module xpb_5_845
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha93ab5f63b7878e531a027b2cf2a0d3d46724fc336972c2d1f28809bcbf440b32de88495cb90a655395928e85d503990fff46fc38d26606767008a01001382c550d5127828fad831c6e386eae33cbef2bc9626cb9be3519620e6848cf052bbe1bfc2576fbff736bc85e5ac8cf919bdd316b6da6e97394de3dfb0cb061c825582;
    5'b00010 : xpb = 1024'ha1c82696b502bd01983ad78e8df9d3291b6e9c5597b6b7e2c07447e1e4e5d45e58888bb2ccface1bd3541289d74262579bceb7a0f799f0831d61d4a3c55490d92d5af041a264b31e7b2d0b332d9db9b4852753feab40761b8c40771f267ad531507d1cb5cf2574eb850b723afa63557cde93d5fade273e9778f21b07b0224499;
    5'b00011 : xpb = 1024'h9a5597372e8d011dfed5876a4cc99914f06ae8e7f8d6439861c00f27fdd76809832892cfce64f5e26d4efc2b51348b1e37a8ff7e620d809ed3c31f468a959eed09e0ce0b1bce8e0b2f768f7b77feb4764db88131ba9d9aa0f79a69b15ca2ee80e137e1fbde53b31a843137e8fbaced26a670d18725152f4b12336b0943c233b0;
    5'b00100 : xpb = 1024'h92e307d7a817453a657037460b995f00c567357a59f5cf4e030bd66e16c8fbb4adc899eccfcf1da90749e5cccb26b3e4d383475bcc8110ba8a2469e94fd6ad00e666abd4953868f7e3c013c3c25faf381649ae64c9fabf2662f45c4392cb07d071f2a741ed81f1498356fd96fcf684d06e4dcd136c031ffeab74bb0ad76222c7;
    5'b00101 : xpb = 1024'h8b70787821a18956cc0ae721ca6924ec9a63820cbb155b03a4579db42fba8f5fd868a109d139456fa144cf6e4518dcab6f5d8f3936f4a0d64085b48c1517bb14c2ec899e0ea243e49809980c0cc0a9f9dedadb97d957e3abce4e4ed5c8f3212002ad6c87fcb02f78827cc344fe401c7a362ac89fb2f110b244b60b0c6b0211de;
    5'b00110 : xpb = 1024'h83fde9189b2bcd7332a596fd8938ead86f5fce9f1c34e6b945a364fa48ac230b0308a826d2a36d363b3fb90fbf0b05720b37d716a16830f1f6e6ff2eda58c9289f726767880c1ed14c531c545721a4bba76c08cae8b5083139a84167ff1b3a6f936831ce0bde6da781a288f2ff89b423fe07c42bf9df0165ddf75b0dfea200f5;
    5'b00111 : xpb = 1024'h7c8b59b914b6118f994046d94808b0c4445c1b317d54726ee6ef2c40619db6b62da8af43d40d94fcd53aa2b138fd2e38a7121ef40bdbc10dad4849d19f99d73c7bf845310175f9be009ca09ca1829f7d6ffd35fdf8122cb6a50233fa354353bf2422f7141b0cabd680c84ea100d34bcdc5e4bfb840ccf2197738ab0f9241f00c;
    5'b01000 : xpb = 1024'h7518ca598e4055abffdaf6b506d876b0195867c3de73fe24883af3867a8f4a615848b660d577bcc36f358c52b2ef56ff42ec66d1764f512963a9947464dae550587e22fa7adfd4aab4e624e4ebe39a3f388e6331076f513c105c268c6b6b6d0eb4ddbc5a2a3aea057fee144f021ce3778dc1bb4487bae2cd1079fb1125e1df23;
    5'b01001 : xpb = 1024'h6da63afa07ca99c86675a690c5a83c9bee54b4563f9389da2986bacc9380de0c82e8bd7dd6e1e48a093075f42ce17fc5dec6aeaee0c2e1451a0adf172a1bf364350400c3f449af97692fa92d36449501011f906416cc75c17bb6191ea193865e459881a0396928347f13d9fd03667b21559eb6d0cea8d380a9bb4b12b981ce3a;
    5'b01010 : xpb = 1024'h6633ab9a8154dde4cd10566c84780287c35100e8a0b3158fcad28212ac7271b7ad88c49ad84c0c50a32b5f95a6d3a88c7aa0f68c4b367160d06c29b9ef5d01781189de8d6db38a841d792d7580a58fc2c9b0bd9726299a46e7100bb0d7bb9fadd65346e6489766637e399fab04b012cb1d7bb25d1596c43442fc9b144d21bd51;
    5'b01011 : xpb = 1024'h5ec11c3afadf220133ab06484347c873984d4d7b01d2a1456c1e4958c5640562d828cbb7d9b634173d26493720c5d153167b3e69b5aa017c86cd745cb49e0f8bee0fbc56e71d6570d1c2b1bdcb068a849241eaca3586becc5269fe430de3b8fd670e0c2c57c5a4927d5f655905f9aa74e558ade95c84b4e7dc3deb15e0c1ac68;
    5'b01100 : xpb = 1024'h574e8cdb7469661d9a45b62402178e5f6d499a0d62f22cfb0d6a109ede55990e02c8d2d4db205bddd72132d89ab7fa19b2558647201d91983d2ebeff79df1d9fca959a206087405d860c3606156785465ad317fd44e3e351bdc3f0d5440bd24cf7c8d17266f3e2c17c852b070743421ead35a975a372a59b757f3b1774619b7f;
    5'b01101 : xpb = 1024'h4fdbfd7bedf3aa3a00e065ffc0e7544b4245e69fc411b8b0aeb5d7e4f7472cb92d68d9f1dc8a83a4711c1c7a14aa22e04e2fce248a9121b3f39009a23f202bb3a71b77e9d9f11b4a3a55ba4e5fc8800823644530544107d7291de3677a33eb9c888396b8762220f07baaf0b5088cd9c87512a501ea60964f0ec08b1908018a96;
    5'b01110 : xpb = 1024'h48696e1c677dee56677b15db7fb71a37174233322531446650019f2b1038c0645808e10eddf4ab6b0b17061b8e9c4ba6ea0a1601f504b1cfa9f15445046139c783a155b3535af636ee9f3e96aa297ac9ebf57263639e2c5c9477d5f9b05c04ec193e5bfe85505f1f7ad0b66309d671723cefa08e314e8702a801db1a9ba179ad;
    5'b01111 : xpb = 1024'h40f6debce1083272ce15c5b73e86e022ec3e7fc48650d01bf14d6671292a540f82a8e82bdf5ed331a511efbd088e746d85e45ddf5f7841eb60529ee7c9a247db6027337cccc4d123a2e8c2def48a758bb4869f9672fb50e1ffd1c88be6841e3ba9f92144947e9d4e79f67c110b20091c04cc9c1a783c77b641432b1c2f4168c4;
    5'b10000 : xpb = 1024'h39844f5d5a92768f34b07592fd56a60ec13acc56e7705bd192992db7421be7baad48ef48e0c8faf83f0cd95e82809d3421bea5bcc9ebd20716b3e98a8ee355ef3cad1146462eac10573247273eeb704d7d17ccc9825875676b2bbb1e1cac378b3ab3e68aa3acdb7d791c41bf0c69a0c5cca997a6bf2a6869da847b1dc2e157db;
    5'b10001 : xpb = 1024'h3211bffdd41cbaab9b4b256ebc266bfa963718e9488fe78733e4f4fd5b0d7b65d7e8f665e23322bed907c2fffc72c5fabd98ed9a345f6222cd15342d542464031932ef0fbf9886fd0b7bcb6f894c6b0f45a8f9fc91b599ecd685adb052d450dacb6eabd0b2db19ac7842076d0db3386f948693330618591d73c5cb1f568146f2;
    5'b10010 : xpb = 1024'h2a9f309e4da6fec801e5d54a7af631e66b33657ba9af733cd530bc4373ff0f110288fd82e39d4a857302aca17664eec1597335779ed2f23e83767ed019657216f5b8ccd9390261e9bfc54fb7d3ad65d10e3a272fa112be7241dfa04288fc6a2a5c297116c20957db7767cd1b0efcd0195c638ebf4d0649d10d071b20ea213609;
    5'b10011 : xpb = 1024'h232ca13ec73142e46880852639c5f7d2402fb20e0acefef2767c83898cf0a2bc2d29049fe507724c0cfd9642f0571787f54d7d550946825a39d7c972dea6802ad23eaaa2b26c3cd6740ed4001e0e6092d6cb5462b06fe2f7ad3992d4bf248379ece4365cd137960a768d92c9104667c324408a4b93f43a84a6486b227dc12520;
    5'b10100 : xpb = 1024'h1bba11df40bb8700cf1b3501f895bdbe152bfea06bee8aa817c84acfa5e2366757c90bbce6719a12a6f87fe46a49404e9127c53273ba1275f0391415a3e78e3eaec4886c2bd617c328585848686f5b549f5c8195bfcd077d18938566f54c9cc97d9efba2e065d43975b35877118fff6cec1d85d7dae22b383f89bb2411611437;
    5'b10101 : xpb = 1024'h1447827fba45cb1d35b5e4ddb76583a9ea284b32cd0e165db9141215bed3ca12826912d9e7dbc1d940f36985e43b69152d020d0fde2da291a69a5eb869289c528b4a6635a53ff2afdca1dc90b2d0561667edaec8cf2a2c0283ed77f92b74b6190e59c0e8ef94126874d91e2512d99716b3fa816421d01bebd8cb0b25a501034e;
    5'b10110 : xpb = 1024'hcd4f32033d00f399c5094b976354995bf2497c52e2da2135a5fd95bd7c55dbdad0919f6e945e99fdaee53275e2d91dbc8dc54ed48a132ad5cfba95b2e69aa6667d043ff1ea9cd9c90eb60d8fd3150d8307edbfbde875087ef476a8b619ccf689f14862efec2509773fee3d314232ec07bd77cf068be0c9f720c5b2738a0f265;
    5'b10111 : xpb = 1024'h56263c0ad5a535602eb449535050f819420e4578f4d2dc8fbaba0a1f0b6f168d7a92113eab0116674e93cc8d81fbaa264b69ccab314c2c9135cf3fdf3aab87a445621c89813a8894534e52147924b99f910092eede4750d5aa15d1d97c4e8b82fcf4b750df08ec67324a981156cc66a43b4787cafabfd530b4dab28cc40e17c;
    5'b11000 : xpb = 1024'hae9d19b6e8d2cc3b348b6c48042f1cbeda93341ac5e459f61ad4213dbcab321c0591a5a9b640b7bbae4265b1356ff43364ab0c8e403b23307a5d7dfef3be3b3f952b3440c10e80bb0c186c0c2acf0a8cb5a62ffa89c7c6a37b87e1aa8817a499ef91a2e4cde7c582f90a560e0e86843d5a6b52eb46e54b36eafe762ee8c336fe;
    5'b11001 : xpb = 1024'ha72a8a57625d10579b261c23c2fee2aaaf8f80ad2703e5abbc1fe883d59cc5c73031acc6b7aadf82483d4f52af621cfa0085546baaaeb34c30bec8a1b8ff495371b1120a3a785ba7c061f0547530054e7e375d2d9924eb28e6e1d43cbe3fbde9804c682add1603b1f8301bbc0fd01be722484e778dd33bea843fc6307c632615;
    5'b11010 : xpb = 1024'h9fb7faf7dbe7547401c0cbff81cea896848bcd3f882371615d6bafc9ee8e59725ad1b3e3b9150748e23838f4295445c09c5f9c4915224367e72013447e4057674e36efd3b3e2369474ab749cbf91001046c88a60a8820fae523bc6cef467d73911072d70ec4441e0f755e16a1119b390ea254a03d4c12c9e1d8116321003152c;
    5'b11011 : xpb = 1024'h98456b9855719890685b7bdb409e6e82598819d1e942fd16feb77710077fed1d8571bb00ba7f2f0f7c332295a3466e873839e4267f95d3839d815de74381657b2abccd9d2d4c118128f4f8e509f1fad20f59b793b7df3433bd95b9612a8ff088a1c1f2b6fb72800ff67ba71812634b3ab20245901baf1d51b6c26633a3a30443;
    5'b11100 : xpb = 1024'h90d2dc38cefbdcaccef62bb6ff6e346e2e8466644a6288cca0033e56207180c8b011c21dbbe956d6162e0c371d38974dd4142c03ea09639f53e2a88a08c2738f0742ab66a6b5ec6ddd3e7d2d5452f593d7eae4c6c73c58b928efabf360b809d8327cb7fd0aa0be3ef5a16cc613ace2e479df411c629d0e055003b6353742f35a;
    5'b11101 : xpb = 1024'h89604cd9488620c93590db92be3dfa5a0380b2f6ab821482414f059c39631473dab1c93abd537e9cb028f5d8972ac0146fee73e1547cf3bb0a43f32cce0381a2e3c88930201fc75a918801759eb3f055a07c11f9d6997d3e94499e8596e02327c3377d4319cefc6df4c7327414f67a8e41bc3ca8a98afeb8e9450636cae2e271;
    5'b11110 : xpb = 1024'h81edbd79c21064e59c2b8b6e7d0dc045d87cff890ca1a037e29acce25254a81f0551d057bebda6634a23df7a111ce8db0bc8bbbebef083d6c0a53dcf93448fb6c04e66f99989a24745d185bde914eb17690d3f2ce5f6a1c3ffa39117cd083c7753f2428928fd3a9cf3ecf8221640123809993834f078ef6c828656385e82d188;
    5'b11111 : xpb = 1024'h7a7b2e1a3b9aa90202c63b4a3bdd8631ad794c1b6dc12bed83e694286b463bca2ff1d774c027ce29e41ec91b8b0f11a1a7a3039c296413f27706887258859dca9cd444c312f37d33fa1b0a063375e5d9319e6c5ff553c6496afd83aa033055c6e4ad07cf382b78cbf312bdd01789a9e1d17633c13766e0201bc7a639f222c09f;
    endcase
end

endmodule

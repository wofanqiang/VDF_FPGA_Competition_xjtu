module xpb_5_980
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3fd27b725d19a509cd2caf1e870be1455749e02de89a94c762f21e7b1550c0c28f3f07210a1261eefa3274fc444c6e3df2297a3979dd15d9e6ddc2ba65d276060ea7cc261f12d605df71e14b79cee6646df5ee4c2d5e25e738919b0fbb7f04b243bdd8fb6d5b7ec4d01f831550840def4443811372be4783a30306aa6c65fbc3;
    5'b00010 : xpb = 1024'h7fa4f6e4ba334a139a595e3d0e17c28aae93c05bd135298ec5e43cf62aa181851e7e0e421424c3ddf464e9f88898dc7be452f472f3ba2bb3cdbb8574cba4ec0c1d4f984c3e25ac0bbee3c296f39dccc8dbebdc985abc4bce7123361f76fe0964877bb1f6dab6fd89a03f062aa1081bde88870226e57c8f0746060d54d8cbf786;
    5'b00011 : xpb = 1024'heca2d01555eba549c80958484c95c7e94679d58e4581ddeaaf9a21b8cef953faa7497ea5410a73e4f391fade98739ef726246c64ae4714203fa08d0f6a4ed60b7a82fc3ada784cc8bbba13fd490eefc55dcd14bfb9444a4f4283f3478526b849c31f8c8974983c0e99ea260f9bc03a47df0a45807ef795aa29998fabc4f8cde;
    5'b00100 : xpb = 1024'h4e9ca873b2785f5e69ad44a30bd53dc3ebb17d86ccf2b2a60debc096a240560239b39f0b5e23092d496b94aa2dd3a82d648bc0ffc4c1871bead7cb8b5c776366c64ffbe9ccba5ad26b2d828b4e5fd560c3d2bf9828f26a8c2cb9da4433d17036dfefd1c404a50285b9be25764a401193c234256b7aadc0de459c9fa528b588a1;
    5'b00101 : xpb = 1024'h8e6f23e60f92046836d9f3c192e11f0942fb5db4b58d476d70dddf11b79116c4c8f2a62c68356b1c439e09a67220166b56b53b393e9e9cf5d1b58e45c249d96cd4f7c80febcd30d84a9f63d6c82ebbc531c8ade456509073654b7553ef5074e923adaabf7200814a89dda88b9ac41f830677a67eed6c0861e89fa64f951b8464;
    5'b00110 : xpb = 1024'h1d945a02aabd74a939012b090992b8fd28cf3ab1c8b03bbd55f3443719df2a7f54e92fd4a8214e7c9e723f5bd30e73dee4c48d8c95c8e28407f411a1ed49dac16f505f875b4f09991777427fa921ddf8abb9a297f7288949e8507e68f0a4d7093863f1912e930781d33d44c1f3780748fbe148b00fdef2b5453331f5789f19bc;
    5'b00111 : xpb = 1024'h5d66d57507d719b3062dda27909e9a4280191adfb14ad084b8e562b22f2feb41e42836f5b233b06b98a4b458175ae21cd6ee07c60fa5f85deed1d45c531c50c77df82bad7a61df9ef6e923cb22f0c45d19af90e42486af3120e21978ac23dbbb7c21ca8c9bee8646a35cc7d743fc15384024c9c3829d3a38e836389fe505157f;
    5'b01000 : xpb = 1024'h9d3950e764f0bebcd35a894617aa7b87d762fb0d99e5654c1bd7812d4480ac0473673e16bc46125a92d729545ba7505ac91781ff89830e37d5af9716b8eec6cd8c9ff7d39974b5a4d65b05169cbfaac187a57f3051e4d5185973b48867a2e06dbfdfa388094a050b737c4aec9480232784684ad6f55b81bc8b393f4a516b1142;
    5'b01001 : xpb = 1024'h2c5e8704001c2efdd581c08d8e5c157bbd36d80aad08599c00ece652a6cebfbeff5dc7befc31f5baedab5f09bc95adce5726d452e0ad53c60bee1a72e3eec82226f88f4b08f68e65a332e3bf7db2ccf5019673e3f2bccdeedc78bd9d68f7428dd495ea59c5dc8b42bcdbe722ed340aed79d1ed0817ce6c0fe7cccaf034eea69a;
    5'b01010 : xpb = 1024'h6c3102765d35d407a2ae6fac1567f6c11480b83895a2ee6363df04cdbc1f80818e9ccee0064457a9e7ddd40600e21c0c49504e8c5a8a699ff2cbdd2d49c13e2835a05b712809646b82a4c50af781b3596f8c6230201af3d6150a58ad247647401853c35533380a078cfb6a383db818dcbe156e1b8a8cb3938acfd19aa154a25d;
    5'b01011 : xpb = 1024'hac037de8ba4f79116fdb1eca9c73d8066bca98667e3d832ac6d12348d17041441ddbd6011056b998e2104902452e8a4a3b79c8c5d4677f79d9a99fe7af93b42e44482797471c3a716216a656715099bddd82507c4d7919bd4d9bf3bcdff54bf25c119c50a09388cc5d1aed4d8e3c26cc0258ef2efd4afb172dd2d8450dba9e20;
    5'b01100 : xpb = 1024'h3b28b405557ae95272025612132571fa519e75639160777aabe6886e33be54fea9d25fa950429cf93ce47eb7a61ce7bdc9891b192b91c5080fe82343da93b582dea0bf0eb69e13322eee84ff5243bbf15773452fee511293d0a0fcd1e149ae1270c7e3225d260f03a67a8983e6f00e91f7c291601fbde56a8a6663eaf13e3378;
    5'b01101 : xpb = 1024'h7afb2f77b2948e5c3f2f05309a31533fa8e8559179fb0c420ed8a6e9490f15c1391166ca5a54fee83716f3b3ea6955fbbbb29552a56edae1f6c5e5fe40662b88ed488b34d5b0e9380e60664acc12a255c569337c1baf387b093297e19cc8b2c4b485bc1dca818dc8769a0c9937741c813c061273927c2cee2d696a955da42f3b;
    5'b01110 : xpb = 1024'ha2065944dbffe9d41563c7810e2ed338ebc328e8d1e0091f3ee0c0eab5d297bc507f0729a40e24891eb29694b57b36f49c1e7a5fc9920702d04695a6b662cdd87a122ac4532c1f8db3844f3ad05c4893f5a282fbc8731518c37a0f69e1d14e4c93c02ef871413ffbff9a8cf90280447316fb4a4b4ef174189fcf63b4127c493;
    5'b01111 : xpb = 1024'h49f2e106aad9a3a70e82eb9697eece78e60612bc75b8955956e02a89c0adea3e5446f793a45344378c1d9e658fa421ad3beb61df7676364a13e22c14d138a2e39648eed2644597febaaa263f26d4aaedad50167be9e55738c4c93c06599c19970cf9dbeaf46f92c490192be4e0ac123675b335b827ad5ec52cfffce5ad8dc056;
    5'b10000 : xpb = 1024'h89c55c7907f348b0dbaf9ab51efaafbe3d4ff2ea5e532a20b9d24904d5feab00e385feb4ae65a62686501361d3f08feb2e14dc18f0534c23fabfeecf370b18e9a4f0baf883586e049a1c078aa0a391521b4604c817437d1ffd5ad716151b1e4950b7b4e661cb11896038aefa31302025b9f6b6cb9a6ba648d003039019f3bc19;
    5'b10001 : xpb = 1024'h18ea9295a31eb8f1ddd6d1fc95ac49b22323cfe771761e709ee7ae2a384cbebb6f7c885cee518986e124491734deed5ebc242e6c477d91b230fe722b620b1a3e3f49526ff2da46c566f3e6338196b3859536f97bb81b75f6805fe02b166f8069656dfbb81e5d97c0a9984b3089e407ebaf6058fcbcde909c2c968f35fd775171;
    5'b10010 : xpb = 1024'h58bd0e0800385dfbab03811b1cb82af77a6db0155a10b33801d9cca54d9d7f7dfebb8f7df863eb75db56be13792b5b9cae4da8a5c15aa78c17dc34e5c7dd90444df11e9611ed1ccb4665c77efb6599ea032ce7c7e5799bddb8f17b3ad1ee851ba92bd4b38bb9168579b7ce45da6815daf3a3da102f9cd81fcf9995e069dd4d34;
    5'b10011 : xpb = 1024'h988f897a5d52030578303039a3c40c3cd1b7904342ab47ff64cbeb2062ee40408dfa969f02764d64d589330fbd77c9daa07722df3b37bd65feb9f7a02db0064a5c98eabc30fff2d125d7a8ca7534804e7122d61412d7c1c4f183164a8d6d89cdece9adaef914954a49d7515b2aec23ca37e75b23a25b1fa3729c9c8ad64348f7;
    5'b10100 : xpb = 1024'h27b4bf96f87d73467a5767811a75a630b78b6d4055ce3c4f49e15045c53c53fb19f12047426230c5305d68c51e66274e2e867532926202f434f87afc58b0079ef6f18233a081cb91f2af87735627a281eb13cac7b3afba9b74881f5f8ec1ebee019ff480b5a71b819336ed9183a00b902d50fd54c4ce09f6cf302830b9c6de4f;
    5'b10101 : xpb = 1024'h67873b09559718504784169fa18187760ed54d6e3e68d116acd36ec0da8d14bda93027684c7492b42a8fddc162b2958c20afef6c0c3f18ce1bd63db6be827da505994e59bf94a197d22168becff688e65909b913e10de082ad19ba6f4a40f0a0455dcd7c23029a46635670a6d424197f71947e68378c517a72332edb262cda12;
    5'b10110 : xpb = 1024'ha759b67bb2b0bd5a14b0c5be288d68bb661f2d9c270365de0fc58d3befddd580386f2e895686f4a324c252bda6ff03ca12d969a5861c2ea802b400712454f3ab14411a7fdea7779db1934a0a49c56f4ac6ffa7600e6c0669e5ab557f05bff552891ba677905e190b3375f3bc24a8276eb5d7ff7baa4a98fe153635859292d5d5;
    5'b10111 : xpb = 1024'h367eec984ddc2d9b16d7fd059f3f02af4bf30a993a265a2df4daf261522be93ac465b8319672d8037f96887307ed613da0e8bbf8dd46743638f283cd4f54f4ffae99b1f74e29505e7e6b28b32ab8917e40f09c13af43ff4068b05e94071457729dd1ed494cf09f427cd58ff27d5c0f34ab41a1acccbd835171c9c12b76166b2d;
    5'b11000 : xpb = 1024'h7651680aaaf5d2a4e404ac24264ae3f4a33ceac722c0eef557cd10dc677ca9fd53a4bf52a08539f279c8fd6f4c39cf7b9312363257238a101fd04687b5276b05bd417e1d6d3c26645ddd09fea48777e2aee68a5fdca22527a141f9a3c2935c24e18fc644ba4c1e074cf51307cde01d23ef8522c03f7bcad514ccc7d5e27c66f0;
    5'b11001 : xpb = 1024'h5769e27462142e5e62be36b9cfc7de88910c7c435e3e3453ce27601c9cabdb7df9b48fae0711d52d49d3324ad282cef21218885ae4dcf9e560ec9e3e0276c5a579a1594dcbdff252ab4e8a7857a9a1628d77f137d7a1dfe244702b8c3e7be44f6460d1676dea43e9654af3e269404e9e4eec4f161eeb5287160537bc5fffc48;
    5'b11010 : xpb = 1024'h45491999a33ae7efb358928a24085f2de05aa7f21e7e780c9fd4947cdf1b7e7a6eda501bea837f41cecfa820f1749b2d134b02bf282ae5783cec8c9e45f9e2606641e1bafbd0d52b0a26c9f2ff49807a96cd6d5faad843e55cd89dc87f66c2f73a03e611e43a230366743253771812d929324604d4acfcac14635a263265f80b;
    5'b11011 : xpb = 1024'h851b950c00548cf9808541a8ab14407337a4882007190cd402c6b2f7f46c3f3cfe19573cf495e130c9021d1d35c1096b05747cf8a207fb5223ca4f58abcc586674e9ade11ae3ab30e998ab3e791866df04c35babd83669cc956a38d83ae5c7a97dc1bf0d5195a1c83693b568c79c20c86d75c718476b442fb76660d09ecbf3ce;
    5'b11100 : xpb = 1024'h1440cb289b7ffd3a82ac78f021c5da671d78651d1a3c0123e7dc181d56ba52f78a0fe0e53481c49123d652d296af66de9383cf4bf93240e05a08d2b4d6cc59bb0f4245588a6583f1b67089e75a0b89127eb4505f790e62a3186f41ed3c3a29c9927805df0e2827ff7ff3519f2050088e62df694969de2e8313f9ec76824f8926;
    5'b11101 : xpb = 1024'h5413469af899a2444fd9280ea8d1bbac74c2454b02d695eb4ace36986c0b13ba194ee8063e9426801e08c7cedafbd51c85ad4985730f56ba40e6956f3c9ecfc11dea117ea97859f795e26b32d3da6f76ecaa3eaba66c888a5100dcfcf7b92e7bd635deda7b83a6c45012d4b470d4167da722ea5cdc9c7606b6fcf320eeb584e9;
    5'b11110 : xpb = 1024'h93e5c20d55b3474e1d05d72d2fdd9cf1cc0c2578eb712ab2adc05513815bd47ca88def2748a6886f183b3ccb1f48435a77d6c3beecec6c9427c45829a27145c72c91dda4c88b2ffd75544c7e4da955db5aa02cf7d3caae718992780cb338332e19f3b7d5e8df2589203257c9c158246ceb666b704f5abd8a59fff9cb5b1b80ac;
    5'b11111 : xpb = 1024'h230af829f0deb78f1f2d0e74a68f36e5b1e00275fe941f0292d5ba38e3a9e837348478cf88926bcf730f72808036a0ce05e616124416b2225e02db85cd71471bc6ea751c380d08be422c2b272e9c780ed49121ab74a2a7480c978121b48c954e2ea9fea7a571abc06991f4001a0c0c32e0d00da171cda7ddb69385713e9f1604;
    endcase
end

endmodule

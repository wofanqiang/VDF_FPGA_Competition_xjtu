module xpb_5_555
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'he59d5dba7328ca6d55533cd683c69f306d3a3c9f6749500fe28ec7755eef669efc0d8a007d61ed2eca344be02ab34a2dd74fc45c115df9aec4c181197521bba6f26434f0fa4a11d4f786c7bc11246c54243d5e5866ddcacd0b78664e1e7fd317917af65226af66b094c0f70a4d60000199f2b751c18d6d6d34da131126f9deb;
    5'b00010 : xpb = 1024'h1cb3abb74e65194daaaa679ad078d3e60da74793ece92a01fc51d8eeabddecd3df81b1400fac3da5d946897c05566945bae9f88b822bbf35d89830232ea43774de4c869e1f49423a9ef0d8f782248d8a8487abcb0cdbb959a16f0cc9c3cffa62f22f5eca44d5ecd612981ee149ac0000333e56ea3831adada69b426224df3bd6;
    5'b00011 : xpb = 1024'h2b0d8192f597a5f47fff9b6838b53dd9147aeb5de35dbf02fa7ac56601cce33dcf4289e017825c78c5e9ce3a08019de8985ef4d143419ed0c4e44834c5f6532f4d72c9ed2eede357ee6945734336d44fc6cb81b0934996067226932ea5b7f7946b470e2f6740e3411be42e51ee8200004cdd825f544a848479e8e393374ed9c1;
    5'b00100 : xpb = 1024'h3967576e9cca329b5554cf35a0f1a7cc1b4e8f27d9d25403f8a3b1dd57bbd9a7bf0362801f587b4bb28d12f80aacd28b75d3f11704577e6bb13060465d486ee9bc990d3c3e9284753de1b1ef04491b15090f579619b772b342de1993879ff4c5e45ebd9489abd9ac25303dc293580000667cadd470635b5b4d3684c449be77ac;
    5'b00101 : xpb = 1024'h47c12d4a43fcbf422aaa0303092e11bf222232f1d046e904f6cc9e54adaad011aec43b20272e9a1e9f3057b60d58072e5348ed5cc56d5e069d7c7857f49a8aa42bbf508b4e3725928d5a1e6ac55b61da4b532d7ba0254f6013959ff86987f1f75d766cf9ac16d0172e7c4d33382e0000801bd9498c7c3232208425f55c2e1597;
    5'b00110 : xpb = 1024'h561b0325eb2f4be8ffff36d0716a7bb228f5d6bbc6bb7e05f4f58acc0399c67b9e8513c02f04b8f18bd39c7410033bd130bde9a286833da189c890698beca65e9ae593da5ddbc6afdcd28ae6866da89f8d97036126932c0ce44d265d4b6fef28d68e1c5ece81c68237c85ca3dd04000099bb04bea8950908f3d1c7266e9db382;
    5'b00111 : xpb = 1024'h6474d9019261d88fd5546a9dd9a6e5a52fc97a85bd301306f31e77435988bce58e45ec6036dad7c47876e13212ae70740e32e5e847991d3c7614a87b233ec2190a0bd7296d8067cd2c4af762477fef64cfdad946ad0108b9b504acc22d57ec5a4fa5cbc3f0ecbced41146c1481da0000b35a3033c4addfdfc71f6857810d516d;
    5'b01000 : xpb = 1024'h72ceaedd39946536aaa99e6b41e34f98369d1e4fb3a4a807f14763baaf77b34f7e06c5003eb0f697651a25f01559a516eba7e22e08aefcd76260c08cba90ddd379321a787d2508ea7bc363de0892362a121eaf2c336ee56685bc33270f3fe98bc8bd7b291357b3584a607b8526b00000ccf95ba8e0c6b6b69a6d0988937cef58;
    5'b01001 : xpb = 1024'h812884b8e0c6f1dd7ffed238aa1fb98b3d70c219aa193d08ef7050320566a9b96dc79da04687156a51bd6aae1804d9b9c91cde73c9c4dc724eacd89e51e2f98de8585dc78cc9aa07cb3bd059c9a47cef54628511b9dcc2135673b98bf127e6bd41d52a8e35c2a9c353ac8af5cb860000e698871dfcdf8d8d6dbaaab9a5ec8d43;
    5'b01010 : xpb = 1024'h8f825a9487f97e8455540606125c237e444465e3a08dd209ed993ca95b55a0235d8876404e5d343d3e60af6c1ab00e5ca691dab98adabc0d3af8f0afe9351548577ea1169c6e4b251ab43cd58ab6c3b496a65af7404a9ec0272b3ff0d30fe3eebaecd9f3582da02e5cf89a66705c00010037b29318f8646441084beab85c2b2e;
    5'b01011 : xpb = 1024'h9ddc30702f2c0b2b2aa939d37a988d714b1809ad9702670aebc22920b144968d4d494ee0563353102b03f42a1d5b42ff8406d6ff4bf09ba8274508c180873102c6a4e465ac12ec426a2ca9514bc90a79d8ea30dcc6b87b6cf7e2c655b4f7e120340489587a9896996644a9d71532000119d6de0835113b3b1455ed1bcacbc919;
    5'b01100 : xpb = 1024'hac36064bd65e97d1fffe6da0e2d4f76451ebad778d76fc0be9eb159807338cf73d0a27805e0971e317a738e8200677a2617bd3450d067b43139120d317d94cbd35cb27b4bbb78d5fb9a515cd0cdb513f1b2e06c24d265819c89a4cba96dfde51ad1c38bd9d038d046f90b947ba0800013376097d512a1211e7a38e4cdd3b6704;
    5'b01101 : xpb = 1024'h9e296d1bba2efb00a4e29973ab71a05e7494e10ae73f0956a3748b9aa1fd659298282a79bb9122764ec3e5f3f539b7adad6a7a4ab698a924f3df9867458f3c630a236551bcb3137f6837fa63511d3d3696ce30f470e07b5e3c54124be9d38f0f72c55f90ea58ae1f21ce1d9670dd9d7fe3b56101cf78bb87481b47966c89e84;
    5'b01110 : xpb = 1024'h183c6cad62d57c56dfa35d64a2f383f8ee1cf1daa4e8859668603531000eccc319435b47a38f30fa518f831d41fed01db84ba3ea6c7f6a2d3b8a11980bab0f809fc879a42b6fd25545fbec21f6241a98abb0b8f4cd7be462b47cc789a08536227044055e3110814cfb68f14a0be3d9d817da81853910628f47cf55aa79383c6f;
    5'b01111 : xpb = 1024'h269642890a0808fdb4f891320b2fedebf4f095a49b5d1a97668921a855fdc32d090433e7ab654fcd3e32c7db44aa04c095c0a0302d9549c827d629a9a2fd2b3b0eeebcf33b1473729574589db736615dedf48eda53e9c10f85344dee826d3353e95bb4c3537b77b804b500bab0b9d9d83179acfa552939661b1cf6db8ba7da5a;
    5'b10000 : xpb = 1024'h34f01864b13a95a48a4dc4ff736c57defbc4396e91d1af9864b20e1fabecb996f8c50c87b33b6ea02ad60c994755396373359c75eeab2963142241bb3a4f46f57e1500424ab9148fe4ecc5197848a823303864bfda579dbc55ebd453645530856273642875e66e230e01102b558fd9d84b18d86f7142103cee6a980c9e177845;
    5'b10001 : xpb = 1024'h4349ee40586d224b5fa2f8ccdba8c1d20297dd388846449962dafa9701dbb000e885e527bb118d73177951574a006e0650aa98bbafc108fe006e59ccd1a162afed3b43915a5db5ad34653195395aeee8727c3aa560c57a6926a35ab8463d2db6db8b138d9851648e174d1f9bfa65d9d864b803e48d5ae713c1b8393db0871630;
    5'b10010 : xpb = 1024'h51a3c41bff9faef234f82c9a43e52bc5096b81027ebad99a6103e70e57caa66ad846bdc7c2e7ac46041c96154caba2a92e1f950170d6e898ecba71de68f37e6a5c6186e06a0256ca83dd9e10fa6d35adb4c0108ae7335715f75ae11d28252ae854a2c2f2babc5af920992f0c9f3bd9d87e572f59a973bdea9505da6ec2f6b41b;
    5'b10011 : xpb = 1024'h5ffd99f7a6d23b990a4d6067ac2195b8103f24cc752f6e9b5f2cd385adb99cd4c8079667cabdcb18f0bfdad34f56d74c0b94914731ecc833d90689f000459a24cb87ca2f79a6f7e7d3560a8cbb7f7c72f703e6706da133c2c81267820a0d2819cdba7257dd27516429e53e7d4411d9d897f65acec58c94c168537b9fd5665206;
    5'b10100 : xpb = 1024'h6e576fd34e04c83fdfa29435145dffab1712c8966ba4039c5d55bffd03a8933eb7c86f07d293e9ebdd631f9152020beee9098d8cf302a7cec552a2019797b5df3aae0d7e894b990522ce77087c91c3383947bc55f40f106f98c9ede6ebf5254b46d221bcff9247cf33314dede8e7d9d8b1958643e1a56b983ba11cd0e7d5eff1;
    5'b10101 : xpb = 1024'h7cb145aef53754e6b4f7c8027c9a699e1de66c606218989d5b7eac74599789a8a78947a7da6a08beca06644f54ad4091c67e89d2b4188769b19eba132ee9d199a9d450cd98f03a227246e3843da409fd7b8b923b7a7ced1c6981744bcddd227cbfe9d12221fd3e3a3c7d5d5e8dbdd9d8cb34b1b8fdbe426f0eeebe01fa458ddc;
    5'b10110 : xpb = 1024'h8b0b1b8a9c69e18d8a4cfbcfe4d6d39124ba102a588d2d9e59a798ebaf868012974a2047e2402791b6a9a90d57587534a3f38618752e67049dead224c63bed5418fa941ca894db3fc1bf4ffffeb650c2bdcf682100eac9c93a38fab0afc51fae39018087446834a545c96ccf3293d9d8e4d3dd2e19d71945e23c5f330cb52bc7;
    5'b10111 : xpb = 1024'h9964f166439c6e345fa22f9d4d133d842b8db3f44f01c29f57d085630575767c870af8e7ea164664a34cedcb5a03a9d78168825e3644469f8a36ea365d8e090e8820d76bb8397c5d1137bc7bbfc8978800133e068758a6760af0811591ad1cdfb2192fec66d32b104f157c3fd769d9d8fe7308a335eff01cb58a00641f24c9b2;
    5'b11000 : xpb = 1024'ha7bec741eacefadb34f7636ab54fa777326157be457657a055f971da5b646ce676cbd187f1ec65378ff032895caede7a5edd7ea3f75a263a76830247f4e024c8f7471abac7de1d7a60b028f780dade4d425713ec0dc68322dba8077a73951a112b30df51893e217b58618bb07c3fd9d9181234185208c6f388d7a1953194679d;
    5'b11001 : xpb = 1024'h56b57c7d01352b93f471f610d31ca18c7bef85766734c29d645a4fbfe50b64863442caf2f9c057bdd3538007bfc0252d838530395bd3589b22fdafb515fcbd1f21e295b27f1c1529d8e92d0a91160e19095f03907ae32bef6d2fbe49b5274b07540fc8cfae01f58daedb4422945b3afe2d780ab1dd6409a15b5c7c1bb219f1d;
    5'b11010 : xpb = 1024'h13c52da37745df60149c532e756e340bce929c215ce7e12ad46e9173543facb25305054f3772244ec9d87cbe7ea736f5b5ad4f4956d315249e7bf30ce8b1e78c61446caa3796626fed06ff4c6a23a7a6d2d9c61e8e1c0f6bc78a82497d3a71e1ee58abf21d4b15c3e439c3b2ce1bb3affc76ac2039ef1770e90368f2cd913d08;
    5'b11011 : xpb = 1024'h221f037f1e786c06e9f186fbddaa9dfed5663feb535c762bd2977deaaa2ea31c42c5ddef3f484321b67bc17c81526b9893224b8f17e8f4bf8ac80b1e80040346d06aaff9473b038d3c7f6bc82b35ee6c151d9c041489ec18984208ae5f226f1367705b573fb60c2eed85d32372f1b3b01615d7955607ee47bc510a23e000daf3;
    5'b11100 : xpb = 1024'h3078d95ac5aaf8adbf46bac945e707f1dc39e3b549d10b2cd0c06a62001d99863286b68f471e61f4a31f063a83fda03b709747d4d8fed45a7714233017561f013f90f34856dfa4aa8bf7d843ec483531576171e99af7c8c568f98f13410a6c44e0880abc62210299f6d1e29417c7b3b02fb5030a7220c51e8f9eab54f27078de;
    5'b11101 : xpb = 1024'h3ed2af366cdd8554949bee96ae2371e4e30d877f4045a02dcee956d9560c8ff022478f2f4ef480c78fc24af886a8d4de4e0c441a9a14b3f563603b41aea83abbaeb73697668445c7db7044bfad5a7bf699a547cf2165a57239b1157822f26976599fba21848bf905001df204bc9db3b049542e7f8e399bf562ec4c8604e016c9;
    5'b11110 : xpb = 1024'h4d2c8512141011fb69f12264165fdbd7e9e12b4936ba352ecd124350abfb865a120867cf56ca9f9a7c658fb6895409812b8140605b2a93904fac535345fa56761ddd79e67628e6e52ae8b13b6e6cc2bbdbe91db4a7d3821f0a689bdd04da66a7d2b76986a6f6ef70096a01756173b3b062f359f4aa5272cc3639edb7174fb4b4;
    5'b11111 : xpb = 1024'h5b865aedbb429ea23f4656317e9c45caf0b4cf132d2eca2fcb3b2fc801ea7cc401c9406f5ea0be6d6908d4748bff3e2408f63ca61c40732b3bf86b64dd4c72308d03bd3585cd88027a611db72f7f09811e2cf39a2e415ecbdb202241e6c263d94bcf18ebc961e5db12b610e60649b3b07c928569c66b49a309878ee829bf529f;
    endcase
end

endmodule

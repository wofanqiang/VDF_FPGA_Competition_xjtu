module xpb_5_520
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7347068c9ac8a597921e9cc3999fdb57ee39d7ee19c26492e8164fcf5e9232ca3b8ad909209191fe1ddca3f1111f6b4b60a755b4152ce2e2944c952854f407aab9367280ad353e590d9f35adf31596101a0fef4a01c5dbcb002834cfc4d2c435c3577d78ab388bbe0d1efefccdbfc1ae1a78b7152b02d50a53c41524090ae715;
    5'b00010 : xpb = 1024'h35e0c7c373a316665937c1b022e56f5e6afdacab5e0d28ae524fe6490a21b88c73cd349976fca56d9c5b089b3ee0c5cc5d34838207a6f57977f9eaf26f159aa3fe1db052aad97f6d08a468b94d4f67ef401ae4fb77058a854ac3d7a4cf7ae5d957a768c7a5a81eee937e171aa3af5d32e6178f4805ba4ce46118af43893367bf;
    5'b00011 : xpb = 1024'ha927ce500e6bbbfdeb565e73bc854ab65937849977cf8d413a66361868b3eb56af580da2978e376bba37ac8c50003117bddbd9361cd3d85c0c46801ac409a24eb75422d3580ebdc616439e674064fdff5a2ad44578cb66504aec0c74944daa0f1afee64050e0aaaca09d1617716f1ee10090465d30bd21eeb4dcc467923e4ed4;
    5'b00100 : xpb = 1024'h6bc18f86e7462cccb26f836045cadebcd5fb5956bc1a515ca49fcc9214437118e79a6932edf94adb38b611367dc18b98ba6907040f4deaf2eff3d5e4de2b3547fc3b60a555b2feda1148d1729a9ecfde8035c9f6ee0b150a9587af499ef5cbb2af4ed18f4b503ddd26fc2e35475eba65cc2f1e900b7499c8c2315e871266cf7e;
    5'b00101 : xpb = 1024'h2e5b50bdc0209d9b7988a84ccf1072c352bf2e14006515780ed9630bbfd2f6db1fdcc4c344645e4ab73475e0ab82e619b6f634d201c7fd89d3a12baef84cc84141229e7753573fee0c4e047df4d8a1bda640bfa8634ac3c4e023521ea99ded56439ebcde45bfd10dad5b46531d4e55ea97cdf6c2e62c11a2cf85f8a6928f5028;
    5'b00110 : xpb = 1024'ha1a2574a5ae943330ba7451068b04e1b40f906021a277a0af6efb2db1e6529a55b679dcc64f5f048d51119d1bca25165179d8a8616f4e06c67edc0d74d40cfebfa5910f8008c7e4719ed3a2be7ee37cdc050aef265109f8fe04b86ee6e70b18c06f63a56f0f85ccbba7a454feb0e1798b246add8112ee6ad234a0dca9b9a373d;
    5'b00111 : xpb = 1024'h643c188133c3b401d2c069fcf1f5e221bdbcdabf5e723e2661294954c9f4af6793a9f95cbb6103b8538f7e7bea63abe6142ab854096ef3034b9b16a1676262e53f404ec9fe30bf5b14f26d37422809ace65ba4a3da504e4a2ae729c37918d32f9b4625a5eb67effc40d95d6dc0fdb31d7de5860aebe65e87309ea7ea1bc2b7e7;
    5'b01000 : xpb = 1024'h26d5d9b80c9e24d099d98ee97b3b76283a80af7ca2bd0241cb62dfce75843529cbec54ed11cc1727d20de3261825066710b7e621fbe9059a2f486c6b8183f5de84278c9bfbd5006f0ff7a0429c61db8c0c669a554f8ffd047582cc9883c0f4d32f9610f4e5d7832cc738758b96ed4ea249845e3dc69dd6613df342099beb3891;
    5'b01001 : xpb = 1024'h9a1ce044a766ca682bf82bad14db518028ba876abc7f66d4b3792f9dd41667f407772df6325da925efea8717294471b2715f3bd61115e87cc3950193d677fd893d5dff1ca90a3ec81d96d5f08f77719c2676899f5155d8cf75ab01684893b908f2ed8e6d91100eead457748864ad105063fd1552f1a0ab6b91b7572da4f61fa6;
    5'b01010 : xpb = 1024'h5cb6a17b80413b36f31150999e20e586a57e5c2800ca2af01db2c6177fa5edb63fb9898688c8bc956e68ebc15705cc336dec69a4038ffb13a742575df099908282453ceea6ae7fdc189c08fbe9b1437b4c817f50c6958789c046a43d533bdaac873d79bc8b7fa21b5ab68ca63a9cabd52f9bed85cc5823459f0bf14d251ea050;
    5'b01011 : xpb = 1024'h1f5062b2591bac05ba2a75862766798d224230e54514ef0b87ec5c912b35737877fbe516df33d004ece7506b84c726b46a799771f60a0daa8aefad280abb237bc72c7ac0a452c0f013a13c0743eb155a728c75023bd536440ae247125de3fc501b8d650b85ef354be115a4c4108c4759fb3ac5b8a70f9b1fac608b6ca54720fa;
    5'b01100 : xpb = 1024'h9297693ef3e4519d4c491249c10654e5107c08d35ed7539e7002ac6089c7a642b386be1fffc562030ac3f45c95e691ffcb20ed260b36f08d1f3c42505faf2b268062ed415187ff49214071b53700ab6a8c9c644c3d9b120f0b0a7be222b6c085dee4e2843127c109ee34a3c0de4c090815b37ccdd212702a0024a090ae52080f;
    5'b01101 : xpb = 1024'h55312a75ccbec26c136237364a4be8eb8d3fdd90a32217b9da3c42da35572c04ebc919b05630757289425906c3a7ec80c7ae1af3fdb1032402e9981a79d0be1fc54a2b134f2c405d1c45a4c0913a7d49b2a759fdb2dac0c955a61eb72d5ee2297334cdd32b97543a7493bbdeb43ba48ce1525500acc9e8040d793ab02e7a88b9;
    5'b01110 : xpb = 1024'h17caebaca599333ada7b5c22d3917cf20a03b24de76cdbd54475d953e0e6b1c7240b7540ac9b88e207c0bdb0f1694701c43b48c1f02b15bae696ede493f251190a3168e54cd08171174ad7cbeb744f28d8b24faf281a6f83a041c18c380703cd0784b9222606e76afaf2d3fc8a2b4011acf12d3387815fde1acdd4cfaea30963;
    5'b01111 : xpb = 1024'h8b11f2394061d8d26c99f8e66d315849f83d8a3c012f40682c8c29233f78e4915f964e49cd2d1ae0259d61a20288b24d24e29e760557f89d7ae3830ce8e658c3c367db65fa05bfca24ea0d79de89e538f2c23ef929e04b4ea069f65bfcd9c802cadc369ad13f73290811d2f957eb01bfc769e448b28434e86e91e9f3b7adf078;
    5'b10000 : xpb = 1024'h4dabb370193c49a133b31dd2f676ec5075015ef9457a048396c5bf9ceb086a5397d8a9da23982e4fa41bc64c304a0cce216fcc43f7d20b345e90d8d70307ebbd084f1937f7aa00de1fef408538c3b71818cd34aa9f1ffa08eb0599310781e9a65f2c21e9cbaf06598e70eb172dda9d449308bc7b8d3bacc27be6841337d67122;
    5'b10001 : xpb = 1024'h104574a6f216ba6ffacc42bf7fbc8056f1c533b689c4c89f00ff56169697f015d01b056a7a0341bf229a2af65e0b674f1dfcfa11ea4c1dcb423e2ea11d297eb64d365709f54e41f21af4739092fd88f73ed82a5c145fa8c335a13c06122a0b49f37c0d38c61e998a14d0033503ca38c95ea794ae67f3249c893b1e32b7fef1cc;
    5'b10010 : xpb = 1024'h838c7b338cdf60078ceadf83195c5baedfff0ba4a3872d31e915a5e5f52a22e00ba5de739a94d3bd4076cee76f2ad29a7ea44fc5ff7900add68ac3c9721d8661066cc98aa283804b2893a93e86131f0758e819a61625848e35c970d5d6fccf7fb6d38ab17157254821ef0231d189fa7779204bc392f5f9a6dcff3356c109d8e1;
    5'b10011 : xpb = 1024'h46263c6a65b9d0d65404046fa2a1efb55cc2e061e7d1f14d534f3c5fa0b9a8a243e83a03f0ffe72cbef533919cec2d1b7b317d93f1f31344ba3819938c3f195a4b54075ca027c15f2398dc49e04cf0e67ef30f578b653348806513aae1a4f1234b2376006bc6b878a84e1a4fa77995fc44bf23f66dad7180ea53cd764132598b;
    5'b10100 : xpb = 1024'h8bffda13e9441a51b1d295c2be783bbd986b51f2c1cb568bd88d2d94c492e647c2a9594476afa9c3d73983bcaad879c77beab61e46d25db9de56f5da660ac53903b452e9dcc02731e9e0f553a86c2c5a4fe050900a4e202cb00b67fec4d12c6df73614f66364ba92ead326d7d693181105dfc294864e95af7a86795c15ada35;
    5'b10101 : xpb = 1024'h7c07042dd95ce73cad3bc61fc5875f13c7c08d0d45df19fba59f22a8aadb612eb7b56e9d67fc8c9a5b503c2cdbccf2e7d8660115f99a08be32320485fb54b3fe4971b7af4b0140cc2c3d45032d9c58d5bf0df453026abdcdcb28eb4fb11fd6fca2cadec8116ed7673bcc316a4b28f32f2ad6b33e7367be654b6c7cb9ca65c14a;
    5'b10110 : xpb = 1024'h3ea0c564b237580b7454eb0c4eccf31a448461ca8a29de170fd8b922566ae6f0eff7ca2dbe67a009d9cea0d7098e4d68d4f32ee3ec141b5515df5a50157646f78e58f58148a581e02742780e87d62ab4e518ea0477aa6c8815c48e24bbc7f8a0371aca170bde6a97c22b498821188eb3f6758b714e1f363f58c116d94a8e41f4;
    5'b10111 : xpb = 1024'h13a869b8b11c8da3b6e0ff8d8128720c1483687ce74a2327a124f9c01fa6cb3283a25be14d2b379584d0581374fa7e9d1805cb1de8e2debf98cb01a2f97d9f0d34033534649c2f42247ab19e20ffc940b23dfb5ecea1b42606030f9c6701a43cb6ab566064dfdc8488a61a5f7082a38c21463a428d6ae196615b0f8cab6c29e;
    5'b11000 : xpb = 1024'h74818d2825da6e71cd8cacbc71b26278af820e75e83706c562289f6b608c9f7d63c4fec7356445777629a972486f13353227b265f3bb10ce8dd94542848be19b8c76a5d3f37f014d2fe6e0c7d52592a42533ceffeeaff70d608865c98b42de798ec232deb186898655a960a2c4c7ebe6dc8d1ab953d98323b9d9c61cd3c1a9b3;
    5'b11001 : xpb = 1024'h371b4e5efeb4df4094a5d1a8faf7f67f2c45e3332c81cae0cc6235e50c1c253f9c075a578bcf58e6f4a80e1c76306db62eb4e033e635236571869b0c9ead7494d15de3a5f12342612aec13d32f5f64834b3ec4b163efa5c7ab24089e95eb001d23121e2dabf61cb6dc0878c09ab7876ba82bf2ec2e90fafdc72e603c53ea2a5d;
    5'b11010 : xpb = 1024'haa6254eb997d84d826c46e6c9497d1d71a7fbb2146442f73b47885b46aae5809d7923360ac60eae51284b20d874fd9018f5c35e7fb62064805d33034f3a17c3f8a9456269e5880ba388b49812274fa93654eb3fb65b58192ab4c3d6e5abdc452e6699ba6572ea874e92777bd68774919c2a4aa015993d0081af275605cf51172;
    5'b11011 : xpb = 1024'h6cfc16227257f5a6eddd93591ddd65dd97438fde8a8ef38f1eb21c2e163dddcc0fd48ef102cbfe54910316b7b51133828be963b5eddc18dee98085ff0dc30f38cf7b93f89bfcc1ce33907c8c7caecc728b59a9acdaf5304cf5e7e0436565e5f67ab986f5519e3ba56f868fdb3e66e49e8e438234344b47e228470f7fdd1d921c;
    5'b11100 : xpb = 1024'h2f95d7594b326675b4f6b845a722f9e41407649bced9b7aa88ebb2a7c1cd638e4816ea81593711c40f817b61e2d28e0388769183e0562b75cd2ddbc927e4a2321462d1ca99a102e22e95af97d6e89e51b1649f5e5034df0740838318700e079a0f0972444c0dced5f5e5a7f91456802359e25a670f02bfbc359ba99f5d4612c6;
    5'b11101 : xpb = 1024'ha2dcdde5e5fb0c0d4715550940c2d53c02413c89e89c1c3d71020277205f965883a1c38a79c8a3c22d5e1f52f3f1f94ee91de737f5830e58617a70f17cd8a9dccd99444b46d6413b3c34e545c9fe3461cb748ea851fabad240abb7e834e0cbcfd260efbcf7465a940304a6f5e21641d1745b117c3a0594c6895fbec36650f9db;
    5'b11110 : xpb = 1024'h65769f1cbed57cdc0e2e79f5ca0869427f0511472ce6e058db3b98f0cbef1c1abbe41f1ad033b731abdc83fd21b353cfe5ab1505e7fd20ef4527c6bb96fa3cd61280821d447a824f373a185124380640f17f8459c73a698c8b475abd3f88ed7366b0db0bf1b5edc48963bf13b805dd563ff9e9af14bd0ca096b458e2e6797a85;
    5'b11111 : xpb = 1024'h2810605397afedaad5479ee2534dfd48fbc8e6047131a47445752f6a777ea1dcf4267aab269ecaa12a5ae8a74f74ae50e23842d3da77338628d51c85b11bcfcf5767bfef421ec363323f4b5c7e71d820178a7a0b3c7a1846d5e2fd924a310f16fb00c65aec2580f50fc2d7318df578db0b98c1e1ef74847aa408f30266a1fb2f;
    endcase
end

endmodule

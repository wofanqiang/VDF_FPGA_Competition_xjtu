module xpb_lut
(
    input logic [16:0] flag[9],
    output logic [1023:0] xpb[27]
);


    always_comb begin
        case(flag[0][5:0])
            6'd0: xpb[0] = 1024'd0;
            6'd1: xpb[0] = 1024'd11454525384925565851030981610095525237135330708387242952012541691402042621681452271329361390848837013342580092128660640518086664281015165389545664756208179145692376357234569976119398356929700888829356807609634068219935781898714912970744491649724942101312076670393225331813467936943319227481230073598687002816;
            6'd2: xpb[0] = 1024'd22909050769851131702061963220191050474270661416774485904025083382804085243362904542658722781697674026685160184257321281036173328562030330779091329512416358291384752714469139952238796713859401777658713615219268136439871563797429825941488983299449884202624153340786450663626935873886638454962460147197374005632;
            6'd3: xpb[0] = 1024'd34363576154776697553092944830286575711405992125161728856037625074206127865044356813988084172546511040027740276385981921554259992843045496168636994268624537437077129071703709928358195070789102666488070422828902204659807345696144738912233474949174826303936230011179675995440403810829957682443690220796061008448;
            6'd4: xpb[0] = 1024'd45818101539702263404123926440382100948541322833548971808050166765608170486725809085317445563395348053370320368514642562072346657124060661558182659024832716582769505428938279904477593427718803555317427230438536272879743127594859651882977966598899768405248306681572901327253871747773276909924920294394748011264;
            6'd5: xpb[0] = 1024'd57272626924627829255154908050477626185676653541936214760062708457010213108407261356646806954244185066712900460643303202590433321405075826947728323781040895728461881786172849880596991784648504444146784038048170341099678909493574564853722458248624710506560383351966126659067339684716596137406150367993435014080;
            6'd6: xpb[0] = 1024'd68727152309553395106185889660573151422811984250323457712075250148412255730088713627976168345093022080055480552771963843108519985686090992337273988537249074874154258143407419856716390141578205332976140845657804409319614691392289477824466949898349652607872460022359351990880807621659915364887380441592122016896;
            6'd7: xpb[0] = 1024'd80181677694478960957216871270668676659947314958710700664087791839814298351770165899305529735941859093398060644900624483626606649967106157726819653293457254019846634500641989832835788498507906221805497653267438477539550473291004390795211441548074594709184536692752577322694275558603234592368610515190809019712;
            6'd8: xpb[0] = 1024'd91636203079404526808247852880764201897082645667097943616100333531216340973451618170634891126790696106740640737029285124144693314248121323116365318049665433165539010857876559808955186855437607110634854460877072545759486255189719303765955933197799536810496613363145802654507743495546553819849840588789496022528;
            6'd9: xpb[0] = 1024'd103090728464330092659278834490859727134217976375485186568112875222618383595133070441964252517639533120083220829157945764662779978529136488505910982805873612311231387215111129785074585212367307999464211268486706613979422037088434216736700424847524478911808690033539027986321211432489873047331070662388183025344;
            6'd10: xpb[0] = 1024'd114545253849255658510309816100955252371353307083872429520125416914020426216814522713293613908488370133425800921286606405180866642810151653895456647562081791456923763572345699761193983569297008888293568076096340682199357818987149129707444916497249421013120766703932253318134679369433192274812300735986870028160;
            6'd11: xpb[0] = 1024'd1933083550056482962541870306236344863790210666523988344006103540445573501186836074607904084679532837325231605957773611119889466249946484729842187301958929668925465360009052399683142734709504055812727275318734904054932750664967269713210838463744913847612939960208420619841619232447878485174840982959962546645;
            6'd12: xpb[0] = 1024'd13387608934982048813572851916331870100925541374911231296018645231847616122868288345937265475528369850667811698086434251637976130530961650119387852058167108814617841717243622375802541091639204944642084082928368972274868532563682182683955330113469855948925016630601645951655087169391197712656071056558649549461;
            6'd13: xpb[0] = 1024'd24842134319907614664603833526427395338060872083298474248031186923249658744549740617266626866377206864010391790215094892156062794811976815508933516814375287960310218074478192351921939448568905833471440890538003040494804314462397095654699821763194798050237093300994871283468555106334516940137301130157336552277;
            6'd14: xpb[0] = 1024'd36296659704833180515634815136522920575196202791685717200043728614651701366231192888595988257226043877352971882343755532674149459092991980898479181570583467106002594431712762328041337805498606722300797698147637108714740096361112008625444313412919740151549169971388096615282023043277836167618531203756023555093;
            6'd15: xpb[0] = 1024'd47751185089758746366665796746618445812331533500072960152056270306053743987912645159925349648074880890695551974472416173192236123374007146288024846326791646251694970788947332304160736162428307611130154505757271176934675878259826921596188805062644682252861246641781321947095490980221155395099761277354710557909;
            6'd16: xpb[0] = 1024'd59205710474684312217696778356713971049466864208460203104068811997455786609594097431254711038923717904038132066601076813710322787655022311677570511082999825397387347146181902280280134519358008499959511313366905245154611660158541834566933296712369624354173323312174547278908958917164474622580991350953397560725;
            6'd17: xpb[0] = 1024'd70660235859609878068727759966809496286602194916847446056081353688857829231275549702584072429772554917380712158729737454228409451936037477067116175839208004543079723503416472256399532876287709388788868120976539313374547442057256747537677788362094566455485399982567772610722426854107793850062221424552084563541;
            6'd18: xpb[0] = 1024'd82114761244535443919758741576905021523737525625234689008093895380259871852957001973913433820621391930723292250858398094746496116217052642456661840595416183688772099860651042232518931233217410277618224928586173381594483223955971660508422280011819508556797476652960997942535894791051113077543451498150771566357;
            6'd19: xpb[0] = 1024'd93569286629461009770789723187000546760872856333621931960106437071661914474638454245242795211470228944065872342987058735264582780498067807846207505351624362834464476217885612208638329590147111166447581736195807449814419005854686573479166771661544450658109553323354223274349362727994432305024681571749458569173;
            6'd20: xpb[0] = 1024'd105023812014386575621820704797096071998008187042009174912118978763063957096319906516572156602319065957408452435115719375782669444779082973235753170107832541980156852575120182184757727947076812055276938543805441518034354787753401486449911263311269392759421629993747448606162830664937751532505911645348145571989;
            6'd21: xpb[0] = 1024'd116478337399312141472851686407191597235143517750396417864131520454465999718001358787901517993167902970751032527244380016300756109060098138625298834864040721125849228932354752160877126304006512944106295351415075586254290569652116399420655754960994334860733706664140673937976298601881070759987141718946832574805;
            6'd22: xpb[0] = 1024'd3866167100112965925083740612472689727580421333047976688012207080891147002373672149215808169359065674650463211915547222239778932499892969459684374603917859337850930720018104799366285469419008111625454550637469808109865501329934539426421676927489827695225879920416841239683238464895756970349681965919925093290;
            6'd23: xpb[0] = 1024'd15320692485038531776114722222568214964715752041435219640024748772293189624055124420545169560207902687993043304044207862757865596780908134849230039360126038483543307077252674775485683826348709000454811358247103876329801283228649452397166168577214769796537956590810066571496706401839076197830912039518612096106;
            6'd24: xpb[0] = 1024'd26775217869964097627145703832663740201851082749822462592037290463695232245736576691874530951056739701335623396172868503275952261061923300238775704116334217629235683434487244751605082183278409889284168165856737944549737065127364365367910660226939711897850033261203291903310174338782395425312142113117299098922;
            6'd25: xpb[0] = 1024'd38229743254889663478176685442759265438986413458209705544049832155097274867418028963203892341905576714678203488301529143794038925342938465628321368872542396774928059791721814727724480540208110778113524973466372012769672847026079278338655151876664653999162109931596517235123642275725714652793372186715986101738;
            6'd26: xpb[0] = 1024'd49684268639815229329207667052854790676121744166596948496062373846499317489099481234533253732754413728020783580430189784312125589623953631017867033628750575920620436148956384703843878897137811666942881781076006080989608628924794191309399643526389596100474186601989742566937110212669033880274602260314673104554;
            6'd27: xpb[0] = 1024'd61138794024740795180238648662950315913257074874984191448074915537901360110780933505862615123603250741363363672558850424830212253904968796407412698384958755066312812506190954679963277254067512555772238588685640149209544410823509104280144135176114538201786263272382967898750578149612353107755832333913360107370;
            6'd28: xpb[0] = 1024'd72593319409666361031269630273045841150392405583371434400087457229303402732462385777191976514452087754705943764687511065348298918185983961796958363141166934212005188863425524656082675610997213444601595396295274217429480192722224017250888626825839480303098339942776193230564046086555672335237062407512047110186;
            6'd29: xpb[0] = 1024'd84047844794591926882300611883141366387527736291758677352099998920705445354143838048521337905300924768048523856816171705866385582466999127186504027897375113357697565220660094632202073967926914333430952203904908285649415974620938930221633118475564422404410416613169418562377514023498991562718292481110734113002;
            6'd30: xpb[0] = 1024'd95502370179517492733331593493236891624663067000145920304112540612107487975825290319850699296149761781391103948944832346384472246748014292576049692653583292503389941577894664608321472324856615222260309011514542353869351756519653843192377610125289364505722493283562643894190981960442310790199522554709421115818;
            6'd31: xpb[0] = 1024'd106956895564443058584362575103332416861798397708533163256125082303509530597506742591180060686998598794733684041073492986902558911029029457965595357409791471649082317935129234584440870681786316111089665819124176422089287538418368756163122101775014306607034569953955869226004449897385630017680752628308108118634;
            6'd32: xpb[0] = 1024'd118411420949368624435393556713427942098933728416920406208137623994911573219188194862509422077847435808076264133202153627420645575310044623355141022165999650794774694292363804560560269038716016999919022626733810490309223320317083669133866593424739248708346646624349094557817917834328949245161982701906795121450;
            6'd33: xpb[0] = 1024'd5799250650169448887625610918709034591370631999571965032018310621336720503560508223823712254038598511975694817873320833359668398749839454189526561905876789006776396080027157199049428204128512167438181825956204712164798251994901809139632515391234741542838819880625261859524857697343635455524522948879887639935;
            6'd34: xpb[0] = 1024'd17253776035095014738656592528804559828505962707959207984030852312738763125241960495153073644887435525318274910001981473877755063030854619579072226662084968152468772437261727175168826561058213056267538633565838780384734033893616722110377007040959683644150896551018487191338325634286954683005753022478574642751;
            6'd35: xpb[0] = 1024'd28708301420020580589687574138900085065641293416346450936043394004140805746923412766482435035736272538660855002130642114395841727311869784968617891418293147298161148794496297151288224917987913945096895441175472848604669815792331635081121498690684625745462973221411712523151793571230273910486983096077261645567;
            6'd36: xpb[0] = 1024'd40162826804946146440718555748995610302776624124733693888055935695542848368604865037811796426585109552003435094259302754913928391592884950358163556174501326443853525151730867127407623274917614833926252248785106916824605597691046548051865990340409567846775049891804937854965261508173593137968213169675948648383;
            6'd37: xpb[0] = 1024'd51617352189871712291749537359091135539911954833120936840068477386944890990286317309141157817433946565346015186387963395432015055873900115747709220930709505589545901508965437103527021631847315722755609056394740985044541379589761461022610481990134509948087126562198163186778729445116912365449443243274635651199;
            6'd38: xpb[0] = 1024'd63071877574797278142780518969186660777047285541508179792081019078346933611967769580470519208282783578688595278516624035950101720154915281137254885686917684735238277866200007079646419988777016611584965864004375053264477161488476373993354973639859452049399203232591388518592197382060231592930673316873322654015;
            6'd39: xpb[0] = 1024'd74526402959722843993811500579282186014182616249895422744093560769748976233649221851799880599131620592031175370645284676468188384435930446526800550443125863880930654223434577055765818345706717500414322671614009121484412943387191286964099465289584394150711279902984613850405665319003550820411903390472009656831;
            6'd40: xpb[0] = 1024'd85980928344648409844842482189377711251317946958282665696106102461151018855330674123129241989980457605373755462773945316986275048716945611916346215199334043026623030580669147031885216702636418389243679479223643189704348725285906199934843956939309336252023356573377839182219133255946870047893133464070696659647;
            6'd41: xpb[0] = 1024'd97435453729573975695873463799473236488453277666669908648118644152553061477012126394458603380829294618716335554902605957504361712997960777305891879955542222172315406937903717008004615059566119278073036286833277257924284507184621112905588448589034278353335433243771064514032601192890189275374363537669383662463;
            6'd42: xpb[0] = 1024'd108889979114499541546904445409568761725588608375057151600131185843955104098693578665787964771678131632058915647031266598022448377278975942695437544711750401318007783295138286984124013416495820166902393094442911326144220289083336025876332940238759220454647509914164289845846069129833508502855593611268070665279;
            6'd43: xpb[0] = 1024'd120344504499425107397935427019664286962723939083444394552143727535357146720375030937117326162526968645401495739159927238540535041559991108084983209467958580463700159652372856960243411773425521055731749902052545394364156070982050938847077431888484162555959586584557515177659537066776827730336823684866757668095;
            6'd44: xpb[0] = 1024'd7732334200225931850167481224945379455160842666095953376024414161782294004747344298431616338718131349300926423831094444479557864999785938919368749207835718675701861440036209598732570938838016223250909101274939616219731002659869078852843353854979655390451759840833682479366476929791513940699363931839850186580;
            6'd45: xpb[0] = 1024'd19186859585151497701198462835040904692296173374483196328036955853184336626428796569760977729566968362643506515959755084997644529280801104308914413964043897821394237797270779574851969295767717112080265908884573684439666784558583991823587845504704597491763836511226907811179944866734833168180594005438537189396;
            6'd46: xpb[0] = 1024'd30641384970077063552229444445136429929431504082870439280049497544586379248110248841090339120415805375986086608088415725515731193561816269698460078720252076967086614154505349550971367652697418000909622716494207752659602566457298904794332337154429539593075913181620133142993412803678152395661824079037224192212;
            6'd47: xpb[0] = 1024'd42095910355002629403260426055231955166566834791257682232062039235988421869791701112419700511264642389328666700217076366033817857842831435088005743476460256112778990511739919527090766009627118889738979524103841820879538348356013817765076828804154481694387989852013358474806880740621471623143054152635911195028;
            6'd48: xpb[0] = 1024'd53550435739928195254291407665327480403702165499644925184074580927390464491473153383749061902113479402671246792345737006551904522123846600477551408232668435258471366868974489503210164366556819778568336331713475889099474130254728730735821320453879423795700066522406583806620348677564790850624284226234598197844;
            6'd49: xpb[0] = 1024'd65004961124853761105322389275423005640837496208032168136087122618792507113154605655078423292962316416013826884474397647069991186404861765867097072988876614404163743226209059479329562723486520667397693139323109957319409912153443643706565812103604365897012143192799809138433816614508110078105514299833285200660;
            6'd50: xpb[0] = 1024'd76459486509779326956353370885518530877972826916419411088099664310194549734836057926407784683811153429356406976603058287588077850685876931256642737745084793549856119583443629455448961080416221556227049946932744025539345694052158556677310303753329307998324219863193034470247284551451429305586744373431972203476;
            6'd51: xpb[0] = 1024'd87914011894704892807384352495614056115108157624806654040112206001596592356517510197737146074659990442698987068731718928106164514966892096646188402501292972695548495940678199431568359437345922445056406754542378093759281475950873469648054795403054250099636296533586259802060752488394748533067974447030659206292;
            6'd52: xpb[0] = 1024'd99368537279630458658415334105709581352243488333193896992124747692998634978198962469066507465508827456041567160860379568624251179247907262035734067257501151841240872297912769407687757794275623333885763562152012161979217257849588382618799287052779192200948373203979485133874220425338067760549204520629346209108;
            6'd53: xpb[0] = 1024'd110823062664556024509446315715805106589378819041581139944137289384400677599880414740395868856357664469384147252989040209142337843528922427425279732013709330986933248655147339383807156151205324222715120369761646230199153039748303295589543778702504134302260449874372710465687688362281386988030434594228033211924;
            6'd54: xpb[0] = 1024'd122277588049481590360477297325900631826514149749968382896149831075802720221561867011725230247206501482726727345117700849660424507809937592814825396769917510132625625012381909359926554508135025111544477177371280298419088821647018208560288270352229076403572526544765935797501156299224706215511664667826720214740;
            6'd55: xpb[0] = 1024'd9665417750282414812709351531181724318951053332619941720030517702227867505934180373039520423397664186626158029788868055599447331249732423649210936509794648344627326800045261998415713673547520279063636376593674520274663753324836348566054192318724569238064699801042103099208096162239392425874204914799812733225;
            6'd56: xpb[0] = 1024'd21119943135207980663740333141277249556086384041007184672043059393629910127615632644368881814246501199968738121917528696117533995530747589038756601266002827490319703157279831974535112030477221167892993184203308588494599535223551261536798683968449511339376776471435328431021564099182711653355434988398499736041;
            6'd57: xpb[0] = 1024'd32574468520133546514771314751372774793221714749394427624055601085031952749297084915698243205095338213311318214046189336635620659811762754428302266022211006636012079514514401950654510387406922056722349991812942656714535317122266174507543175618174453440688853141828553762835032036126030880836665061997186738857;
            6'd58: xpb[0] = 1024'd44028993905059112365802296361468300030357045457781670576068142776433995370978537187027604595944175226653898306174849977153707324092777919817847930778419185781704455871748971926773908744336622945551706799422576724934471099020981087478287667267899395542000929812221779094648499973069350108317895135595873741673;
            6'd59: xpb[0] = 1024'd55483519289984678216833277971563825267492376166168913528080684467836037992659989458356965986793012239996478398303510617671793988373793085207393595534627364927396832228983541902893307101266323834381063607032210793154406880919696000449032158917624337643313006482615004426461967910012669335799125209194560744489;
            6'd60: xpb[0] = 1024'd66938044674910244067864259581659350504627706874556156480093226159238080614341441729686327377641849253339058490432171258189880652654808250596939260290835544073089208586218111879012705458196024723210420414641844861374342662818410913419776650567349279744625083153008229758275435846955988563280355282793247747305;
            6'd61: xpb[0] = 1024'd78392570059835809918895241191754875741763037582943399432105767850640123236022894001015688768490686266681638582560831898707967316935823415986484925047043723218781584943452681855132103815125725612039777222251478929594278444717125826390521142217074221845937159823401455090088903783899307790761585356391934750121;
            6'd62: xpb[0] = 1024'd89847095444761375769926222801850400978898368291330642384118309542042165857704346272345050159339523280024218674689492539226053981216838581376030589803251902364473961300687251831251502172055426500869134029861112997814214226615840739361265633866799163947249236493794680421902371720842627018242815429990621752937;
            6'd63: xpb[0] = 1024'd101301620829686941620957204411945926216033698999717885336130851233444208479385798543674411550188360293366798766818153179744140645497853746765576254559460081510166337657921821807370900528985127389698490837470747066034150008514555652332010125516524106048561313164187905753715839657785946245724045503589308755753;
        endcase
    end

    always_comb begin
        case(flag[0][11:6])
            6'd0: xpb[1] = 1024'd0;
            6'd1: xpb[1] = 1024'd112756146214612507471988186022041451453169029708105128288143392924846251101067250815003772941037197306709378858946813820262227309778868912155121919315668260655858714015156391783490298885914828278527847645080381134254085790413270565302754617166249048149873389834581131085529307594729265473205275577187995758569;
            6'd2: xpb[1] = 1024'd101445596745100273545177444639268470161639632290474572448154930784715606864825362719992474667416720303975608310436134205945390778716517489755083713615005480378026753460741566229350358580312450835745497681773522422143810730605644357640530664649268647032926876255045204140952087115529897929291861327750397032807;
            6'd3: xpb[1] = 1024'd90135047275588039618366703256495488870110234872844016608166468644584962628583474624981176393796243301241837761925454591628554247654166067355045507914342700100194792906326740675210418274710073392963147718466663710033535670798018149978306712132288245915980362675509277196374866636330530385378447078312798307045;
            6'd4: xpb[1] = 1024'd78824497806075805691555961873722507578580837455213460768178006504454318392341586529969878120175766298508067213414774977311717716591814644955007302213679919822362832351911915121070477969107695950180797755159804997923260610990391942316082759615307844799033849095973350251797646157131162841465032828875199581283;
            6'd5: xpb[1] = 1024'd67513948336563571764745220490949526287051440037582904928189544364323674156099698434958579846555289295774296664904095362994881185529463222554969096513017139544530871797497089566930537663505318507398447791852946285812985551182765734653858807098327443682087335516437423307220425677931795297551618579437600855521;
            6'd6: xpb[1] = 1024'd56203398867051337837934479108176544995522042619952349088201082224193029919857810339947281572934812293040526116393415748678044654467111800154930890812354359266698911243082264012790597357902941064616097828546087573702710491375139526991634854581347042565140821936901496362643205198732427753638204330000002129759;
            6'd7: xpb[1] = 1024'd44892849397539103911123737725403563703992645202321793248212620084062385683615922244935983299314335290306755567882736134361208123404760377754892685111691578988866950688667438458650657052300563621833747865239228861592435431567513319329410902064366641448194308357365569418065984719533060209724790080562403403997;
            6'd8: xpb[1] = 1024'd33582299928026869984312996342630582412463247784691237408224157943931741447374034149924685025693858287572985019372056520044371592342408955354854479411028798711034990134252612904510716746698186179051397901932370149482160371759887111667186949547386240331247794777829642473488764240333692665811375831124804678235;
            6'd9: xpb[1] = 1024'd22271750458514636057502254959857601120933850367060681568235695803801097211132146054913386752073381284839214470861376905727535061280057532954816273710366018433203029579837787350370776441095808736269047938625511437371885311952260904004962997030405839214301281198293715528911543761134325121897961581687205952473;
            6'd10: xpb[1] = 1024'd10961200989002402130691513577084619829404452949430125728247233663670452974890257959902088478452904282105443922350697291410698530217706110554778068009703238155371069025422961796230836135493431293486697975318652725261610252144634696342739044513425438097354767618757788584334323281934957577984547332249607226711;
            6'd11: xpb[1] = 1024'd123717347203614909602679699599126071282573482657535254016390626588516704075957508774905861419490101588814822781297511111672925839996575022709899987325371498811229783040579353579721135021408259572014545620399033859515696042557905261645493661679674486247228157453338919669863630876664223051189822909437602985280;
            6'd12: xpb[1] = 1024'd112406797734102675675868958216353089991044085239904698176402164448386059839715620679894563145869624586081052232786831497356089308934223600309861781624708718533397822486164528025581194715805882129232195657092175147405420982750279053983269709162694085130281643873802992725286410397464855507276408660000004259518;
            6'd13: xpb[1] = 1024'd101096248264590441749058216833580108699514687822274142336413702308255415603473732584883264872249147583347281684276151883039252777871872177909823575924045938255565861931749702471441254410203504686449845693785316435295145922942652846321045756645713684013335130294267065780709189918265487963362994410562405533756;
            6'd14: xpb[1] = 1024'd89785698795078207822247475450807127407985290404643586496425240168124771367231844489871966598628670580613511135765472268722416246809520755509785370223383157977733901377334876917301314104601127243667495730478457723184870863135026638658821804128733282896388616714731138836131969439066120419449580161124806807994;
            6'd15: xpb[1] = 1024'd78475149325565973895436734068034146116455892987013030656436778027994127130989956394860668325008193577879740587254792654405579715747169333109747164522720377699901940822920051363161373798998749800885145767171599011074595803327400430996597851611752881779442103135195211891554748959866752875536165911687208082232;
            6'd16: xpb[1] = 1024'd67164599856053739968625992685261164824926495569382474816448315887863482894748068299849370051387716575145970038744113040088743184684817910709708958822057597422069980268505225809021433493396372358102795803864740298964320743519774223334373899094772480662495589555659284946977528480667385331622751662249609356470;
            6'd17: xpb[1] = 1024'd55854050386541506041815251302488183533397098151751918976459853747732838658506180204838071777767239572412199490233433425771906653622466488309670753121394817144238019714090400254881493187793994915320445840557881586854045683712148015672149946577792079545549075976123358002400308001468017787709337412812010630708;
            6'd18: xpb[1] = 1024'd44543500917029272115004509919715202241867700734121363136471391607602194422264292109826773504146762569678428941722753811455070122560115065909632547420732036866406059159675574700741552882191617472538095877251022874743770623904521808009925994060811678428602562396587431057823087522268650243795923163374411904946;
            6'd19: xpb[1] = 1024'd33232951447517038188193768536942220950338303316490807296482929467471550186022404014815475230526285566944658393212074197138233591497763643509594341720069256588574098605260749146601612576589240029755745913944164162633495564096895600347702041543831277311656048817051504113245867043069282699882508913936813179184;
            6'd20: xpb[1] = 1024'd21922401978004804261383027154169239658808905898860251456494467327340905949780515919804176956905808564210887844701394582821397060435412221109556136019406476310742138050845923592461672270986862586973395950637305450523220504289269392685478089026850876194709535237515577168668646563869915155969094664499214453422;
            6'd21: xpb[1] = 1024'd10611852508492570334572285771396258367279508481229695616506005187210261713538627824792878683285331561477117296190714968504560529373060798709517930318743696032910177496431098038321731965384485144191045987330446738412945444481643185023254136509870475077763021657979650224091426084670547612055680415061615727660;
            6'd22: xpb[1] = 1024'd123367998723105077806560471793437709820448538189334823904649398112056512814605878639796651624322528868186496155137528788766787839151929710864639849634411956688768891511587489821812030851299313422718893632410827872667031234894913750326008753676119523227636411492560781309620733679399813085260955992249611486229;
            6'd23: xpb[1] = 1024'd112057449253592843879749730410664728528919140771704268064660935971925868578363990544785353350702051865452725606626849174449951308089578288464601643933749176410936930957172664267672090545696935979936543669103969160556756175087287542663784801159139122110689897913024854365043513200200445541347541742812012760467;
            6'd24: xpb[1] = 1024'd100746899784080609952938989027891747237389743354073712224672473831795224342122102449774055077081574862718955058116169560133114777027226866064563438233086396133104970402757838713532150240094558537154193705797110448446481115279661335001560848642158720993743384333488927420466292721001077997434127493374414034705;
            6'd25: xpb[1] = 1024'd89436350314568376026128247645118765945860345936443156384684011691664580105880214354762756803461097859985184509605489945816278245964875443664525232532423615855273009848343013159392209934492181094371843742490251736336206055472035127339336896125178319876796870753953000475889072241801710453520713243936815308943;
            6'd26: xpb[1] = 1024'd78125800845056142099317506262345784654330948518812600544695549551533935869638326259751458529840620857251413961094810331499441714902524021264487026831760835577441049293928187605252269628889803651589493779183393024225930995664408919677112943608197918759850357174417073531311851762602342909607298994499216583181;
            6'd27: xpb[1] = 1024'd66815251375543908172506764879572803362801551101182044704707087411403291633396438164740160256220143854517643412584130717182605183840172598864448821131098055299609088739513362051112329323287426208807143815876534312115655935856782712014888991091217517642903843594881146586734631283402975365693884745061617857419;
            6'd28: xpb[1] = 1024'd55504701906031674245696023496799822071272153683551488864718625271272647397154550069728861982599666851783872864073451102865768652777821176464410615430435275021777128185098536496972389017685048766024793852569675600005380876049156504352665038574237116525957330015345219642157410804203607821780470495624019131657;
            6'd29: xpb[1] = 1024'd44194152436519440318885282114026840779742756265920933024730163131142003160912661974717563708979189849050102315562771488548932121715469754064372409729772494743945167630683710942832448712082671323242443889262816887895105816241530296690441086057256715409010816435809292697580190325004240277867056246186420405895;
            6'd30: xpb[1] = 1024'd32883602967007206392074540731253859488213358848290377184741700991011358924670773879706265435358712846316331767052091874232095590653118331664334204029109714466113207076268885388692508406480293880460093925955958175784830756433904089028217133540276314292064302856273365753002969845804872733953641996748821680133;
            6'd31: xpb[1] = 1024'd21573053497494972465263799348480878196683961430659821344753238850880714688428885784694967161738235843582561218541412259915259059590766909264295998328446934188281246521854059834552568100877916437677743962649099463674555696626277881365993181023295913175117789276737438808425749366605505190040227747311222954371;
            6'd32: xpb[1] = 1024'd10262504027982738538453057965707896905154564013029265504764776710750070452186997689683668888117758840848790670030732645598422528528415486864257792627784153910449285967439234280412627795275538994895393999342240751564280636818651673703769228506315512058171275697201511863848528887406137646126813497873624228609;
            6'd33: xpb[1] = 1024'd123018650242595246010441243987749348358323593721134393792908169635596321553254248504687441829154956147558169528977546465860649838307284399019379711943452414566307999982595626063902926681190367273423241644422621885818366427231922239006523845672564560208044665531782642949377836482135403119332089075061619987178;
            6'd34: xpb[1] = 1024'd111708100773083012083630502604976367066794196303503837952919707495465677317012360409676143555534479144824398980466866851543813307244932976619341506242789634288476039428180800509762986375587989830640891681115763173708091367424296031344299893155584159091098151952246716004800616002936035575418674825624021261416;
            6'd35: xpb[1] = 1024'd100397551303570778156819761222203385775264798885873282112931245355335033080770472314664845281914002142090628431956187237226976776182581554219303300542126854010644078873765974955623046069985612387858541717808904461597816307616669823682075940638603757974151638372710789060223395523736668031505260576186422535654;
            6'd36: xpb[1] = 1024'd89087001834058544230009019839430404483735401468242726272942783215204388844528584219653547008293525139356857883445507622910140245120230131819265094841464073732812118319351149401483105764383234945076191754502045749487541247809043616019851988121623356857205124793174862115646175044537300487591846326748823809892;
            6'd37: xpb[1] = 1024'd77776452364546310303198278456657423192206004050612170432954321075073744608286696124642248734673048136623087334934828008593303714057878709419226889140801293454980157764936323847343165458780857502293841791195187037377266188001417408357628035604642955740258611213638935171068954565337932943678432077311225084130;
            6'd38: xpb[1] = 1024'd66465902895034076376387537073884441900676606632981614592965858934943100372044808029630950461052571133889316786424148394276467182995527287019188683440138513177148197210521498293203225153178480059511491827888328325266991128193791200695404083087662554623312097634103008226491734086138565399765017827873626358368;
            6'd39: xpb[1] = 1024'd55155353425521842449576795691111460609147209215351058752977396794812456135802919934619652187432094131155546237913468779959630651933175864619150477739475732899316236656106672739063284847576102616729141864581469613156716068386164993033180130570682153506365584054567081281914513606939197855851603578436027632606;
            6'd40: xpb[1] = 1024'd43844803956009608522766054308338479317617811797720502912988934654681811899561031839608353913811617128421775689402789165642794120870824442219112272038812952621484276101691847184923344541973725173946791901274610901046441008578538785370956178053701752389419070475031154337337293127739830311938189328998428906844;
            6'd41: xpb[1] = 1024'd32534254486497374595955312925565498026088414380089947073000472514551167663319143744597055640191140125688005140892109551325957589808473019819074066338150172343652315547277021630783404236371347731164441937967752188936165948770912577708732225536721351272472556895495227392760072648540462768024775079560830181082;
            6'd42: xpb[1] = 1024'd21223705016985140669144571542792516734559016962459391233012010374420523427077255649585757366570663122954234592381429937009121058746121597419035860637487392065820354992862196076643463930768970288382091974660893476825890888963286370046508273019740950155526043315959300448182852169341095224111360830123231455320;
            6'd43: xpb[1] = 1024'd9913155547472906742333830160019535443029619544828835393023548234289879190835367554574459092950186120220464043870750322692284527683770175018997654936824611787988394438447370522503523625166592845599742011354034764715615829155660162384284320502760549038579529736423373503605631690141727680197946580685632729558;
            6'd44: xpb[1] = 1024'd122669301762085414214322016182060986896198649252933963681166941159136130291902618369578232033987383426929842902817564142954511837462639087174119574252492872443847108453603762305993822511081421124127589656434415898969701619568930727687038937669009597188452919571004504589134939284870993153403222157873628488127;
            6'd45: xpb[1] = 1024'd111358752292573180287511274799288005604669251835303407841178479019005486055660730274566933760366906424196072354306884528637675306400287664774081368551830092166015147899188936751853882205479043681345239693127557186859426559761304520024814985152029196071506405991468577644557718805671625609489807908436029762365;
            6'd46: xpb[1] = 1024'd100048202823060946360700533416515024313139854417672852001190016878874841819418842179555635486746429421462301805796204914320838775337936242374043162851167311888183187344774111197713941899876666238562889729820698474749151499953678312362591032635048794954559892411932650699980498326472258065576393658998431036603;
            6'd47: xpb[1] = 1024'd88737653353548712433889792033742043021610457000042296161201554738744197583176954084544337213125952418728531257285525300004002244275584819974004957150504531610351226790359285643574001594274288795780539766513839762638876440146052104700367080118068393837613378832396723755403277847272890521662979409560832310841;
            6'd48: xpb[1] = 1024'd77427103884036478507079050650969061730081059582411740321213092598613553346935065989533038939505475415994760708774845685687165713213233397573966751449841751332519266235944460089434061288671911352998189803206981050528601380338425897038143127601087992720666865252860796810826057368073522977749565160123233585079;
            6'd49: xpb[1] = 1024'd66116554414524244580268309268196080438551662164781184481224630458482909110693177894521740665884998413260990160264166071370329182150881975173928545749178971054687305681529634535294120983069533910215839839900122338418326320530799689375919175084107591603720351673324869866248836888874155433836150910685634859317;
            6'd50: xpb[1] = 1024'd54806004945012010653457567885423099147022264747150628641236168318352264874451289799510442392264521410527219611753486457053492651088530552773890340048516190776855345127114808981154180677467156467433489876593263626308051260723173481713695222567127190486773838093788942921671616409674787889922736661248036133555;
            6'd51: xpb[1] = 1024'd43495455475499776726646826502650117855492867329520072801247706178221620638209401704499144118644044407793449063242806842736656120026179130373852134347853410499023384572699983427014240371864779024651139913286404914197776200915547274051471270050146789369827324514253015977094395930475420346009322411810437407793;
            6'd52: xpb[1] = 1024'd32184906005987542799836085119877136563963469911889516961259244038090976401967513609487845845023567405059678514732127228419819588963827707973813928647190630221191424018285157872874300066262401581868789949979546202087501141107921066389247317533166388252880810934717089032517175451276052802095908162372838682031;
            6'd53: xpb[1] = 1024'd20874356536475308873025343737104155272434072494258961121270781897960332165725625514476547571403090402325907966221447614102983057901476285573775722946527849943359463463870332318734359760660024139086439986672687489977226081300294858727023365016185987135934297355181162087939954972076685258182493912935239956269;
            6'd54: xpb[1] = 1024'd9563807066963074946214602354331173980904675076628405281282319757829687929483737419465249297782613399592137417710767999786146526839124863173737517245865069665527502909455506764594419455057646696304090023365828777866951021492668651064799412499205586018987783775645235143362734492877317714269079663497641230507;
            6'd55: xpb[1] = 1024'd122319953281575582418202788376372625434073704784733533569425712682675939030550988234469022238819810706301516276657581820048373836617993775328859436561533330321386216924611898548084718340972474974831937668446209912121036811905939216367554029665454634168861173610226366228892042087606583187474355240685636989076;
            6'd56: xpb[1] = 1024'd111009403812063348491392046993599644142544307367102977729437250542545294794309100139457723965199333703567745728146902205731537305555642352928821230860870550043554256370197072993944778035370097532049587705139351200010761752098313008705330077148474233051914660030690439284314821608407215643560940991248038263314;
            6'd57: xpb[1] = 1024'd99698854342551114564581305610826662851014909949472421889448788402414650558067212044446425691578856700833975179636222591414700774493290930528783025160207769765722295815782247439804837729767720089267237741832492487900486692290686801043106124631493831934968146451154512339737601129207848099647526741810439537552;
            6'd58: xpb[1] = 1024'd88388304873038880637770564228053681559485512531841866049460326262284006321825323949435127417958379698100204631125542977097864243430939508128744819459544989487890335261367421885664897424165342646484887778525633775790211632483060593380882172114513430818021632871618585395160380650008480555734112492372840811790;
            6'd59: xpb[1] = 1024'd77077755403526646710959822845280700267956115114211310209471864122153362085583435854423829144337902695366434082614863362781027712368588085728706613758882209210058374706952596331524957118562965203702537815218775063679936572675434385718658219597533029701075119292082658450583160170809113011820698242935242086028;
            6'd60: xpb[1] = 1024'd65767205934014412784149081462507718976426717696580754369483401982022717849341547759412530870717425692632663534104183748464191181306236663328668408058219428932226414152537770777385016812960587760920187851911916351569661512867808178056434267080552628584128605712546731506005939691609745467907283993497643360266;
            6'd61: xpb[1] = 1024'd54456656464502178857338340079734737684897320278950198529494939841892073613099659664401232597096948689898892985593504134147354650243885240928630202357556648654394453598122945223245076507358210318137837888605057639459386453060181970394210314563572227467182092133010804561428719212410377923993869744060044634504;
            6'd62: xpb[1] = 1024'd43146106994989944930527598696961756393367922861319642689506477701761429376857771569389934323476471687165122437082824519830518119181533818528591996656893868376562493043708119669105136201755832875355487925298198927349111393252555762731986362046591826350235578553474877616851498733211010380080455494622445908742;
            6'd63: xpb[1] = 1024'd31835557525477711003716857314188775101838525443689086849518015561630785140615883474378636049855994684431351888572144905513681588119182396128553790956231088098730532489293294114965195896153455432573137961991340215238836333444929555069762409529611425233289064973938950672274278254011642836167041245184847182980;
        endcase
    end

    always_comb begin
        case(flag[0][16:12])
            5'd0: xpb[2] = 1024'd0;
            5'd1: xpb[2] = 1024'd20525008055965477076906115931415793810309128026058531009529553421500140904373995379367337776235517681697581340061465291196845057056830973728515585255568307820898571934878468560825255590551077989790787998684481503128561273637303347407538457012631024116342551394403023727697057774812275292253626995747248457218;
            5'd2: xpb[2] = 1024'd41050016111930954153812231862831587620618256052117062019059106843000281808747990758734675552471035363395162680122930582393690114113661947457031170511136615641797143869756937121650511181102155979581575997368963006257122547274606694815076914025262048232685102788806047455394115549624550584507253991494496914436;
            5'd3: xpb[2] = 1024'd61575024167896431230718347794247381430927384078175593028588660264500422713121986138102013328706553045092744020184395873590535171170492921185546755766704923462695715804635405682475766771653233969372363996053444509385683820911910042222615371037893072349027654183209071183091173324436825876760880987241745371654;
            5'd4: xpb[2] = 1024'd82100032223861908307624463725663175241236512104234124038118213686000563617495981517469351104942070726790325360245861164787380228227323894914062341022273231283594287739513874243301022362204311959163151994737926012514245094549213389630153828050524096465370205577612094910788231099249101169014507982988993828872;
            5'd5: xpb[2] = 1024'd102625040279827385384530579657078969051545640130292655047647767107500704521869976896836688881177588408487906700307326455984225285284154868642577926277841539104492859674392342804126277952755389948953939993422407515642806368186516737037692285063155120581712756972015118638485288874061376461268134978736242286090;
            5'd6: xpb[2] = 1024'd123150048335792862461436695588494762861854768156351186057177320529000845426243972276204026657413106090185488040368791747181070342340985842371093511533409846925391431609270811364951533543306467938744727992106889018771367641823820084445230742075786144698055308366418142366182346648873651753521761974483490743308;
            5'd7: xpb[2] = 1024'd19608360707633598139543884115096123927465469056674032938575018885524090993308828745556293218990949462439919972972763603798851558556596481544448971772647113812599328974578062588146549942340340207225318382404130675535568065240226658887790629405187719547577956346704108063772876349757294028656699143605144716195;
            5'd8: xpb[2] = 1024'd40133368763599075216450000046511917737774597082732563948104572307024231897682824124923630995226467144137501313034228894995696615613427455272964557028215421633497900909456531148971805532891418197016106381088612178664129338877530006295329086417818743663920507741107131791469934124569569320910326139352393173413;
            5'd9: xpb[2] = 1024'd60658376819564552293356115977927711548083725108791094957634125728524372802056819504290968771461984825835082653095694186192541672670258429001480142283783729454396472844334999709797061123442496186806894379773093681792690612514833353702867543430449767780263059135510155519166991899381844613163953135099641630631;
            5'd10: xpb[2] = 1024'd81183384875530029370262231909343505358392853134849625967163679150024513706430814883658306547697502507532663993157159477389386729727089402729995727539352037275295044779213468270622316713993574176597682378457575184921251886152136701110406000443080791896605610529913179246864049674194119905417580130846890087849;
            5'd11: xpb[2] = 1024'd101708392931495506447168347840759299168701981160908156976693232571524654610804810263025644323933020189230245333218624768586231786783920376458511312794920345096193616714091936831447572304544652166388470377142056688049813159789440048517944457455711816012948161924316202974561107449006395197671207126594138545067;
            5'd12: xpb[2] = 1024'd122233400987460983524074463772175092979011109186966687986222785993024795515178805642392982100168537870927826673280090059783076843840751350187026898050488652917092188648970405392272827895095730156179258375826538191178374433426743395925482914468342840129290713318719226702258165223818670489924834122341387002285;
            5'd13: xpb[2] = 1024'd18691713359301719202181652298776454044621810087289534867620484349548041082243662111745248661746381243182258605884061916400858060056361989360382358289725919804300086014277656615467844294129602424659848766123779847942574856843149970368042801797744414978813361299005192399848694924702312765059771291463040975172;
            5'd14: xpb[2] = 1024'd39216721415267196279087768230192247854930938113348065877150037771048181986617657491112586437981898924879839945945527207597703117113192963088897943545294227625198657949156125176293099884680680414450636764808261351071136130480453317775581258810375439095155912693408216127545752699514588057313398287210289432390;
            5'd15: xpb[2] = 1024'd59741729471232673355993884161608041665240066139406596886679591192548322890991652870479924214217416606577421286006992498794548174170023936817413528800862535446097229884034593737118355475231758404241424763492742854199697404117756665183119715823006463211498464087811239855242810474326863349567025282957537889608;
            5'd16: xpb[2] = 1024'd80266737527198150432900000093023835475549194165465127896209144614048463795365648249847261990452934288275002626068457789991393231226854910545929114056430843266995801818913062297943611065782836394032212762177224357328258677755060012590658172835637487327841015482214263582939868249139138641820652278704786346826;
            5'd17: xpb[2] = 1024'd100791745583163627509806116024439629285858322191523658905738698035548604699739643629214599766688451969972583966129923081188238288283685884274444699311999151087894373753791530858768866656333914383823000760861705860456819951392363359998196629848268511444183566876617287310636926023951413934074279274452034804044;
            5'd18: xpb[2] = 1024'd121316753639129104586712231955855423096167450217582189915268251457048745604113639008581937542923969651670165306191388372385083345340516858002960284567567458908792945688669999419594122246884992373613788759546187363585381225029666707405735086860899535560526118271020311038333983798763689226327906270199283261262;
            5'd19: xpb[2] = 1024'd17775066010969840264819420482456784161778151117905036796665949813571991171178495477934204104501813023924597238795360229002864561556127497176315744806804725796000843053977250642789138645918864642094379149843429020349581648446073281848294974190301110410048766251306276735924513499647331501462843439320937234149;
            5'd20: xpb[2] = 1024'd38300074066935317341725536413872577972087279143963567806195503235072132075552490857301541880737330705622178578856825520199709618612958470904831330062373033616899414988855719203614394236469942631885167148527910523478142922083376629255833431202932134526391317645709300463621571274459606793716470435068185691367;
            5'd21: xpb[2] = 1024'd58825082122900794418631652345288371782396407170022098815725056656572272979926486236668879656972848387319759918918290811396554675669789444633346915317941341437797986923734187764439649827021020621675955147212392026606704195720679976663371888215563158642733869040112324191318629049271882085970097430815434148585;
            5'd22: xpb[2] = 1024'd79350090178866271495537768276704165592705535196080629825254610078072413884300481616036217433208366069017341258979756102593399732726620418361862500573509649258696558858612656325264905417572098611466743145896873529735265469357983324070910345228194182759076420434515347919015686824084157378223724426562682605803;
            5'd23: xpb[2] = 1024'd99875098234831748572443884208119959403014663222139160834784163499572554788674476995403555209443883750714922599041221393790244789783451392090378085829077957079595130793491124886090161008123176601257531144581355032863826742995286671478448802240825206875418971828918371646712744598896432670477351422309931063021;
            5'd24: xpb[2] = 1024'd120400106290797225649350000139535753213323791248197691844313716921072695693048472374770892985679401432412503939102686684987089846840282365818893671084646264900493702728369593446915416598674254591048319143265836535992388016632590018885987259253456230991761523223321395374409802373708707962730978418057179520239;
            5'd25: xpb[2] = 1024'd16858418662637961327457188666137114278934492148520538725711415277595941260113328844123159547257244804666935871706658541604871063055893004992249131323883531787701600093676844670110432997708126859528909533563078192756588440048996593328547146582857805841284171203607361072000332074592350237865915587178833493126;
            5'd26: xpb[2] = 1024'd37383426718603438404363304597552908089243620174579069735240968699096082164487324223490497323492762486364517211768123832801716120112723978720764716579451839608600172028555313230935688588259204849319697532247559695885149713686299940736085603595488829957626722598010384799697389849404625530119542582926081950344;
            5'd27: xpb[2] = 1024'd57908434774568915481269420528968701899552748200637600744770522120596223068861319602857835099728280168062098551829589123998561177169554952449280301835020147429498743963433781791760944178810282839110485530932041199013710987323603288143624060608119854073969273992413408527394447624216900822373169578673330407562;
            5'd28: xpb[2] = 1024'd78433442830534392558175536460384495709861876226696131754300075542096363973235314982225172875963797849759679891891054415195406234226385926177795887090588455250397315898312250352586199769361360828901273529616522702142272260960906635551162517620750878190311825386816432255091505399029176114626796574420578864780;
            5'd29: xpb[2] = 1024'd98958450886499869635081652391800289520171004252754662763829628963596504877609310361592510652199315531457261231952519706392251291283216899906311472346156763071295887833190718913411455359912438818692061528301004205270833534598209982958700974633381902306654376781219455982788563173841451406880423570167827321998;
            5'd30: xpb[2] = 1024'd119483458942465346711987768323216083330480132278813193773359182385096645781983305740959848428434833213154842572013984997589096348340047873634827057601725070892194459768069187474236710950463516808482849526985485708399394808235513330366239431646012926422996928175622479710485620948653726699134050565915075779216;
            5'd31: xpb[2] = 1024'd15941771314306082390094956849817444396090833179136040654756880741619891349048162210312114990012676585409274504617956854206877564555658512808182517840962337779402357133376438697431727349497389076963439917282727365163595231651919904808799318975414501272519576155908445408076150649537368974268987735036729752103;
        endcase
    end

    always_comb begin
        case(flag[1][5:0])
            6'd0: xpb[3] = 1024'd0;
            6'd1: xpb[3] = 1024'd80266737527198150432900000093023835475549194165465127896209144614048463795365648249847261990452934288275002626068457789991393231226854910545929114056430843266995801818913062297943611065782836394032212762177224357328258677755060012590658172835637487327841015482214263582939868249139138641820652278704786346826;
            6'd2: xpb[3] = 1024'd36466779370271559467001072781233238206399961205194571664286434163120032253422157589679452766248194267106855844679422145403722621612489486536698103096530645600300929068254907258256982940048467066754227915967208868292156505289223252216337775988045525388862127550311469135773208424349644266522614730783978209321;
            6'd3: xpb[3] = 1024'd116733516897469709899901072874257073681949155370659699560495578777168496048787805839526714756701128555381858470747879935395115852839344397082627217152961488867296730887167969556200594005831303460786440678144433225620415183044283264806995948823683012716703143032525732718713076673488782908343267009488764556147;
            6'd4: xpb[3] = 1024'd72933558740543118934002145562466476412799922410389143328572868326240064506844315179358905532496388534213711689358844290807445243224978973073396206193061291200601858136509814516513965880096934133508455831934417736584313010578446504432675551976091050777724255100622938271546416848699288533045229461567956418642;
            6'd5: xpb[3] = 1024'd29133600583616527968103218250675879143650689450118587096650157875311632964900824519191096308291648513045564907969808646219774633610613549064165195233161093533906985385851659476827337754362564806230470985724402247548210838112609744058355155128499088838745367168720143824379757023909794157747191913647148281137;
            6'd6: xpb[3] = 1024'd109400338110814678401003218343699714619199883615583714992859302489360096760266472769038358298744582801320567534038266436211167864837468459610094309289591936800902787204764721774770948820145401200262683747901626604876469515867669756649013327964136576166586382650934407407319625273048932799567844192351934627963;
            6'd7: xpb[3] = 1024'd65600379953888087435104291031909117350050650655313158760936592038431665218322982108870549074539842780152420752649230791623497255223103035600863298329691739134207914454106566735084320694411031872984698901691611115840367343401832996274692931116544614227607494719031612960152965448259438424269806644431126490458;
            6'd8: xpb[3] = 1024'd21800421796961496469205363720118520080901417695042602529013881587503233676379491448702739850335102758984273971260195147035826645608737611591632287369791541467513041703448411695397692568676662545706714055481595626804265170935996235900372534268952652288628606787128818512986305623469944048971769096510318352953;
            6'd9: xpb[3] = 1024'd102067159324159646902105363813142355556450611860507730425223026201551697471745139698550001840788037047259276597328652937027219876835592522137561401426222384734508843522361473993341303634459498939738926817658819984132523848691056248491030707104590139616469622269343082095926173872609082690792421375215104699779;
            6'd10: xpb[3] = 1024'd58267201167233055936206436501351758287301378900237174193300315750623265929801649038382192616583297026091129815939617292439549267221227098128330390466322187067813970771703318953654675508725129612460941971448804495096421676225219488116710310256998177677490734337440287648759514047819588315494383827294296562274;
            6'd11: xpb[3] = 1024'd14467243010306464970307509189561161018152145939966617961377605299694834387858158378214383392378557004922983034550581647851878657606861674119099379506421989401119098021045163913968047382990760285182957125238789006060319503759382727742389913409406215738511846405537493201592854223030093940196346279373488424769;
            6'd12: xpb[3] = 1024'd94733980537504615403207509282584996493701340105431745857586749913743298183223806628061645382831491293197985660619039437843271888833716584665028493562852832668114899839958226211911658448773596679215169887416013363388578181514442740333048086245043703066352861887751756784532722472169232582016998558078274771595;
            6'd13: xpb[3] = 1024'd50934022380578024437308581970794399224552107145161189625664039462814866641280315967893836158626751272029838879230003793255601279219351160655797482602952635001420027089300071172225030323039227351937185041205997874352476009048605979958727689397451741127373973955848962337366062647379738206718961010157466634090;
            6'd14: xpb[3] = 1024'd7134064223651433471409654659003801955402874184890633393741329011886435099336825307726026934422011250861692097840968148667930669604985736646566471643052437334725154338641916132538402197304858024659200194995982385316373836582769219584407292549859779188395086023946167890199402822590243831420923462236658496585;
            6'd15: xpb[3] = 1024'd87400801750849583904309654752027637430952068350355761289950473625934898894702473557573288924874945539136694723909425938659323900831840647192495585699483280601720956157554978430482013263087694418691412957173206742644632514337829232175065465385497266516236101506160431473139271071729382473241575740941444843411;
            6'd16: xpb[3] = 1024'd43600843593922992938410727440237040161802835390085205058027763175006467352758982897405479700670205517968547942520390294071653291217475223183264574739583082935026083406896823390795385137353325091413428110963191253608530341871992471800745068537905304577257213574257637025972611246939888097943538193020636705906;
            6'd17: xpb[3] = 1024'd123867581121121143371310727533260875637352029555550332954236907789054931148124631147252741691123139806243550568588848084063046522444330133729193688796013926202021885225809885688738996203136161485445640873140415610936789019627052484391403241373542791905098229056471900608912479496079026739764190471725423052732;
            6'd18: xpb[3] = 1024'd80067622964194552405411800221470278368202796595279776722314197338126499606181140487084932466918399785075403787199812439475375912829964709719962677836113728535327012475151730649052368077401792158167656026930400121900686847161215724017082844525950829966119341124569106161745819671289532364466152923804614915227;
            6'd19: xpb[3] = 1024'd36267664807267961439512872909679681099053563635009220490391486887198068064237649826917123242713659763907257005810776794887705303215599285710731666876213530868632139724493575609365739951667422830889671180720384632864584674695378963642762447678358868027140453192666311714579159846500037989168115375883806777722;
            6'd20: xpb[3] = 1024'd116534402334466111872412873002703516574602757800474348386600631501246531859603298076764385233166594052182259631879234584879098534442454196256660780932644374135627941543406637907309351017450259224921883942897608990192843352450438976233420620513996355354981468674880575297519028095639176630988767654588593124548;
            6'd21: xpb[3] = 1024'd72734444177539520906513945690912919305453524840203792154677921050318100317659807416596576008961854031014112850490198940291427924828088772247429769972744176468933068792748482867622722891715889897643899096687593501156741179984602215859100223666404393416002580742977780850352368270849682255690730106667784987043;
            6'd22: xpb[3] = 1024'd28934486020612929940615018379122322036304291879933235922755210599389668775716316756428766784757114009845966069101163295703757315213723348238198759012843978802238196042090327827936094765981520570365914250477578012120639007518765455484779826818812431477023692811074986403185708446060187880392692558746976849538;
            6'd23: xpb[3] = 1024'd109201223547811080373515018472146157511853486045398363818964355213438132571081965006276028775210048298120968695169621085695150546440578258784127873069274822069233997861003390125879705831764356964398127012654802369448897685273825468075437999654449918804864708293289249986125576695199326522213344837451763196364;
            6'd24: xpb[3] = 1024'd65401265390884489407616091160355560242704253085127807587041644762509701029138474346108219551005308276952821913780585441107479936826212834774896862109374624402539125110345235086193077706029987637120142166444786880412795512807988707701117602806857956865885820361386455538958916870409832146915307289530955058859;
            6'd25: xpb[3] = 1024'd21601307233957898441717163848564962973555020124857251355118934311581269487194983685940410326800568255784675132391549796519809327211847410765665851149474426735844252359687080046506449580295618309842157320234771391376693340342151947326797205959265994926906932429483661091792257045620337771617269741610146921354;
            6'd26: xpb[3] = 1024'd101868044761156048874617163941588798449104214290322379251328078925629733282560631935787672317253502544059677758460007586511202558438702321311594965205905270002840054178600142344450060646078454703874370082411995748704952018097211959917455378794903482254747947911697924674732125294759476413437922020314933268180;
            6'd27: xpb[3] = 1024'd58068086604229457908718236629798201179954981330051823019405368474701301740617141275619863093048762522891530977070971941923531948824336897302363954246005072336145181427941987304763432520344085376596385236201980259668849845631375199543134981947311520315769059979795130227565465469969982038139884472394125130675;
            6'd28: xpb[3] = 1024'd14268128447302866942819309318007603910805748369781266787482658023772870198673650615452053868844022501723384195681936297335861339209971473293132943286104874669450308677283832265076804394609716049318400389991964770632747673165538439168814585099719558376790172047892335780398805645180487662841846924473316993170;
            6'd29: xpb[3] = 1024'd94534865974501017375719309411031439386354942535246394683691802637821333994039298865299315859296956789998386821750394087327254570436826383839062057342535717936446110496196894563020415460392552443350613152169189127961006350920598451759472757935357045704631187530106599363338673894319626304662499203178103339996;
            6'd30: xpb[3] = 1024'd50734907817574426409820382099240842117205709574975838451769092186892902452095808205131506635092216768830240040361358442739583960822460959829831046382635520269751237745538739523333787334658183116072628305959173638924904178454761691385152361087765083765652299598203804916172014069530131929364461655257295202491;
            6'd31: xpb[3] = 1024'd6934949660647835443921454787450244848056476614705282219846381735964470910152317544963697410887476747662093258972322798151913351208095535820600035422735322603056364994880584483647159208923813788794643459749158149888802005988924931010831964240173121826673411666301010469005354244740637554066424107336487064986;
            6'd32: xpb[3] = 1024'd87201687187845985876821454880474080323605670780170410116055526350012934705517965794810959401340411035937095885040780588143306582434950446366529149479166165870052166813793646781590770274706650182826856221926382507217060683743984943601490137075810609154514427148515274051945222493879776195887076386041273411812;
            6'd33: xpb[3] = 1024'd43401729030919394910922527568683483054456437819899853884132815899084503163574475134643150177135671014768949103651744943555635972820585022357298138519265968203357294063135491741904142148972280855548871375716367018180958511278148183227169740228218647215535539216612479604778562669090281820589038838120465274307;
            6'd34: xpb[3] = 1024'd123668466558117545343822527661707318530005631985364981780341960513132966958940123384490412167588605303043951729720202733547029204047439932903227252575696811470353095882048554039847753214755117249581084137893591375509217189033208195817827913063856134543376554698826743187718430918229420462409691116825251621133;
            6'd35: xpb[3] = 1024'd79868508401190954377923600349916721260856399025094425548419250062204535416996632724322602943383865281875804948331167088959358594433074508893996241615796613803658223131390399000161125089020747922303099291683575886473115016567371435443507516216264172604397666766923948740551771093439926087111653568904443483628;
            6'd36: xpb[3] = 1024'd36068550244264363412024673038126123991707166064823869316496539611276103875053142064154793719179125260707658166942131444371687984818709084884765230655896416136963350380732243960474496963286378595025114445473560397437012844101534675069187119368672210665418778835021154293385111268650431711813616020983635346123;
            6'd37: xpb[3] = 1024'd116335287771462513844924673131149959467256360230288997212705684225324567670418790314002055709632059548982660793010589234363081216045563995430694344712327259403959152199645306258418108029069214989057327207650784754765271521856594687659845292204309697993259794317235417876324979517789570353634268299688421692949;
            6'd38: xpb[3] = 1024'd72535329614535922879025745819359362198107127270018440980782973774396136128475299653834246485427319527814514011621553589775410606431198571421463333752427061737264279448987151218731479903334845661779342361440769265729169349390757927285524895356717736054280906385332623429158319693000075978336230751767613555444;
            6'd39: xpb[3] = 1024'd28735371457609331913126818507568764928957894309747884748860263323467704586531808993666437261222579506646367230232517945187739996816833147412232322792526864070569406698328996179044851777600476334501357515230753776693067176924921166911204498509125774115302018453429828981991659868210581603038193203846805417939;
            6'd40: xpb[3] = 1024'd109002108984807482346026818600592600404507088475213012645069407937516168381897457243513699251675513794921369856300975735179133228043688057958161436848957707337565208517242058476988462843383312728533570277407978134021325854679981179501862671344763261443143033935644092564931528117349720244858845482551591764765;
            6'd41: xpb[3] = 1024'd65202150827880891380127891288802003135357855514942456413146697486587736839953966583345890027470773773753223074911940090591462618429322633948930425889057509670870335766583903437301834717648943401255585431197962644985223682214144419127542274497171299504164146003741298117764868292560225869560807934630783627260;
            6'd42: xpb[3] = 1024'd21402192670954300414228963977011405866208622554671900181223987035659305298010475923178080803266033752585076293522904446003792008814957209939699414929157312004175463015925748397615206591914574073977600584987947155949121509748307658753221877649579337565185258071838503670598208467770731494262770386709975489755;
            6'd43: xpb[3] = 1024'd101668930198152450847128964070035241341757816720137028077433131649707769093376124173025342793718968040860078919591362235995185240041812120485628528985588155271171264834838810695558817657697410468009813347165171513277380187503367671343880050485216824893026273554052767253538076716909870136083422665414761836581;
            6'd44: xpb[3] = 1024'd57868972041225859881230036758244644072608583759866471845510421198779337551432633512857533569514228019691932138202326591407514630427446696476397518025687957604476392084180655655872189531963041140731828500955156024241278015037530910969559653637624862954047385622149972806371416892120375760785385117493953699076;
            6'd45: xpb[3] = 1024'd14069013884299268915331109446454046803459350799595915613587710747850906009489142852689724345309487998523785356813290946819844020813081272467166507065787759937781519333522500616185561406228671813453843654745140535205175842571694150595239256790032901015068497690247178359204757067330881385487347569573145561571;
            6'd46: xpb[3] = 1024'd94335751411497419348231109539477882279008544965061043509796855361899369804854791102536986335762422286798787982881748736811237252039936183013095621122218603204777321152435562914129172472011508207486056416922364892533434520326754163185897429625670388342909513172461441942144625316470020027307999848277931908397;
            6'd47: xpb[3] = 1024'd50535793254570828382332182227687285009859312004790487277874144910970938262911300442369177111557682265630641201492713092223566642425570759003864610162318405538082448401777407874442544346277138880208071570712349403497332347860917402811577032778078426403930625240558647494977965491680525652009962300357123770892;
            6'd48: xpb[3] = 1024'd6735835097644237416433254915896687740710079044519931045951434460042506720967809782201367887352942244462494420103677447635896032811205334994633599202418207871387575651119252834755916220542769552930086724502333914461230175395080642437256635930486464464951737308655853047811305666891031276711924752436315633387;
            6'd49: xpb[3] = 1024'd87002572624842387849333255008920523216259273209985058942160579074090970516333458032048629877805876532737497046172135237627289264038060245540562713258849051138383377470032315132699527286325605946962299486679558271789488853150140655027914808766123951792792752790870116630751173916030169918532577031141101980213;
            6'd50: xpb[3] = 1024'd43202614467915796883434327697129925947110040249714502710237868623162538974389967371880820653601136511569350264783099593039618654423694821531331702298948853471688504719374160093012899160591236619684314640469542782753386680684303894653594411918531989853813864858967322183584514091240675543234539483220293842708;
            6'd51: xpb[3] = 1024'd123469351995113947316334327790153761422659234415179630606447013237211002769755615621728082644054070799844352890851557383031011885650549732077260816355379696738684306538287222390956510226374073013716527402646767140081645358439363907244252584754169477181654880341181585766524382340379814185055191761925080189534;
            6'd52: xpb[3] = 1024'd79669393838187356350435400478363164153510001454909074374524302786282571227812124961560273419849330778676206109462521738443341276036184308068029805395479499071989433787629067351269882100639703686438542556436751651045543185973527146869932187906577515242675992409278791319357722515590319809757154214004272052029;
            6'd53: xpb[3] = 1024'd35869435681260765384536473166572566884360768494638518142601592335354139685868634301392464195644590757508059328073486093855670666421818884058798794435579301405294561036970912311583253974905334359160557710226736162009441013507690386495611791058985553303697104477375996872191062690800825434459116666083463914524;
            6'd54: xpb[3] = 1024'd116136173208458915817436473259596402359909962660103646038810736949402603481234282551239726186097525045783061954141943883847063897648673794604727908492010144672290362855883974609526865040688170753192770472403960519337699691262750399086269963894623040631538119959590260455130930939939964076279768944788250261350;
            6'd55: xpb[3] = 1024'd72336215051532324851537545947805805090760729699833089806888026498474171939290791891071916961892785024614915172752908239259393288034308370595496897532109947005595490105225819569840236914953801425914785626193945030301597518796913638711949567047031078692559232027687466007964271115150469700981731396867442123845;
            6'd56: xpb[3] = 1024'd28536256894605733885638618636015207821611496739562533574965316047545740397347301230904107737688045003446768391363872594671722678419942946586265886572209749338900617354567664530153608789219432098636800779983929541265495346331076878337629170199439116753580344095784671560797611290360975325683693848946633986340;
            6'd57: xpb[3] = 1024'd108802994421803884318538618729039043297160690905027661471174460661594204192712949480751369728140979291721771017432330384663115909646797857132195000628640592605896419173480726828097219855002268492669013542161153898593754024086136890928287343035076604081421359577998935143737479539500113967504346127651420333166;
            6'd58: xpb[3] = 1024'd65003036264877293352639691417248446028011457944757105239251750210665772650769458820583560503936239270553624236043294740075445300032432433122963989668740394939201546422822571788410591729267899165391028695951138409557651851620300130553966946187484642142442471646096140696570819714710619592206308579730612195661;
            6'd59: xpb[3] = 1024'd21203078107950702386740764105457848758862224984486549007329039759737341108825968160415751279731499249385477454654259095487774690418067009113732978708840197272506673672164416748723963603533529838113043849741122920521549679154463370179646549339892680203463583714193346249404159889921125216908271031809804058156;
            6'd60: xpb[3] = 1024'd101469815635148852819640764198481684234411419149951676903538184373785804904191616410263013270184433537660480080722716885479167921644921919659662092765271040539502475491077479046667574669316366232145256611918347277849808356909523382770304722175530167531304599196407609832344028139060263858728923310514590404982;
            6'd61: xpb[3] = 1024'd57669857478222261853741836886691086965262186189681120671615473922857373362248125750095204045979693516492333299333681240891497312030556495650431081805370842872807602740419324006980946543581996904867271765708331788813706184443686622395984325327938205592325711264504815385177368314270769483430885762593782267477;
            6'd62: xpb[3] = 1024'd13869899321295670887842909574900489696112953229410564439692763471928941820304635089927394821774953495324186517944645596303826702416191071641200070845470645206112729989761168967294318417847627577589286919498316299777604011977849862021663928480346243653346823332602020938010708489481275108132848214672974129972;
            6'd63: xpb[3] = 1024'd94136636848493821320742909667924325171662147394875692335901908085977405615670283339774656812227887783599189144013103386295219933643045982187129184901901488473108531808674231265237929483630463971621499681675540657105862689732909874612322101315983730981187838814816284520950576738620413749953500493377760476798;
        endcase
    end

    always_comb begin
        case(flag[1][11:6])
            6'd0: xpb[4] = 1024'd0;
            6'd1: xpb[4] = 1024'd50336678691567230354843982356133727902512914434605136103979197635048974073726792679606847588023147762431042362624067741707549324028680558177898173942001290806413659058016076225551301357896094644343514835465525168069760517267073114238001704468391769042208950882913490073783916913830919374655462945456952339293;
            6'd2: xpb[4] = 1024'd100673357383134460709687964712267455805025828869210272207958395270097948147453585359213695176046295524862084725248135483415098648057361116355796347884002581612827318116032152451102602715792189288687029670931050336139521034534146228476003408936783538084417901765826980147567833827661838749310925890913904678586;
            6'd3: xpb[4] = 1024'd26943340390576949665733019663586750962840316178079724183805737840170026883871239128805471549411768977849977680414709790543584131244821339978534396809672831485550302604477011339023664882171078211720346898009335657844920701580322569749026543721945857859806949234623412191245222667564125106847699009745262533548;
            6'd4: xpb[4] = 1024'd77280019082144180020577002019720478865353230612684860287784935475219000957598031808412319137434916740281020043038777532251133455273501898156432570751674122291963961662493087564574966240067172856063861733474860825914681218847395683987028248190337626902015900117536902265029139581395044481503161955202214872841;
            6'd5: xpb[4] = 1024'd3550002089586668976622056971039774023167717921554312263632278045291079694015685578004095510800390193268912998205351839379618938460962121779170619677344372164686946150937946452496028406446061779097178960553146147620080885893572025260051382975499946677404947586333334308706528421297330839039935074033572727803;
            6'd6: xpb[4] = 1024'd53886680781153899331466039327173501925680632356159448367611475680340053767742478257610943098823537955699955360829419581087168262489642679957068793619345662971100605208954022678047329764342156423440693796018671315689841403160645139498053087443891715719613898469246824382490445335128250213695398019490525067096;
            6'd7: xpb[4] = 1024'd104223359472721129686310021683307229828193546790764584471590673315389027841469270937217790686846685718130997723453487322794717586518323238134966967561346953777514264266970098903598631122238251067784208631484196483759601920427718253736054791912283484761822849352160314456274362248959169588350860964947477406389;
            6'd8: xpb[4] = 1024'd30493342480163618642355076634626524986008034099634036447438015885461106577886924706809567060212159171118890678620061629923203069705783461757705016487017203650237248755414957791519693288617139990817525858562481805465001587473894595009077926697445804537211896820956746499951751088861455945887634083778835261351;
            6'd9: xpb[4] = 1024'd80830021171730848997199058990760252888520948534239172551417213520510080651613717386416414648235306933549933041244129371630752393734464019935603190429018494456650907813431034017070994646513234635161040694028006973534762104740967709247079631165837573579420847703870236573735668002692375320543097029235787600644;
            6'd10: xpb[4] = 1024'd7100004179173337953244113942079548046335435843108624527264556090582159388031371156008191021600780386537825996410703678759237876921924243558341239354688744329373892301875892904992056812892123558194357921106292295240161771787144050520102765950999893354809895172666668617413056842594661678079870148067145455606;
            6'd11: xpb[4] = 1024'd57436682870740568308088096298213275948848350277713760631243753725631133461758163835615038609623928148968868359034771420466787200950604801736239413296690035135787551359891969130543358170788218202537872756571817463309922289054217164758104470419391662397018846055580158691196973756425581052735333093524097794899;
            6'd12: xpb[4] = 1024'd107773361562307798662932078654347003851361264712318896735222951360680107535484956515221886197647075911399910721658839162174336524979285359914137587238691325942201210417908045356094659528684312846881387592037342631379682806321290278996106174887783431439227796938493648764980890670256500427390796038981050134192;
            6'd13: xpb[4] = 1024'd34043344569750287618977133605666299009175752021188348711070293930752186271902610284813662571012549364387803676825413469302822008166745583536875636164361575814924194906352904244015721695063201769914704819115627953085082473367466620269129309672945751214616844407290080808658279510158786784927569157812407989154;
            6'd14: xpb[4] = 1024'd84380023261317517973821115961800026911688666455793484815049491565801160345629402964420510159035697126818846039449481211010371332195426141714773810106362866621337853964368980469567023052959296414258219654581153121154842990634539734507131014141337520256825795290203570882442196423989706159583032103269360328447;
            6'd15: xpb[4] = 1024'd10650006268760006929866170913119322069503153764662936790896834135873239082047056734012286532401170579806738994616055518138856815382886365337511859032033116494060838452813839357488085219338185337291536881659438442860242657680716075780154148926499840032214842759000002926119585263891992517119805222100718183409;
            6'd16: xpb[4] = 1024'd60986684960327237284710153269253049972016068199268072894876031770922213155773849413619134120424318342237781357240123259846406139411566923515410032974034407300474497510829915583039386577234279981635051717124963610930003174947789190018155853394891609074423793641913492999903502177722911891775268167557670522702;
            6'd17: xpb[4] = 1024'd111323363651894467639554135625386777874528982633873208998855229405971187229500642093225981708447466104668823719864191001553955463440247481693308206916035698106888156568845991808590687935130374625978566552590488778999763692214862304256157557863283378116632744524826983073687419091553831266430731113014622861995;
            6'd18: xpb[4] = 1024'd37593346659336956595599190576706073032343469942742660974702571976043265965918295862817758081812939557656716675030765308682440946627707705316046255841705947979611141057290850696511750101509263549011883779668774100705163359261038645529180692648445697892021791993623415117364807931456117623967504231845980716957;
            6'd19: xpb[4] = 1024'd87930025350904186950443172932839800934856384377347797078681769611092240039645088542424605669836087320087759037654833050389990270656388263493944429783707238786024800115306926922063051459405358193355398615134299268774923876528111759767182397116837466934230742876536905191148724845287036998622967177302933056250;
            6'd20: xpb[4] = 1024'd14200008358346675906488227884159096092670871686217249054529112181164318776062742312016382043201560773075651992821407357518475753843848487116682478709377488658747784603751785809984113625784247116388715842212584590480323543574288101040205531901999786709619790345333337234826113685189323356159740296134290911212;
            6'd21: xpb[4] = 1024'd64536687049913906261332210240292823995183786120822385158508309816213292849789534991623229631224708535506694355445475099226025077872529045294580652651378779465161443661767862035535414983680341760732230677678109758550084060841361215278207236370391555751828741228246827308610030599020242730815203241591243250505;
            6'd22: xpb[4] = 1024'd114873365741481136616176192596426551897696700555427521262487507451262266923516327671230077219247856297937736718069542840933574401901209603472478826593380070271575102719783938261086716341576436405075745513143634926619844578108434329516208940838783324794037692111160317382393947512851162105470666187048195589798;
            6'd23: xpb[4] = 1024'd41143348748923625572221247547745847055511187864296973238334850021334345659933981440821853592613329750925629673236117148062059885088669827095216875519050320144298087208228797149007778507955325328109062740221920248325244245154610670789232075623945644569426739579956749426071336352753448463007439305879553444760;
            6'd24: xpb[4] = 1024'd91480027440490855927065229903879574958024102298902109342314047656383319733660774120428701180636477513356672035860184889769609209117350385273115049461051610950711746266244873374559079865851419972452577575687445416395004762421683785027233780092337413611635690462870239499855253266584367837662902251336505784053;
            6'd25: xpb[4] = 1024'd17750010447933344883110284855198870115838589607771561318161390226455398470078427890020477554001950966344564991026759196898094692304810608895853098386721860823434730754689732262480142032230308895485894802765730738100404429467860126300256914877499733387024737931666671543532642106486654195199675370167863639015;
            6'd26: xpb[4] = 1024'd68086689139500575237954267211332598018351504042376697422140587861504372543805220569627325142025098728775607353650826938605644016333491167073751272328723151629848389812705808488031443390126403539829409638231255906170164946734933240538258619345891502429233688814580161617316559020317573569855138315624815978308;
            6'd27: xpb[4] = 1024'd118423367831067805592798249567466325920864418476981833526119785496553346617532013249234172730048246491206649716274894680313193340362171725251649446270724442436262048870721884713582744748022498184172924473696781074239925464002006354776260323814283271471442639697493651691100475934148492944510601261081768317601;
            6'd28: xpb[4] = 1024'd44693350838510294548843304518785621078678905785851285501967128066625425353949667018825949103413719944194542671441468987441678823549631948874387495196394692308985033359166743601503806914401387107206241700775066395945325131048182696049283458599445591246831687166290083734777864774050779302047374379913126172563;
            6'd29: xpb[4] = 1024'd95030029530077524903687286874919348981191820220456421605946325701674399427676459698432796691436867706625585034065536729149228147578312507052285669138395983115398692417182819827055108272297481751549756536240591564015085648315255810287285163067837360289040638049203573808561781687881698676702837325370078511856;
            6'd30: xpb[4] = 1024'd21300012537520013859732341826238644139006307529325873581793668271746478164094113468024573064802341159613477989232111036277713630765772730675023718064066232988121676905627678714976170438676370674583073763318876885720485315361432151560308297852999680064429685518000005852239170527783985034239610444201436366818;
            6'd31: xpb[4] = 1024'd71636691229087244214576324182372372041519221963931009685772865906795452237820906147631420652825488922044520351856178777985262954794453288852921892006067523794535335963643754940527471796572465318926588598784402053790245832628505265798310002321391449106638636400913495926023087441614904408895073389658388706111;
            6'd32: xpb[4] = 1024'd121973369920654474569420306538506099944032136398536145789752063541844426311547698827238268240848636684475562714480246519692812278823133847030820065948068814600948995021659831166078773154468559963270103434249927221860006349895578380036311706789783218148847587283826985999807004355445823783550536335115341045404;
            6'd33: xpb[4] = 1024'd48243352928096963525465361489825395101846623707405597765599406111916505047965352596830044614214110137463455669646820826821297762010594070653558114873739064473671979510104690053999835320847448886303420661328212543565406016941754721309334841574945537924236634752623418043484393195348110141087309453946698900366;
            6'd34: xpb[4] = 1024'd98580031619664193880309343845959123004359538142010733869578603746965479121692145276436892202237257899894498032270888568528847086039274628831456288815740355280085638568120766279551136678743543530646935496793737711635166534208827835547336546043337306966445585635536908117268310109179029515742772399403651239659;
            6'd35: xpb[4] = 1024'd24850014627106682836354398797278418162174025450880185845425946317037557858109799046028668575602731352882390987437462875657332569226734852454194337741410605152808623056565625167472198845122432453680252723872023033340566201255004176820359680828499626741834633104333340160945698949081315873279545518235009094621;
            6'd36: xpb[4] = 1024'd75186693318673913191198381153412146064686939885485321949405143952086531931836591725635516163625879115313433350061530617364881893255415410632092511683411895959222282114581701393023500203018527098023767559337548201410326718522077291058361385296891395784043583987246830234729615862912235247935008463691961433914;
            6'd37: xpb[4] = 1024'd1456676326116402147243436104731441222501427194354773925252486522158610668254245495227292536991352568301326305228104924493367376442875634254830560609082145831945266603026560280944562369397416021057084786415833523115726385568253632331384520082053715559432631456043262278407004702814521605471781582523319288876;
            6'd38: xpb[4] = 1024'd51793355017683632502087418460865169125014341628959910029231684157207584741981038174834140125014500330732368667852172666200916700471556192432728734551083436638358925661042636506495863727293510665400599621881358691185486902835326746569386224550445484601641582338956752352190921616645440980127244527980271628169;
            6'd39: xpb[4] = 1024'd102130033709250862856931400816998897027527256063565046133210881792256558815707830854440987713037648093163411030476240407908466024500236750610626908493084727444772584719058712732047165085189605309744114457346883859255247420102399860807387929018837253643850533221870242425974838530476360354782707473437223967462;
            6'd40: xpb[4] = 1024'd28400016716693351812976455768318192185341743372434498109058224362328637552125484624032764086403121546151303985642814715036951507687696974233364957418754977317495569207503571619968227251568494232777431684425169180960647087148576202080411063803999573419239580690666674469652227370378646712319480592268581822424;
            6'd41: xpb[4] = 1024'd78736695408260582167820438124451920087854657807039634213037421997377611625852277303639611674426269308582346348266882456744500831716377532411263131360756268123909228265519647845519528609464588877120946519890694349030407604415649316318412768272391342461448531573580164543436144284209566086974943537725534161717;
            6'd42: xpb[4] = 1024'd5006678415703071123865493075771215245669145115909086188884764567449690362269931073231388047791742761570239303433456763872986314903837756034001180286426517996632212753964506733440590775843477800154263746968979670735807271461825657591435903057553662236837579042376596587113533124111852444511716656556892016679;
            6'd43: xpb[4] = 1024'd55343357107270301478709475431904943148182059550514222292863962202498664435996723752838235635814890524001281666057524505580535638932518314211899354228427808803045871811980582958991892133739572444497778582434504838805567788728898771829437607525945431279046529925290086660897450037942771819167179602013844355972;
            6'd44: xpb[4] = 1024'd105680035798837531833553457788038671050694973985119358396843159837547638509723516432445083223838038286432324028681592247288084962961198872389797528170429099609459530869996659184543193491635667088841293417900030006875328305995971886067439311994337200321255480808203576734681366951773691193822642547470796695265;
            6'd45: xpb[4] = 1024'd31950018806280020789598512739357966208509461293988810372690502407619717246141170202036859597203511739420216983848166554416570446148659096012535577096099349482182515358441518072464255658014556011874610644978315328580727973042148227340462446779499520096644528277000008778358755791675977551359415666302154550227;
            6'd46: xpb[4] = 1024'd82286697497847251144442495095491694111022375728593946476669700042668691319867962881643707185226659501851259346472234296124119770177339654190433751038100640288596174416457594298015557015910650656218125480443840496650488490309221341578464151247891289138853479159913498852142672705506896926014878611759106889520;
            6'd47: xpb[4] = 1024'd8556680505289740100487550046810989268836863037463398452517042612740770056285616651235483558592132954839152301638808603252605253364799877813171799963770890161319158904902453185936619182289539579251442707522125818355888157355397682851487286033053608914242526628709930895820061545409183283551651730590464744482;
            6'd48: xpb[4] = 1024'd58893359196856970455331532402944717171349777472068534556496240247789744130012409330842331146615280717270194664262876344960154577393480435991069973905772180967732817962918529411487920540185634223594957542987650986425648674622470797089488990501445377956451477511623420969603978459240102658207114676047417083775;
            6'd49: xpb[4] = 1024'd109230037888424200810175514759078445073862691906673670660475437882838718203739202010449178734638428479701237026886944086667703901422160994168968147847773471774146477020934605637039221898081728867938472378453176154495409191889543911327490694969837146998660428394536911043387895373071022032862577621504369423068;
            6'd50: xpb[4] = 1024'd35500020895866689766220569710397740231677179215543122636322780452910796940156855780040955108003901932689129982053518393796189384609621217791706196773443721646869461509379464524960284064460617790971789605531461476200808858935720252600513829754999466774049475863333343087065284212973308390399350740335727278030;
            6'd51: xpb[4] = 1024'd85836699587433920121064552066531468134190093650148258740301978087959771013883648459647802696027049695120172344677586135503738708638301775969604370715445012453283120567395540750511585422356712435315304440996986644270569376202793366838515534223391235816258426746246833160849201126804227765054813685792679617323;
            6'd52: xpb[4] = 1024'd12106682594876409077109607017850763292004580959017710716149320658031849750301302229239579069392523148108065299844160442632224191825761999592342419641115262326006105055840399638432647588735601358348621668075271965975969043248969708111538669008553555591647474215043265204526589966706514122591586804624037472285;
            6'd53: xpb[4] = 1024'd62443361286443639431953589373984491194517495393622846820128518293080823824028094908846426657415670910539107662468228184339773515854442557770240593583116553132419764113856475863983948946631696002692136503540797134045729560516042822349540373476945324633856425097956755278310506880537433497247049750080989811578;
            6'd54: xpb[4] = 1024'd112780039978010869786797571730118219097030409828227982924107715928129797897754887588453274245438818672970150025092295926047322839883123115948138767525117843938833423171872552089535250304527790647035651339006322302115490077783115936587542077945337093676065375980870245352094423794368352871902512695537942150871;
            6'd55: xpb[4] = 1024'd39050022985453358742842626681437514254844897137097434899955058498201876634172541358045050618804292125958042980258870233175808323070583339570876816450788093811556407660317410977456312470906679570068968566084607623820889744829292277860565212730499413451454423449666677395771812634270639229439285814369300005833;
            6'd56: xpb[4] = 1024'd89386701677020589097686609037571242157357811571702571003934256133250850707899334037651898206827439888389085342882937974883357647099263897748774990392789384617970066718333487203007613828802774214412483401550132791890650262096365392098566917198891182493663374332580167469555729548101558604094748759826252345126;
            6'd57: xpb[4] = 1024'd15656684684463078053731663988890537315172298880572022979781598703322929444316987807243674580192913341376978298049512282011843130286724121371513039318459634490693051206778346090928675995181663137445800628628418113596049929142541733371590051984053502269052421801376599513233118388003844961631521878657610200088;
            6'd58: xpb[4] = 1024'd65993363376030308408575646345024265217685213315177159083760796338371903518043780486850522168216061103808020660673580023719392454315404679549411213260460925297106710264794422316479977353077757781789315464093943281665810446409614847609591756452445271311261372684290089587017035301834764336286984824114562539381;
            6'd59: xpb[4] = 1024'd116330042067597538763419628701157993120198127749782295187739993973420877591770573166457369756239208866239063023297647765426941778344085237727309387202462216103520369322810498542031278710973852426132830299559468449735570963676687961847593460920837040353470323567203579660800952215665683710942447769571514878674;
            6'd60: xpb[4] = 1024'd42600025075040027719464683652477288278012615058651747163587336543492956328188226936049146129604682319226955978464222072555427261531545461350047436128132465976243353811255357429952340877352741349166147526637753771440970630722864303120616595705999360128859371036000011704478341055567970068479220888402872733636;
            6'd61: xpb[4] = 1024'd92936703766607258074308666008611016180525529493256883267566534178541930401915019615655993717627830081657998341088289814262976585560226019527945610070133756782657012869271433655503642235248835993509662362103278939510731147989937417358618300174391129171068321918913501778262257969398889443134683833859825072929;
            6'd62: xpb[4] = 1024'd19206686774049747030353720959930311338340016802126335243413876748614009138332673385247770090993303534645891296254864121391462068747686243150683658995804006655379997357716292543424704401627724916542979589181564261216130815036113758631641434959553448946457369387709933821939646809301175800671456952691182927891;
            6'd63: xpb[4] = 1024'd69543365465616977385197703316064039240852931236731471347393074383662983212059466064854617679016451297076933658878931863099011392776366801328581832937805297461793656415732368768976005759523819560886494424647089429285891332303186872869643139427945217988666320270623423895723563723132095175326919898148135267184;
        endcase
    end

    always_comb begin
        case(flag[1][16:12])
            5'd0: xpb[5] = 1024'd0;
            5'd1: xpb[5] = 1024'd119880044157184207740041685672197767143365845671336607451372272018711957285786258744461465267039599059507976021502999604806560716805047359506480006879806588268207315473748444994527307117419914205230009260112614597355651849570259987107644843896336987030875271153536913969507480636963014549982382843605087606477;
            5'd2: xpb[5] = 1024'd115693392630243674081284443939581101542033264216937530774612688972447019234263378578907859319421523809572802635548505775034057592768874384457799888743282135602723956377925672651424375043322622689149820911837989348346942848919623201250311118109444524794930638892956769908908433199997396082846075860584580728623;
            5'd3: xpb[5] = 1024'd111506741103303140422527202206964435940700682762538454097853105926182081182740498413354253371803448559637629249594011945261554468732701409409119770606757682937240597282102900308321442969225331173069632563563364099338233848268986415392977392322552062558986006632376625848309385763031777615709768877564073850769;
            5'd4: xpb[5] = 1024'd107320089576362606763769960474347770339368101308139377421093522879917143131217618247800647424185373309702455863639518115489051344696528434360439652470233230271757238186280127965218510895128039656989444215288738850329524847618349629535643666535659600323041374371796481787710338326066159148573461894543566972915;
            5'd5: xpb[5] = 1024'd103133438049422073105012718741731104738035519853740300744333939833652205079694738082247041476567298059767282477685024285716548220660355459311759534333708777606273879090457355622115578821030748140909255867014113601320815846967712843678309940748767138087096742111216337727111290889100540681437154911523060095061;
            5'd6: xpb[5] = 1024'd98946786522481539446255477009114439136702938399341224067574356787387267028171857916693435528949222809832109091730530455944045096624182484263079416197184324940790519994634583279012646746933456624829067518739488352312106846317076057820976214961874675851152109850636193666512243452134922214300847928502553217207;
            5'd7: xpb[5] = 1024'd94760134995541005787498235276497773535370356944942147390814773741122328976648977751139829581331147559896935705776036626171541972588009509214399298060659872275307160898811810935909714672836165108748879170464863103303397845666439271963642489174982213615207477590056049605913196015169303747164540945482046339353;
            5'd8: xpb[5] = 1024'd90573483468600472128740993543881107934037775490543070714055190694857390925126097585586223633713072309961762319821542796399038848551836534165719179924135419609823801802989038592806782598738873592668690822190237854294688845015802486106308763388089751379262845329475905545314148578203685280028233962461539461499;
            5'd9: xpb[5] = 1024'd86386831941659938469983751811264442332705194036143994037295607648592452873603217420032617686094997060026588933867048966626535724515663559117039061787610966944340442707166266249703850524641582076588502473915612605285979844365165700248975037601197289143318213068895761484715101141238066812891926979441032583645;
            5'd10: xpb[5] = 1024'd82200180414719404811226510078647776731372612581744917360536024602327514822080337254479011738476921810091415547912555136854032600479490584068358943651086514278857083611343493906600918450544290560508314125640987356277270843714528914391641311814304826907373580808315617424116053704272448345755619996420525705791;
            5'd11: xpb[5] = 1024'd78013528887778871152469268346031111130040031127345840683776441556062576770557457088925405790858846560156242161958061307081529476443317609019678825514562061613373724515520721563497986376446999044428125777366362107268561843063892128534307586027412364671428948547735473363517006267306829878619313013400018827937;
            5'd12: xpb[5] = 1024'd73826877360838337493712026613414445528707449672946764007016858509797638719034576923371799843240771310221068776003567477309026352407144633970998707378037608947890365419697949220395054302349707528347937429091736858259852842413255342676973860240519902435484316287155329302917958830341211411483006030379511950083;
            5'd13: xpb[5] = 1024'd69640225833897803834954784880797779927374868218547687330257275463532700667511696757818193895622696060285895390049073647536523228370971658922318589241513156282407006323875176877292122228252416012267749080817111609251143841762618556819640134453627440199539684026575185242318911393375592944346699047359005072229;
            5'd14: xpb[5] = 1024'd65453574306957270176197543148181114326042286764148610653497692417267762615988816592264587948004620810350722004094579817764020104334798683873638471104988703616923647228052404534189190154155124496187560732542486360242434841111981770962306408666734977963595051765995041181719863956409974477210392064338498194375;
            5'd15: xpb[5] = 1024'd61266922780016736517440301415564448724709705309749533976738109371002824564465936426710982000386545560415548618140085987991516980298625708824958352968464250951440288132229632191086258080057832980107372384267861111233725840461344985104972682879842515727650419505414897121120816519444356010074085081317991316521;
            5'd16: xpb[5] = 1024'd57080271253076202858683059682947783123377123855350457299978526324737886512943056261157376052768470310480375232185592158219013856262452733776278234831939798285956929036406859847983326005960541464027184035993235862225016839810708199247638957092950053491705787244834753060521769082478737542937778098297484438667;
            5'd17: xpb[5] = 1024'd52893619726135669199925817950331117522044542400951380623218943278472948461420176095603770105150395060545201846231098328446510732226279758727598116695415345620473569940584087504880393931863249947946995687718610613216307839160071413390305231306057591255761154984254608999922721645513119075801471115276977560813;
            5'd18: xpb[5] = 1024'd48706968199195135541168576217714451920711960946552303946459360232208010409897295930050164157532319810610028460276604498674007608190106783678917998558890892954990210844761315161777461857765958431866807339443985364207598838509434627532971505519165129019816522723674464939323674208547500608665164132256470682959;
            5'd19: xpb[5] = 1024'd44520316672254601882411334485097786319379379492153227269699777185943072358374415764496558209914244560674855074322110668901504484153933808630237880422366440289506851748938542818674529783668666915786618991169360115198889837858797841675637779732272666783871890463094320878724626771581882141528857149235963805105;
            5'd20: xpb[5] = 1024'd40333665145314068223654092752481120718046798037754150592940194139678134306851535598942952262296169310739681688367616839129001360117760833581557762285841987624023492653115770475571597709571375399706430642894734866190180837208161055818304053945380204547927258202514176818125579334616263674392550166215456927251;
            5'd21: xpb[5] = 1024'd36147013618373534564896851019864455116714216583355073916180611093413196255328655433389346314678094060804508302413123009356498236081587858532877644149317534958540133557292998132468665635474083883626242294620109617181471836557524269960970328158487742311982625941934032757526531897650645207256243183194950049397;
            5'd22: xpb[5] = 1024'd31960362091433000906139609287247789515381635128955997239421028047148258203805775267835740367060018810869334916458629179583995112045414883484197526012793082293056774461470225789365733561376792367546053946345484368172762835906887484103636602371595280076037993681353888696927484460685026740119936200174443171543;
            5'd23: xpb[5] = 1024'd27773710564492467247382367554631123914049053674556920562661445000883320152282895102282134419441943560934161530504135349811491988009241908435517407876268629627573415365647453446262801487279500851465865598070859119164053835256250698246302876584702817840093361420773744636328437023719408272983629217153936293689;
            5'd24: xpb[5] = 1024'd23587059037551933588625125822014458312716472220157843885901861954618382100760014936728528471823868310998988144549641520038988863973068933386837289739744176962090056269824681103159869413182209335385677249796233870155344834605613912388969150797810355604148729160193600575729389586753789805847322234133429415835;
            5'd25: xpb[5] = 1024'd19400407510611399929867884089397792711383890765758767209142278908353444049237134771174922524205793061063814758595147690266485739936895958338157171603219724296606697174001908760056937339084917819305488901521608621146635833954977126531635425010917893368204096899613456515130342149788171338711015251112922537981;
            5'd26: xpb[5] = 1024'd15213755983670866271110642356781127110051309311359690532382695862088505997714254605621316576587717811128641372640653860493982615900722983289477053466695271631123338078179136416954005264987626303225300553246983372137926833304340340674301699224025431132259464639033312454531294712822552871574708268092415660127;
            5'd27: xpb[5] = 1024'd11027104456730332612353400624164461508718727856960613855623112815823567946191374440067710628969642561193467986686160030721479491864550008240796935330170818965639978982356364073851073190890334787145112204972358123129217832653703554816967973437132968896314832378453168393932247275856934404438401285071908782273;
            5'd28: xpb[5] = 1024'd6840452929789798953596158891547795907386146402561537178863529769558629894668494274514104681351567311258294600731666200948976367828377033192116817193646366300156619886533591730748141116793043271064923856697732874120508832003066768959634247650240506660370200117873024333333199838891315937302094302051401904419;
            5'd29: xpb[5] = 1024'd2653801402849265294838917158931130306053564948162460502103946723293691843145614108960498733733492061323121214777172371176473243792204058143436699057121913634673260790710819387645209042695751754984735508423107625111799831352429983102300521863348044424425567857292880272734152401925697470165787319030895026565;
            5'd30: xpb[5] = 1024'd122533845560033473034880602831128897449419410619499067953476218742005649128931872853421964000773091120831097236280171975983033960597251417649916705936928501902880576264459264382172516160115665960214744768535722222467451680922689970209945365759685031455300839010829794242241633038888712020148170162635982633042;
            5'd31: xpb[5] = 1024'd118347194033092939376123361098512231848086829165099991276716635695740711077408992687868358053155015870895923850325678146210530836561078442601236587800404049237397217168636492039069584086018374444134556420261096973458742680272053184352611639972792569219356206750249650181642585601923093553011863179615475755188;
        endcase
    end

    always_comb begin
        case(flag[2][5:0])
            6'd0: xpb[6] = 1024'd0;
            6'd1: xpb[6] = 1024'd57080271253076202858683059682947783123377123855350457299978526324737886512943056261157376052768470310480375232185592158219013856262452733776278234831939798285956929036406859847983326005960541464027184035993235862225016839810708199247638957092950053491705787244834753060521769082478737542937778098297484438667;
            6'd2: xpb[6] = 1024'd114160542506152405717366119365895566246754247710700914599957052649475773025886112522314752105536940620960750464371184316438027712524905467552556469663879596571913858072813719695966652011921082928054368071986471724450033679621416398495277914185900106983411574489669506121043538164957475085875556196594968877334;
            6'd3: xpb[6] = 1024'd47174118075103867177250251644028916625432944440315687771803723909236764201520029873457056943647736621997976289099283040077977727946137866773674579479488353924180112539649362206319738826364418670771354499592467740310689669211227824777938301595620711208297458320387201151458779173507579611694644468266858831670;
            6'd4: xpb[6] = 1024'd104254389328180070035933311326976699748810068295666145071782250233974650714463086134614432996416206932478351521284875198296991584208590600549952814311428152210137041576056222054303064832324960134798538535585703602535706509021936024025577258688570764700003245565221954211980548255986317154632422566564343270337;
            6'd5: xpb[6] = 1024'd37267964897131531495817443605110050127488765025280918243628921493735641890097003485756737834527002933515577346012973921936941599629822999771070924127036909562403296042891864564656151646768295877515524963191699618396362498611747450308237646098291368924889129395939649242395789264536421680451510838236233224673;
            6'd6: xpb[6] = 1024'd94348236150207734354500503288057833250865888880631375543607447818473528403040059746914113887295473243995952578198566080155955455892275733547349158958976707848360225079298724412639477652728837341542708999184935480621379338422455649555876603191241422416594916640774402302917558347015159223389288936533717663340;
            6'd7: xpb[6] = 1024'd27361811719159195814384635566191183629544585610246148715454119078234519578673977098056418725406269245033178402926664803795905471313508132768467268774585465200626479546134366922992564467172173084259695426790931496482035328012267075838536990600962026641480800471492097333332799355565263749208377208205607617676;
            6'd8: xpb[6] = 1024'd84442082972235398673067695249138966752921709465596606015432645402972406091617033359213794778174739555513553635112256962014919327575960866544745503606525263486583408582541226770975890473132714548286879462784167358707052167822975275086175947693912080133186587716326850393854568438044001292146155306503092056343;
            6'd9: xpb[6] = 1024'd17455658541186860132951827527272317131600406195211379187279316662733397267250950710356099616285535556550779459840355685654869342997193265765863613422134020838849663049376869281328977287576050291003865890390163374567708157412786701368836335103632684358072471547044545424269809446594105817965243578174982010679;
            6'd10: xpb[6] = 1024'd74535929794263062991634887210220100254977530050561836487257842987471283780194006971513475669054005867031154692025947843873883199259645999542141848254073819124806592085783729129312303293536591755031049926383399236792724997223494900616475292196582737849778258791879298484791578529072843360903021676472466449346;
            6'd11: xpb[6] = 1024'd7549505363214524451519019488353450633656226780176609659104514247232274955827924322655780507164801868068380516754046567513833214680878398763259958069682576477072846552619371639665390107979927497748036353989395252653380986813306326899135679606303342074664142622596993515206819537622947886722109948144356403682;
            6'd12: xpb[6] = 1024'd64629776616290727310202079171301233757033350635527066959083040571970161468770980583813156559933272178548755748939638725732847070943331132539538192901622374763029775589026231487648716113940468961775220389982631114878397826624014526146774636699253395566369929867431746575728588620101685429659888046441840842349;
            6'd13: xpb[6] = 1024'd121710047869366930168885138854249016880410474490877524259061566896708047981714036844970532612701742489029130981125230883951860927205783866315816427733562173048986704625433091335632042119901010425802404425975866977103414666434722725394413593792203449058075717112266499636250357702580422972597666144739325281016;
            6'd14: xpb[6] = 1024'd54723623438318391628769271132382367259089171220492297430908238156469039157347954196112837450812538490066356805853329607591810942627016265536934537549170930401252959092268733845985128934344346168519390853581862992964070656024534151677073981201924053282961600942984194666665598711130527498416754416411215235352;
            6'd15: xpb[6] = 1024'd111803894691394594487452330815330150382466295075842754730886764481206925670291010457270213503581008800546732038038921765810824798889468999313212772381110728687209888128675593693968454940304887632546574889575098855189087495835242350924712938294874106774667388187818947727187367793609265041354532514708699674019;
            6'd16: xpb[6] = 1024'd44817470260346055947336463093463500761144991805457527902733435740967916845924927808412518341691804801583957862767020489450774814310701398534330882196719486039476142595511236204321541754748223375263561317181094871049743485425053777207373325704594710999553272018536642757602608802159369567173620786380589628355;
            6'd17: xpb[6] = 1024'd101897741513422258806019522776411283884522115660807985202711962065705803358867984069569894394460275112064333094952612647669788670573154132310609117028659284325433071631918096052304867760708764839290745353174330733274760325235761976455012282797544764491259059263371395818124377884638107110111398884678074067022;
            6'd18: xpb[6] = 1024'd34911317082373720265903655054544634263200812390422758374558633325466794534501901420712199232571071113101558919680711371309738685994386531531727226844268041677699326098753738562657954575152100582007731780780326749135416314825573402737672670207265368716144943094089090848539618893188211635930487156349964021358;
            6'd19: xpb[6] = 1024'd91991588335449923124586714737492417386577936245773215674537159650204681047444957681869575285339541423581934151866303529528752542256839265308005461676207839963656255135160598410641280581112642046034915816773562611360433154636281601985311627300215422207850730338923843909061387975666949178868265254647448460025;
            6'd20: xpb[6] = 1024'd25005163904401384584470847015625767765256632975387988846383830909965672223078875033011880123450337424619159976594402253168702557678071664529123571491816597315922509601996240920994367395555977788751902244379558627221089144226093028267972014709936026432736614169641538939476628984217053704687353526319338414361;
            6'd21: xpb[6] = 1024'd82085435157477587443153906698573550888633756830738446146362357234703558736021931294169256176218807735099535208779994411387716413940524398305401806323756395601879438638403100768977693401516519252779086280372794489446105984036801227515610971802886079924442401414476291999998398066695791247625131624616822853028;
            6'd22: xpb[6] = 1024'd15099010726429048903038038976706901267312453560353219318209028494464549911655848645311561014329603736136761033508093135027666429361756797526519916139365152954145693105238743279330780215959854995496072707978790505306761973626612653798271359212606684149328285245193987030413639075245895773444219896288712807364;
            6'd23: xpb[6] = 1024'd72179281979505251761721098659654684390689577415703676618187554819202436424598904906468937067098074046617136265693685293246680285624209531302798150971304951240102622141645603127314106221920396459523256743972026367531778813437320853045910316305556737641034072490028740090935408157724633316381997994586197246031;
            6'd24: xpb[6] = 1024'd5192857548456713221605230937788034769368274145318449790034226078963427600232822257611241905208870047654362090421784016886630301045441930523916260786913708592368876608481245637667193036363732202240243171578022383392434803027132279328570703715277341865919956320746435121350649166274737842201086266258087200367;
            6'd25: xpb[6] = 1024'd62273128801532916080288290620735817892745398000668907090012752403701314113175878518768617957977340358134737322607376175105644157307894664300194495618853506878325805644888105485650519042324273666267427207571258245617451642837840478576209660808227395357625743565581188181872418248753475385138864364555571639034;
            6'd26: xpb[6] = 1024'd119353400054609118938971350303683601016122521856019364389991278728439200626118934779925994010745810668615112554792968333324658013570347398076472730450793305164282734681294965333633845048284815130294611243564494107842468482648548677823848617901177448849331530810415941242394187331232212928076642462853056077701;
            6'd27: xpb[6] = 1024'd52366975623560580398855482581816951394801218585634137561837949988200191801752852131068298848856606669652338379521067056964608028991579797297590840266402062516548989148130607843986931862728150873011597671170490123703124472238360104106509005310898053074217414641133636272809428339782317453895730734524946032037;
            6'd28: xpb[6] = 1024'd109447246876636783257538542264764734518178342440984594861816476312938078314695908392225674901625076980132713611706659215183621885254032531073869075098341860802505918184537467691970257868688692337038781707163725985928141312049068303354147962403848106565923201885968389333331197422261054996833508832822430470704;
            6'd29: xpb[6] = 1024'd42460822445588244717422674542898084896857039170599368033663147572699069490329825743367979739735872981169939436434757938823571900675264930294987184913950618154772172651373110202323344683132028079755768134769722001788797301638879729636808349813568710790809085716686084363746438430811159522652597104494320425040;
            6'd30: xpb[6] = 1024'd99541093698664447576105734225845868020234163025949825333641673897436956003272882004525355792504343291650314668620350097042585756937717664071265419745890416440729101687779970050306670689092569543782952170762957864013814141449587928884447306906518764282514872961520837424268207513289897065590375202791804863707;
            6'd31: xpb[6] = 1024'd32554669267615909035989866503979218398912859755564598505488345157197947178906799355667660630615139292687540493348448820682535772358950063292383529561499173792995356154615612560659757503535905286499938598368953879874470131039399355167107694316239368507400756792238532454683448521840001591409463474463694818043;
            6'd32: xpb[6] = 1024'd89634940520692111894672926186927001522289983610915055805466871481935833691849855616825036683383609603167915725534040978901549628621402797068661764393438972078952285191022472408643083509496446750527122634362189742099486970850107554414746651409189421999106544037073285515205217604318739134347241572761179256710;
            6'd33: xpb[6] = 1024'd22648516089643573354557058465060351900968680340529828977313542741696824867483772967967341521494405604205141550262139702541499644042635196289779874209047729431218539657858114918996170323939782493244109061968185757960142960439918980697407038818910026223992427867790980545620458612868843660166329844433069211046;
            6'd34: xpb[6] = 1024'd79728787342719776213240118148008135024345804195880286277292069066434711380426829229124717574262875914685516782447731860760513500305087930066058109040987527717175468694264974766979496329900323957271293097961421620185159800250627179945045995911860079715698215112625733606142227695347581203104107942730553649713;
            6'd35: xpb[6] = 1024'd12742362911671237673124250426141485403024500925495059449138740326195702556060746580267022412373671915722742607175830584400463515726320329287176218856596285069441723161100617277332583144343659699988279525567417636045815789840438606227706383321580683940584098943343428636557468703897685728923196214402443604049;
            6'd36: xpb[6] = 1024'd69822634164747440531807310109089268526401624780845516749117266650933589069003802841424398465142142226203117839361422742619477371988773063063454453688536083355398652197507477125315909150304201164015463561560653498270832629651146805475345340414530737432289886188178181697079237786376423271860974312699928042716;
            6'd37: xpb[6] = 1024'd2836209733698901991691442387222618905080321510460289920963937910694580244637720192566703303252938227240343664089521466259427387410005462284572563504144840707664906664343119635668995964747536906732449989166649514131488619240958231758005727824251341657175770018895876727494478794926527797680062584371817997052;
            6'd38: xpb[6] = 1024'd59916480986775104850374502070170402028457445365810747220942464235432466757580776453724079356021408537720718896275113624478441243672458196060850798336084638993621835700749979483652321970708078370759634025159885376356505459051666431005644684917201395148881557263730629788016247877405265340617840682669302435719;
            6'd39: xpb[6] = 1024'd116996752239851307709057561753118185151834569221161204520920990560170353270523832714881455408789878848201094128460705782697455099934910929837129033168024437279578764737156839331635647976668619834786818061153121238581522298862374630253283642010151448640587344508565382848538016959884002883555618780966786874386;
            6'd40: xpb[6] = 1024'd50010327808802769168941694031251535530513265950775977692767661819931344446157750066023760246900674849238319953188804506337405115356143329058247142983633194631845019203992481841988734791111955577503804488759117254442178288452186056535944029419872052865473228339283077878953257968434107409374707052638676828722;
            6'd41: xpb[6] = 1024'd107090599061878972027624753714199318653890389806126434992746188144669230959100806327181136299669145159718695185374396664556418971618596062834525377815572992917801948240399341689972060797072497041530988524752353116667195128262894255783582986512822106357179015584117830939475027050912844952312485150936161267389;
            6'd42: xpb[6] = 1024'd40104174630830433487508885992332669032569086535741208164592859404430222134734723678323441137779941160755921010102495388196368987039828462055643487631181750270068202707234984200325147611515832784247974952358349132527851117852705682066243373922542710582064899414835525969890268059462949478131573422608051221725;
            6'd43: xpb[6] = 1024'd97184445883906636346191945675280452155946210391091665464571385729168108647677779939480817190548411471236296242288087546415382843302281195831921722463121548556025131743641844048308473617476374248275158988351584994752867957663413881313882331015492764073770686659670279030412037141941687021069351520905535660392;
            6'd44: xpb[6] = 1024'd30198021452858097806076077953413802534624907120706438636418056988929099823311697290623122028659207472273522067016186270055332858723513595053039832278730305908291386210477486558661560431919709990992145415957581010613523947253225307596542718425213368298656570490387974060827278150491791546888439792577425614728;
            6'd45: xpb[6] = 1024'd87278292705934300664759137636361585658002030976056895936396583313666986336254753551780498081427677782753897299201778428274346714985966328829318067110670104194248315246884346406644886437880251455019329451950816872838540787063933506844181675518163421790362357735222727121349047232970529089826217890874910053395;
            6'd46: xpb[6] = 1024'd20291868274885762124643269914494936036680727705671669108243254573427977511888670902922802919538473783791123123929877151914296730407198728050436176926278861546514569713719988916997973252323587197736315879556812888699196776653744933126842062927884026015248241565940422151764288241520633615645306162546800007731;
            6'd47: xpb[6] = 1024'd77372139527961964983326329597442719160057851561022126408221780898165864024831727164080178972306944094271498356115469310133310586669651461826714411758218659832471498750126848764981299258284128661763499915550048750924213616464453132374481020020834079506954028810775175212286057323999371158583084260844284446398;
            6'd48: xpb[6] = 1024'd10385715096913426443210461875576069538736548290636899580068452157926855200465644515222483810417740095308724180843568033773260602090883861047832521573827417184737753216962491275334386072727464404480486343156044766784869606054264558657141407430554683731839912641492870242701298332549475684402172532516174400734;
            6'd49: xpb[6] = 1024'd67465986349989629301893521558523852662113672145987356880046978482664741713408700776379859863186210405789099413029160191992274458353336594824110756405767215470694682253369351123317712078688005868507670379149280629009886445864972757904780364523504737223545699886327623303223067415028213227339950630813658839401;
            6'd50: xpb[6] = 1024'd479561918941090761777653836657203040792368875602130051893649742425732889042618127522164701297006406826325237757258915632224473774568994045228866221375972822960936720204993633670798893131341611224656806755276644870542435454784184187440751933225341448431583717045318333638308423578317753159038902485548793737;
            6'd51: xpb[6] = 1024'd57559833172017293620460713519604986164169492730952587351872176067163619401985674388679540754065476717306700469942851073851238330037021727821507101053315771108917865756611853481654124899091883075251840842748512507095559275265492383435079709026175394940137370961880071394160077506057055296096817000783033232404;
            6'd52: xpb[6] = 1024'd114640104425093496479143773202552769287546616586303044651850702391901505914928730649836916806833947027787075702128443232070252186299474461597785335885255569394874794793018713329637450905052424539279024878741748369320576115076200582682718666119125448431843158206714824454681846588535792839034595099080517671071;
            6'd53: xpb[6] = 1024'd47653679994044957939027905480686119666225313315917817823697373651662497090562648000979221644944743028824301526856541955710202201720706860818903445700864326747141049259854355839990537719495760281996011306347744385181232104666012008965379053528846052656729042037432519485097087597085897364853683370752407625407;
            6'd54: xpb[6] = 1024'd104733951247121160797710965163633902789602437171268275123675899976400383603505704262136597697713213339304676759042134113929216057983159594595181680532804125033097978296261215687973863725456301746023195342340980247406248944476720208213018010621796106148434829282267272545618856679564634907791461469049892064074;
            6'd55: xpb[6] = 1024'd37747526816072622257595097441767253168281133900883048295522571236161374779139621613278902535824009340341902583770232837569166073404391993816299790348412882385364232763096858198326950539899637488740181769946976263266904934066531634495678398031516710373320713112984967576034097688114739433610549740721782018410;
            6'd56: xpb[6] = 1024'd94827798069148825116278157124715036291658257756233505595501097560899261292082677874436278588592479650822277815955824995788179929666844727592578025180352680671321161799503718046310276545860178952767365805940212125491921773877239833743317355124466763865026500357819720636555866770593476976548327839019266457077;
            6'd57: xpb[6] = 1024'd27841373638100286576162289402848386670336954485848278767347768820660252467716595225578583426703275651859503640683923719428129945088077126813696134995961438023587416266339360556663363360303514695484352233546208141352577763467051260025977742534187368089912384188537415666971107779143581502367416110691156411413;
            6'd58: xpb[6] = 1024'd84921644891176489434845349085796169793714078341198736067326295145398138980659651486735959479471745962339878872869515877647143801350529860589974369827901236309544345302746220404646689366264056159511536269539444003577594603277759459273616699627137421581618171433372168727492876861622319045305194208988640850080;
            6'd59: xpb[6] = 1024'd17935220460127950894729481363929520172392775070813509239172966405159130156293568837878264317582541963377104697597614601287093816771762259811092479643509993661810599769581862914999776180707391902228522697145440019438250592867570885556277087036858025806504055264089863757908117870172423571124282480660530804416;
            6'd60: xpb[6] = 1024'd75015491713204153753412541046877303295769898926163966539151492729897016669236625099035640370351012273857479929783206759506107673034214993587370714475449791947767528805988722762983102186667933366255706733138675881663267432678279084803916044129808079298209842508924616818429886952651161114062060578958015243083;
            6'd61: xpb[6] = 1024'd8029067282155615213296673325010653674448595655778739710998163989658007844870542450177945208461808274894705754511305483146057688455447392808488824291058549300033783272824365273336189001111269108972693160744671897523923422268090511086576431539528683523095726339642311848845127961201265639881148850629905197419;
            6'd62: xpb[6] = 1024'd65109338535231818071979733007958436797825719511129197010976690314395894357813598711335321261230278585375080986696897641365071544717900126584767059122998347585990712309231225121319515007071810572999877196737907759748940262078798710334215388632478737014801513584477064909366897043680003182818926948927389636086;
            6'd63: xpb[6] = 1024'd122189609788308020930662792690906219921202843366479654310955216639133780870756654972492697313998748895855456218882489799584085400980352860361045293954938145871947641345638084969302841013032352037027061232731143621973957101889506909581854345725428790506507300829311817969888666126158740725756705047224874074753;
        endcase
    end

    always_comb begin
        case(flag[2][11:6])
            6'd0: xpb[7] = 1024'd0;
            6'd1: xpb[7] = 1024'd55203185357259482390546924969039570299881540096094427482801887898894772046390572323635002152109544896892682043610588523224035416401585259582163403770546903224213895812473727479655927827475687779744047660337139637834613091479318335864514733135149394731393184660029513000303907134708845251575793318896764029089;
            6'd2: xpb[7] = 1024'd110406370714518964781093849938079140599763080192188854965603775797789544092781144647270004304219089793785364087221177046448070832803170519164326807541093806448427791624947454959311855654951375559488095320674279275669226182958636671729029466270298789462786369320059026000607814269417690503151586637793528058178;
            6'd3: xpb[7] = 1024'd41542860387653705772841847502304278154946193162547598320273808631707420801862578060889935241670960381234896723374272135093042408363535444191330086295309668738951012867849965101337544290909857617921945372624179067139478424217058234628565629722218734927359650565971480970805193330197902737608690130064697602936;
            6'd4: xpb[7] = 1024'd96746045744913188163388772471343848454827733258642025803075696530602192848253150384524937393780505278127578766984860658317077824765120703773493490065856571963164908680323692580993472118385545397665993032961318704974091515696376570493080362857368129658752835226000993971109100464906747989184483448961461632025;
            6'd5: xpb[7] = 1024'd27882535418047929155136770035568986010010846229000769157745729364520069557334583798144868331232375865577111403137955746962049400325485628800496768820072434253688129923226202723019160754344027456099843084911218496444343756954798133392616526309288075123326116471913448941306479525686960223641586941232631176783;
            6'd6: xpb[7] = 1024'd83085720775307411545683695004608556309892386325095196640547617263414841603725156121779870483341920762469793446748544270186084816727070888382660172590619337477902025735699930202675088581819715235843890745248358134278956848434116469257131259444437469854719301131942961941610386660395805475217380260129395205872;
            6'd7: xpb[7] = 1024'd14222210448442152537431692568833693865075499295453939995217650097332718312806589535399801420793791349919326082901639358831056392287435813409663451344835199768425246978602440344700777217778197294277740797198257925749209089692538032156667422896357415319292582377855416911807765721176017709674483752400564750630;
            6'd8: xpb[7] = 1024'd69425395805701634927978617537873264164957039391548367478019537996227490359197161859034803572903336246812008126512227882055091808689021072991826855115382102992639142791076167824356705045253885074021788457535397563583822181171856368021182156031506810050685767037884929912111672855884862961250277071297328779719;
            6'd9: xpb[7] = 1024'd561885478836375919726615102098401720140152361907110832689570830145367068278595272654734510355206834261540762665322970700063384249385998018830133869597965283162364033978677966382393681212367132455638509485297355054074422430277930920718319483426755515259048283797384882309051916665075195707380563568498324477;
            6'd10: xpb[7] = 1024'd55765070836095858310273540071137972020021692458001538315491458729040139114669167596289736662464751731154222806275911493924098800650971257600993537640144868507376259846452405446038321508688054912199686169822436992888687513909596266785233052618576150246652232943826897882612959051373920447283173882465262353566;
            6'd11: xpb[7] = 1024'd110968256193355340700820465040177542319903232554095965798293346627934911161059739919924738814574296628046904849886500017148134217052556517183156941410691771731590155658926132925694249336163742691943733830159576630723300605388914602649747785753725544978045417603856410882916866186082765698858967201362026382655;
            6'd12: xpb[7] = 1024'd42104745866490081692568462604402679875086345524454709152963379461852787870141173333544669752026167215496437486039595105793105792612921442210160220164907634022113376901828643067719937972122224750377583882109476422193552846647336165549283949205645490442618698849768865853114245246862977933316070693633195927413;
            6'd13: xpb[7] = 1024'd97307931223749564083115387573442250174967885620549136635765267360747559916531745657179671904135712112389119529650183629017141209014506701792323623935454537246327272714302370547375865799597912530121631542446616060028165938126654501413798682340794885174011883509798378853418152381571823184891864012529959956502;
            6'd14: xpb[7] = 1024'd28444420896884305074863385137667387730150998590907879990435300194665436625613179070799602841587582699838652165803278717662112784574871626819326902689670399536850493957204880689401554435556394588555481594396515851498418179385076064313334845792714830638585164755710833823615531442352035419348967504801129501260;
            6'd15: xpb[7] = 1024'd83647606254143787465410310106706958030032538687002307473237188093560208672003751394434604993697127596731334209413867240886148200976456886401490306460217302761064389769678608169057482263032082368299529254733655489333031270864394400177849578927864225369978349415740346823919438577060880670924760823697893530349;
            6'd16: xpb[7] = 1024'd14784095927278528457158307670932095585215651657361050827907220927478085381085184808054535931148998184180866845566962329531119776536821811428493585214433165051587611012581118311083170898990564426733379306683555280803283512122815963077385742379784170834551630661652801794116817637841092905381864315969063075107;
            6'd17: xpb[7] = 1024'd69987281284538010847705232639971665885097191753455478310709108826372857427475757131689538083258543081073548889177550852755155192938407071010656988984980068275801506825054845790739098726466252206477426967020694918637896603602134298941900475514933565565944815321682314794420724772549938156957657634865827104196;
            6'd18: xpb[7] = 1024'd1123770957672751839453230204196803440280304723814221665379141660290734136557190545309469020710413668523081525330645941400126768498771996037660267739195930566324728067957355932764787362424734264911277018970594710108148844860555861841436638966853511030518096567594769764618103833330150391414761127136996648954;
            6'd19: xpb[7] = 1024'd56326956314932234230000155173236373740161844819908649148181029559185506182947762868944471172819958565415763568941234464624162184900357255619823671509742833790538623880431083412420715189900422044655324679307734347942761936339874197705951372102002905761911281227624282764922010968038995642990554446033760678043;
            6'd20: xpb[7] = 1024'd111530141672191716620547080142275944040043384916003076630982917458080278229338335192579473324929503462308445612551822987848197601301942515201987075280289737014752519692904810892076643017376109824399372339644873985777375027819192533570466105237152300493304465887653795765225918102747840894566347764930524707132;
            6'd21: xpb[7] = 1024'd42666631345326457612295077706501081595226497886361819985652950291998154938419768606199404262381374049757978248704918076493169176862307440228990354034505599305275740935807321034102331653334591882833222391594773777247627269077614096470002268689072245957877747133566250735423297163528053129023451257201694251890;
            6'd22: xpb[7] = 1024'd97869816702585940002842002675540651895108037982456247468454838190892926984810340929834406414490918946650660292315506599717204593263892699811153757805052502529489636748281048513758259480810279662577270051931913415082240360556932432334517001824221640689270931793595763735727204298236898380599244576098458280979;
            6'd23: xpb[7] = 1024'd29006306375720680994590000239765789450291150952814990823124871024810803693891774343454337351942789534100192928468601688362176168824257624838157036559268364820012857991183558655783948116768761721011120103881813206552492601815353995234053165276141586153844213039508218705924583359017110615056348068369627825737;
            6'd24: xpb[7] = 1024'd84209491732980163385136925208805359750172691048909418305926758923705575740282346667089339504052334430992874972079190211586211585225842884420320440329815268044226753803657286135439875944244449500755167764218952844387105693294672331098567898411290980885237397699537731706228490493725955866632141387266391854826;
            6'd25: xpb[7] = 1024'd15345981406114904376884922773030497305355804019268161660596791757623452449363780080709270441504205018442407608232285300231183160786207809447323719084031130334749975046559796277465564580202931559189017816168852635857357934553093893998104061863210926349810678945450186676425869554506168101089244879537561399584;
            6'd26: xpb[7] = 1024'd70549166763374386767431847742070067605237344115362589143398679656518224495754352404344272593613749915335089651842873823455218577187793069029487122854578033558963870859033523757121492407678619338933065476505992273691971026032412229862618794998360321081203863605479699676729776689215013352665038198434325428673;
            6'd27: xpb[7] = 1024'd1685656436509127759179845306295205160420457085721332498068712490436101204835785817964203531065620502784622287995968912100190152748157994056490401608793895849487092101936033899147181043637101397366915528455892065162223267290833792762154958450280266545777144851392154646927155749995225587122141690705494973431;
            6'd28: xpb[7] = 1024'd56888841793768610149726770275334775460301997181815759980870600389330873251226358141599205683175165399677304331606557435324225569149743253638653805379340799073700987914409761378803108871112789177110963188793031702996836358770152128626669691585429661277170329511421667647231062884704070838697935009602259002520;
            6'd29: xpb[7] = 1024'd112092027151028092540273695244374345760183537277910187463672488288225645297616930465234207835284710296569986375217145958548260985551328513220817209149887702297914883726883488858459036698588476956855010849130171340831449450249470464491184424720579056008563514171451180647534970019412916090273728328499023031609;
            6'd30: xpb[7] = 1024'd43228516824162833532021692808599483315366650248268930818342521122143522006698363878854138772736580884019519011370241047193232561111693438247820487904103564588438104969785999000484725334546959015288860901080071132301701691507892027390720588172499001473136795417363635617732349080193128324730831820770192576367;
            6'd31: xpb[7] = 1024'd98431702181422315922568617777639053615248190344363358301144409021038294053088936202489140924846125780912201054980829570417267977513278697829983891674650467812652000782259726480140653162022646795032908561417210770136314782987210363255235321307648396204529980077393148618036256214901973576306625139666956605456;
            6'd32: xpb[7] = 1024'd29568191854557056914316615341864191170431303314722101655814441854956170762170369616109071862297996368361733691133924659062239553073643622856987170428866330103175222025162236622166341797981128853466758613367110561606567024245631926154771484759568341669103261323305603588233635275682185810763728631938126150214;
            6'd33: xpb[7] = 1024'd84771377211816539304863540310903761470312843410816529138616329753850942808560941939744074014407541265254415734744513182286274969475228882439150574199413233327389117837635964101822269625456816633210806273704250199441180115724950262019286217894717736400496445983335116588537542410391031062339521950834890179303;
            6'd34: xpb[7] = 1024'd15907866884951280296611537875128899025495956381175272493286362587768819517642375353364004951859411852703948370897608270931246545035593807466153852953629095617912339080538474243847958261415298691644656325654149990911432356983371824918822381346637681865069727229247571558734921471171243296796625443106059724061;
            6'd35: xpb[7] = 1024'd71111052242210762687158462844168469325377496477269699976088250486663591564032947676999007103968956749596630414508196794155281961437179067048317256724175998842126234893012201723503886088890986471388703985991289628746045448462690160783337114481787076596462911889277084559038828605880088548372418762002823753150;
            6'd36: xpb[7] = 1024'd2247541915345503678906460408393606880560609447628443330758283320581468273114381090618938041420827337046163050661291882800253536997543992075320535478391861132649456135914711865529574724849468529822554037941189420216297689721111723682873277933707022061036193135189539529236207666660300782829522254273993297908;
            6'd37: xpb[7] = 1024'd57450727272604986069453385377433177180442149543722870813560171219476240319504953414253940193530372233938845094271880406024288953399129251657483939248938764356863351948388439345185502552325156309566601698278329058050910781200430059547388011068856416792429377795219052529540114801369146034405315573170757326997;
            6'd38: xpb[7] = 1024'd112653912629864468460000310346472747480323689639817298296362059118371012365895525737888942345639917130831527137882468929248324369800714511239647343019485667581077247760862166824841430379800844089310649358615468695885523872679748395411902744204005811523822562455248565529844021936077991285981108892067521356086;
            6'd39: xpb[7] = 1024'd43790402302999209451748307910697885035506802610176041651032091952288889074976959151508873283091787718281059774035564017893295945361079436266650621773701529871600469003764676966867119015759326147744499410565368487355776113938169958311438907655925756988395843701161020500041400996858203520438212384338690900844;
            6'd40: xpb[7] = 1024'd98993587660258691842295232879737455335388342706270469133833979851183661121367531475143875435201332615173741817646152541117331361762664695848814025544248433095814364816238404446523046843235013927488547070902508125190389205417488294175953640791075151719789028361190533500345308131567048772014005703235454929933;
            6'd41: xpb[7] = 1024'd30130077333393432834043230443962592890571455676629212488504012685101537830448964888763806372653203202623274453799247629762302937323029620875817304298464295386337586059140914588548735479193495985922397122852407916660641446675909857075489804242995097184362309607102988470542687192347261006471109195506624474691;
            6'd42: xpb[7] = 1024'd85333262690652915224590155413002163190452995772723639971305900583996309876839537212398808524762748099515956497409836152986338353724614880457980708069011198610551481871614642068204663306669183765666444783189547554495254538155228192940004537378144491915755494267132501470846594327056106258046902514403388503780;
            6'd43: xpb[7] = 1024'd16469752363787656216338152977227300745636108743082383325975933417914186585920970626018739462214618686965489133562931241631309929284979805484983986823227060901074703114517152210230351942627665824100294835139447345965506779413649755839540700830064437380328775513044956441043973387836318492504006006674558048538;
            6'd44: xpb[7] = 1024'd71672937721047138606885077946266871045517648839176810808777821316808958632311542949653741614324163583858171177173519764855345345686565065067147390593773964125288598926990879689886279770103353603844342495476586983800119870892968091704055433965213832111721960173074469441347880522545163744079799325571322077627;
            6'd45: xpb[7] = 1024'd2809427394181879598633075510492008600700761809535554163447854150726835341392976363273672551776034171307703813326614853500316921246929990094150669347989826415811820169893389831911968406061835662278192547426486775270372112151389654603591597417133777576295241418986924411545259583325375978536902817842491622385;
            6'd46: xpb[7] = 1024'd58012612751441361989180000479531578900582301905629981646249742049621607387783548686908674703885579068200385856937203376724352337648515249676314073118536729640025715982367117311567896233537523442022240207763626413104985203630707990468106330552283172307688426079016437411849166718034221230112696136739255651474;
            6'd47: xpb[7] = 1024'd113215798108700844379726925448571149200463842001724409129051629948516379434174121010543676855995123965093067900547791899948387754050100509258477476889083632864239611794840844791223824061013211221766287868100766050939598295110026326332621063687432567039081610739045950412153073852743066481688489455636019680563;
            6'd48: xpb[7] = 1024'd44352287781835585371474923012796286755646954972083152483721662782434256143255554424163607793446994552542600536700886988593359329610465434285480755643299495154762833037743354933249512696971693280200137920050665842409850536368447889232157227139352512503654891984958405382350452913523278716145592947907189225321;
            6'd49: xpb[7] = 1024'd99555473139095067762021847981835857055528495068177579966523550681329028189646126747798609945556539449435282580311475511817394746012050693867644159413846398378976728850217082412905440524447381059944185580387805480244463627847766225096671960274501907235048076644987918382654360048232123967721386266803953254410;
            6'd50: xpb[7] = 1024'd30691962812229808753769845546060994610711608038536323321193583515246904898727560161418540883008410036884815216464570600462366321572415618894647438168062260669499950093119592554931129160405863118378035632337705271714715869106187787996208123726421852699621357890900373352851739109012336202178489759075122799168;
            6'd51: xpb[7] = 1024'd85895148169489291144316770515100564910593148134630750803995471414141676945118132485053543035117954933777497260075159123686401737974000878476810841938609163893713845905593320034587056987881550898122083292674844909549328960585506123860722856861571247431014542550929886353155646243721181453754283077971886828257;
            6'd52: xpb[7] = 1024'd17031637842624032136064768079325702465776261104989494158665504248059553654199565898673473972569825521227029896228254212331373313534365803503814120692825026184237067148495830176612745623840032956555933344624744701019581201843927686760259020313491192895587823796842341323353025304501393688211386570243056373015;
            6'd53: xpb[7] = 1024'd72234823199883514526611693048365272765657801201083921641467392146954325700590138222308476124679370418119711939838842735555408729935951063085977524463371929408450962960969557656268673451315720736299981004961884338854194293323246022624773753448640587626981008456871854323656932439210238939787179889139820402104;
            6'd54: xpb[7] = 1024'd3371312873018255518359690612590410320840914171442664996137424980872202409671571635928407062131241005569244575991937824200380305496315988112980803217587791698974184203872067798294362087274202794733831056911784130324446534581667585524309916900560533091554289702784309293854311499990451174244283381410989946862;
            6'd55: xpb[7] = 1024'd58574498230277737908906615581629980620722454267537092478939312879766974456062143959563409214240785902461926619602526347424415721897901247695144206988134694923188080016345795277950289914749890574477878717248923768159059626060985921388824650035709927822947474362813822294158218634699296425820076700307753975951;
            6'd56: xpb[7] = 1024'd113777683587537220299453540550669550920603994363631519961741200778661746502452716283198411366350330799354608663213114870648451138299486507277307610758681598147401975828819522757606217742225578354221926377586063405993672717540304257253339383170859322554340659022843335294462125769408141677395870019204518005040;
            6'd57: xpb[7] = 1024'd44914173260671961291201538114894688475787107333990263316411233612579623211534149696818342303802201386804141299366209959293422713859851432304310889512897460437925197071722032899631906378184060412655776429535963197463924958798725820152875546622779268018913940268755790264659504830188353911852973511475687549798;
            6'd58: xpb[7] = 1024'd100117358617931443681748463083934258775668647430084690799213121511474395257924722020453344455911746283696823342976798482517458130261436691886474293283444363662139092884195760379287834205659748192399824089873102835298538050278044156017390279757928662750307124928785303264963411964897199163428766830372451578887;
            6'd59: xpb[7] = 1024'd31253848291066184673496460648159396330851760400443434153883154345392271967006155434073275393363616871146355979129893571162429705821801616913477572037660225952662314127098270521313522841618230250833674141823002626768790291536465718916926443209848608214880406174697758235160791025677411397885870322643621123645;
            6'd60: xpb[7] = 1024'd86457033648325667064043385617198966630733300496537861636685042244287044013396727757708277545473161768039038022740482094386465122223386876495640975808207129176876209939571998000969450669093918030577721802160142264603403383015784054781441176344998002946273590834727271235464698160386256649461663641540385152734;
            6'd61: xpb[7] = 1024'd17593523321460408055791383181424104185916413466896604991355075078204920722478161171328208482925032355488570658893577183031436697783751801522644254562422991467399431182474508142995139305052400089011571854110042056073655624274205617680977339796917948410846872080639726205662077221166468883918767133811554697492;
            6'd62: xpb[7] = 1024'd72796708678719890446338308150463674485797953562991032474156962977099692768868733494963210635034577252381252702504165706255472114185337061104807658332969894691613326994948235622651067132528087868755619514447181693908268715753523953545492072932067343142240056740669239205965984355875314135494560452708318726581;
            6'd63: xpb[7] = 1024'd3933198351854631438086305714688812040981066533349775828826995811017569477950166908583141572486447839830785338657260794900443689745701986131810937087185756982136548237850745764676755768486569927189469566397081485378520957011945516445028236383987288606813337986581694176163363416655526369951663944979488271339;
        endcase
    end

    always_comb begin
        case(flag[2][16:12])
            5'd0: xpb[8] = 1024'd0;
            5'd1: xpb[8] = 1024'd59136383709114113828633230683728382340862606629444203311628883709912341524340739232218143724595992736723467382267849318124479106147287245713974340857732660206350444050324473244332683595962257706933517226734221123213134048491263852309542969519136683338206522646611207176467270551364371621527457263876252300428;
            5'd2: xpb[8] = 1024'd118272767418228227657266461367456764681725213258888406623257767419824683048681478464436287449191985473446934764535698636248958212294574491427948681715465320412700888100648946488665367191924515413867034453468442246426268096982527704619085939038273366676413045293222414352934541102728743243054914527752504600856;
            5'd3: xpb[8] = 1024'd53342455443217600087100764646370714277889392762596925806754796064760129235713078786639359959130303900727252739346054519794373477600641402586762897556866939685360657581402202395367811596369567399490354071815423523275041295252894783963650338874180600747799664525716563499295283580164481847463681965003162416953;
            5'd4: xpb[8] = 1024'd112478839152331713915733995330099096618751999392041129118383679774672470760053818018857503683726296637450720121613903837918852583747928648300737238414599599891711101631726675639700495192331825106423871298549644646488175343744158636273193308393317284086006187172327770675762554131528853468991139228879414717381;
            5'd5: xpb[8] = 1024'd47548527177321086345568298609013046214916178895749648301880708419607916947085418341060576193664615064731038096424259721464267849053995559459551454256001219164370871112479931546402939596776877092047190916896625923336948542014525715617757708229224518157392806404821919822123296608964592073399906666130072533478;
            5'd6: xpb[8] = 1024'd106684910886435200174201529292741428555778785525193851613509592129520258471426157573278719918260607801454505478692109039588746955201282805173525795113733879370721315162804404790735623192739134798980708143630847046550082590505789567927300677748361201495599329051433126998590567160328963694927363930006324833906;
            5'd7: xpb[8] = 1024'd41754598911424572604035832571655378151942965028902370797006620774455704658457757895481792428198926228734823453502464923134162220507349716332340010955135498643381084643557660697438067597184186784604027761977828323398855788776156647271865077584268435566985948283927276144951309637764702299336131367256982650003;
            5'd8: xpb[8] = 1024'd100890982620538686432669063255383760492805571658346574108635504484368046182798497127699936152794918965458290835770314241258641326654636962046314351812868158849731528693882133941770751193146444491537544988712049446611989837267420499581408047103405118905192470930538483321418580189129073920863588631133234950431;
            5'd9: xpb[8] = 1024'd35960670645528058862503366534297710088969751162055093292132533129303492369830097449903008662733237392738608810580670124804056591960703873205128567654269778122391298174635389848473195597591496477160864607059030723460763035537787578925972446939312352976579090163032632467779322666564812525272356068383892766528;
            5'd10: xpb[8] = 1024'd95097054354642172691136597218026092429832357791499296603761416839215833894170836682121152387329230129462076192848519442928535698107991118919102908512002438328741742224959863092805879193553754184094381833793251846673897084029051431235515416458449036314785612809643839644246593217929184146799813332260145066956;
            5'd11: xpb[8] = 1024'd30166742379631545120970900496940042025996537295207815787258445484151280081202437004324224897267548556742394167658875326473950963414058030077917124353404057601401511705713118999508323597998806169717701452140233123522670282299418510580079816294356270386172232042137988790607335695364922751208580769510802883053;
            5'd12: xpb[8] = 1024'd89303126088745658949604131180668424366859143924652019098887329194063621605543176236542368621863541293465861549926724644598430069561345275791891465211136717807751955756037592243841007193961063876651218678874454246735804330790682362889622785813492953724378754688749195967074606246729294372736038033387055183481;
            5'd13: xpb[8] = 1024'd24372814113735031379438434459582373963023323428360538282384357838999067792574776558745441131801859720746179524737080528143845334867412186950705681052538337080411725236790848150543451598406115862274538297221435523584577529061049442234187185649400187795765373921243345113435348724165032977144805470637712999578;
            5'd14: xpb[8] = 1024'd83509197822849145208071665143310756303885930057804741594013241548911409316915515790963584856397852457469646907004929846268324441014699432664680021910270997286762169287115321394876135194368373569208055523955656646797711577552313294543730155168536871133971896567854552289902619275529404598672262734513965300006;
            5'd15: xpb[8] = 1024'd18578885847838517637905968422224705900050109561513260777510270193846855503947116113166657366336170884749964881815285729813739706320766343823494237751672616559421938767868577301578579598813425554831375142302637923646484775822680373888294555004444105205358515800348701436263361752965143203081030171764623116103;
            5'd16: xpb[8] = 1024'd77715269556952631466539199105953088240912716190957464089139153903759197028287855345384801090932163621473432264083135047938218812468053589537468578609405276765772382818193050545911263194775683261764892369036859046859618824313944226197837524523580788543565038446959908612730632304329514824608487435640875416531;
            5'd17: xpb[8] = 1024'd12784957581942003896373502384867037837076895694665983272636182548694643215319455667587873600870482048753750238893490931483634077774120500696282794450806896038432152298946306452613707599220735247388211987383840323708392022584311305542401924359488022614951657679454057759091374781765253429017254872891533232628;
            5'd18: xpb[8] = 1024'd71921341291056117725006733068595420177939502324110186584265066258606984739660194899806017325466474785477217621161340249608113183921407746410257135308539556244782596349270779696946391195182992954321729214118061446921526071075575157851944893878624705953158180326065264935558645333129625050544712136767785533056;
            5'd19: xpb[8] = 1024'd6991029316045490154841036347509369774103681827818705767762094903542430926691795222009089835404793212757535595971696133153528449227474657569071351149941175517442365830024035603648835599628044939945048832465042723770299269345942237196509293714531940024544799558559414081919387810565363654953479574018443349153;
            5'd20: xpb[8] = 1024'd66127413025159603983474267031237752114966288457262909079390978613454772451032534454227233560000785949481002978239545451278007555374761903283045692007673835723792809880348508847981519195590302646878566059199263846983433317837206089506052263233668623362751322205170621258386658361929735276480936837894695649581;
            5'd21: xpb[8] = 1024'd1197101050148976413308570310151701711130467960971428262888007258390218638064134776430306069939104376761320953049901334823422820680828814441859907849075454996452579361101764754683963600035354632501885677546245123832206516107573168850616663069575857434137941437664770404747400839365473880889704275145353465678;
            5'd22: xpb[8] = 1024'd60333484759263090241941800993880084051993074590415631574516890968302560162404874008648449794535097113484788335317750652947901926828116060155834248706808115202803023411426237999016647195997612339435402904280466247045340564598837021160159632588712540772344464084275977581214671390729845502417161539021605766106;
            5'd23: xpb[8] = 1024'd119469868468377204070575031677608466392855681219859834886145774678214901686745613240866593519131089850208255717585599971072381032975403305869808589564540775409153467461750711243349330791959870046368920131014687370258474613090100873469702602107849224110550986730887184757681941942094217123944618802897858066534;
            5'd24: xpb[8] = 1024'd54539556493366576500409334956522415989019860723568354069642803323150347873777213563069666029069408277488573692395955854617796298281470217028622805405942394681813236942503967150051775196404922031992239749361668647107247811360467952814267001943756458181937605963381333904042684419529955728353386240148515882631;
            5'd25: xpb[8] = 1024'd113675940202480690329042565640250798329882467353012557381271687033062689398117952795287809753665401014212041074663805172742275404428757462742597146263675054888163680992828440394384458792367179738925756976095889770320381859851731805123809971462893141520144128609992541080509954970894327349880843504024768183059;
            5'd26: xpb[8] = 1024'd48745628227470062758876868919164747926046646856721076564768715677998135585149553117490882263603719441492359049474161056287690669734824373901411362105076674160823450473581696301086903196812231724549076594442871047169155058122098884468374371298800375591530747842486690226870697448330065954289610941275425999156;
            5'd27: xpb[8] = 1024'd107882011936584176587510099602893130266909253486165279876397599387910477109490292349709025988199712178215826431742010374412169775882111619615385702962809334367173894523906169545419586792774489431482593821177092170382289106613362736777917340817937058929737270489097897403337967999694437575817068205151678299584;
            5'd28: xpb[8] = 1024'd42951699961573549017344402881807079863073432989873799059894628032845923296521892671912098498138030605496144406552366257957585041188178530774199918804210953639833664004659425452122031197219541417105913439524073447231062304883729816122481740653844293001123889721592046549698710477130176180225835642402336115681;
            5'd29: xpb[8] = 1024'd102088083670687662845977633565535462203936039619318002371523511742758264820862631904130242222734023342219611788820215576082064147335465776488174259661943613846184108054983898696454714793181799124039430666258294570444196353374993668432024710172980976339330412368203253726165981028494547801753292906278588416109;
            5'd30: xpb[8] = 1024'd37157771695677035275811936844449411800100219123026521555020540387693711007894232226333314732672341769499929763630571459627479412641532687646988475503345233118843877535737154603157159197626851109662750284605275847292969551645360747776589110008888210410717031600697402872526723505930286406162060343529246232206;
            5'd31: xpb[8] = 1024'd96294155404791149104445167528177794140962825752470724866649424097606052532234971458551458457268334506223397145898420777751958518788819933360962816361077893325194321586061627847489842793589108816596267511339496970506103600136624600086132079528024893748923554247308610048993994057294658027689517607405498532634;
        endcase
    end

    always_comb begin
        case(flag[3][5:0])
            6'd0: xpb[9] = 1024'd0;
            6'd1: xpb[9] = 1024'd77715269556952631466539199105953088240912716190957464089139153903759197028287855345384801090932163621473432264083135047938218812468053589537468578609405276765772382818193050545911263194775683261764892369036859046859618824313944226197837524523580788543565038446959908612730632304329514824608487435640875416531;
            6'd2: xpb[9] = 1024'd31363843429780521534279470807091743737127005256179244050146452742541498719266571780754530967206652933503715120708776661297373784094886844519777032202479512597854091066814883754192287198034160802219587129686478247354876798406991679430696479363932127820310173479802759195354736534730396632098285044656156348731;
            6'd3: xpb[9] = 1024'd109079112986733153000818669913044831978039721447136708139285606646300695747554427126139332058138816554977147384791911709235592596562940434057245610811884789363626473885007934300103550392809844063984479498723337294214495622720935905628534003887512916363875211926762667808085368839059911456706772480297031765262;
            6'd4: xpb[9] = 1024'd62727686859561043068558941614183487474254010512358488100292905485082997438533143561509061934413305867007430241417553322594747568189773689039554064404959025195708182133629767508384574396068321604439174259372956494709753596813983358861392958727864255640620346959605518390709473069460793264196570089312312697462;
            6'd5: xpb[9] = 1024'd16376260732388933136299213315322142970468299577580268061300204323865299129511859996878791810687795179037713098043194935953902539816606944021862517998033261027789890382251600716665598399326799144893869020022575695205011570907030812094251913568215594917365481992448368973333577299861675071686367698327593629662;
            6'd6: xpb[9] = 1024'd94091530289341564602838412421275231211381015768537732150439358227624496157799715342263592901619958800511145362126329983892121352284660533559331096607438537793562273200444651262576861594102482406658761389059434742064630395220975038292089438091796383460930520439408277586064209604191189896294855133968469046193;
            6'd7: xpb[9] = 1024'd47740104162169454670578684122413886707595304833759512111446657066406797848778431777633322777894448112541428218751971597251276323911493788541639550200512773625643981449066484470857885597360959947113456149709053942559888369314022491524948392932147722737675655472251128168688313834592071703784652742983749978393;
            6'd8: xpb[9] = 1024'd1388678034997344738318955823552542203809593898981292072453955905189099539757148213003052654168937424571711075377613210610431295538327043523948003793587009457725689697688317679138909600619437487568150910358673143055146343407069944757807347772499062014420790505093978751312418064992953511274450351999030910593;
            6'd9: xpb[9] = 1024'd79103947591949976204858154929505630444722310089938756161593109808948296568045003558387853745101101046045143339460748258548650108006380633061416582402992286223498072515881368225050172795395120749333043279395532189914765167721014170955644872296079850557985828952053887364043050369322468335882937787639906327124;
            6'd10: xpb[9] = 1024'd32752521464777866272598426630644285940936599155160536122600408647730598259023719993757583621375590358075426196086389871907805079633213888043725035996066522055579780764503201433331196798653598289787738040045151390410023141814061624188503827136431189834730963984896737946667154599723350143372735396655187259324;
            6'd11: xpb[9] = 1024'd110467791021730497739137625736597374181849315346118000211739562551489795287311575339142384712307753979548858460169524919846023892101267477581193614605471798821352163582696251979242459993429281551552630409082010437269641966128005850386341351660011978378296002431856646559397786904052864967981222832296062675855;
            6'd12: xpb[9] = 1024'd64116364894558387806877897437736029678063604411339780172746861390272096978290291774512114588582243291579141316795166533205178863728100732563502068198546034653433871831318085187523483996687759092007325169731629637764899940221053303619200306500363317655041137464699497142021891134453746775471020441311343608055;
            6'd13: xpb[9] = 1024'd17764938767386277874618169138874685174277893476561560133754160229054398669269008209881844464856732603609424173420808146564333835354933987545810521791620270485515580079939918395804507999946236632462019930381248838260157914314100756852059261340714656931786272497542347724645995364854628582960818050326624540255;
            6'd14: xpb[9] = 1024'd95480208324338909341157368244827773415190609667519024222893314132813595697556863555266645555788896225082856437503943194502552647822987577083279100401025547251287962898132968941715771194721919894226912299418107885119776738628044983049896785864295445475351310944502256337376627669184143407569305485967499956786;
            6'd15: xpb[9] = 1024'd49128782197166799408897639945966428911404898732740804183900612971595897388535579990636375432063385537113139294129584807861707619449820832065587553994099783083369671146754802149996795197980397434681607060067727085615034712721092436282755740704646784752096445977345106920000731899585025215059103094982780888986;
            6'd16: xpb[9] = 1024'd2777356069994689476637911647105084407619187797962584144907911810378199079514296426006105308337874849143422150755226421220862591076654087047896007587174018915451379395376635358277819201238874975136301820717346286110292686814139889515614695544998124028841581010187957502624836129985907022548900703998061821186;
            6'd17: xpb[9] = 1024'd80492625626947320943177110753058172648531903988920048234047065714137396107802151771390906399270038470616854414838361469159081403544707676585364586196579295681223762213569685904189082396014558236901194189754205332969911511128084115713452220068578912572406619457147866115355468434315421847157388139638937237717;
            6'd18: xpb[9] = 1024'd34141199499775211010917382454196828144746193054141828195054364552919697798780868206760636275544527782647137271464003082518236375171540931567673039789653531513305470462191519112470106399273035777355888950403824533465169485221131568946311174908930251849151754489990716697979572664716303654647185748654218169917;
            6'd19: xpb[9] = 1024'd111856469056727842477456581560149916385658909245099292284193518456678894827068723552145437366476691404120569535547138130456455187639594521105141618399058808279077853280384569658381369594048719039120781319440683580324788309535075795144148699432511040392716792936950625310710204969045818479255673184295093586448;
            6'd20: xpb[9] = 1024'd65505042929555732545196853261288571881873198310321072245200817295461196518047439987515167242751180716150852392172779743815610159266427776087450071992133044111159561529006402866662393597307196579575476080090302780820046283628123248377007654272862379669461927969793475893334309199446700286745470793310374518648;
            6'd21: xpb[9] = 1024'd19153616802383622612937124962427227378087487375542852206208116134243498209026156422884897119025670028181135248798421357174765130893261031069758525585207279943241269777628236074943417600565674120030170840739921981315304257721170701609866609113213718946207063002636326475958413429847582094235268402325655450848;
            6'd22: xpb[9] = 1024'd96868886359336254079476324068380315619000203566500316295347270038002695237314011768269698209957833649654567512881556405112983943361314620607227104194612556709013652595821286620854680795341357381795063209776781028174923082035114927807704133636794507489772101449596235088689045734177096918843755837966530867379;
            6'd23: xpb[9] = 1024'd50517460232164144147216595769518971115214492631722096256354568876784996928292728203639428086232322961684850369507198018472138914988147875589535557787686792541095360844443119829135704798599834922249757970426400228670181056128162381040563088477145846766517236482439085671313149964577978726333553446981811799579;
            6'd24: xpb[9] = 1024'd4166034104992034214956867470657626611428781696943876217361867715567298619271444639009157962506812273715133226132839631831293886614981130571844011380761028373177069093064953037416728801858312462704452731076019429165439030221209834273422043317497186043262371515281936253937254194978860533823351055997092731779;
            6'd25: xpb[9] = 1024'd81881303661944665681496066576610714852341497887901340306501021619326495647559299984393959053438975895188565490215974679769512699083034720109312589990166305138949451911258003583327991996633995724469345100112878476025057854535154060471259567841077974586827409962241844866667886499308375358431838491637968148310;
            6'd26: xpb[9] = 1024'd35529877534772555749236338277749370348555786953123120267508320458108797338538016419763688929713465207218848346841616293128667670709867975091621043583240540971031160159879836791609015999892473264924039860762497676520315828628201513704118522681429313863572544995084695449291990729709257165921636100653249080510;
            6'd27: xpb[9] = 1024'd113245147091725187215775537383702458589468503144080584356647474361867994366825871765148490020645628828692280610924751341066886483177921564629089622192645817736803542978072887337520279194668156526688932229799356723379934652942145739901956047205010102407137583442044604062022623034038771990530123536294124497041;
            6'd28: xpb[9] = 1024'd66893720964553077283515809084841114085682792209302364317654773200650296057804588200518219896920118140722563467550392954426041454804754819611398075785720053568885251226694720545801303197926634067143626990448975923875192627035193193134815002045361441683882718474887454644646727264439653798019921145309405429241;
            6'd29: xpb[9] = 1024'd20542294837380967351256080785979769581897081274524144278662072039432597748783304635887949773194607452752846324176034567785196426431588074593706529378794289400966959475316553754082327201185111607598321751098595124370450601128240646367673956885712780960627853507730305227270831494840535605509718754324686361441;
            6'd30: xpb[9] = 1024'd98257564394333598817795279891932857822809797465481608367801225943191794777071159981272750864126771074226278588259169615723415238899641664131175107988199566166739342293509604299993590395960794869363214120135454171230069425442184872565511481409293569504192891954690213840001463799170050430118206189965561777972;
            6'd31: xpb[9] = 1024'd51906138267161488885535551593071513319024086530703388328808524781974096468049876416642480740401260386256561444884811229082570210526474919113483561581273801998821050542131437508274614399219272409817908880785073371725327399535232325798370436249644908780938026987533064422625568029570932237608003798980842710172;
            6'd32: xpb[9] = 1024'd5554712139989378953275823294210168815238375595925168289815823620756398159028592852012210616675749698286844301510452842441725182153308174095792015174348037830902758790753270716555638402477749950272603641434692572220585373628279779031229391089996248057683162020375915005249672259971814045097801407996123642372;
            6'd33: xpb[9] = 1024'd83269981696942010419815022400163257056151091786882632378954977524515595187316448197397011707607913319760276565593587890379943994621361763633260593783753314596675141608946321262466901597253433212037496010471551619080204197942224005229066915613577036601248200467335823617980304564301328869706288843636999058903;
            6'd34: xpb[9] = 1024'd36918555569769900487555294101301912552365380852104412339962276363297896878295164632766741583882402631790559422219229503739098966248195018615569047376827550428756849857568154470747925600511910752492190771121170819575462172035271458461925870453928375877993335500178674200604408794702210677196086452652279991103;
            6'd35: xpb[9] = 1024'd114633825126722531954094493207255000793278097043061876429101430267057093906583019978151542674814566253263991686302364551677317778716248608153037625986232827194529232675761205016659188795287594014257083140158029866435080996349215684659763394977509164421558373947138582813335041099031725501804573888293155407634;
            6'd36: xpb[9] = 1024'd68282398999550422021834764908393656289492386108283656390108729105839395597561736413521272551089055565294274542928006165036472750343081863135346079579307063026610940924383038224940212798546071554711777900807649066930338970442263137892622349817860503698303508979981433395959145329432607309294371497308436339834;
            6'd37: xpb[9] = 1024'd21930972872378312089575036609532311785706675173505436351116027944621697288540452848891002427363544877324557399553647778395627721969915118117654533172381298858692649173004871433221236801804549095166472661457268267425596944535310591125481304658211842975048644012824283978583249559833489116784169106323717272034;
            6'd38: xpb[9] = 1024'd99646242429330943556114235715485400026619391364462900440255181848380894316828308194275803518295708498797989663636782826333846534437968707655123111781786575624465031991197921979132499996580232356931365030494127314285215768849254817323318829181792631518613682459784192591313881864163003941392656541964592688565;
            6'd39: xpb[9] = 1024'd53294816302158833623854507416624055522833680429684680401262480687163196007807024629645533394570197810828272520262424439693001506064801962637431565374860811456546740239819755187413523999838709897386059791143746514780473742942302270556177784022143970795358817492627043173937986094563885748882454150979873620765;
            6'd40: xpb[9] = 1024'd6943390174986723691594779117762711019047969494906460362269779525945497698785741065015263270844687122858555376888066053052156477691635217619740018967935047288628448488441588395694548003097187437840754551793365715275731717035349723789036738862495310072103952525469893756562090324964767556372251759995154552965;
            6'd41: xpb[9] = 1024'd84658659731939355158133978223715799259960685685863924451408933429704694727073596410400064361776850744331987640971201100990375290159688807157208597577340324054400831306634638941605811197872870699605646920830224762135350541349293949986874263386076098615668990972429802369292722629294282380980739195636029969496;
            6'd42: xpb[9] = 1024'd38307233604767245225874249924854454756174974751085704412416232268486996418052312845769794238051340056362270497596842714349530261786522062139517051170414559886482539555256472149886835201131348240060341681479843962630608515442341403219733218226427437892414126005272652951916826859695164188470536804651310901696;
            6'd43: xpb[9] = 1024'd116022503161719876692413449030807542997087690942043168501555386172246193446340168191154595328983503677835702761679977762287749074254575651676985629779819836652254922373449522695798098395907031501825234050516703009490227339756285629417570742750008226435979164452232561564647459164024679013079024240292186318227;
            6'd44: xpb[9] = 1024'd69671077034547766760153720731946198493301980007264948462562685011028495137318884626524325205257992989865985618305619375646904045881408906659294083372894072484336630622071355904079122399165509042279928811166322209985485313849333082650429697590359565712724299485075412147271563394425560820568821849307467250427;
            6'd45: xpb[9] = 1024'd23319650907375656827893992433084853989516269072486728423569983849810796828297601061894055081532482301896268474931260989006059017508242161641602536965968308316418338870693189112360146402423986582734623571815941410480743287942380535883288652430710904989469434517918262729895667624826442628058619458322748182627;
            6'd46: xpb[9] = 1024'd101034920464328288294433191539037942230428985263444192512709137753569993856585456407278856172464645923369700739014396036944277829976295751179071115575373585082190721688886239658271409597199669844499515940852800457340362112256324762081126176954291693533034472964878171342626299929155957452667106893963623599158;
            6'd47: xpb[9] = 1024'd54683494337156178362173463240176597726643274328665972473716436592352295547564172842648586048739135235399983595640037650303432801603129006161379569168447820914272429937508072866552433600458147384954210701502419657835620086349372215313985131794643032809779607997721021925250404159556839260156904502978904531358;
            6'd48: xpb[9] = 1024'd8332068209984068429913734941315253222857563393887752434723735431134597238542889278018315925013624547430266452265679263662587773229962261143688022761522056746354138186129906074833457603716624925408905462152038858330878060442419668546844086634994372086524743030563872507874508389957721067646702111994185463558;
            6'd49: xpb[9] = 1024'd86047337766936699896452934047268341463770279584845216523862889334893794266830744623403117015945788168903698716348814311600806585698015850681156601370927333512126521004322956620744720798492308187173797831188897905190496884756363894744681611158575160630089781477523781120605140694287235892255189547635060880089;
            6'd50: xpb[9] = 1024'd39695911639764589964193205748406996959984568650066996484870188173676095957809461058772846892220277480933981572974455924959961557324849105663465054964001569344208229252944789829025744801750785727628492591838517105685754858849411347977540565998926499906834916510366631703229244924688117699744987156650341812289;
            6'd51: xpb[9] = 1024'd117411181196717221430732404854360085200897284841024460574009342077435292986097316404157647983152441102407413837057590972898180369792902695200933633573406846109980612071137840374937007996526468989393384960875376152545373683163355574175378090522507288450399954957326540315959877229017632524353474592291217228820;
            6'd52: xpb[9] = 1024'd71059755069545111498472676555498740697111573906246240535016640916217594677076032839527377859426930414437696693683232586257335341419735950183242087166481081942062320319759673583218031999784946529848079721524995353040631657256403027408237045362858627727145089990169390898583981459418514331843272201306498161020;
            6'd53: xpb[9] = 1024'd24708328942373001566212948256637396193325862971468020496023939754999896368054749274897107735701419726467979550308874199616490313046569205165550540759555317774144028568381506791499056003043424070302774482174614553535889631349450480641096000203209967003890225023012241481208085689819396139333069810321779093220;
            6'd54: xpb[9] = 1024'd102423598499325633032752147362590484434238579162425484585163093658759093396342604620281908826633583347941411814392009247554709125514622794703019119368960594539916411386574557337410319197819107332067666851211473600395508455663394706838933524726790755547455263469972150093938717994148910963941557245962654509751;
            6'd55: xpb[9] = 1024'd56072172372153523100492419063729139930452868227647264546170392497541395087321321055651638702908072659971694671017650860913864097141456049685327572962034830371998119635196390545691343201077584872522361611861092800890766429756442160071792479567142094824200398502815000676562822224549792771431354854977935441951;
            6'd56: xpb[9] = 1024'd9720746244981413168232690764867795426667157292869044507177691336323696778300037491021368579182561972001977527643292474273019068768289304667636026555109066204079827883818223753972367204336062412977056372510712001386024403849489613304651434407493434100945533535657851259186926454950674578921152463993216374151;
            6'd57: xpb[9] = 1024'd87436015801934044634771889870820883667579873483826508596316845240082893806587892836406169670114725593475409791726427522211237881236342894205104605164514342969852210702011274299883630399111745674741948741547571048245643228163433839502488958931074222644510571982617759871917558759280189403529639899634091790682;
            6'd58: xpb[9] = 1024'd41084589674761934702512161571959539163794162549048288557324144078865195497566609271775899546389214905505692648352069135570392852863176149187413058757588578801933918950633107508164654402370223215196643502197190248740901202256481292735347913771425561921255707015460610454541662989681071211019437508649372722882;
            6'd59: xpb[9] = 1024'd118799859231714566169051360677912627404706878740005752646463297982624392525854464617160700637321378526979124912435204183508611665331229738724881637366993855567706301768826158054075917597145906476961535871234049295600520026570425518933185438295006350464820745462420519067272295294010586035627924944290248139413;
            6'd60: xpb[9] = 1024'd72448433104542456236791632379051282900921167805227532607470596821406694216833181052530430513595867839009407769060845796867766636958062993707190090960068091399788010017447991262356941600404384017416230631883668496095778000663472972166044393135357689741565880495263369649896399524411467843117722553305529071613;
            6'd61: xpb[9] = 1024'd26097006977370346304531904080189938397135456870449312568477895660188995907811897487900160389870357151039690625686487410226921608584896248689498544553142327231869718266069824470637965603662861557870925392533287696591035974756520425398903347975709029018311015528106220232520503754812349650607520162320810003813;
            6'd62: xpb[9] = 1024'd103812276534322977771071103186143026638048173061406776657617049563948192936099752833284961480802520772513122889769622458165140421052949838226967123162547603997642101084262875016549228798438544819635817761570146743450654799070464651596740872499289817561876053975066128845251136059141864475216007597961685420344;
            6'd63: xpb[9] = 1024'd57460850407150867838811374887281682134262462126628556618624348402730494627078469268654691357077010084543405746395264071524295392679783093209275576755621839829723809332884708224830252801697022360090512522219765943945912773163512104829599827339641156838621189007908979427875240289542746282705805206976966352544;
        endcase
    end

    always_comb begin
        case(flag[3][11:6])
            6'd0: xpb[10] = 1024'd0;
            6'd1: xpb[10] = 1024'd11109424279978757906551646588420337630476751191850336579631647241512796318057185704024421233351499396573688603020905684883450364306616348191584030348696075661805517581506541433111276804955499900545207282869385144441170747256559558062458782179992496115366324040751830010499344519943628090195602815992247284744;
            6'd2: xpb[10] = 1024'd22218848559957515813103293176840675260953502383700673159263294483025592636114371408048842466702998793147377206041811369766900728613232696383168060697392151323611035163013082866222553609910999801090414565738770288882341494513119116124917564359984992230732648081503660020998689039887256180391205631984494569488;
            6'd3: xpb[10] = 1024'd33328272839936273719654939765261012891430253575551009738894941724538388954171557112073263700054498189721065809062717054650351092919849044574752091046088226985416552744519624299333830414866499701635621848608155433323512241769678674187376346539977488346098972122255490031498033559830884270586808447976741854232;
            6'd4: xpb[10] = 1024'd44437697119915031626206586353681350521907004767401346318526588966051185272228742816097684933405997586294754412083622739533801457226465392766336121394784302647222070326026165732445107219821999602180829131477540577764682989026238232249835128719969984461465296163007320041997378079774512360782411263968989138976;
            6'd5: xpb[10] = 1024'd55547121399893789532758232942101688152383755959251682898158236207563981590285928520122106166757496982868443015104528424417251821533081740957920151743480378309027587907532707165556384024777499502726036414346925722205853736282797790312293910899962480576831620203759150052496722599718140450978014079961236423720;
            6'd6: xpb[10] = 1024'd66656545679872547439309879530522025782860507151102019477789883449076777908343114224146527400108996379442131618125434109300702185839698089149504182092176453970833105489039248598667660829732999403271243697216310866647024483539357348374752693079954976692197944244510980062996067119661768541173616895953483708464;
            6'd7: xpb[10] = 1024'd77765969959851305345861526118942363413337258342952356057421530690589574226400299928170948633460495776015820221146339794184152550146314437341088212440872529632638623070545790031778937634688499303816450980085696011088195230795916906437211475259947472807564268285262810073495411639605396631369219711945730993208;
            6'd8: xpb[10] = 1024'd88875394239830063252413172707362701043814009534802692637053177932102370544457485632195369866811995172589508824167245479067602914452930785532672242789568605294444140652052331464890214439643999204361658262955081155529365978052476464499670257439939968922930592326014640083994756159549024721564822527937978277952;
            6'd9: xpb[10] = 1024'd99984818519808821158964819295783038674290760726653029216684825173615166862514671336219791100163494569163197427188151163951053278759547133724256273138264680956249658233558872898001491244599499104906865545824466299970536725309036022562129039619932465038296916366766470094494100679492652811760425343930225562696;
            6'd10: xpb[10] = 1024'd111094242799787579065516465884203376304767511918503365796316472415127963180571857040244212333514993965736886030209056848834503643066163481915840303486960756618055175815065414331112768049554999005452072828693851444411707472565595580624587821799924961153663240407518300104993445199436280901956028159922472847440;
            6'd11: xpb[10] = 1024'd122203667079766336972068112472623713935244263110353702375948119656640759498629042744268633566866493362310574633229962533717954007372779830107424333835656832279860693396571955764224044854510498905997280111563236588852878219822155138687046603979917457269029564448270130115492789719379908992151630975914720132184;
            6'd12: xpb[10] = 1024'd9246395675620353479820831656229618821022587176468354827447911833176660479377089538277983585560318449441113828793374784022340530838175843743848239168021867007975536408507279859705082467948793085232289786045381886929688116857817923784526816476680504117575985074904902095885606165394904065228543965281372932597;
            6'd13: xpb[10] = 1024'd20355819955599111386372478244649956451499338368318691407079559074689456797434275242302404818911817846014802431814280468905790895144792191935432269516717942669781053990013821292816359272904292985777497068914767031370858864114377481846985598656673000232942309115656732106384950685338532155424146781273620217341;
            6'd14: xpb[10] = 1024'd31465244235577869292924124833070294081976089560169027986711206316202253115491460946326826052263317242588491034835186153789241259451408540127016299865414018331586571571520362725927636077859792886322704351784152175812029611370937039909444380836665496348308633156408562116884295205282160245619749597265867502085;
            6'd15: xpb[10] = 1024'd42574668515556627199475771421490631712452840752019364566342853557715049433548646650351247285614816639162179637856091838672691623758024888318600330214110093993392089153026904159038912882815292786867911634653537320253200358627496597971903163016657992463674957197160392127383639725225788335815352413258114786829;
            6'd16: xpb[10] = 1024'd53684092795535385106027418009910969342929591943869701145974500799227845751605832354375668518966316035735868240876997523556141988064641236510184360562806169655197606734533445592150189687770792687413118917522922464694371105884056156034361945196650488579041281237912222137882984245169416426010955229250362071573;
            6'd17: xpb[10] = 1024'd64793517075514143012579064598331306973406343135720037725606148040740642069663018058400089752317815432309556843897903208439592352371257584701768390911502245317003124316039987025261466492726292587958326200392307609135541853140615714096820727376642984694407605278664052148382328765113044516206558045242609356317;
            6'd18: xpb[10] = 1024'd75902941355492900919130711186751644603883094327570374305237795282253438387720203762424510985669314828883245446918808893323042716677873932893352421260198320978808641897546528458372743297681792488503533483261692753576712600397175272159279509556635480809773929319415882158881673285056672606402160861234856641061;
            6'd19: xpb[10] = 1024'd87012365635471658825682357775171982234359845519420710884869442523766234705777389466448932219020814225456934049939714578206493080984490281084936451608894396640614159479053069891484020102637292389048740766131077898017883347653734830221738291736627976925140253360167712169381017805000300696597763677227103925805;
            6'd20: xpb[10] = 1024'd98121789915450416732234004363592319864836596711271047464501089765279031023834575170473353452372313622030622652960620263089943445291106629276520481957590472302419677060559611324595296907592792289593948049000463042459054094910294388284197073916620473040506577400919542179880362324943928786793366493219351210549;
            6'd21: xpb[10] = 1024'd109231214195429174638785650952012657495313347903121384044132737006791827341891760874497774685723813018604311255981525947973393809597722977468104512306286547964225194642066152757706573712548292190139155331869848186900224842166853946346655856096612969155872901441671372190379706844887556876988969309211598495293;
            6'd22: xpb[10] = 1024'd120340638475407932545337297540432995125790099094971720623764384248304623659948946578522195919075312415177999859002431632856844173904339325659688542654982623626030712223572694190817850517503792090684362614739233331341395589423413504409114638276605465271239225482423202200879051364831184967184572125203845780037;
            6'd23: xpb[10] = 1024'd7383367071261949053090016724038900011568423161086373075264176424840524640696993372531545937769137502308539054565843883161230697369735339296112447987347658354145555235508018286298888130942086269919372289221378629418205486459076289506594850773368512119785646109057974181271867810846180040261485114570498580450;
            6'd24: xpb[10] = 1024'd18492791351240706959641663312459237642045174352936709654895823666353320958754179076555967171120636898882227657586749568044681061676351687487696478336043734015951072817014559719410164935897586170464579572090763773859376233715635847569053632953361008235151970149809804191771212330789808130457087930562745865194;
            6'd25: xpb[10] = 1024'd29602215631219464866193309900879575272521925544787046234527470907866117276811364780580388404472136295455916260607655252928131425982968035679280508684739809677756590398521101152521441740853086071009786854960148918300546980972195405631512415133353504350518294190561634202270556850733436220652690746554993149938;
            6'd26: xpb[10] = 1024'd40711639911198222772744956489299912902998676736637382814159118149378913594868550484604809637823635692029604863628560937811581790289584383870864539033435885339562107980027642585632718545808585971554994137829534062741717728228754963693971197313346000465884618231313464212769901370677064310848293562547240434682;
            6'd27: xpb[10] = 1024'd51821064191176980679296603077720250533475427928487719393790765390891709912925736188629230871175135088603293466649466622695032154596200732062448569382131961001367625561534184018743995350764085872100201420698919207182888475485314521756429979493338496581250942272065294223269245890620692401043896378539487719426;
            6'd28: xpb[10] = 1024'd62930488471155738585848249666140588163952179120338055973422412632404506230982921892653652104526634485176982069670372307578482518902817080254032599730828036663173143143040725451855272155719585772645408703568304351624059222741874079818888761673330992696617266312817124233768590410564320491239499194531735004170;
            6'd29: xpb[10] = 1024'd74039912751134496492399896254560925794428930312188392553054059873917302549040107596678073337878133881750670672691277992461932883209433428445616630079524112324978660724547266884966548960675085673190615986437689496065229969998433637881347543853323488811983590353568954244267934930507948581435102010523982288914;
            6'd30: xpb[10] = 1024'd85149337031113254398951542842981263424905681504038729132685707115430098867097293300702494571229633278324359275712183677345383247516049776637200660428220187986784178306053808318077825765630585573735823269307074640506400717254993195943806326033315984927349914394320784254767279450451576671630704826516229573658;
            6'd31: xpb[10] = 1024'd96258761311092012305503189431401601055382432695889065712317354356942895185154479004726915804581132674898047878733089362228833611822666124828784690776916263648589695887560349751189102570586085474281030552176459784947571464511552754006265108213308481042716238435072614265266623970395204761826307642508476858402;
            6'd32: xpb[10] = 1024'd107368185591070770212054836019821938685859183887739402291949001598455691503211664708751337037932632071471736481753995047112283976129282473020368721125612339310395213469066891184300379375541585374826237835045844929388742211768112312068723890393300977158082562475824444275765968490338832852021910458500724143146;
            6'd33: xpb[10] = 1024'd118477609871049528118606482608242276316335935079589738871580648839968487821268850412775758271284131468045425084774900731995734340435898821211952751474308414972200731050573432617411656180497085275371445117915230073829912959024671870131182672573293473273448886516576274286265313010282460942217513274492971427890;
            6'd34: xpb[10] = 1024'd5520338466903544626359201791848181202114259145704391323080441016504388802016897206785108289977956555175964280338312982300120863901294834848376656806673449700315574062508756712892693793935379454606454792397375371906722856060334655228662885070056520121995307143211046266658129456297456015294426263859624228303;
            6'd35: xpb[10] = 1024'd16629762746882302532910848380268518832591010337554727902712088258017185120074082910809529523329455951749652883359218667183571228207911183039960687155369525362121091644015298146003970598890879355151662075266760516347893603316894213291121667250049016237361631183962876277157473976241084105490029079851871513047;
            6'd36: xpb[10] = 1024'd27739187026861060439462494968688856463067761529405064482343735499529981438131268614833950756680955348323341486380124352067021592514527531231544717504065601023926609225521839579115247403846379255696869358136145660789064350573453771353580449430041512352727955224714706287656818496184712195685631895844118797791;
            6'd37: xpb[10] = 1024'd38848611306839818346014141557109194093544512721255401061975382741042777756188454318858371990032454744897030089401030036950471956821143879423128747852761676685732126807028381012226524208801879156242076641005530805230235097830013329416039231610034008468094279265466536298156163016128340285881234711836366082535;
            6'd38: xpb[10] = 1024'd49958035586818576252565788145529531724021263913105737641607029982555574074245640022882793223383954141470718692421935721833922321127760227614712778201457752347537644388534922445337801013757379056787283923874915949671405845086572887478498013790026504583460603306218366308655507536071968376076837527828613367279;
            6'd39: xpb[10] = 1024'd61067459866797334159117434733949869354498015104956074221238677224068370392302825726907214456735453538044407295442841406717372685434376575806296808550153828009343161970041463878449077818712878957332491206744301094112576592343132445540956795970019000698826927346970196319154852056015596466272440343820860652023;
            6'd40: xpb[10] = 1024'd72176884146776092065669081322370206984974766296806410800870324465581166710360011430931635690086952934618095898463747091600823049740992923997880838898849903671148679551548005311560354623668378857877698489613686238553747339599692003603415578150011496814193251387722026329654196575959224556468043159813107936767;
            6'd41: xpb[10] = 1024'd83286308426754849972220727910790544615451517488656747380501971707093963028417197134956056923438452331191784501484652776484273414047609272189464869247545979332954197133054546744671631428623878758422905772483071382994918086856251561665874360330003992929559575428473856340153541095902852646663645975805355221511;
            6'd42: xpb[10] = 1024'd94395732706733607878772374499210882245928268680507083960133618948606759346474382838980478156789951727765473104505558461367723778354225620381048899596242054994759714714561088177782908233579378658968113055352456527436088834112811119728333142509996489044925899469225686350652885615846480736859248791797602506255;
            6'd43: xpb[10] = 1024'd105505156986712365785324021087631219876405019872357420539765266190119555664531568543004899390141451124339161707526464146251174142660841968572632929944938130656565232296067629610894185038534878559513320338221841671877259581369370677790791924689988985160292223509977516361152230135790108827054851607789849790999;
            6'd44: xpb[10] = 1024'd116614581266691123691875667676051557506881771064207757119396913431632351982588754247029320623492950520912850310547369831134624506967458316764216960293634206318370749877574171044005461843490378460058527621091226816318430328625930235853250706869981481275658547550729346371651574655733736917250454423782097075743;
            6'd45: xpb[10] = 1024'd3657309862545140199628386859657462392660095130322409570896705608168252963336801041038670642186775608043389506110782081439011030432854330400640865625999241046485592889509495139486499456928672639293537295573372114395240225661593020950730919366744528124204968177364118352044391101748731990327367413148749876156;
            6'd46: xpb[10] = 1024'd14766734142523898106180033448077800023136846322172746150528352849681049281393986745063091875538275004617078109131687766322461394739470678592224895974695316708291110471016036572597776261884172539838744578442757258836410972918152579013189701546737024239571292218115948362543735621692360080522970229140997160900;
            6'd47: xpb[10] = 1024'd25876158422502656012731680036498137653613597514023082730160000091193845599451172449087513108889774401190766712152593451205911759046087026783808926323391392370096628052522578005709053066839672440383951861312142403277581720174712137075648483726729520354937616258867778373043080141635988170718573045133244445644;
            6'd48: xpb[10] = 1024'd36985582702481413919283326624918475284090348705873419309791647332706641917508358153111934342241273797764455315173499136089362123352703374975392956672087468031902145634029119438820329871795172340929159144181527547718752467431271695138107265906722016470303940299619608383542424661579616260914175861125491730388;
            6'd49: xpb[10] = 1024'd48095006982460171825834973213338812914567099897723755889423294574219438235565543857136355575592773194338143918194404820972812487659319723166976987020783543693707663215535660871931606676750672241474366427050912692159923214687831253200566048086714512585670264340371438394041769181523244351109778677117739015132;
            6'd50: xpb[10] = 1024'd59204431262438929732386619801759150545043851089574092469054941815732234553622729561160776808944272590911832521215310505856262851965936071358561017369479619355513180797042202305042883481706172142019573709920297836601093961944390811263024830266707008701036588381123268404541113701466872441305381493109986299876;
            6'd51: xpb[10] = 1024'd70313855542417687638938266390179488175520602281424429048686589057245030871679915265185198042295771987485521124236216190739713216272552419550145047718175695017318698378548743738154160286661672042564780992789682981042264709200950369325483612446699504816402912421875098415040458221410500531500984309102233584620;
            6'd52: xpb[10] = 1024'd81423279822396445545489912978599825805997353473274765628318236298757827189737100969209619275647271384059209727257121875623163580579168767741729078066871770679124215960055285171265437091617171943109988275659068125483435456457509927387942394626692000931769236462626928425539802741354128621696587125094480869364;
            6'd53: xpb[10] = 1024'd92532704102375203452041559567020163436474104665125102207949883540270623507794286673234040508998770780632898330278027560506613944885785115933313108415567846340929733541561826604376713896572671843655195558528453269924606203714069485450401176806684497047135560503378758436039147261297756711892189941086728154108;
            6'd54: xpb[10] = 1024'd103642128382353961358593206155440501066950855856975438787581530781783419825851472377258461742350270177206586933298933245390064309192401464124897138764263922002735251123068368037487990701528171744200402841397838414365776950970629043512859958986676993162501884544130588446538491781241384802087792757078975438852;
            6'd55: xpb[10] = 1024'd114751552662332719265144852743860838697427607048825775367213178023296216143908658081282882975701769573780275536319838930273514673499017812316481169112959997664540768704574909470599267506483671644745610124267223558806947698227188601575318741166669489277868208584882418457037836301185012892283395573071222723596;
            6'd56: xpb[10] = 1024'd1794281258186735772897571927466743583205931114940427818712970199832117124656704875292232994395594660910814731883251180577901196964413825952905074445325032392655611716510233566080305119921965823980619798749368856883757595262851386672798953663432536126414629211517190437430652747200007965360308562437875524009;
            6'd57: xpb[10] = 1024'd12903705538165493679449218515887081213682682306790764398344617441344913442713890579316654227747094057484503334904156865461351561271030174144489104794021108054461129298016774999191581924877465724525827081618754001324928342519410944735257735843425032241780953252269020447929997267143636055555911378430122808753;
            6'd58: xpb[10] = 1024'd24013129818144251586000865104307418844159433498641100977976264682857709760771076283341075461098593454058191937925062550344801925577646522336073135142717183716266646879523316432302858729832965625071034364488139145766099089775970502797716518023417528357147277293020850458429341787087264145751514194422370093497;
            6'd59: xpb[10] = 1024'd35122554098123009492552511692727756474636184690491437557607911924370506078828261987365496694450092850631880540945968235228252289884262870527657165491413259378072164461029857865414135534788465525616241647357524290207269837032530060860175300203410024472513601333772680468928686307030892235947117010414617378241;
            6'd60: xpb[10] = 1024'd46231978378101767399104158281148094105112935882341774137239559165883302396885447691389917927801592247205569143966873920111702654190879218719241195840109335039877682042536399298525412339743965426161448930226909434648440584289089618922634082383402520587879925374524510479428030826974520326142719826406864662985;
            6'd61: xpb[10] = 1024'd57341402658080525305655804869568431735589687074192110716871206407396098714942633395414339161153091643779257746987779604995153018497495566910825226188805410701683199624042940731636689144699465326706656213096294579089611331545649176985092864563395016703246249415276340489927375346918148416338322642399111947729;
            6'd62: xpb[10] = 1024'd68450826938059283212207451457988769366066438266042447296502853648908895032999819099438760394504591040352946350008685289878603382804111915102409256537501486363488717205549482164747965949654965227251863495965679723530782078802208735047551646743387512818612573456028170500426719866861776506533925458391359232473;
            6'd63: xpb[10] = 1024'd79560251218038041118759098046409106996543189457892783876134500890421691351057004803463181627856090436926634953029590974762053747110728263293993286886197562025294234787056023597859242754610465127797070778835064867971952826058768293110010428923380008933978897496780000510926064386805404596729528274383606517217;
        endcase
    end

    always_comb begin
        case(flag[3][16:12])
            5'd0: xpb[11] = 1024'd0;
            5'd1: xpb[11] = 1024'd90669675498016799025310744634829444627019940649743120455766148131934487669114190507487602861207589833500323556050496659645504111417344611485577317234893637687099752368562565030970519559565965028342278061704450012413123573315327851172469211103372505049345221537531830521425408906749032686925131090375853801961;
            5'd2: xpb[11] = 1024'd57272655311908856651822561864844456509341454173750556783400441198892080000919242104960134507757505357557497704643499884711944381993468888415994509453456234440508830167553912724310799927614724335374358515021660178461886296409758929379959852523515560831870539660946603012744289739569432356731572354126113119591;
            5'd3: xpb[11] = 1024'd23875635125800914278334379094859468391662967697757993111034734265849672332724293702432666154307420881614671853236503109778384652569593165346411701672018831193917907966545260417651080295663483642406438968338870344510649019504190007587450493943658616614395857784361375504063170572389832026538013617876372437221;
            5'd4: xpb[11] = 1024'd114545310623817713303645123729688913018682908347501113566800882397784160001838484209920269015515010715114995409286999769423888763986937776831989018906912468881017660335107825448621599855229448670748717030043320356923772592819517858759919705047031121663741079321893206025488579479138864713463144708252226239182;
            5'd5: xpb[11] = 1024'd81148290437709770930156940959703924901004421871508549894435175464741752333643535807392800662064926239172169557880002994490329034563062053762406211125475065634426738134099173141961880223278207977780797483360530522972535315913948936967410346467174177446266397445307978516807460311959264383269585972002485556812;
            5'd6: xpb[11] = 1024'd47751270251601828556668758189718936783325935395515986222069468531699344665448587404865332308614841763229343706473006219556769305139186330692823403344037662387835815933090520835302160591326967284812877936677740689021298039008380015174900987887317233228791715568722751008126341144779664053076027235752744874442;
            5'd7: xpb[11] = 1024'd14354250065493886183180575419733948665647448919523422549703761598656936997253639002337863955164757287286517855066009444623209575715310607623240595562600259141244893732081868528642440959375726591844958389994950855070060762102811093382391629307460289011317033692137523499445221977600063722882468499503004192072;
            5'd8: xpb[11] = 1024'd105023925563510685208491320054563393292667389569266543005469909730591424666367829509825466816372347120786841411116506104268713687132655219108817912797493896828344646100644433559612960518941691620187236451699400867483184335418138944554860840410832794060662255229669354020870630884349096409807599589878857994033;
            5'd9: xpb[11] = 1024'd71626905377402742835003137284578405174988903093273979333104202797549016998172881107297998462922262644844015559709509329335153957708779496039235105016056493581753723899635781252953240886990450927219316905016611033531947058512570022762351481830975849843187573353084126512189511717169496079614040853629117311663;
            5'd10: xpb[11] = 1024'd38229885191294800461514954514593417057310416617281415660738495864506609329977932704770530109472178168901189708302512554401594228284903772969652297234619090335162801698627128946293521255039210234251397358333821199580709781607001100969842123251118905625712891476498899003508392549989895749420482117379376629293;
            5'd11: xpb[11] = 1024'd4832865005186858088026771744608428939631930141288851988372788931464201661782984302243061756022093692958363856895515779468034498861028049900069489453181687088571879497618476639633801623087969541283477811651031365629472504701432179177332764671261961408238209599913671494827273382810295419226923381129635946923;
            5'd12: xpb[11] = 1024'd95502540503203657113337516379437873566651870791031972444138937063398689330897174809730664617229683526458687412946012439113538610278372661385646806688075324775671631866181041670604321182653934569625755873355481378042596078016760030349801975774634466457583431137445502016252682289559328106152054471505489748884;
            5'd13: xpb[11] = 1024'd62105520317095714739849333609452885448973384315039408771773230130356281662702226407203196263779599050515861561539015664179978880854496938316063998906637921529080709665172389363944601550702693876657836326672691544091358801111191108557292617194777522240108749260860274507571563122379727775958495735255749066514;
            5'd14: xpb[11] = 1024'd28708500130987772366361150839467897331294897839046845099407523197313873994507278004675727910329514574573035710132018889246419151430621215246481191125200518282489787464163737057284881918751453183689916779989901710140121524205622186764783258614920578022634067384275046998890443955200127445764936999006008384144;
            5'd15: xpb[11] = 1024'd119378175629004571391671895474297341958314838488789965555173671329248361663621468512163330771537104408073359266182515548891923262847965826732058508360094155969589539832726302088255401478317418212032194841694351722553245097520950037937252469718293083071979288921806877520315852861949160132690068089381862186105;
            5'd16: xpb[11] = 1024'd85981155442896629018183712704312353840636352012797401882807964396205953995426520109635862418087019932130533414775518773958363533424090103662475700578656752722998617631717649781595681846366177519064275295011561888602007820615381116144743111138436138854504607045221650011634733694769559802496509353132121503735;
            5'd17: xpb[11] = 1024'd52584135256788686644695529934327365722957865536804838210442257463163546327231571707108394064636935456187707563368521999024803804000214380592892892797219349476407695430708997474935962214414936826096355748328772054650770543709812194352233752558579194637029925168636422502953614527589959472302950616882380821365;
            5'd18: xpb[11] = 1024'd19187115070680744271207347164342377605279379060812274538076550530121138659036623304580925711186850980244881711961525224091244074576338657523310085015781946229816773229700345168276242582463696133128436201645982220699533266804243272559724393978722250419555243292051194994272495360410359142109391880632640138995;
            5'd19: xpb[11] = 1024'd109856790568697543296518091799171822232299319710555394993842698662055626328150813812068528572394440813745205268012021883736748185993683269008887402250675583916916525598262910199246762142029661161470714263350432233112656840119571123732193605082094755468900464829583025515697904267159391829034522971008493940956;
            5'd20: xpb[11] = 1024'd76459770382589600923029909029186834114620833234562831321476991729013218659955865409541060218944356337802379416605025108803188456569807545939304594469238180670325603397254257892587042510078420468502794716667642399161419563214002201939684246502237811251425782952997798007016785099979791498840964234758753258586;
            5'd21: xpb[11] = 1024'd43062750196481658549541726259201845996942346758570267649111284795970810991760917007013591865494271861859553565198028333869628727145931822869721786687800777423734681196245605585927322878127179775534875169984852565210182286308433280147174887922380867033951101076412570498335665932800191168647405498509012576216;
            5'd22: xpb[11] = 1024'd9665730010373716176053543489216857879263860282577703976745577862928403323565968604486123512044187385916727713791031558936068997722056099800138978906363374177143758995236953279267603246175939082566955623302062731258945009402864358354665529342523922816476419199827342989654546765620590838453846762259271893846;
            5'd23: xpb[11] = 1024'd100335405508390515201364288124046302506283800932320824432511725994862890992680159111973726373251777219417051269841528218581573109139400711285716296141257011864243511363799518310238122805741904110909233685006512743672068582718192209527134740445896427865821640737359173511079955672369623525378977852635125695807;
            5'd24: xpb[11] = 1024'd66938385322282572827876105354061314388605314456328260760146019061820483324485210709446258019801692743474225418434531443648013379715524988216133488359819608617652589162790866003578403173790663417941314138323722909720831305812623287734625381866039483648346958860773946002398836505190023195185419116385385013437;
            5'd25: xpb[11] = 1024'd33541365136174630454387922584076326270926827980335697087780312128778075656290262306918789666351608267531399567027534668714453650291649265146550680578382205371061666961782213696918683541839422724973394591640933075769594028907054365942116023286182539430872276984188718493717717338010422864991860380135644331067;
            5'd26: xpb[11] = 1024'd144344950066688080899739814091338153248341504343133415414605195735667988095313904391321312901523791588573715620537893780893920867773542076967872796944802124470744760773561390258963909888182032005475044958143241818356752001485444149606664706325595213397595107603490985036598170830822534798301643885903648697;
            5'd27: xpb[11] = 1024'd90814020448083487106210484448920782780268282154086253871180753327670155657209504411878924174109113625088897271671034553426398032285118153562545190031838439811570497129336126421229483469454147060347753106662593254231480325316813295322075875809698100262742816645135321506462007077579855221723432734261757450658;
            5'd28: xpb[11] = 1024'd57417000261975544732722301678935794662589795678093690198815046394627747989014556009351455820659029149146071420264037778492838302861242430492962382250401036564979574928327474114569763837502906367379833559979803420280243048411244373529566517229841156045268134768550093997780887910400254891529873998012016768288;
            5'd29: xpb[11] = 1024'd24019980075867602359234118908950806544911309202101126526449339461585340320819607606823987467208944673203245568857041003559278573437366707423379574468963633318388652727318821807910044205551665674411914013297013586329005771505675451737057158649984211827793452891964866489099768743220654561336315261762276085918;
            5'd30: xpb[11] = 1024'd114689655573884401384544863543780251171931249851844246982215487593519827989933798114311590328416534506703569124907537663204782684854711318908956891703857271005488405095881386838880563765117630702754192075001463598742129344821003302909526369753356716877138674429496697010525177649969687248261446352138129887879;
            5'd31: xpb[11] = 1024'd81292635387776459011056680773795263054252763375851683309849780660477420321738849711784121974966450030760743273500540888271222955430835595839374083922419867758897482894872734532220844133166390009786272528318673764790892067915434381117017011173499772659663992552911469501844058482790086918067887615888389205509;
        endcase
    end

    always_comb begin
        case(flag[4][5:0])
            6'd0: xpb[12] = 1024'd0;
            6'd1: xpb[12] = 1024'd85981155442896629018183712704312353840636352012797401882807964396205953995426520109635862418087019932130533414775518773958363533424090103662475700578656752722998617631717649781595681846366177519064275295011561888602007820615381116144743111138436138854504607045221650011634733694769559802496509353132121503735;
            6'd2: xpb[12] = 1024'd47895615201668516637568498003810274936574276899859119637484073727435012653543901309256653621516365554817917422093544113337663226006959872769791276140982464512306560693864082225561124501215149316818352981635883930839654791009865459324507652593642828442189310676326241993162939315610486587874328879638648523139;
            6'd3: xpb[12] = 1024'd9810074960440404256953283303308196032512201786920837392160183058664071311661282508877444824945711177505301429411569452716962918589829641877106851703308176301614503756010514669526567156064121114572430668260205973077301761404349802504272194048849518029874014307430833974691144936451413373252148406145175542543;
            6'd4: xpb[12] = 1024'd95791230403337033275136996007620549873148553799718239274968147454870025307087802618513307243032731109635834844187088226675326452013919745539582552281964929024613121387728164451122249002430298633636705963271767861679309582019730918649015305187285656884378621352652483986325878631220973175748657759277297046278;
            6'd5: xpb[12] = 1024'd57705690162108920894521781307118470969086478686779957029644256786099083965205183818134098446462076732323218851505113566054626144596789514646898127844290640813921064449874596895087691657279270431390783649896089903916956552414215261828779846642492346472063324983757075967854084252061899961126477285783824065682;
            6'd6: xpb[12] = 1024'd19620149920880808513906566606616392065024403573841674784320366117328142623322565017754889649891422355010602858823138905433925837179659283754213703406616352603229007512021029339053134312128242229144861336520411946154603522808699605008544388097699036059748028614861667949382289872902826746504296812290351085086;
            6'd7: xpb[12] = 1024'd105601305363777437532090279310928745905660755586639076667128330513534096618749085127390752067978442287141136273598657679392289370603749387416689403985273105326227625143738679120648816158494419748209136631531973834756611343424080721153287499236135174914252635660083317961017023567672386549000806165422472588821;
            6'd8: xpb[12] = 1024'd67515765122549325151475064610426667001598680473700794421804439844763155276866466327011543271407787909828520280916683018771589063186619156524004979547598817115535568205885111564614258813343391545963214318156295876994258313818565064333052040691341864501937339291187909942545229188513313334378625691928999608225;
            6'd9: xpb[12] = 1024'd29430224881321212770859849909924588097536605360762512176480549175992213934983847526632334474837133532515904288234708358150888755769488925631320555109924528904843511268031544008579701468192363343717292004780617919231905284213049407512816582146548554089622042922292501924073434809354240119756445218435526627629;
            6'd10: xpb[12] = 1024'd115411380324217841789043562614236941938172957373559914059288513572198167930410367636268196892924153464646437703010227132109252289193579029293796255688581281627842128899749193790175383314558540862781567299792179807833913104828430523657559693284984692944126649967514151935708168504123799922252954571567648131364;
            6'd11: xpb[12] = 1024'd77325840082989729408428347913734863034110882260621631813964622903427226588527748835888988096353499087333821710328252471488551981776448798401111831250906993417150071961895626234140825969407512660535644986416501850071560075222914866837324234740191382531811353598618743917236374124964726707630774098074175150768;
            6'd12: xpb[12] = 1024'd39240299841761617027813133213232784130048807147683349568640732234656285246645130035509779299782844710021205717646277810867851674359318567508427406813232705206458015024042058678106268624256484458289722673040823892309207045617399210017088776195398072119496057229723335898764579745805653493008593624580702170172;
            6'd13: xpb[12] = 1024'd1154759600533504647197918512730705225986732034745067323316841565885343904762511235130570503212190332708589724964303150247151366942188336615742982375558416995765958086188491122071711279105456256043800359665145934546854016011883553196853317650604761707180760860827927880292785366646580278386413151087229189576;
            6'd14: xpb[12] = 1024'd87135915043430133665381631217043059066623084047542469206124805962091297900189031344766432921299210264839123139739821924205514900366278440278218682954215169718764575717906140903667393125471633775108075654676707823148861836627264669341596428789040900561685367906049577891927519061416140080882922504219350693311;
            6'd15: xpb[12] = 1024'd49050374802202021284766416516540980162561008934604186960800915293320356558306412544387224124728555887526507147057847263584814592949148209385534258516540881508072518780052573347632835780320605572862153341301029865386508807021749012521360970244247590149370071537154169873455724682257066866260742030725877712715;
            6'd16: xpb[12] = 1024'd10964834560973908904151201816038901258498933821665904715477024624549415216423793744008015328157901510213891154375872602964114285532017978492849834078866593297380461842199005791598278435169577370616231027925351907624155777416233355701125511699454279737054775168258761854983930303097993651638561557232404732119;
            6'd17: xpb[12] = 1024'd96945990003870537922334914520351255099135285834463306598284989020755369211850313853643877746244921442344424569151391376922477818956108082155325534657523346020379079473916655573193960281535754889680506322936913796226163598031614471845868622837890418591559382213480411866618663997867553454135070910364526235854;
            6'd18: xpb[12] = 1024'd58860449762642425541719699819849176195073210721525024352961098351984427869967695053264668949674267065031808576469416716301777511538977851262641110219849057809687022536063088017159402936384726687434584009561235838463810568426098815025633164293097108179244085844585003848146869618708480239512890436871053255258;
            6'd19: xpb[12] = 1024'd20774909521414313161104485119347097291011135608586742107637207683213486528085076252885460153103612687719192583787442055681077204121847620369956685782174769598994965598209520461124845591233698485188661696185557880701457538820583158205397705748303797766928789475689595829675075239549407024890709963377580274662;
            6'd20: xpb[12] = 1024'd106756064964310942179288197823659451131647487621384143990445172079419440523511596362521322571190632619849725998562960829639440737545937724032432386360831522321993583229927170242720527437599876004252936991197119769303465359435964274350140816886739936621433396520911245841309808934318966827387219316509701778397;
            6'd21: xpb[12] = 1024'd68670524723082829798672983123157372227585412508445861745121281410648499181628977562142113774619978242537110005880986169018740430128807493139747961923157234111301526292073602686685970092448847802007014677821441811541112329830448617529905358341946626209118100152015837822838014555159893612765038843016228797801;
            6'd22: xpb[12] = 1024'd30584984481854717418057768422655293323523337395507579499797390741877557839746358761762904978049323865224494013199011508398040122711677262247063537485482945900609469354220035130651412747297819599761092364445763853778759300224932960709669899797153315796802803783120429804366220176000820398142858369522755817205;
            6'd23: xpb[12] = 1024'd116566139924751346436241481126967647164159689408304981382605355138083511835172878871398767396136343797355027427974530282356403656135767365909539238064139698623608086985937684912247094593663997118825367659457325742380767120840314076854413010935589454651307410828342079816000953870770380200639367722654877320940;
            6'd24: xpb[12] = 1024'd78480599683523234055626266426465568260097614295366699137281464469312570493290260071019558599565689420042411435292555621735703348718637135016854813626465410412916030048084117356212537248512968916579445346081647784618414091234798420034177552390796144238992114459446671797529159491611306986017187249161404340344;
            6'd25: xpb[12] = 1024'd40395059442295121675011051725963489356035539182428416891957573800541629151407641270640349802995035042729795442610580961115003041301506904124170389188791122202223973110230549800177979903361940714333523032705969826856061061629282763213942093846002833826676818090551263779057365112452233771395006775667931359748;
            6'd26: xpb[12] = 1024'd2309519201067009294395837025461410451973464069490134646633683131770687809525022470261141006424380665417179449928606300494302733884376673231485964751116833991531916172376982244143422558210912512087600719330291869093708032023767106393706635301209523414361521721655855760585570733293160556772826302174458379152;
            6'd27: xpb[12] = 1024'd88290674643963638312579549729773764292609816082287536529441647527976641804951542579897003424511400597547712864704125074452666267308466776893961665329773586714530533804094632025739104404577090031151876014341853757695715852639148222538449746439645662268866128766877505772220304428062720359269335655306579882887;
            6'd28: xpb[12] = 1024'd50205134402735525931964335029271685388547740969349254284117756859205700463068923779517794627940746220235096872022150413831965959891336546001277240892099298503838476866241064469704547059426061828905953700966175799933362823033632565718214287894852351856550832397982097753748510048903647144647155181813106902291;
            6'd29: xpb[12] = 1024'd12119594161507413551349120328769606484485665856410972038793866190434759121186304979138585831370091842922480879340175753211265652474206315108592816454425010293146419928387496913669989714275033626660031387590497842171009793428116908897978829350059041444235536029086689735276715669744573930024974708319633921695;
            6'd30: xpb[12] = 1024'd98100749604404042569532833033081960325122017869208373921601830586640713116612825088774448249457111775053014294115694527169629185898296418771068517033081763016145037560105146695265671560641211145724306682602059730773017614043498025042721940488495180298740143074308339746911449364514133732521484061451755425430;
            6'd31: xpb[12] = 1024'd60015209363175930188917618332579881421059942756270091676277939917869771774730206288395239452886457397740398301433719866548928878481166187878384092595407474805452980622251579139231114215490182943478384369226381773010664584437982368222486481943701869886424846705412931728439654985355060517899303587958282444834;
            6'd32: xpb[12] = 1024'd21929669121947817808302403632077802516997867643331809430954049249098830432847587488016030656315803020427782308751745205928228571064035956985699668157733186594760923684398011583196556870339154741232462055850703815248311554832466711402251023398908559474109550336517523709967860606195987303277123114464809464238;
            6'd33: xpb[12] = 1024'd107910824564844446826486116336390156357634219656129211313762013645304784428274107597651893074402822952558315723527263979886592104488126060648175368736389939317759541316115661364792238716705332260296737350862265703850319375447847827546994134537344698328614157381739173721602594300965547105773632467596930967973;
            6'd34: xpb[12] = 1024'd69825284323616334445870901635888077453572144543190929068438122976533843086391488797272684277832168575245699730845289319265891797070995829755490944298715651107067484378262093808757681371554304058050815037486587746087966345842332170726758675992551387916298861012843765703130799921806473891151451994103457987377;
            6'd35: xpb[12] = 1024'd31739744082388222065255686935385998549510069430252646823114232307762901744508869996893475481261514197933083738163314658645191489653865598862806519861041362896375427440408526252723124026403275855804892724110909788325613316236816513906523217447758077503983564643948357684659005542647400676529271520609985006781;
            6'd36: xpb[12] = 1024'd117720899525284851083439399639698352390146421443050048705922196703968855739935390106529337899348534130063617152938833432603555023077955702525282220439698115619374045072126176034318805872769453374869168019122471676927621136852197630051266328586194216358488171689170007696293739237416960479025780873742106510516;
            6'd37: xpb[12] = 1024'd79635359284056738702824184939196273486084346330111766460598306035197914398052771306150129102777879752751001160256858771982854715660825471632597796002023827408681988134272608478284248527618425172623245705746793719165268107246681973231030870041400905946172875320274599677821944858257887264403600400248633529920;
            6'd38: xpb[12] = 1024'd41549819042828626322208970238694194582022271217173484215274415366426973056170152505770920306207225375438385167574884111362154408243695240739913371564349539197989931196419040922249691182467396970377323392371115761402915077641166316410795411496607595533857578951379191659350150479098814049781419926755160549324;
            6'd39: xpb[12] = 1024'd3464278801600513941593755538192115677960196104235201969950524697656031714287533705391711509636570998125769174892909450741454100826565009847228947126675250987297874258565473366215133837316368768131401078995437803640562048035650659590559952951814285121542282582483783640878356099939740835159239453261687568728;
            6'd40: xpb[12] = 1024'd89445434244497142959777468242504469518596548117032603852758489093861985709714053815027573927723590930256302589668428224699817634250655113509704647705332003710296491890283123147810815683682546287195676374006999692242569868651031775735303064090250423976046889627705433652513089794709300637655748806393809072463;
            6'd41: xpb[12] = 1024'd51359894003269030579162253542002390614534473004094321607434598425091044367831435014648365131152936552943686596986453564079117326833524882617020223267657715499604434952429555591776258338531518084949754060631321734480216839045516118915067605545457113563731593258810025634041295415550227423033568332900336091867;
            6'd42: xpb[12] = 1024'd13274353762040918198547038841500311710472397891156039362110707756320103025948816214269156334582282175631070604304478903458417019416394651724335798829983427288912378014575988035741700993380489882703831747255643776717863809440000462094832147000663803151416296889914617615569501036391154208411387859406863111271;
            6'd43: xpb[12] = 1024'd99255509204937547216730751545812665551108749903953441244918672152526057021375336323905018752669302107761604019079997677416780552840484755386811499408640180011910995646293637817337382839746667401768107042267205665319871630055381578239575258139099942005920903935136267627204234731160714010907897212538984615006;
            6'd44: xpb[12] = 1024'd61169968963709434836115536845310586647046674791015158999594781483755115679492717523525809956098647730448988026398023016796080245423354524494127074970965891801218938708440070261302825494595639199522184728891527707557518600449865921419339799594306631593605607566240859608732440352001640796285716739045511634410;
            6'd45: xpb[12] = 1024'd23084428722481322455500322144808507742984599678076876754270890814984174337610098723146601159527993353136372033716048356175379938006224293601442650533291603590526881770586502705268268149444610997276262415515849749795165570844350264599104341049513321181290311197345451590260645972842567581663536265552038653814;
            6'd46: xpb[12] = 1024'd109065584165377951473684034849120861583620951690874278637078855211190128333036618832782463577615013285266905448491567130133743471430314397263918351111948356313525499402304152486863949995810788516340537710527411638397173391459731380743847452187949460035794918242567101601895379667612127384160045618684160157549;
            6'd47: xpb[12] = 1024'd70980043924149839093068820148618782679558876577935996391754964542419186991154000032403254781044358907954289455809592469513043164013184166371233926674274068102833442464450584930829392650659760314094615397151733680634820361854215723923611993643156149623479621873671693583423585288453054169537865145190687176953;
            6'd48: xpb[12] = 1024'd32894503682921726712453605448116703775496801464997714146431073873648245649271381232024045984473704530641673463127617808892342856596053935478549502236599779892141385526597017374794835305508732111848693083776055722872467332248700067103376535098362839211164325504776285564951790909293980954915684671697214196357;
            6'd49: xpb[12] = 1024'd118875659125818355730637318152429057616133153477795116029239038269854199644697901341659908402560724462772206877903136582850706390020144039141025202815256532615140003158314667156390517151874909630912968378787617611474475152864081183248119646236798978065668932549997935576586524604063540757412194024829335700092;
            6'd50: xpb[12] = 1024'd80790118884590243350022103451926978712071078364856833783915147601083258302815282541280699605990070085459590885221161922230006082603013808248340778377582244404447946220461099600355959806723881428667046065411939653712122123258565526427884187692005667653353636181102527558114730224904467542790013551335862719496;
            6'd51: xpb[12] = 1024'd42704578643362130969406888751424899808009003251918551538591256932312316960932663740901490809419415708146974892539187261609305775185883577355656353939907956193755889282607532044321402461572853226421123752036261695949769093653049869607648729147212357241038339812207119539642935845745394328167833077842389738900;
            6'd52: xpb[12] = 1024'd4619038402134018588791674050922820903946928138980269293267366263541375619050044940522282012848761330834358899857212600988605467768753346462971929502233667983063832344753964488286845116421825024175201438660583738187416064047534212787413270602419046828723043443311711521171141466586321113545652604348916758304;
            6'd53: xpb[12] = 1024'd90600193845030647606975386755235174744583280151777671176075330659747329614476565050158144430935781262964892314632731374946969001192843450125447630080890420706062449976471614269882526962788002543239476733672145626789423884662915328932156381740855185683227650488533361532805875161355880916042161957481038262039;
            6'd54: xpb[12] = 1024'd52514653603802535226360172054733095840521205038839388930751439990976388272593946249778935634365126885652276321950756714326268693775713219232763205643216132495370393038618046713847969617636974340993554420296467669027070855057399672111920923196061875270912354119637953514334080782196807701419981483987565281443;
            6'd55: xpb[12] = 1024'd14429113362574422845744957354231016936459129925901106685427549322205446930711327449399726837794472508339660329268782053705568386358582988340078781205541844284678336100764479157813412272485946138747632106920789711264717825451884015291685464651268564858597057750742545495862286403037734486797801010494092300847;
            6'd56: xpb[12] = 1024'd100410268805471051863928670058543370777095481938698508568235513718411400926137847559035589255881492440470193744044300827663931919782673092002554481784198597007676953732482128939409094118852123657811907401932351599866725646067265131436428575789704703713101664795964195507497020097807294289294310363626213804582;
            6'd57: xpb[12] = 1024'd62324728564242939483313455358041291873033406825760226322911623049640459584255228758656380459310838063157577751362326167043231612365542861109870057346524308796984896794628561383374536773701095455565985088556673642104372616461749474616193117244911393300786368427068787489025225718648221074672129890132740823986;
            6'd58: xpb[12] = 1024'd24239188323014827102698240657539212968971331712821944077587732380869518242372609958277171662740183685844961758680351506422531304948412630217185632908850020586292839856774993827339979428550067253320062775180995684342019586856233817795957658700118082888471072058173379470553431339489147860049949416639267843390;
            6'd59: xpb[12] = 1024'd110220343765911456120881953361851566809607683725619345960395696777075472237799130067913034080827203617975495173455870280380894838372502733879661333487506773309291457488492643608935661274916244772384338070192557572944027407471614933940700769838554221742975679103395029482188165034258707662546458769771389347125;
            6'd60: xpb[12] = 1024'd72134803524683343740266738661349487905545608612681063715071806108304530895916511267533825284256549240662879180773895619760194530955372502986976909049832485098599400550639076052901103929765216570138415756816879615181674377866099277120465311293760911330660382734499621463716370655099634447924278296277916366529;
            6'd61: xpb[12] = 1024'd34049263283455231359651523960847409001483533499742781469747915439533589554033892467154616487685894863350263188091920959139494223538242272094292484612158196887907343612785508496866546584614188367892493443441201657419321348260583620300229852748967600918345086365604213445244576275940561233302097822784443385933;
            6'd62: xpb[12] = 1024'd120030418726351860377835236665159762842119885512540183352555879835739543549460412576790478905772914795480796602867439733097857756962332375756768185190814949610905961244503158278462228430980365886956768738452763546021329168875964736444972963887403739772849693410825863456879309970710121035798607175916564889668;
            6'd63: xpb[12] = 1024'd81944878485123747997220021964657683938057810399601901107231989166968602207577793776411270109202260418168180610185465072477157449545202144864083760753140661400213904306649590722427671085829337684710846425077085588258976139270449079624737505342610429360534397041930455438407515591551047821176426702423091909072;
        endcase
    end

    always_comb begin
        case(flag[4][11:6])
            6'd0: xpb[13] = 1024'd0;
            6'd1: xpb[13] = 1024'd43859338243895635616604807264155605033995735286663618861908098498197660865695174976032061312631606040855564617503490411856457142128071913971399336315466373189521847368796023166393113740678309482464924111701407630496623109664933422804502046797817118948219100673035047419935721212391974606554246228929618928476;
            6'd2: xpb[13] = 1024'd87718676487791271233209614528311210067991470573327237723816196996395321731390349952064122625263212081711129235006980823712914284256143827942798672630932746379043694737592046332786227481356618964929848223402815260993246219329866845609004093595634237896438201346070094839871442424783949213108492457859237856952;
            6'd3: xpb[13] = 1024'd7511319047562165451015494387652382357288778734255172457592440429616087259776386018081112723237143813123544445052977800990307585542995407359037883930068078634874867536816852161549102030517722726084574726716983045125508478773903495448527570710221907577837398604988084229700635563247290802544048860163262301097;
            6'd4: xpb[13] = 1024'd51370657291457801067620301651807987391284514020918791319500538927813748125471560994113174035868749853979109062556468212846764727671067321330437220245534451824396714905612875327942215771196032208549498838418390675622131588438836918253029617508039026526056499278023131649636356775639265409098295089092881229573;
            6'd5: xpb[13] = 1024'd95229995535353436684225108915963592425280249307582410181408637426011408991166735970145235348500355894834673680059958624703221869799139235301836556561000825013918562274408898494335329511874341691014422950119798306118754698103770341057531664305856145474275599951058179069572077988031240015652541318022500158049;
            6'd6: xpb[13] = 1024'd15022638095124330902030988775304764714577557468510344915184880859232174519552772036162225446474287626247088890105955601980615171085990814718075767860136157269749735073633704323098204061035445452169149453433966090251016957547806990897055141420443815155674797209976168459401271126494581605088097720326524602194;
            6'd7: xpb[13] = 1024'd58881976339019966518635796039460369748573292755173963777092979357429835385247947012194286759105893667102653507609446013837072313214062728689475104175602530459271582442429727489491317801713754934634073565135373720747640067212740413701557188218260934103893897883011215879336992338886556211642343949256143530670;
            6'd8: xpb[13] = 1024'd102741314582915602135240603303615974782569028041837582639001077855627496250943121988226348071737499707958218125112936425693529455342134642660874440491068903648793429811225750655884431542392064417098997676836781351244263176877673836506059235016078053052112998556046263299272713551278530818196590178185762459146;
            6'd9: xpb[13] = 1024'd22533957142686496353046483162957147071866336202765517372777321288848261779329158054243338169711431439370633335158933402970922756628986222077113651790204235904624602610450556484647306091553168178253724180150949135376525436321710486345582712130665722733512195814964252689101906689741872407632146580489786903291;
            6'd10: xpb[13] = 1024'd66393295386582131969651290427112752105862071489429136234685419787045922645024333030275399482343037480226197952662423814827379898757058136048512988105670609094146449979246579651040419832231477660718648291852356765873148545986643909150084758928482841681731296487999300109037627902133847014186392809419405831767;
            6'd11: xpb[13] = 1024'd110252633630477767586256097691268357139857806776092755096593518285243583510719508006307460794974643521081762570165914226683837040885130050019912324421136982283668297348042602817433533572909787143183572403553764396369771655651577331954586805726299960629950397161034347528973349114525821620740639038349024760243;
            6'd12: xpb[13] = 1024'd30045276190248661804061977550609529429155114937020689830369761718464349039105544072324450892948575252494177780211911203961230342171981629436151535720272314539499470147267408646196408122070890904338298906867932180502033915095613981794110282840887630311349594419952336918802542252989163210176195440653049204388;
            6'd13: xpb[13] = 1024'd73904614434144297420666784814765134463150850223684308692277860216662009904800719048356512205580181293349742397715401615817687484300053543407550872035738687729021317516063431812589521862749200386803223018569339810998657024760547404598612329638704749259568695092987384338738263465381137816730441669582668132864;
            6'd14: xpb[13] = 1024'd117763952678039933037271592078920739497146585510347927554185958714859670770495894024388573518211787334205307015218892027674144626428125457378950208351205060918543164884859454978982635603427509869268147130270747441495280134425480827403114376436521868207787795766022431758673984677773112423284687898512287061340;
            6'd15: xpb[13] = 1024'd37556595237810827255077471938261911786443893671275862287962202148080436298881930090405563616185719065617722225264889004951537927714977036795189419650340393174374337684084260807745510152588613630422873633584915225627542393869517477242637853551109537889186993024940421148503177816236454012720244300816311505485;
            6'd16: xpb[13] = 1024'd81415933481706462871682279202417516820439628957939481149870300646278097164577105066437624928817325106473286842768379416807995069843048950766588755965806766363896185052880283974138623893266923112887797745286322856124165503534450900047139900348926656837406093697975468568438899028628428619274490529745930433961;
            6'd17: xpb[13] = 1024'd1208576041477357089488159061758689109736937118867415883646544079498862692963141132454615026791256837885702052814376394085388371129900530182827967264942098619727357852105089802901498442428026874042524248600490640256427762978487549886663377463514326518805290956893457958268092167091770208710046932049954878106;
            6'd18: xpb[13] = 1024'd45067914285372992706092966325914294143732672405531034745554642577696523558658316108486676339422862878741266670317866805941845513257972444154227303580408471809249205220901112969294612183106336356507448360301898270753050872643420972691165424261331445467024391629928505378203813379483744815264293160979573806582;
            6'd19: xpb[13] = 1024'd88927252529268628322697773590069899177728407692194653607462741075894184424353491084518737652054468919596831287821357217798302655386044358125626639895874844998771052589697136135687725923784645838972372472003305901249673982308354395495667471059148564415243492302963552798139534591875719421818539389909192735058;
            6'd20: xpb[13] = 1024'd8719895089039522540503653449411071467025715853122588341238984509114949952739527150535727750028400651009246497867354195075695956672895937541865851195010177254602225388921941964450600472945749600127098975317473685381936241752391045335190948173736234096642689561881542187968727730339061011254095792213217179203;
            6'd21: xpb[13] = 1024'd52579233332935158157108460713566676501021451139786207203147083007312610818434702126567789062660006691864811115370844606932153098800967851513265187510476550444124072757717965130843714213624059082592023087018881315878559351417324468139692994971553353044861790234916589607904448942731035617808342021142836107679;
            6'd22: xpb[13] = 1024'd96438571576830793773713267977722281535017186426449826065055181505510271684129877102599850375291612732720375732874335018788610240929039765484664523825942923633645920126513988297236827954302368565056947198720288946375182461082257890944195041769370471993080890907951637027840170155123010224362588250072455036155;
            6'd23: xpb[13] = 1024'd16231214136601687991519147837063453824314494587377760798831424938731037212515913168616840473265544464132790942920331996066003542215891344900903735125078255889477092925738794125999702503463472326211673702034456730507444720526294540783718518883958141674480088166869626417669363293586351813798144652376479480300;
            6'd24: xpb[13] = 1024'd60090552380497323608123955101219058858310229874041379660739523436928698078211088144648901785897150504988355560423822407922460684343963258872303071440544629078998940294534817292392816244141781808676597813735864361004067830191227963588220565681775260622699188839904673837605084505978326420352390881306098408776;
            6'd25: xpb[13] = 1024'd103949890624392959224728762365374663892305965160704998522647621935126358943906263120680963098528756545843920177927312819778917826472035172843702407756011002268520787663330840458785929984820091291141521925437271991500690939856161386392722612479592379570918289512939721257540805718370301026906637110235717337252;
            6'd26: xpb[13] = 1024'd23742533184163853442534642224715836181603273321632933256423865368347124472292299186697953196502688277256335387973309797056311127758886752259941619055146334524351960462555646287548804533981195052296248428751439775632953199300198036232246089594180049252317486771857710647369998856833642616342193512539741781397;
            6'd27: xpb[13] = 1024'd67601871428059489059139449488871441215599008608296552118331963866544785337987474162730014509134294318111900005476800208912768269886958666231340955370612707713873807831351669453941918274659504534761172540452847406129576308965131459036748136391997168200536587444892758067305720069225617222896439741469360709873;
            6'd28: xpb[13] = 1024'd111461209671955124675744256753027046249594743894960170980240062364742446203682649138762075821765900358967464622980290620769225412015030580202740291686079080903395655200147692620335032015337814017226096652154255036626199418630064881841250183189814287148755688117927805487241441281617591829450685970398979638349;
            6'd29: xpb[13] = 1024'd31253852231726018893550136612368218538892052055888105714016305797963211732068685204779065919739832090379879833026287598046618713301882159618979502985214413159226827999372498449097906564498917778380823155468422820758461678074101531680773660304401956830154885376845794877070634420080933418886242372703004082494;
            6'd30: xpb[13] = 1024'd75113190475621654510154943876523823572887787342551724575924404296160872597763860180811127232371438131235444450529778009903075855429954073590378839300680786348748675368168521615491020305177227260845747267169830451255084787739034954485275707102219075778373986049880842297006355632472908025440488601632623010970;
            6'd31: xpb[13] = 1024'd118972528719517290126759751140679428606883522629215343437832502794358533463459035156843188545003044172091009068033268421759532997558025987561778175616147159538270522736964544781884134045855536743310671378871238081751707897403968377289777753900036194726593086722915889716942076844864882631994734830562241939446;
            6'd32: xpb[13] = 1024'd38765171279288184344565631000020600896180830790143278171608746227579298991845071222860178642976975903503424278079265399036926298844877566978017386915282491794101695536189350610647008595016640504465397882185405865883970156848005027129301231014623864407992283981833879106771269983328224221430291232866266383591;
            6'd33: xpb[13] = 1024'd82624509523183819961170438264176205930176566076806897033516844725776959857540246198892239955608581944358988895582755810893383440972949480949416723230748864983623542904985373777040122335694949986930321993886813496380593266512938449933803277812440983356211384654868926526706991195720198827984537461795885312067;
            6'd34: xpb[13] = 1024'd2417152082954714178976318123517378219473874237734831767293088158997725385926282264909230053582513675771404105628752788170776742259801060365655934529884197239454715704210179605802996884856053748085048497200981280512855525956975099773326754927028653037610581913786915916536184334183540417420093864099909756212;
            6'd35: xpb[13] = 1024'd46276490326850349795581125387672983253469609524398450629201186657195386251621457240941291366214119716626968723132243200027233884387872974337055270845350570428976563073006202772196110625534363230549972608902388911009478635621908522577828801724845771985829682586821963336471905546575515023974340093029528684688;
            6'd36: xpb[13] = 1024'd90135828570745985412185932651828588287465344811062069491109285155393047117316632216973352678845725757482533340635733611883691026515944888308454607160816943618498410441802225938589224366212672713014896720603796541506101745286841945382330848522662890934048783259857010756407626758967489630528586321959147613164;
            6'd37: xpb[13] = 1024'd9928471130516879629991812511169760576762652971990004224885528588613812645702668282990342776819657488894948550681730589161084327802796467724693818459952275874329583241027031767352098915373776474169623223917964325638364004730878595221854325637250560615447980518775000146236819897430831219964142724263172057309;
            6'd38: xpb[13] = 1024'd53787809374412515246596619775325365610758388258653623086793627086811473511397843259022404089451263529750513168185221001017541469930868381696093154775418649063851430609823054933745212656052085956634547335619371956134987114395812018026356372435067679563667081191810047566172541109822805826518388953192790985785;
            6'd39: xpb[13] = 1024'd97647147618308150863201427039480970644754123545317241948701725585009134377093018235054465402082869570606077785688711412873998612058940295667492491090885022253373277978619078100138326396730395439099471447320779586631610224060745440830858419232884798511886181864845094986108262322214780433072635182122409914261;
            6'd40: xpb[13] = 1024'd17439790178079045081007306898822142934051431706245176682477969018229899905479054301071455500056801302018492995734708390151391913345791875083731702390020354509204450777843883928901200945891499200254197950634947370763872483504782090670381896347472468193285379123763084375937455460678122022508191584426434358406;
            6'd41: xpb[13] = 1024'd61299128421974680697612114162977747968047166992908795544386067516427560771174229277103516812688407342874057613238198802007849055473863789055131038705486727698726298146639907095294314686569808682719122062336355001260495593169715513474883943145289587141504479796798131795873176673070096629062437813356053286882;
            6'd42: xpb[13] = 1024'd105158466665870316314216921427133353002042902279572414406294166014625221636869404253135578125320013383729622230741689213864306197601935703026530375020953100888248145515435930261687428427248118165184046174037762631757118702834648936279385989943106706089723580469833179215808897885462071235616684042285672215358;
            6'd43: xpb[13] = 1024'd24951109225641210532022801286474525291340210440500349140070409447845987165255440319152568223293945115142037440787686191141699498888787282442769586320088433144079318314660736090450302976409221926338772677351930415889380962278685586118909467057694375771122777728751168605638091023925412825052240444589696659503;
            6'd44: xpb[13] = 1024'd68810447469536846148627608550630130325335945727163968001978507946043648030950615295184629535925551155997602058291176602998156641016859196414168922635554806333601165683456759256843416717087531408803696789053338046386004071943619008923411513855511494719341878401786216025573812236317387431606486673519315587979;
            6'd45: xpb[13] = 1024'd112669785713432481765232415814785735359331681013827586863886606444241308896645790271216690848557157196853166675794667014854613783144931110385568258951021179523123013052252782423236530457765840891268620900754745676882627181608552431727913560653328613667560979074821263445509533448709362038160732902448934516455;
            6'd46: xpb[13] = 1024'd32462428273203375983038295674126907648628989174755521597662849877462074425031826337233680946531088928265581885840663992132007084431782689801807470250156511778954185851477588251999405006926944652423347404068913461014889441052589081567437037767916283348960176333739252835338726587172703627596289304752958960600;
            6'd47: xpb[13] = 1024'd76321766517099011599643102938282512682624724461419140459570948375659735290727001313265742259162694969121146503344154403988464226559854603773206806565622884968476033220273611418392518747605254134888271515770321091511512550717522504371939084565733402297179277006774300255274447799564678234150535533682577889076;
            6'd48: xpb[13] = 1024'd120181104760994647216247910202438117716620459748082759321479046873857396156422176289297803571794301009976711120847644815844921368687926517744606142881089258157997880589069634584785632488283563617353195627471728722008135660382455927176441131363550521245398377679809347675210169011956652840704781762612196817552;
            6'd49: xpb[13] = 1024'd39973747320765541434053790061779290005917767909010694055255290307078161684808212355314793669768232741389126330893641793122314669974778097160845354180224590413829053388294440413548507037444667378507922130785896506140397919826492577015964608478138190926797574938727337065039362150419994430140338164916221261697;
            6'd50: xpb[13] = 1024'd83833085564661177050658597325934895039913503195674312917163388805275822550503387331346854982399838782244690948397132204978771812102850011132244690495690963603350900757090463579941620778122976860972846242487304136637021029491425999820466655275955309875016675611762384484975083362811969036694584393845840190173;
            6'd51: xpb[13] = 1024'd3625728124432071268464477185276067329210811356602247650939632238496588078889423397363845080373770513657106158443129182256165113389701590548483901794826295859182073556315269408704495327284080622127572745801471920769283288935462649659990132390542979556415872870680373874804276501275310626130140796149864634318;
            6'd52: xpb[13] = 1024'd47485066368327706885069284449431672363206546643265866512847730736694248944584598373395906393005376554512670775946619594112622255517773504519883238110292669048703920925111292575097609067962390104592496857502879551265906398600396072464492179188360098504634973543715421294739997713667285232684387025079483562794;
            6'd53: xpb[13] = 1024'd91344404612223342501674091713587277397202281929929485374755829234891909810279773349427967705636982595368235393450110005969079397645845418491282574425759042238225768293907315741490722808640699587057420969204287181762529508265329495268994225986177217452854074216750468714675718926059259839238633254009102491270;
            6'd54: xpb[13] = 1024'd11137047171994236719479971572928449686499590090857420108532072668112675338665809415444957803610914326780650603496106983246472698932696997907521785724894374494056941093132121570253597357801803348212147472518454965894791767709366145108517703100764887134253271475668458104504912064522601428674189656313126935415;
            6'd55: xpb[13] = 1024'd54996385415889872336084778837084054720495325377521038970440171166310336204360984391477019116242520367636215220999597395102929841060768911878921122040360747683578788461928144736646711098480112830677071584219862596391414877374299567913019749898582006082472372148703505524440633276914576035228435885242745863891;
            6'd56: xpb[13] = 1024'd98855723659785507952689586101239659754491060664184657832348269664507997070056159367509080428874126408491779838503087806959386983188840825850320458355827120873100635830724167903039824839158422313141995695921270226888037987039232990717521796696399125030691472821738552944376354489306550641782682114172364792367;
            6'd57: xpb[13] = 1024'd18648366219556402170495465960580832043788368825112592566124513097728762598442195433526070526848058139904195048549084784236780284475692405266559669654962453128931808629948973731802699388319526074296722199235438011020300246483269640557045273810986794712090670080656542334205547627769892231218238516476389236512;
            6'd58: xpb[13] = 1024'd62507704463452037787100273224736437077784104111776211428032611595926423464137370409558131839479664180759759666052575196093237426603764319237959005970428826318453655998744996898195813128997835556761646310936845641516923356148203063361547320608803913660309770753691589754141268840161866837772484745406008164988;
            6'd59: xpb[13] = 1024'd106367042707347673403705080488892042111779839398439830289940710094124084329832545385590193152111270221615324283556065607949694568731836233209358342285895199507975503367541020064588926869676145039226570422638253272013546465813136486166049367406621032608528871426726637174076990052553841444326730974335627093464;
            6'd60: xpb[13] = 1024'd26159685267118567621510960348233214401077147559367765023716953527344849858218581451607183250085201953027739493602062585227087870018687812625597553585030531763806676166765825893351801418837248800381296925952421056145808725257173136005572844521208702289928068685644626563906183191017183033762287376639651537609;
            6'd61: xpb[13] = 1024'd70019023511014203238115767612388819435072882846031383885625052025542510723913756427639244562716807993883304111105552997083545012146759726596996889900496904953328523535561849059744915159515558282846221037653828686642431834922106558810074891319025821238147169358679673983841904403409157640316533605569270466085;
            6'd62: xpb[13] = 1024'd113878361754909838854720574876544424469068618132695002747533150523740171589608931403671305875348414034738868728609043408940002154274831640568396226215963278142850370904357872226138028900193867765311145149355236317139054944587039981614576938116842940186366270031714721403777625615801132246870779834498889394561;
            6'd63: xpb[13] = 1024'd33671004314680733072526454735885596758365926293622937481309393956960937117994967469688295973322345766151283938655040386217395455561683219984635437515098610398681543703582678054900903449354971526465871652669404101271317204031076631454100415231430609867765467290632710793606818754264473836306336236802913838706;
        endcase
    end

    always_comb begin
        case(flag[4][16:12])
            5'd0: xpb[14] = 1024'd0;
            5'd1: xpb[14] = 1024'd77530342558576368689131262000041201792361661580286556343217492455158597983690142445720357285953951807006848556158530798073852597689755133956034773830564983588203391072378701221294017190033281008930795764370811731767940313696010054258602462029247728815984567963667758213542539966656448442860582465732532767182;
            5'd2: xpb[14] = 1024'd30993989433027995979463596595267970840024896034837428558303129845340300630071145981425643357250229304570547704859568161568641354538289933356909422644798926242716107575186185104957795188549356296551393920354383617171519777171123335552226354375266008365149232513218458396978551859384263868602475104839471050033;
            5'd3: xpb[14] = 1024'd108524331991604364668594858595309172632386557615123984901520622300498898613761288427146000643204181111577396261018098959642493952228045067312944196475363909830919498647564886326251812378582637305482189684725195348939460090867133389810828816404513737181133800476886216610521091826040712311463057570572003817215;
            5'd4: xpb[14] = 1024'd61987978866055991958927193190535941680049792069674857116606259690680601260142291962851286714500458609141095409719136323137282709076579866713818845289597852485432215150372370209915590377098712593102787840708767234343039554342246671104452708750532016730298465026436916793957103718768527737204950209678942100066;
            5'd5: xpb[14] = 1024'd15451625740507619249259527785762710727713026524225729331691897080862303906523295498556572785796736106704794558420173686632071465925114666114693494103831795139944931653179854093579368375614787880723385996692339119746619017817359952398076601096550296279463129575987616977393115611496343162946842848785880382917;
            5'd6: xpb[14] = 1024'd92981968299083987938390789785803912520074688104512285674909389536020901890213437944276930071750687913711643114578704484705924063614869800070728267934396778728148322725558555314873385565648068889654181761063150851514559331513370006656679063125798025095447697539655375190935655578152791605807425314518413150099;
            5'd7: xpb[14] = 1024'd46445615173535615228723124381030681567737922559063157889995026926202604536594441479982216143046965411275342263279741848200712820463404599471602916748630721382661039228366039198537163564164144177274779917046722736918138794988483287950302955471816304644612362089206075374371667470880607031549317953625351432950;
            5'd8: xpb[14] = 1024'd123975957732111983917854386381071883360099584139349714233212519381361202520284583925702573429000917218282190819438272646274565418153159733427637690579195704970864430300744740419831180754197425186205575681417534468686079108684493342208905417501064033460596930052873833587914207437537055474409900419357884200132;
            5'd9: xpb[14] = 1024'd77439604606563611208186720976298652407762818593900586448298156771542905166665587461407859500297194715845889968139310009769354175001694532828512339393429647625377146803552224303494958752713500473826173837401106354089658572159606623502529309847082313009761594602424533771350219330264870900151793058464822482983;
            5'd10: xpb[14] = 1024'd30903251481015238498519055571525421455426053048451458663383794161724607813046590997113145571593472213409589116840347373264142931850229332229386988207663590279889863306359708187158736751229575761446771993384678239493238035634719904796153202193100592558926259151975233954786231222992686325893685697571760765834;
            5'd11: xpb[14] = 1024'd108433594039591607187650317571566623247787714628738015006601286616883205796736733442833502857547424020416437672998878171337995529539984466185421762038228573868093254378738409408452753941262856770377567757755489971261178349330729959054755664222348321374910827115642992168328771189649134768754268163304293533016;
            5'd12: xpb[14] = 1024'd61897240914043234477982652166793392295450949083288887221686924007064908443117736978538788928843701517980136821699915534832784286388519265586296410852462516522605970881545893292116531939778932057998165913739061856664757812805843240348379556568366600924075491665193692351764783082376950194496160802411231815867;
            5'd13: xpb[14] = 1024'd15360887788494861768314986762020161343114183537839759436772561397246611089498740514244075000139979015543835970400952898327573043237054064987171059666696459177118687384353377175780309938295007345618764069722633742068337276280956521642003448914384880473240156214744392535200794975104765620238053441518170098718;
            5'd14: xpb[14] = 1024'd92891230347071230457446248762061363135475845118126315779990053852405209073188882959964432286093930822550684526559483696401425640926809198943205833497261442765322078456732078397074327128328288354549559834093445473836277589976966575900605910943632609289224724178412150748743334941761214063098635907250702865900;
            5'd15: xpb[14] = 1024'd46354877221522857747778583357288132183139079572677187995075691242586911719569886495669718357390208320114383675260521059896214397775343998344080482311495385419834794959539562280738105126844363642170157990077017359239857053452079857194229803289650888838389388727962850932179346834489029488840528546357641148751;
            5'd16: xpb[14] = 1024'd123885219780099226436909845357329333975500741152963744338293183697745509703260028941390075643344160127121232231419051857970066995465099132300115256142060369008038186031918263502032122316877644651100953754447829091007797367148089911452832265318898617654373956691630609145721886801145477931701111012090173915933;
            5'd17: xpb[14] = 1024'd77348866654550853727242179952556103023163975607514616553378821087927212349641032477095361714640437624684931380120089221464855752313633931700989904956294311662550902534725747385695900315393719938721551910431400976411376830623203192746456157664916897203538621241181309329157898693873293357443003651197112198784;
            5'd18: xpb[14] = 1024'd30812513529002481017574514547782872070827210062065488768464458478108914996022036012800647785936715122248630528821126584959644509162168731101864553770528254317063619037533231269359678313909795226342150066414972861814956294098316474040080050010935176752703285790732009512593910586601108783184896290304050481635;
            5'd19: xpb[14] = 1024'd108342856087578849706705776547824073863188871642352045111681950933267512979712178458521005071890666929255479084979657383033497106851923865057899327601093237905267010109911932490653695503943076235272945830785784593582896607794326528298682512040182905568687853754399767726136450553257557226045478756036583248817;
            5'd20: xpb[14] = 1024'd61806502962030476997038111143050842910852106096902917326767588323449215626093181994226291143186944426819178233680694746528285863700458664458773976415327180559779726612719416374317473502459151522893543986769356478986476071269439809592306404386201185117852518303950467909572462445985372651787371395143521531668;
            5'd21: xpb[14] = 1024'd15270149836482104287370445738277611958515340551453789541853225713630918272474185529931577214483221924382877382381732110023074620548993463859648625229561123214292443115526900257981251500975226810514142142752928364390055534744553090885930296732219464667017182853501168093008474338713188077529264034250459814519;
            5'd22: xpb[14] = 1024'd92800492395058472976501707738318813750877002131740345885070718168789516256164327975651934500437173731389725938540262908096927218238748597815683399060126106802495834187905601479275268691008507819444937907123740096157995848440563145144532758761467193483001750817168926306551014305369636520389846499982992581701;
            5'd23: xpb[14] = 1024'd46264139269510100266834042333545582798540236586291218100156355558971218902545331511357220571733451228953425087241300271591715975087283397216558047874360049457008550690713085362939046689524583107065536063107311981561575311915676426438156651107485473032166415366719626489987026198097451946131739139089930864552;
            5'd24: xpb[14] = 1024'd123794481828086468955965304333586784590901898166577774443373848014129816886235473957077577857687403035960273643399831069665568572777038531172592821704925033045211941763091786584233063879557864115996331827478123713329515625611686480696759113136733201848150983330387384703529566164753900388992321604822463631734;
            5'd25: xpb[14] = 1024'd77258128702538096246297638928813553638565132621128646658459485404311519532616477492782863928983680533523972792100868433160357329625573330573467470519158975699724658265899270467896841878073939403616929983461695598733095089086799761990383005482751481397315647879938084886965578057481715814734214243929401914585;
            5'd26: xpb[14] = 1024'd30721775576989723536629973524040322686228367075679518873545122794493222178997481028488150000279958031087671940801905796655146086474108129974342119333392918354237374768706754351560619876590014691237528139445267484136674552561913043284006897828769760946480312429488785070401589950209531240476106883036340197436;
            5'd27: xpb[14] = 1024'd108252118135566092225761235524081524478590028655966075216762615249651820162687623474208507286233909838094520496960436594728998684163863263930376893163957901942440765841085455572854637066623295700168323903816079215904614866257923097542609359858017489762464880393156543283944129916865979683336689348768872964618;
            5'd28: xpb[14] = 1024'd61715765010017719516093570119308293526253263110516947431848252639833522809068627009913793357530187335658219645661473958223787441012398063331251541978191844596953482343892939456518415065139370987788922059799651101308194329733036378836233252204035769311629544942707243467380141809593795109078581987875811247469;
            5'd29: xpb[14] = 1024'd15179411884469346806425904714535062573916497565067819646933890030015225455449630545619079428826464833221918794362511321718576197860932862732126190792425787251466198846700423340182193063655446275409520215783222986711773793208149660129857144550054048860794209492257943650816153702321610534820474626982749530320;
            5'd30: xpb[14] = 1024'd92709754443045715495557166714576264366278159145354375990151382485173823439139772991339436714780416640228767350521042119792428795550687996688160964622990770839669589919079124561476210253688727284340315980154034718479714106904159714388459606579301777676778777455925701864358693668978058977681057092715282297502;
            5'd31: xpb[14] = 1024'd46173401317497342785889501309803033413941393599905248205237019875355526085520776527044722786076694137792466499222079483287217552399222796089035613437224713494182306421886608445139988252204802571960914136137606603883293570379272995682083498925320057225943442005476402047794705561705874403422949731822220580353;
        endcase
    end

    always_comb begin
        case(flag[5][5:0])
            6'd0: xpb[15] = 1024'd0;
            6'd1: xpb[15] = 1024'd123885219780099226436909845357329333975500741152963744338293183697745509703260028941390075643344160127121232231419051857970066995465099132300115256142060369008038186031918263502032122316877644651100953754447829091007797367148089911452832265318898617654373956691630609145721886801145477931701111012090173915933;
            6'd2: xpb[15] = 1024'd123703743876073711475020763309844235206303055180191804548454512330514124069210918972765080072030645944799315055380610281361070150088977930045070387267789697082385697494265309666434005442238083580891709900508418335651233884075283049940685960954567786041928009969144160261337245528362322846283532197554753347535;
            6'd3: xpb[15] = 1024'd123522267972048196513131681262359136437105369207419864758615840963282738435161809004140084500717131762477397879342168704752073304712856727790025518393519025156733208956612355830835888567598522510682466046569007580294670401002476188428539656590236954429482063246657711376952604255579167760865953383019332779137;
            6'd4: xpb[15] = 1024'd123340792068022681551242599214874037667907683234647924968777169596051352801112699035515088929403617580155480703303727128143076459336735525534980649519248353231080720418959401995237771692958961440473222192629596824938106917929669326916393352225906122817036116524171262492567962982796012675448374568483912210739;
            6'd5: xpb[15] = 1024'd123159316163997166589353517167388938898709997261875985178938498228819967167063589066890093358090103397833563527265285551534079613960614323279935780644977681305428231881306448159639654818319400370263978338690186069581543434856862465404247047861575291204590169801684813608183321710012857590030795753948491642341;
            6'd6: xpb[15] = 1024'd122977840259971651627464435119903840129512311289104045389099826861588581533014479098265097786776589215511646351226843974925082768584493121024890911770707009379775743343653494324041537943679839300054734484750775314224979951784055603892100743497244459592144223079198364723798680437229702504613216939413071073943;
            6'd7: xpb[15] = 1024'd122796364355946136665575353072418741360314625316332105599261155494357195898965369129640102215463075033189729175188402398316085923208371918769846042896436337454123254806000540488443421069040278229845490630811364558868416468711248742379954439132913627979698276356711915839414039164446547419195638124877650505545;
            6'd8: xpb[15] = 1024'd122614888451920621703686271024933642591116939343560165809422484127125810264916259161015106644149560850867811999149960821707089077832250716514801174022165665528470766268347586652845304194400717159636246776871953803511852985638441880867808134768582796367252329634225466955029397891663392333778059310342229937147;
            6'd9: xpb[15] = 1024'd122433412547895106741797188977448543821919253370788226019583812759894424630867149192390111072836046668545894823111519245098092232456129514259756305147894993602818277730694632817247187319761156089427002922932543048155289502565635019355661830404251964754806382911739018070644756618880237248360480495806809368749;
            6'd10: xpb[15] = 1024'd122251936643869591779908106929963445052721567398016286229745141392663038996818039223765115501522532486223977647073077668489095387080008312004711436273624321677165789193041678981649070445121595019217759068993132292798726019492828157843515526039921133142360436189252569186260115346097082162942901681271388800351;
            6'd11: xpb[15] = 1024'd122070460739844076818019024882478346283523881425244346439906470025431653362768929255140119930209018303902060471034636091880098541703887109749666567399353649751513300655388725146050953570482033949008515215053721537442162536420021296331369221675590301529914489466766120301875474073313927077525322866735968231953;
            6'd12: xpb[15] = 1024'd121888984835818561856129942834993247514326195452472406650067798658200267728719819286515124358895504121580143294996194515271101696327765907494621698525082977825860812117735771310452836695842472878799271361114310782085599053347214434819222917311259469917468542744279671417490832800530771992107744052200547663555;
            6'd13: xpb[15] = 1024'd121707508931793046894240860787508148745128509479700466860229127290968882094670709317890128787581989939258226118957752938662104850951644705239576829650812305900208323580082817474854719821202911808590027507174900026729035570274407573307076612946928638305022596021793222533106191527747616906690165237665127095157;
            6'd14: xpb[15] = 1024'd121526033027767531932351778740023049975930823506928527070390455923737496460621599349265133216268475756936308942919311362053108005575523502984531960776541633974555835042429863639256602946563350738380783653235489271372472087201600711794930308582597806692576649299306773648721550254964461821272586423129706526759;
            6'd15: xpb[15] = 1024'd121344557123742016970462696692537951206733137534156587280551784556506110826572489380640137644954961574614391766880869785444111160199402300729487091902270962048903346504776909803658486071923789668171539799296078516015908604128793850282784004218266975080130702576820324764336908982181306735855007608594285958361;
            6'd16: xpb[15] = 1024'd121163081219716502008573614645052852437535451561384647490713113189274725192523379412015142073641447392292474590842428208835114314823281098474442223028000290123250857967123955968060369197284228597962295945356667760659345121055986988770637699853936143467684755854333875879952267709398151650437428794058865389963;
            6'd17: xpb[15] = 1024'd120981605315690987046684532597567753668337765588612707700874441822043339558474269443390146502327933209970557414803986632226117469447159896219397354153729618197598369429471002132462252322644667527753052091417257005302781637983180127258491395489605311855238809131847426995567626436614996565019849979523444821565;
            6'd18: xpb[15] = 1024'd120800129411665472084795450550082654899140079615840767911035770454811953924425159474765150931014419027648640238765545055617120624071038693964352485279458946271945880891818048296864135448005106457543808237477846249946218154910373265746345091125274480242792862409360978111182985163831841479602271164988024253167;
            6'd19: xpb[15] = 1024'd120618653507639957122906368502597556129942393643068828121197099087580568290376049506140155359700904845326723062727103479008123778694917491709307616405188274346293392354165094461266018573365545387334564383538435494589654671837566404234198786760943648630346915686874529226798343891048686394184692350452603684769;
            6'd20: xpb[15] = 1024'd120437177603614442161017286455112457360744707670296888331358427720349182656326939537515159788387390663004805886688661902399126933318796289454262747530917602420640903816512140625667901698725984317125320529599024739233091188764759542722052482396612817017900968964388080342413702618265531308767113535917183116371;
            6'd21: xpb[15] = 1024'd120255701699588927199128204407627358591547021697524948541519756353117797022277829568890164217073876480682888710650220325790130087942675087199217878656646930494988415278859186790069784824086423246916076675659613983876527705691952681209906178032281985405455022241901631458029061345482376223349534721381762547973;
            6'd22: xpb[15] = 1024'd120074225795563412237239122360142259822349335724753008751681084985886411388228719600265168645760362298360971534611778749181133242566553884944173009782376258569335926741206232954471667949446862176706832821720203228519964222619145819697759873667951153793009075519415182573644420072699221137931955906846341979575;
            6'd23: xpb[15] = 1024'd119892749891537897275350040312657161053151649751981068961842413618655025754179609631640173074446848116039054358573337172572136397190432682689128140908105586643683438203553279118873551074807301106497588967780792473163400739546338958185613569303620322180563128796928733689259778799916066052514377092310921411177;
            6'd24: xpb[15] = 1024'd119711273987512382313460958265172062283953963779209129172003742251423640120130499663015177503133333933717137182534895595963139551814311480434083272033834914718030949665900325283275434200167740036288345113841381717806837256473532096673467264939289490568117182074442284804875137527132910967096798277775500842779;
            6'd25: xpb[15] = 1024'd119529798083486867351571876217686963514756277806437189382165070884192254486081389694390181931819819751395220006496454019354142706438190278179038403159564242792378461128247371447677317325528178966079101259901970962450273773400725235161320960574958658955671235351955835920490496254349755881679219463240080274381;
            6'd26: xpb[15] = 1024'd119348322179461352389682794170201864745558591833665249592326399516960868852032279725765186360506305569073302830458012442745145861062069075923993534285293570866725972590594417612079200450888617895869857405962560207093710290327918373649174656210627827343225288629469387036105854981566600796261640648704659705983;
            6'd27: xpb[15] = 1024'd119166846275435837427793712122716765976360905860893309802487728149729483217983169757140190789192791386751385654419570866136149015685947873668948665411022898941073484052941463776481083576249056825660613552023149451737146807255111512137028351846296995730779341906982938151721213708783445710844061834169239137585;
            6'd28: xpb[15] = 1024'd118985370371410322465904630075231667207163219888121370012649056782498097583934059788515195217879277204429468478381129289527152170309826671413903796536752227015420995515288509940882966701609495755451369698083738696380583324182304650624882047481966164118333395184496489267336572436000290625426483019633818569187;
            6'd29: xpb[15] = 1024'd118803894467384807504015548027746568437965533915349430222810385415266711949884949819890199646565763022107551302342687712918155324933705469158858927662481555089768506977635556105284849826969934685242125844144327941024019841109497789112735743117635332505887448462010040382951931163217135540008904205098398000789;
            6'd30: xpb[15] = 1024'd118622418563359292542126465980261469668767847942577490432971714048035326315835839851265204075252248839785634126304246136309158479557584266903814058788210883164116018439982602269686732952330373615032881990204917185667456358036690927600589438753304500893441501739523591498567289890433980454591325390562977432391;
            6'd31: xpb[15] = 1024'd118440942659333777580237383932776370899570161969805550643133042680803940681786729882640208503938734657463716950265804559700161634181463064648769189913940211238463529902329648434088616077690812544823638136265506430310892874963884066088443134388973669280995555017037142614182648617650825369173746576027556863993;
            6'd32: xpb[15] = 1024'd118259466755308262618348301885291272130372475997033610853294371313572555047737619914015212932625220475141799774227362983091164788805341862393724321039669539312811041364676694598490499203051251474614394282326095674954329391891077204576296830024642837668549608294550693729798007344867670283756167761492136295595;
            6'd33: xpb[15] = 1024'd118077990851282747656459219837806173361174790024261671063455699946341169413688509945390217361311706292819882598188921406482167943429220660138679452165398867387158552827023740762892382328411690404405150428386684919597765908818270343064150525660312006056103661572064244845413366072084515198338588946956715727197;
            6'd34: xpb[15] = 1024'd117896514947257232694570137790321074591977104051489731273617028579109783779639399976765221789998192110497965422150479829873171098053099457883634583291128195461506064289370786927294265453772129334195906574447274164241202425745463481552004221295981174443657714849577795961028724799301360112921010132421295158799;
            6'd35: xpb[15] = 1024'd117715039043231717732681055742835975822779418078717791483778357211878398145590290008140226218684677928176048246112038253264174252676978255628589714416857523535853575751717833091696148579132568263986662720507863408884638942672656620039857916931650342831211768127091347076644083526518205027503431317885874590401;
            6'd36: xpb[15] = 1024'd117533563139206202770791973695350877053581732105945851693939685844647012511541180039515230647371163745854131070073596676655177407300857053373544845542586851610201087214064879256098031704493007193777418866568452653528075459599849758527711612567319511218765821404604898192259442253735049942085852503350454022003;
            6'd37: xpb[15] = 1024'd117352087235180687808902891647865778284384046133173911904101014477415626877492070070890235076057649563532213894035155100046180561924735851118499976668316179684548598676411925420499914829853446123568175012629041898171511976527042897015565308202988679606319874682118449307874800980951894856668273688815033453605;
            6'd38: xpb[15] = 1024'd117170611331155172847013809600380679515186360160401972114262343110184241243442960102265239504744135381210296717996713523437183716548614648863455107794045507758896110138758971584901797955213885053358931158689631142814948493454236035503419003838657847993873927959632000423490159708168739771250694874279612885207;
            6'd39: xpb[15] = 1024'd116989135427129657885124727552895580745988674187630032324423671742952855609393850133640243933430621198888379541958271946828186871172493446608410238919774835833243621601106017749303681080574323983149687304750220387458385010381429173991272699474327016381427981237145551539105518435385584685833116059744192316809;
            6'd40: xpb[15] = 1024'd116807659523104142923235645505410481976790988214858092534585000375721469975344740165015248362117107016566462365919830370219190025796372244353365370045504163907591133063453063913705564205934762912940443450810809632101821527308622312479126395109996184768982034514659102654720877162602429600415537245208771748411;
            6'd41: xpb[15] = 1024'd116626183619078627961346563457925383207593302242086152744746329008490084341295630196390252790803592834244545189881388793610193180420251042098320501171233491981938644525800110078107447331295201842731199596871398876745258044235815450966980090745665353156536087792172653770336235889819274514997958430673351180013;
            6'd42: xpb[15] = 1024'd116444707715053112999457481410440284438395616269314212954907657641258698707246520227765257219490078651922628013842947217001196335044129839843275632296962820056286155988147156242509330456655640772521955742931988121388694561163008589454833786381334521544090141069686204885951594617036119429580379616137930611615;
            6'd43: xpb[15] = 1024'd116263231811027598037568399362955185669197930296542273165068986274027313073197410259140261648176564469600710837804505640392199489668008637588230763422692148130633667450494202406911213582016079702312711888992577366032131078090201727942687482017003689931644194347199756001566953344252964344162800801602510043217;
            6'd44: xpb[15] = 1024'd116081755907002083075679317315470086900000244323770333375230314906795927439148300290515266076863050287278793661766064063783202644291887435333185894548421476204981178912841248571313096707376518632103468035053166610675567595017394866430541177652672858319198247624713307117182312071469809258745221987067089474819;
            6'd45: xpb[15] = 1024'd115900280002976568113790235267984988130802558350998393585391643539564541805099190321890270505549536104956876485727622487174205798915766233078141025674150804279328690375188294735714979832736957561894224181113755855319004111944588004918394873288342026706752300902226858232797670798686654173327643172531668906421;
            6'd46: xpb[15] = 1024'd115718804098951053151901153220499889361604872378226453795552972172333156171050080353265274934236021922634959309689180910565208953539645030823096156799880132353676201837535340900116862958097396491684980327174345099962440628871781143406248568924011195094306354179740409348413029525903499087910064357996248338023;
            6'd47: xpb[15] = 1024'd115537328194925538190012071173014790592407186405454514005714300805101770537000970384640279362922507740313042133650739333956212108163523828568051287925609460428023713299882387064518746083457835421475736473234934344605877145798974281894102264559680363481860407457253960464028388253120344002492485543460827769625;
            6'd48: xpb[15] = 1024'd115355852290900023228122989125529691823209500432682574215875629437870384902951860416015283791608993557991124957612297757347215262787402626313006419051338788502371224762229433228920629208818274351266492619295523589249313662726167420381955960195349531869414460734767511579643746980337188917074906728925407201227;
            6'd49: xpb[15] = 1024'd115174376386874508266233907078044593054011814459910634426036958070638999268902750447390288220295479375669207781573856180738218417411281424057961550177068116576718736224576479393322512334178713281057248765356112833892750179653360558869809655831018700256968514012281062695259105707554033831657327914389986632829;
            6'd50: xpb[15] = 1024'd114992900482848993304344825030559494284814128487138694636198286703407613634853640478765292648981965193347290605535414604129221572035160221802916681302797444651066247686923525557724395459539152210848004911416702078536186696580553697357663351466687868644522567289794613810874464434770878746239749099854566064431;
            6'd51: xpb[15] = 1024'd114811424578823478342455742983074395515616442514366754846359615336176228000804530510140297077668451011025373429496973027520224726659039019547871812428526772725413759149270571722126278584899591140638761057477291323179623213507746835845517047102357037032076620567308164926489823161987723660822170285319145496033;
            6'd52: xpb[15] = 1024'd114629948674797963380566660935589296746418756541594815056520943968944842366755420541515301506354936828703456253458531450911227881282917817292826943554256100799761270611617617886528161710260030070429517203537880567823059730434939974333370742738026205419630673844821716042105181889204568575404591470783724927635;
            6'd53: xpb[15] = 1024'd114448472770772448418677578888104197977221070568822875266682272601713456732706310572890305935041422646381539077420089874302231035906796615037782074679985428874108782073964664050930044835620469000220273349598469812466496247362133112821224438373695373807184727122335267157720540616421413489987012656248304359237;
            6'd54: xpb[15] = 1024'd114266996866746933456788496840619099208023384596050935476843601234482071098657200604265310363727908464059621901381648297693234190530675412782737205805714756948456293536311710215331927960980907930011029495659059057109932764289326251309078134009364542194738780399848818273335899343638258404569433841712883790839;
            6'd55: xpb[15] = 1024'd114085520962721418494899414793134000438825698623278995687004929867250685464608090635640314792414394281737704725343206721084237345154554210527692336931444085022803804998658756379733811086341346859801785641719648301753369281216519389796931829645033710582292833677362369388951258070855103319151855027177463222441;
            6'd56: xpb[15] = 1024'd113904045058695903533010332745648901669628012650507055897166258500019299830558980667015319221100880099415787549304765144475240499778433008272647468057173413097151316461005802544135694211701785789592541787780237546396805798143712528284785525280702878969846886954875920504566616798071948233734276212642042654043;
            6'd57: xpb[15] = 1024'd113722569154670388571121250698163802900430326677735116107327587132787914196509870698390323649787365917093870373266323567866243654402311806017602599182902741171498827923352848708537577337062224719383297933840826791040242315070905666772639220916372047357400940232389471620181975525288793148316697398106622085645;
            6'd58: xpb[15] = 1024'd113541093250644873609232168650678704131232640704963176317488915765556528562460760729765328078473851734771953197227881991257246809026190603762557730308632069245846339385699894872939460462422663649174054079901416035683678831998098805260492916552041215744954993509903022735797334252505638062899118583571201517247;
            6'd59: xpb[15] = 1024'd113359617346619358647343086603193605362034954732191236527650244398325142928411650761140332507160337552450036021189440414648249963650069401507512861434361397320193850848046941037341343587783102578964810225962005280327115348925291943748346612187710384132509046787416573851412692979722482977481539769035780948849;
            6'd60: xpb[15] = 1024'd113178141442593843685454004555708506592837268759419296737811573031093757294362540792515336935846823370128118845150998838039253118273948199252467992560090725394541362310393987201743226713143541508755566372022594524970551865852485082236200307823379552520063100064930124967028051706939327892063960954500360380451;
            6'd61: xpb[15] = 1024'd112996665538568328723564922508223407823639582786647356947972901663862371660313430823890341364533309187806201669112557261430256272897826996997423123685820053468888873772741033366145109838503980438546322518083183769613988382779678220724054003459048720907617153342443676082643410434156172806646382139964939812053;
            6'd62: xpb[15] = 1024'd112815189634542813761675840460738309054441896813875417158134230296630986026264320855265345793219795005484284493074115684821259427521705794742378254811549381543236385235088079530546992963864419368337078664143773014257424899706871359211907699094717889295171206619957227198258769161373017721228803325429519243655;
            6'd63: xpb[15] = 1024'd112633713730517298799786758413253210285244210841103477368295558929399600392215210886640350221906280823162367317035674108212262582145584592487333385937278709617583896697435125694948876089224858298127834810204362258900861416634064497699761394730387057682725259897470778313874127888589862635811224510894098675257;
        endcase
    end

    always_comb begin
        case(flag[5][11:6])
            6'd0: xpb[16] = 1024'd0;
            6'd1: xpb[16] = 1024'd112452237826491783837897676365768111516046524868331537578456887562168214758166100918015354650592766640840450140997232531603265736769463390232288517063008037691931408159782171859350759214585297227918590956264951503544297933561257636187615090366056226070279313174984329429489486615806707550393645696358678106859;
            6'd2: xpb[16] = 1024'd100837779968858826276996425326721790287394622610927391028781920059359534179023062926015638086527858972237750874536971628627467632697706445909416909109685034450172141749993126381071279237653388734526984304142663160724235016901618499410251611048883002873738722935851600828872445157684782083668601566091761729387;
            6'd3: xpb[16] = 1024'd89223322111225868716095174287675469058742720353523244479106952556550853599880024934015921522462951303635051608076710725651669528625949501586545301156362031208412875340204080902791799260721480241135377652020374817904172100241979362632888131731709779677198132696718872228255403699562856616943557435824845351915;
            6'd4: xpb[16] = 1024'd77608864253592911155193923248629147830090818096119097929431985053742173020736986942016204958398043635032352341616449822675871424554192557263673693203039027966653608930415035424512319283789571747743770999898086475084109183582340225855524652414536556480657542457586143627638362241440931150218513305557928974443;
            6'd5: xpb[16] = 1024'd65994406395959953594292672209582826601438915838714951379757017550933492441593948950016488394333135966429653075156188919700073320482435612940802085249716024724894342520625989946232839306857663254352164347775798132264046266922701089078161173097363333284116952218453415027021320783319005683493469175291012596971;
            6'd6: xpb[16] = 1024'd54379948538326996033391421170536505372787013581310804830082050048124811862450910958016771830268228297826953808695928016724275216410678668617930477296393021483135076110836944467953359329925754760960557695653509789443983350263061952300797693780190110087576361979320686426404279325197080216768425045024096219499;
            6'd7: xpb[16] = 1024'd42765490680694038472490170131490184144135111323906658280407082545316131283307872966017055266203320629224254542235667113748477112338921724295058869343070018241375809701047898989673879352993846267568951043531221446623920433603422815523434214463016886891035771740187957825787237867075154750043380914757179842027;
            6'd8: xpb[16] = 1024'd31151032823061080911588919092443862915483209066502511730732115042507450704164834974017338702138412960621555275775406210772679008267164779972187261389747014999616543291258853511394399376061937774177344391408933103803857516943783678746070735145843663694495181501055229225170196408953229283318336784490263464555;
            6'd9: xpb[16] = 1024'd19536574965428123350687668053397541686831306809098365181057147539698770125021796982017622138073505292018856009315145307796880904195407835649315653436424011757857276881469808033114919399130029280785737739286644760983794600284144541968707255828670440497954591261922500624553154950831303816593292654223347087083;
            6'd10: xpb[16] = 1024'd7922117107795165789786417014351220458179404551694218631382180036890089545878758990017905574008597623416156742854884404821082800123650891326444045483101008516098010471680762554835439422198120787394131087164356418163731683624505405191343776511497217301414001022789772023936113492709378349868248523956430709611;
            6'd11: xpb[16] = 1024'd120374354934286949627684093380119331974225929420025756209839067599058304304044859908033260224601364264256606883852116936424348536893114281558732562546109046208029418631462934414186198636783418015312722043429307921708029617185763041378958866877553443371693314197774101453425600108516085900261894220315108816470;
            6'd12: xpb[16] = 1024'd108759897076653992066782842341073010745574027162621609660164100096249623724901821916033543660536456595653907617391856033448550432821357337235860954592786042966270152221673888935906718659851509521921115391307019578887966700526123904601595387560380220175152723958641372852808558650394160433536850090048192438998;
            6'd13: xpb[16] = 1024'd97145439219021034505881591302026689516922124905217463110489132593440943145758783924033827096471548927051208350931595130472752328749600392912989346639463039724510885811884843457627238682919601028529508739184731236067903783866484767824231908243206996978612133719508644252191517192272234966811805959781276061526;
            6'd14: xpb[16] = 1024'd85530981361388076944980340262980368288270222647813316560814165090632262566615745932034110532406641258448509084471334227496954224677843448590117738686140036482751619402095797979347758705987692535137902087062442893247840867206845631046868428926033773782071543480375915651574475734150309500086761829514359684054;
            6'd15: xpb[16] = 1024'd73916523503755119384079089223934047059618320390409170011139197587823581987472707940034393968341733589845809818011073324521156120606086504267246130732817033240992352992306752501068278729055784041746295434940154550427777950547206494269504949608860550585530953241243187050957434276028384033361717699247443306582;
            6'd16: xpb[16] = 1024'd62302065646122161823177838184887725830966418133005023461464230085014901408329669948034677404276825921243110551550812421545358016534329559944374522779494029999233086582517707022788798752123875548354688782817866207607715033887567357492141470291687327388990363002110458450340392817906458566636673568980526929110;
            6'd17: xpb[16] = 1024'd50687607788489204262276587145841404602314515875600876911789262582206220829186631956034960840211918252640411285090551518569559912462572615621502914826171026757473820172728661544509318775191967054963082130695577864787652117227928220714777990974514104192449772762977729849723351359784533099911629438713610551638;
            6'd18: xpb[16] = 1024'd39073149930856246701375336106795083373662613618196730362114295079397540250043593964035244276147010584037712018630290615593761808390815671298631306872848023515714553762939616066229838798260058561571475478573289521967589200568289083937414511657340880995909182523845001249106309901662607633186585308446694174166;
            6'd19: xpb[16] = 1024'd27458692073223289140474085067748762145010711360792583812439327576588859670900555972035527712082102915435012752170029712617963704319058726975759698919525020273955287353150570587950358821328150068179868826451001179147526283908649947160051032340167657799368592284712272648489268443540682166461541178179777796694;
            6'd20: xpb[16] = 1024'd15844234215590331579572834028702440916358809103388437262764360073780179091757517980035811148017195246832313485709768809642165600247301782652888090966202017032196020943361525109670878844396241574788262174328712836327463367249010810382687553022994434602828002045579544047872226985418756699736497047912861419222;
            6'd21: xpb[16] = 1024'd4229776357957374018671582989656119687706906845984290713089392570971498512614479988036094583952287578229614219249507906666367496175544838330016483012879013790436754533572479631391398867464333081396655522206424493507400450589371673605324073705821211406287411806446815447255185527296831233011452917645945041750;
            6'd22: xpb[16] = 1024'd116682014184449157856569259355424231203753431714315828291546280133139713270780580906051449234545054219070064360246740438269633232945008228562305000075887051482368162693354651490742158082049630309315246478471375997051698384150629309792939164071877437476566724981431144876744672143103538783405098614004623148609;
            6'd23: xpb[16] = 1024'd105067556326816200295668008316377909975101529456911681741871312630331032691637542914051732670480146550467365093786479535293835128873251284239433392122564048240608896283565606012462678105117721815923639826349087654231635467490990173015575684754704214280026134742298416276127630684981613316680054483737706771137;
            6'd24: xpb[16] = 1024'd93453098469183242734766757277331588746449627199507535192196345127522352112494504922052016106415238881864665827326218632318037024801494339916561784169241044998849629873776560534183198128185813322532033174226799311411572550831351036238212205437530991083485544503165687675510589226859687849955010353470790393665;
            6'd25: xpb[16] = 1024'd81838640611550285173865506238285267517797724942103388642521377624713671533351466930052299542350331213261966560865957729342238920729737395593690176215918041757090363463987515055903718151253904829140426522104510968591509634171711899460848726120357767886944954264032959074893547768737762383229966223203874016193;
            6'd26: xpb[16] = 1024'd70224182753917327612964255199238946289145822684699242092846410121904990954208428938052582978285423544659267294405696826366440816657980451270818568262595038515331097054198469577624238174321996335748819869982222625771446717512072762683485246803184544690404364024900230474276506310615836916504922092936957638721;
            6'd27: xpb[16] = 1024'd58609724896284370052063004160192625060493920427295095543171442619096310375065390946052866414220515876056568027945435923390642712586223506947946960309272035273571830644409424099344758197390087842357213217859934282951383800852433625906121767486011321493863773785767501873659464852493911449779877962670041261249;
            6'd28: xpb[16] = 1024'd46995267038651412491161753121146303831842018169890948993496475116287629795922352954053149850155608207453868761485175020414844608514466562625075352355949032031812564234620378621065278220458179348965606565737645940131320884192794489128758288168838098297323183546634773273042423394371985983054833832403124883777;
            6'd29: xpb[16] = 1024'd35380809181018454930260502082099982603190115912486802443821507613478949216779314962053433286090700538851169495024914117439046504442709618302203744402626028790053297824831333142785798243526270855573999913615357597311257967533155352351394808851664875100782593307502044672425381936250060516329789702136208506305;
            6'd30: xpb[16] = 1024'd23766351323385497369359251043053661374538213655082655894146540110670268637636276970053716722025792870248470228564653214463248400370952673979332136449303025548294031415042287664506318266594362362182393261493069254491195050873516215574031329534491651904242003068369316071808340478128135049604745571869292128833;
            6'd31: xpb[16] = 1024'd12151893465752539808458000004007340145886311397678509344471572607861588058493238978054000157960885201645770962104392311487450296299195729656460528495980022306534765005253242186226838289662453868790786609370780911671132134213877078796667850217318428707701412829236587471191299020006209582879701441602375751361;
            6'd32: xpb[16] = 1024'd537435608119582247556748964961018917234409140274362794796605105052907479350200986054283593895977533043071695644131408511652192227438785333588920542657019064775498595464196707947358312730545375399179957248492568851069217554237942019304370900145205511160822590103858870574257561884284116154657311335459373889;
            6'd33: xpb[16] = 1024'd112989673434611366085454425330729130433280934008605900373253492667221122237516301904069638244488744173883521836641363940114917928996902175565877437605665056756706906755246368567298117527315842603317770913513444072395367151115495578206919461266201431581440135765088188300063744177690991666548303007694137480748;
            6'd34: xpb[16] = 1024'd101375215576978408524553174291682809204629031751201753823578525164412441658373263912069921680423836505280822570181103037139119824925145231243005829652342053514947640345457323089018637550383934109926164261391155729575304234455856441429555981949028208384899545525955459699446702719569066199823258877427221103276;
            6'd35: xpb[16] = 1024'd89760757719345450963651923252636487975977129493797607273903557661603761079230225920070205116358928836678123303720842134163321720853388286920134221699019050273188373935668277610739157573452025616534557609268867386755241317796217304652192502631854985188358955286822731098829661261447140733098214747160304725804;
            6'd36: xpb[16] = 1024'd78146299861712493402750672213590166747325227236393460724228590158795080500087187928070488552294021168075424037260581231187523616781631342597262613745696047031429107525879232132459677596520117123142950957146579043935178401136578167874829023314681761991818365047690002498212619803325215266373170616893388348332;
            6'd37: xpb[16] = 1024'd66531842004079535841849421174543845518673324978989314174553622655986399920944149936070771988229113499472724770800320328211725512709874398274391005792373043789669841116090186654180197619588208629751344305024290701115115484476939031097465543997508538795277774808557273897595578345203289799648126486626471970860;
            6'd38: xpb[16] = 1024'd54917384146446578280948170135497524290021422721585167624878655153177719341801111944071055424164205830870025504340059425235927408638117453951519397839050040547910574706301141175900717642656300136359737652902002358295052567817299894320102064680335315598737184569424545296978536887081364332923082356359555593388;
            6'd39: xpb[16] = 1024'd43302926288813620720046919096451203061369520464181021075203687650369038762658073952071338860099298162267326237879798522260129304566360509628647789885727037306151308296512095697621237665724391642968131000779714015474989651157660757542738585363162092402196594330291816696361495428959438866198038226092639215916;
            6'd40: xpb[16] = 1024'd31688468431180663159145668057404881832717618206776874525528720147560358183515035960071622296034390493664626971419537619284331200494603565305776181932404034064392041886723050219341757688792483149576524348657425672654926734498021620765375106045988869205656004091159088095744453970837513399472994095825722838444;
            6'd41: xpb[16] = 1024'd20074010573547705598244417018358560604065715949372727975853752644751677604371997968071905731969482825061927704959276716308533096422846620982904573979081030822632775476934004741062277711860574656184917696535137329834863817838382483988011626728815646009115413852026359495127412512715587932747949965558806460972;
            6'd42: xpb[16] = 1024'd8459552715914748037343165979312239375413813691968581426178785141942997025228959976072189167904575156459228438499015813332734992351089676660032966025758027580873509067144959262782797734928666162793311044412848987014800901178743347210648147411642422812574823612893630894510371054593662466022905835291890083500;
            6'd43: xpb[16] = 1024'd120911790542406531875240842345080350891460338560300119004635672704111211783395060894087543818497341797299678579496248344936000729120553066892321483088766065272804917226927131122133556949513963390711902000677800490559098834740000983398263237777698648882854136787877960323999857670400370016416551531650568190359;
            6'd44: xpb[16] = 1024'd109297332684773574314339591306034029662808436302895972454960705201302531204252022902087827254432434128696979313035987441960202625048796122569449875135443062031045650817138085643854076972582054897320295348555512147739035918080361846620899758460525425686313546548745231723382816212278444549691507401383651812887;
            6'd45: xpb[16] = 1024'd97682874827140616753438340266987708434156534045491825905285737698493850625108984910088110690367526460094280046575726538984404520977039178246578267182120058789286384407349040165574596995650146403928688696433223804918973001420722709843536279143352202489772956309612503122765774754156519082966463271116735435415;
            6'd46: xpb[16] = 1024'd86068416969507659192537089227941387205504631788087679355610770195685170045965946918088394126302618791491580780115465636008606416905282233923706659228797055547527117997559994687295117018718237910537082044310935462098910084761083573066172799826178979293232366070479774522148733296034593616241419140849819057943;
            6'd47: xpb[16] = 1024'd74453959111874701631635838188895065976852729530683532805935802692876489466822908926088677562237711122888881513655204733032808312833525289600835051275474052305767851587770949209015637041786329417145475392188647119278847168101444436288809320509005756096691775831347045921531691837912668149516375010582902680471;
            6'd48: xpb[16] = 1024'd62839501254241744070734587149848744748200827273279386256260835190067808887679870934088960998172803454286182247194943830057010208761768345277963443322151049064008585177981903730736157064854420923753868740066358776458784251441805299511445841191832532900151185592214317320914650379790742682791330880315986302999;
            6'd49: xpb[16] = 1024'd51225043396608786509833336110802423519548925015875239706585867687259128308536832942089244434107895785683482980734682927081212104690011400955091835368828045822249318768192858252456677087922512430362262087944070433638721334782166162734082361874659309703610595353081588720297608921668817216066286750049069925527;
            6'd50: xpb[16] = 1024'd39610585538975828948932085071756102290897022758471093156910900184450447729393794950089527870042988117080783714274422024105414000618254456632220227415505042580490052358403812774177197110990603936970655435821782090818658418122527025956718882557486086507070005113948860119680567463546891749341242619782153548055;
            6'd51: xpb[16] = 1024'd27996127681342871388030834032709781062245120501066946607235932681641767150250756958089811305978080448478084447814161121129615896546497512309348619462182039338730785948614767295897717134058695443579048783699493747998595501462887889179355403240312863310529414874816131519063526005424966282616198489515237170583;
            6'd52: xpb[16] = 1024'd16381669823709913827129582993663459833593218243662800057560965178833086571107718966090094741913172779875385181353900218153817792474740567986477011508859036096971519538825721817618237157126786950187442131577205405178532584803248752401991923923139640113988824635683402918446484547303040815891154359248320793111;
            6'd53: xpb[16] = 1024'd4767211966076956266228331954617138604941315986258653507885997676024405991964680974090378177848265111272685914893639315178019688402983623663605403555536032855212253129036676339338757180194878456795835479454917062358469668143609615624628444605966416917448234396550674317829443089181115349166110228981404415639;
            6'd54: xpb[16] = 1024'd117219449792568740104126008320385250120987840854590191086342885238192620750130781892105732828441031752113136055890871846781285425172447013895893920618544070547143661288818848198689516394780175684714426435719868565902767601704867251812243534972022642987727547571535003747318929704987822899559755925340082522498;
            6'd55: xpb[16] = 1024'd105604991934935782543224757281338928892335938597186044536667917735383940170987743900106016264376124083510436789430610943805487321100690069573022312665221067305384394879029802720410036417848267191322819783597580223082704685045228115034880055654849419791186957332402275146701888246865897432834711795073166145026;
            6'd56: xpb[16] = 1024'd93990534077302824982323506242292607663684036339781897986992950232575259591844705908106299700311216414907737522970350040829689217028933125250150704711898064063625128469240757242130556440916358697931213131475291880262641768385588978257516576337676196594646367093269546546084846788743971966109667664806249767554;
            6'd57: xpb[16] = 1024'd82376076219669867421422255203246286435032134082377751437317982729766579012701667916106583136246308746305038256510089137853891112957176180927279096758575060821865862059451711763851076463984450204539606479353003537442578851725949841480153097020502973398105776854136817945467805330622046499384623534539333390082;
            6'd58: xpb[16] = 1024'd70761618362036909860521004164199965206380231824973604887643015226957898433558629924106866572181401077702338990049828234878093008885419236604407488805252057580106595649662666285571596487052541711147999827230715194622515935066310704702789617703329750201565186615004089344850763872500121032659579404272417012610;
            6'd59: xpb[16] = 1024'd59147160504403952299619753125153643977728329567569458337968047724149217854415591932107150008116493409099639723589567331902294904813662292281535880851929054338347329239873620807292116510120633217756393175108426851802453018406671567925426138386156527005024596375871360744233722414378195565934535274005500635138;
            6'd60: xpb[16] = 1024'd47532702646770994738718502086107322749076427310165311788293080221340537275272553940107433444051585740496940457129306428926496800741905347958664272898606051096588062830084575329012636533188724724364786522986138508982390101747032431148062659068983303808484006136738632143616680956256270099209491143738584257666;
            6'd61: xpb[16] = 1024'd35918244789138037177817251047061001520424525052761165238618112718531856696129515948107716879986678071894241190669045525950698696670148403635792664945283047854828796420295529850733156556256816230973179870863850166162327185087393294370699179751810080611943415897605903542999639498134344632484447013471667880194;
            6'd62: xpb[16] = 1024'd24303786931505079616916000008014680291772622795357018688943145215723176116986477956108000315921770403291541924208784622974900592598391459312921056991960044613069530010506484372453676579324907737581573218741561823342264268427754157593335700434636857415402825658473174942382598040012419165759402883204751502722;
            6'd63: xpb[16] = 1024'd12689329073872122056014748968968359063120720537952872139268177712914495537843439964108283751856862734688842657748523719999102488526634514990049449038637041371310263600717438894174196602392999244189966566619273480522201351768115020815972221117463634218862235419340446341765556581890493699034358752937835125250;
        endcase
    end

    always_comb begin
        case(flag[5][16:12])
            5'd0: xpb[17] = 1024'd0;
            5'd1: xpb[17] = 1024'd1074871216239164495113497929922037834468818280548725589593210210105814958700401972108567187791955066086143391288262817023304384454877570667177841085314038129550997190928393415894716625461090750798359914496985137702138435108475884038608741800290411022321645180207717741148515123768568232309314622670918747778;
            5'd2: xpb[17] = 1024'd2149742432478328990226995859844075668937636561097451179186420420211629917400803944217134375583910132172286782576525634046608768909755141334355682170628076259101994381856786831789433250922181501596719828993970275404276870216951768077217483600580822044643290360415435482297030247537136464618629245341837495556;
            5'd3: xpb[17] = 1024'd3224613648717493485340493789766113503406454841646176768779630630317444876101205916325701563375865198258430173864788451069913153364632712001533523255942114388652991572785180247684149876383272252395079743490955413106415305325427652115826225400871233066964935540623153223445545371305704696927943868012756243334;
            5'd4: xpb[17] = 1024'd4299484864956657980453991719688151337875273122194902358372840840423259834801607888434268751167820264344573565153051268093217537819510282668711364341256152518203988763713573663578866501844363003193439657987940550808553740433903536154434967201161644089286580720830870964594060495074272929237258490683674991112;
            5'd5: xpb[17] = 1024'd5374356081195822475567489649610189172344091402743627947966051050529074793502009860542835938959775330430716956441314085116521922274387853335889205426570190647754985954641967079473583127305453753991799572484925688510692175542379420193043709001452055111608225901038588705742575618842841161546573113354593738890;
            5'd6: xpb[17] = 1024'd6449227297434986970680987579532227006812909683292353537559261260634889752202411832651403126751730396516860347729576902139826306729265424003067046511884228777305983145570360495368299752766544504790159486981910826212830610650855304231652450801742466133929871081246306446891090742611409393855887736025512486668;
            5'd7: xpb[17] = 1024'd7524098513674151465794485509454264841281727963841079127152471470740704710902813804759970314543685462603003739017839719163130691184142994670244887597198266906856980336498753911263016378227635255588519401478895963914969045759331188270261192602032877156251516261454024188039605866379977626165202358696431234446;
            5'd8: xpb[17] = 1024'd8598969729913315960907983439376302675750546244389804716745681680846519669603215776868537502335640528689147130306102536186435075639020565337422728682512305036407977527427147327157733003688726006386879315975881101617107480867807072308869934402323288178573161441661741929188120990148545858474516981367349982224;
            5'd9: xpb[17] = 1024'd9673840946152480456021481369298340510219364524938530306338891890952334628303617748977104690127595594775290521594365353209739460093898136004600569767826343165958974718355540743052449629149816757185239230472866239319245915976282956347478676202613699200894806621869459670336636113917114090783831604038268730002;
            5'd10: xpb[17] = 1024'd10748712162391644951134979299220378344688182805487255895932102101058149587004019721085671877919550660861433912882628170233043844548775706671778410853140381295509971909283934158947166254610907507983599144969851377021384351084758840386087418002904110223216451802077177411485151237685682323093146226709187477780;
            5'd11: xpb[17] = 1024'd11823583378630809446248477229142416179157001086035981485525312311163964545704421693194239065711505726947577304170890987256348229003653277338956251938454419425060969100212327574841882880071998258781959059466836514723522786193234724424696159803194521245538096982284895152633666361454250555402460849380106225558;
            5'd12: xpb[17] = 1024'd12898454594869973941361975159064454013625819366584707075118522521269779504404823665302806253503460793033720695459153804279652613458530848006134093023768457554611966291140720990736599505533089009580318973963821652425661221301710608463304901603484932267859742162492612893782181485222818787711775472051024973336;
            5'd13: xpb[17] = 1024'd13973325811109138436475473088986491848094637647133432664711732731375594463105225637411373441295415859119864086747416621302956997913408418673311934109082495684162963482069114406631316130994179760378678888460806790127799656410186492501913643403775343290181387342700330634930696608991387020021090094721943721114;
            5'd14: xpb[17] = 1024'd15048197027348302931588971018908529682563455927682158254304942941481409421805627609519940629087370925206007478035679438326261382368285989340489775194396533813713960672997507822526032756455270511177038802957791927829938091518662376540522385204065754312503032522908048376079211732759955252330404717392862468892;
            5'd15: xpb[17] = 1024'd16123068243587467426702468948830567517032274208230883843898153151587224380506029581628507816879325991292150869323942255349565766823163560007667616279710571943264957863925901238420749381916361261975398717454777065532076526627138260579131127004356165334824677703115766117227726856528523484639719340063781216670;
            5'd16: xpb[17] = 1024'd17197939459826631921815966878752605351501092488779609433491363361693039339206431553737075004671281057378294260612205072372870151278041130674845457365024610072815955054854294654315466007377452012773758631951762203234214961735614144617739868804646576357146322883323483858376241980297091716949033962734699964448;
            5'd17: xpb[17] = 1024'd18272810676065796416929464808674643185969910769328335023084573571798854297906833525845642192463236123464437651900467889396174535732918701342023298450338648202366952245782688070210182632838542763572118546448747340936353396844090028656348610604936987379467968063531201599524757104065659949258348585405618712226;
            5'd18: xpb[17] = 1024'd19347681892304960912042962738596681020438729049877060612677783781904669256607235497954209380255191189550581043188730706419478920187796272009201139535652686331917949436711081486104899258299633514370478460945732478638491831952565912694957352405227398401789613243738919340673272227834228181567663208076537460004;
            5'd19: xpb[17] = 1024'd20422553108544125407156460668518718854907547330425786202270993992010484215307637470062776568047146255636724434476993523442783304642673842676378980620966724461468946627639474901999615883760724265168838375442717616340630267061041796733566094205517809424111258423946637081821787351602796413876977830747456207782;
            5'd20: xpb[17] = 1024'd21497424324783289902269958598440756689376365610974511791864204202116299174008039442171343755839101321722867825765256340466087689097551413343556821706280762591019943818567868317894332509221815015967198289939702754042768702169517680772174836005808220446432903604154354822970302475371364646186292453418374955560;
            5'd21: xpb[17] = 1024'd22572295541022454397383456528362794523845183891523237381457414412222114132708441414279910943631056387809011217053519157489392073552428984010734662791594800720570941009496261733789049134682905766765558204436687891744907137277993564810783577806098631468754548784362072564118817599139932878495607076089293703338;
            5'd22: xpb[17] = 1024'd23647166757261618892496954458284832358314002172071962971050624622327929091408843386388478131423011453895154608341781974512696458007306554677912503876908838850121938200424655149683765760143996517563918118933673029447045572386469448849392319606389042491076193964569790305267332722908501110804921698760212451116;
            5'd23: xpb[17] = 1024'd24722037973500783387610452388206870192782820452620688560643834832433744050109245358497045319214966519981297999630044791536000842462184125345090344962222876979672935391353048565578482385605087268362278033430658167149184007494945332888001061406679453513397839144777508046415847846677069343114236321431131198894;
            5'd24: xpb[17] = 1024'd25796909189739947882723950318128908027251638733169414150237045042539559008809647330605612507006921586067441390918307608559305226917061696012268186047536915109223932582281441981473199011066178019160637947927643304851322442603421216926609803206969864535719484324985225787564362970445637575423550944102049946672;
            5'd25: xpb[17] = 1024'd26871780405979112377837448248050945861720457013718139739830255252645373967510049302714179694798876652153584782206570425582609611371939266679446027132850953238774929773209835397367915636527268769958997862424628442553460877711897100965218545007260275558041129505192943528712878094214205807732865566772968694450;
            5'd26: xpb[17] = 1024'd27946651622218276872950946177972983696189275294266865329423465462751188926210451274822746882590831718239728173494833242605913995826816837346623868218164991368325926964138228813262632261988359520757357776921613580255599312820372985003827286807550686580362774685400661269861393217982774040042180189443887442228;
            5'd27: xpb[17] = 1024'd29021522838457441368064444107895021530658093574815590919016675672857003884910853246931314070382786784325871564783096059629218380281694408013801709303479029497876924155066622229157348887449450271555717691418598717957737747928848869042436028607841097602684419865608379011009908341751342272351494812114806190006;
            5'd28: xpb[17] = 1024'd30096394054696605863177942037817059365126911855364316508609885882962818843611255219039881258174741850412014956071358876652522764736571978680979550388793067627427921345995015645052065512910541022354077605915583855659876183037324753081044770408131508625006065045816096752158423465519910504660809434785724937784;
            5'd29: xpb[17] = 1024'd31171265270935770358291439967739097199595730135913042098203096093068633802311657191148448445966696916498158347359621693675827149191449549348157391474107105756978918536923409060946782138371631773152437520412568993362014618145800637119653512208421919647327710226023814493306938589288478736970124057456643685562;
            5'd30: xpb[17] = 1024'd32246136487174934853404937897661135034064548416461767687796306303174448761012059163257015633758651982584301738647884510699131533646327120015335232559421143886529915727851802476841498763832722523950797434909554131064153053254276521158262254008712330669649355406231532234455453713057046969279438680127562433340;
            5'd31: xpb[17] = 1024'd33321007703414099348518435827583172868533366697010493277389516513280263719712461135365582821550607048670445129936147327722435918101204690682513073644735182016080912918780195892736215389293813274749157349406539268766291488362752405196870995809002741691971000586439249975603968836825615201588753302798481181118;
        endcase
    end

    always_comb begin
        case(flag[6][5:0])
            6'd0: xpb[18] = 1024'd0;
            6'd1: xpb[18] = 1024'd17197939459826631921815966878752605351501092488779609433491363361693039339206431553737075004671281057378294260612205072372870151278041130674845457365024610072815955054854294654315466007377452012773758631951762203234214961735614144617739868804646576357146322883323483858376241980297091716949033962734699964448;
            6'd2: xpb[18] = 1024'd34395878919653263843631933757505210703002184977559218866982726723386078678412863107474150009342562114756588521224410144745740302556082261349690914730049220145631910109708589308630932014754904025547517263903524406468429923471228289235479737609293152714292645766646967716752483960594183433898067925469399928896;
            6'd3: xpb[18] = 1024'd51593818379479895765447900636257816054503277466338828300474090085079118017619294661211225014013843172134882781836615217118610453834123392024536372095073830218447865164562883962946398022132356038321275895855286609702644885206842433853219606413939729071438968649970451575128725940891275150847101888204099893344;
            6'd4: xpb[18] = 1024'd68791757839306527687263867515010421406004369955118437733965453446772157356825726214948300018685124229513177042448820289491480605112164522699381829460098440291263820219417178617261864029509808051095034527807048812936859846942456578470959475218586305428585291533293935433504967921188366867796135850938799857792;
            6'd5: xpb[18] = 1024'd85989697299133159609079834393763026757505462443898047167456816808465196696032157768685375023356405286891471303061025361864350756390205653374227286825123050364079775274271473271577330036887260063868793159758811016171074808678070723088699344023232881785731614416617419291881209901485458584745169813673499822240;
            6'd6: xpb[18] = 1024'd103187636758959791530895801272515632109006554932677656600948180170158236035238589322422450028027686344269765563673230434237220907668246784049072744190147660436895730329125767925892796044264712076642551791710573219405289770413684867706439212827879458142877937299940903150257451881782550301694203776408199786688;
            6'd7: xpb[18] = 1024'd120385576218786423452711768151268237460507647421457266034439543531851275374445020876159525032698967401648059824285435506610091058946287914723918201555172270509711685383980062580208262051642164089416310423662335422639504732149299012324179081632526034500024260183264387008633693862079642018643237739142899751136;
            6'd8: xpb[18] = 1024'd13516819994488313975728807625206410067310312784501191339799051828567419376342313519881528822712574149583204677440147144403897369383108710843603533903865839648836965869263139896893488867502410380879871447226857779509358843664016383976940380753943161590350679652470812836903407768448100718473581875252005231253;
            6'd9: xpb[18] = 1024'd30714759454314945897544774503959015418811405273280800773290415190260458715548745073618603827383855206961498938052352216776767520661149841518448991268890449721652920924117434551208954874879862393653630079178619982743573805399630528594680249558589737947497002535794296695279649748745192435422615837986705195701;
            6'd10: xpb[18] = 1024'd47912698914141577819360741382711620770312497762060410206781778551953498054755176627355678832055136264339793198664557289149637671939190972193294448633915059794468875978971729205524420882257314406427388711130382185977788767135244673212420118363236314304643325419117780553655891729042284152371649800721405160149;
            6'd11: xpb[18] = 1024'd65110638373968209741176708261464226121813590250840019640273141913646537393961608181092753836726417321718087459276762361522507823217232102868139905998939669867284831033826023859839886889634766419201147343082144389212003728870858817830159987167882890661789648302441264412032133709339375869320683763456105124597;
            6'd12: xpb[18] = 1024'd82308577833794841662992675140216831473314682739619629073764505275339576733168039734829828841397698379096381719888967433895377974495273233542985363363964279940100786088680318514155352897012218431974905975033906592446218690606472962447899855972529467018935971185764748270408375689636467586269717726190805089045;
            6'd13: xpb[18] = 1024'd99506517293621473584808642018969436824815775228399238507255868637032616072374471288566903846068979436474675980501172506268248125773314364217830820728988890012916741143534613168470818904389670444748664606985668795680433652342087107065639724777176043376082294069088232128784617669933559303218751688925505053493;
            6'd14: xpb[18] = 1024'd116704456753448105506624608897722042176316867717178847940747231998725655411580902842303978850740260493852970241113377578641118277051355494892676278094013500085732696198388907822786284911767122457522423238937430998914648614077701251683379593581822619733228616952411715987160859650230651020167785651660205017941;
            6'd15: xpb[18] = 1024'd9835700529149996029641648371660214783119533080222773246106740295441799413478195486025982640753867241788115094268089216434924587488176291012361610442707069224857976683671985139471511727627368748985984262501953355784502725592418623336140892703239746823555036421618141815430573556599109719998129787769310498058;
            6'd16: xpb[18] = 1024'd27033639988976627951457615250412820134620625569002382679598103657134838752684627039763057645425148299166409354880294288807794738766217421687207067807731679297673931738526279793786977735004820761759742894453715559018717687328032767953880761507886323180701359304941625673806815536896201436947163750504010462506;
            6'd17: xpb[18] = 1024'd44231579448803259873273582129165425486121718057781992113089467018827878091891058593500132650096429356544703615492499361180664890044258552362052525172756289370489886793380574448102443742382272774533501526405477762252932649063646912571620630312532899537847682188265109532183057517193293153896197713238710426954;
            6'd18: xpb[18] = 1024'd61429518908629891795089549007918030837622810546561601546580830380520917431097490147237207654767710413922997876104704433553535041322299683036897982537780899443305841848234869102417909749759724787307260158357239965487147610799261057189360499117179475894994005071588593390559299497490384870845231675973410391402;
            6'd19: xpb[18] = 1024'd78627458368456523716905515886670636189123903035341210980072193742213956770303921700974282659438991471301292136716909505926405192600340813711743439902805509516121796903089163756733375757137176800081018790309002168721362572534875201807100367921826052252140327954912077248935541477787476587794265638708110355850;
            6'd20: xpb[18] = 1024'd95825397828283155638721482765423241540624995524120820413563557103906996109510353254711357664110272528679586397329114578299275343878381944386588897267830119588937751957943458411048841764514628812854777422260764371955577534270489346424840236726472628609286650838235561107311783458084568304743299601442810320298;
            6'd21: xpb[18] = 1024'd113023337288109787560537449644175846892126088012900429847054920465600035448716784808448432668781553586057880657941319650672145495156423075061434354632854729661753707012797753065364307771892080825628536054212526575189792496006103491042580105531119204966432973721559044965688025438381660021692333564177510284746;
            6'd22: xpb[18] = 1024'd6154581063811678083554489118114019498928753375944355152414428762316179450614077452170436458795160333993025511096031288465951805593243871181119686981548298800878987498080830382049534587752327117092097077777048932059646607520820862695341404652536332056759393190765470793957739344750118721522677700286615764863;
            6'd23: xpb[18] = 1024'd23352520523638310005370455996866624850429845864723964585905792124009218789820509005907511463466441391371319771708236360838821956871285001855965144346572908873694942552935125036365000595129779129865855709728811135293861569256435007313081273457182908413905716074088954652333981325047210438471711663021315729311;
            6'd24: xpb[18] = 1024'd40550459983464941927186422875619230201930938353503574019397155485702258129026940559644586468137722448749614032320441433211692108149326132530810601711597518946510897607789419690680466602507231142639614341680573338528076530992049151930821142261829484771052038957412438510710223305344302155420745625756015693759;
            6'd25: xpb[18] = 1024'd57748399443291573849002389754371835553432030842283183452888518847395297468233372113381661472809003506127908292932646505584562259427367263205656059076622129019326852662643714344995932609884683155413372973632335541762291492727663296548561011066476061128198361840735922369086465285641393872369779588490715658207;
            6'd26: xpb[18] = 1024'd74946338903118205770818356633124440904933123331062792886379882209088336807439803667118736477480284563506202553544851577957432410705408393880501516441646739092142807717498008999311398617262135168187131605584097744996506454463277441166300879871122637485344684724059406227462707265938485589318813551225415622655;
            6'd27: xpb[18] = 1024'd92144278362944837692634323511877046256434215819842402319871245570781376146646235220855811482151565620884496814157056650330302561983449524555346973806671349164958762772352303653626864624639587180960890237535859948230721416198891585784040748675769213842491007607382890085838949246235577306267847513960115587103;
            6'd28: xpb[18] = 1024'd109342217822771469614450290390629651607935308308622011753362608932474415485852666774592886486822846678262791074769261722703172713261490655230192431171695959237774717827206598307942330632017039193734648869487622151464936377934505730401780617480415790199637330490706373944215191226532669023216881476694815551551;
            6'd29: xpb[18] = 1024'd2473461598473360137467329864567824214737973671665937058722117229190559487749959418314890276836453426197935927923973360496979023698311451349877763520389528376899998312489675624627557447877285485198209893052144508334790489449223102054541916601832917289963749959912799772484905132901127723047225612803921031668;
            6'd30: xpb[18] = 1024'd19671401058299992059283296743320429566239066160445546492213480590883598826956390972051965281507734483576230188536178432869849174976352582024723220885414138449715953367343970278943023455254737497971968525003906711569005451184837246672281785406479493647110072843236283630861147113198219439996259575538620996116;
            6'd31: xpb[18] = 1024'd36869340518126623981099263622073034917740158649225155925704843952576638166162822525789040286179015540954524449148383505242719326254393712699568678250438748522531908422198264933258489462632189510745727156955668914803220412920451391290021654211126070004256395726559767489237389093495311156945293538273320960564;
            6'd32: xpb[18] = 1024'd54067279977953255902915230500825640269241251138004765359196207314269677505369254079526115290850296598332818709760588577615589477532434843374414135615463358595347863477052559587573955470009641523519485788907431118037435374656065535907761523015772646361402718609883251347613631073792402873894327501008020925012;
            6'd33: xpb[18] = 1024'd71265219437779887824731197379578245620742343626784374792687570675962716844575685633263190295521577655711112970372793649988459628810475974049259592980487968668163818531906854241889421477387093536293244420859193321271650336391679680525501391820419222718549041493206735205989873054089494590843361463742720889460;
            6'd34: xpb[18] = 1024'd88463158897606519746547164258330850972243436115563984226178934037655756183782117187000265300192858713089407230984998722361329780088517104724105050345512578740979773586761148896204887484764545549067003052810955524505865298127293825143241260625065799075695364376530219064366115034386586307792395426477420853908;
            6'd35: xpb[18] = 1024'd105661098357433151668363131137083456323744528604343593659670297399348795522988548740737340304864139770467701491597203794734199931366558235398950507710537188813795728641615443550520353492141997561840761684762717727740080259862907969760981129429712375432841687259853702922742357014683678024741429389212120818356;
            6'd36: xpb[18] = 1024'd122859037817259783590179098015836061675245621093123203093161660761041834862194980294474415309535420827845995752209408867107070082644599366073795965075561798886611683696469738204835819499519449574614520316714479930974295221598522114378720998234358951789988010143177186781118598994980769741690463351946820782804;
            6'd37: xpb[18] = 1024'd15990281592961674113196137489774234282048286456167128398521169057757978864092272938196419099549027575781140605364120504900876393081420162193481297424255368025736964181752815521521046315379695866078081340279002287844149333113239486031482297355776078880314429612383612609388312901349228441520807488055926262921;
            6'd38: xpb[18] = 1024'd33188221052788306035012104368526839633549378944946737832012532419451018203298704491933494104220308633159434865976325577273746544359461292868326754789279978098552919236607110175836512322757147878851839972230764491078364294848853630649222166160422655237460752495707096467764554881646320158469841450790626227369;
            6'd39: xpb[18] = 1024'd50386160512614937956828071247279444985050471433726347265503895781144057542505136045670569108891589690537729126588530649646616695637502423543172212154304588171368874291461404830151978330134599891625598604182526694312579256584467775266962034965069231594607075379030580326140796861943411875418875413525326191817;
            6'd40: xpb[18] = 1024'd67584099972441569878644038126032050336551563922505956698995259142837096881711567599407644113562870747916023387200735722019486846915543554218017669519329198244184829346315699484467444337512051904399357236134288897546794218320081919884701903769715807951753398262354064184517038842240503592367909376260026156265;
            6'd41: xpb[18] = 1024'd84782039432268201800460005004784655688052656411285566132486622504530136220917999153144719118234151805294317647812940794392356998193584684892863126884353808317000784401169994138782910344889503917173115868086051100781009180055696064502441772574362384308899721145677548042893280822537595309316943338994726120713;
            6'd42: xpb[18] = 1024'd101979978892094833722275971883537261039553748900065175565977985866223175560124430706881794122905432862672611908425145866765227149471625815567708584249378418389816739456024288793098376352266955929946874500037813304015224141791310209120181641379008960666046044029001031901269522802834687026265977301729426085161;
            6'd43: xpb[18] = 1024'd119177918351921465644091938762289866391054841388844784999469349227916214899330862260618869127576713920050906169037350939138097300749666946242554041614403028462632694510878583447413842359644407942720633131989575507249439103526924353737921510183655537023192366912324515759645764783131778743215011264464126049609;
            6'd44: xpb[18] = 1024'd12309162127623356167108978236228038997857506751888710304828857524632358901228154904340872917590320667986051022192062576931903611186487742362239373963096597601757974996161660764099069175504654234184194155554097864119293215041641725390682809305072664113518786381530941587915478689500237443045355400573231529726;
            6'd45: xpb[18] = 1024'd29507101587449988088924945114980644349358599240668319738320220886325398240434586458077947922261601725364345282804267649304773762464528873037084831328121207674573930051015955418414535182882106246957952787505860067353508176777255870008422678109719240470665109264854425446291720669797329159994389363307931494174;
            6'd46: xpb[18] = 1024'd46705041047276620010740911993733249700859691729447929171811584248018437579641018011815022926932882782742639543416472721677643913742570003711930288693145817747389885105870250072730001190259558259731711419457622270587723138512870014626162546914365816827811432148177909304667962650094420876943423326042631458622;
            6'd47: xpb[18] = 1024'd63902980507103251932556878872485855052360784218227538605302947609711476918847449565552097931604163840120933804028677794050514065020611134386775746058170427820205840160724544727045467197637010272505470051409384473821938100248484159243902415719012393184957755031501393163044204630391512593892457288777331423070;
            6'd48: xpb[18] = 1024'd81100919966929883854372845751238460403861876707007148038794310971404516258053881119289172936275444897499228064640882866423384216298652265061621203423195037893021795215578839381360933205014462285279228683361146677056153061984098303861642284523658969542104077914824877021420446610688604310841491251512031387518;
            6'd49: xpb[18] = 1024'd98298859426756515776188812629991065755362969195786757472285674333097555597260312673026247940946725954877522325253087938796254367576693395736466660788219647965837750270433134035676399212391914298052987315312908880290368023719712448479382153328305545899250400798148360879796688590985696027790525214246731351966;
            6'd50: xpb[18] = 1024'd115496798886583147698004779508743671106864061684566366905777037694790594936466744226763322945618007012255816585865293011169124518854734526411312118153244258038653705325287428689991865219769366310826745947264671083524582985455326593097122022132952122256396723681471844738172930571282787744739559176981431316414;
            6'd51: xpb[18] = 1024'd8628042662285038221021818982681843713666727047610292211136545991506738938364036870485326735631613760190961439020004648962930829291555322530997450501937827177778985810570506006677092035629612602290306970829193440394437096970043964749883321254369249346723143150678270566442644477651246444569903313090536796531;
            6'd52: xpb[18] = 1024'd25825982122111670142837785861434449065167819536389901644627909353199778277570468424222401740302894817569255699632209721335800980569596453205842907866962437250594940865424800660992558043007064615064065602780955643628652058705658109367623190059015825703869466034001754424818886457948338161518937275825236760979;
            6'd53: xpb[18] = 1024'd43023921581938302064653752740187054416668912025169511078119272714892817616776899977959476744974175874947549960244414793708671131847637583880688365231987047323410895920279095315308024050384516627837824234732717846862867020441272253985363058863662402061015788917325238283195128438245429878467971238559936725427;
            6'd54: xpb[18] = 1024'd60221861041764933986469719618939659768170004513949120511610636076585856955983331531696551749645456932325844220856619866081541283125678714555533822597011657396226850975133389969623490057761968640611582866684480050097081982176886398603102927668308978418162111800648722141571370418542521595417005201294636689875;
            6'd55: xpb[18] = 1024'd77419800501591565908285686497692265119671097002728729945101999438278896295189763085433626754316737989704138481468824938454411434403719845230379279962036267469042806029987684623938956065139420653385341498636242253331296943912500543220842796472955554775308434683972205999947612398839613312366039164029336654323;
            6'd56: xpb[18] = 1024'd94617739961418197830101653376444870471172189491508339378593362799971935634396194639170701758988019047082432742081030010827281585681760975905224737327060877541858761084841979278254422072516872666159100130588004456565511905648114687838582665277602131132454757567295689858323854379136705029315073126764036618771;
            6'd57: xpb[18] = 1024'd111815679421244829751917620255197475822673281980287948812084726161664974973602626192907776763659300104460727002693235083200151736959802106580070194692085487614674716139696273932569888079894324678932858762539766659799726867383728832456322534082248707489601080450619173716700096359433796746264107089498736583219;
            6'd58: xpb[18] = 1024'd4946923196946720274934659729135648429475947343331874117444234458381118975499918836629780553672906852395871855847946720993958047396622902699755527040779056753799996624979351249255114895754570970396419786104289016669580978898446204109083833203665834579927499919825599544969810265802255446094451225607842063336;
            6'd59: xpb[18] = 1024'd22144862656773352196750626607888253780977039832111483550935597820074158314706350390366855558344187909774166116460151793366828198674664033374600984405803666826615951679833645903570580903132022983170178418056051219903795940634060348726823702008312410937073822803149083403346052246099347163043485188342542027784;
            6'd60: xpb[18] = 1024'd39342802116599984118566593486640859132478132320891092984426961181767197653912781944103930563015468967152460377072356865739698349952705164049446441770828276899431906734687940557886046910509474995943937050007813423138010902369674493344563570812958987294220145686472567261722294226396438879992519151077241992232;
            6'd61: xpb[18] = 1024'd56540741576426616040382560365393464483979224809670702417918324543460236993119213497841005567686750024530754637684561938112568501230746294724291899135852886972247861789542235212201512917886927008717695681959575626372225864105288637962303439617605563651366468569796051120098536206693530596941553113811941956680;
            6'd62: xpb[18] = 1024'd73738681036253247962198527244146069835480317298450311851409687905153276332325645051578080572358031081909048898296767010485438652508787425399137356500877497045063816844396529866516978925264379021491454313911337829606440825840902782580043308422252140008512791453119534978474778186990622313890587076546641921128;
            6'd63: xpb[18] = 1024'd90936620496079879884014494122898675186981409787229921284901051266846315671532076605315155577029312139287343158908972082858308803786828556073982813865902107117879771899250824520832444932641831034265212945863100032840655787576516927197783177226898716365659114336443018836851020167287714030839621039281341885576;
        endcase
    end

    always_comb begin
        case(flag[6][11:6])
            6'd0: xpb[19] = 1024'd0;
            6'd1: xpb[19] = 1024'd108134559955906511805830461001651280538482502276009530718392414628539355010738508159052230581700593196665637419521177155231178955064869686748828271230926717190695726954105119175147910940019283047038971577814862236074870749312131071815523046031545292722805437219766502695227262147584805747788655002016041850024;
            6'd2: xpb[19] = 1024'd92202424227688282212861994598488128332266577426283377308652974192101814684167877408089389948743512083888125431584860875883294069288519038942496417445522393447700779338639021012665582688521360372767745547242484625785380648403365370666067522379861136178790971025415947360347996221240978478458620177406489215717;
            6'd3: xpb[19] = 1024'd76270288499470052619893528195324976126050652576557223898913533755664274357597246657126549315786430971110613443648544596535409183512168391136164563660118069704705831723172922850183254437023437698496519516670107015495890547494599669516611998728176979634776504831065392025468730294897151209128585352796936581410;
            6'd4: xpb[19] = 1024'd60338152771251823026925061792161823919834727726831070489174093319226734031026615906163708682829349858333101455712228317187524297735817743329832709874713745961710884107706824687700926185525515024225293486097729405206400446585833968367156475076492823090762038636714836690589464368553323939798550528187383947103;
            6'd5: xpb[19] = 1024'd44406017043033593433956595388998671713618802877104917079434652882789193704455985155200868049872268745555589467775912037839639411959467095523500856089309422218715936492240726525218597934027592349954067455525351794916910345677068267217700951424808666546747572442364281355710198442209496670468515703577831312796;
            6'd6: xpb[19] = 1024'd28473881314815363840988128985835519507402878027378763669695212446351653377885354404238027416915187632778077479839595758491754526183116447717169002303905098475720988876774628362736269682529669675682841424952974184627420244768302566068245427773124510002733106248013726020830932515865669401138480878968278678489;
            6'd7: xpb[19] = 1024'd12541745586597134248019662582672367301186953177652610259955772009914113051314723653275186783958106520000565491903279479143869640406765799910837148518500774732726041261308530200253941431031747001411615394380596574337930143859536864918789904121440353458718640053663170685951666589521842131808446054358726044182;
            6'd8: xpb[19] = 1024'd120676305542503646053850123584323647839669455453662140978348186638453468062053231812327417365658699716666202911424456634375048595471635486659665419749427491923421768215413649375401852371051030048450586972195458810412800893171667936734312950152985646181524077273429673381178928737106647879597101056374767894206;
            6'd9: xpb[19] = 1024'd104744169814285416460881657181160495633453530603935987568608746202015927735482601061364576732701618603888690923488140355027163709695284838853333565964023168180426820599947551212919524119553107374179360941623081200123310792262902235584857426501301489637509611079079118046299662810762820610267066231765215259899;
            6'd10: xpb[19] = 1024'd88812034086067186867913190777997343427237605754209834158869305765578387408911970310401736099744537491111178935551824075679278823918934191047001712178618844437431872984481453050437195868055184699908134911050703589833820691354136534435401902849617333093495144884728562711420396884418993340937031407155662625592;
            6'd11: xpb[19] = 1024'd72879898357848957274944724374834191221021680904483680749129865329140847082341339559438895466787456378333666947615507796331393938142583543240669858393214520694436925369015354887954867616557262025636908880478325979544330590445370833285946379197933176549480678690378007376541130958075166071606996582546109991285;
            6'd12: xpb[19] = 1024'd56947762629630727681976257971671039014805756054757527339390424892703306755770708808476054833830375265556154959679191516983509052366232895434338004607810196951441977753549256725472539365059339351365682849905948369254840489536605132136490855546249020005466212496027452041661865031731338802276961757936557356978;
            6'd13: xpb[19] = 1024'd41015626901412498089007791568507886808589831205031373929650984456265766429200078057513214200873294152778642971742875237635624166589882247628006150822405873208447030138083158562990211113561416677094456819333570758965350388627839430987035331894564863461451746301676896706782599105387511532946926933327004722671;
            6'd14: xpb[19] = 1024'd25083491173194268496039325165344734602373906355305220519911544019828226102629447306550373567916213040001130983806558958287739280813531599821674297037001549465452082522617060400507882862063494002823230788761193148675860287719073729837579808242880706917437280107326341371903333179043684263616892108717452088364;
            6'd15: xpb[19] = 1024'd9151355444976038903070858762181582396157981505579067110172103583390685776058816555587532934959131927223618995870242678939854395037180952015342443251597225722457134907150962238025554610565571328552004758188815538386370186810308028688124284591196550373422813912975786037024067252699856994286857284107899454057;
            6'd16: xpb[19] = 1024'd117285915400882550708901319763832862934640483781588597828564518211930040786797324714639763516659725123889256415391419834171033350102050638764170714482523942913152861861256081413173465550584854375590976336003677774461240936122439100503647330622741843096228251132742288732251329400284662742075512286123941304081;
            6'd17: xpb[19] = 1024'd101353779672664321115932853360669710728424558931862444418825077775492500460226693963676922883702644011111744427455103554823148464325699990957838860697119619170157914245789983250691137299086931701319750305431300164171750835213673399354191806971057686552213784938391733397372063473940835472745477461514388669774;
            6'd18: xpb[19] = 1024'd85421643944446091522964386957506558522208634082136291009085637339054960133656063212714082250745562898334232439518787275475263578549349343151507006911715295427162966630323885088208809047589009027048524274858922553882260734304907698204736283319373530008199318744041178062492797547597008203415442636904836035467;
            6'd19: xpb[19] = 1024'd69489508216227861929995920554343406315992709232410137599346196902617419807085432461751241617788481785556720451582470996127378692772998695345175153126310971684168019014857786925726480796091086352777298244286544943592770633396141997055280759667689373464184852549690622727613531621253180934085407812295283401160;
            6'd20: xpb[19] = 1024'd53557372488009632337027454151180254109776784382683984189606756466179879480514801710788400984831400672779208463646154716779493806996648047538843299340906647941173071399391688763244152544593163678506072213714167333303280532487376295905825236016005216920170386355340067392734265694909353664755372987685730766853;
            6'd21: xpb[19] = 1024'd37625236759791402744058987748017101903560859532957830779867316029742339153944170959825560351874319560001696475709838437431608921220297399732511445555502324198178123783925590600761824293095241004234846183141789723013790431578610594756369712364321060376155920160989512057854999768565526395425338163076178132546;
            6'd22: xpb[19] = 1024'd21693101031573173151090521344853949697344934683231677370127875593304798827373540208862719718917238447224184487773522158083724035443946751926179591770098000455183176168459492438279496041597318329963620152569412112724300330669844893606914188712636903832141453966638956722975733842221699126095303338466625498239;
            6'd23: xpb[19] = 1024'd5760965303354943558122054941690797491129009833505523960388435156867258500802909457899879085960157334446672499837205878735839149667596104119847737984693676712188228552993394275797167790099395655692394121997034502434810229761079192457458665060952747288126987772288401388096467915877871856765268513857072863932;
            6'd24: xpb[19] = 1024'd113895525259261455363952515943342078029611512109515054678780849785406613511541417616952109667660750531112309919358383033967018104732465790868676009215620393902883955507098513450945078730118678702731365699811896738509680979073210264272981711092498040010932424992054904083323730063462677604553923515873114713956;
            6'd25: xpb[19] = 1024'd97963389531043225770984049540178925823395587259788901269041409348969073184970786865989269034703669418334797931422066754619133218956115143062344155430216070159889007891632415288462750478620756028460139669239519128220190878164444563123526187440813883466917958797704348748444464137118850335223888691263562079649;
            6'd26: xpb[19] = 1024'd82031253802824996178015583137015773617179662410062747859301968912531532858400156115026428401746588305557285943485750475271248333179764495256012301644811746416894060276166317125980422227122833354188913638667141517930700777255678861974070663789129726922903492603353793413565198210775023065893853866654009445342;
            6'd27: xpb[19] = 1024'd66099118074606766585047116733852621410963737560336594449562528476093992531829525364063587768789507192779773955549434195923363447403413847449680447859407422673899112660700218963498093975624910679917687608094763907641210676346913160824615140137445570378889026409003238078685932284431195796563819042044456811035;
            6'd28: xpb[19] = 1024'd50166982346388536992078650330689469204747812710610441039823088039656452205258894613100747135832426080002261967613117916575478561627063199643348594074003098930904165045234120801015765724126988005646461577522386297351720575438147459675159616485761413834874560214652682743806666358087368527233784217434904176728;
            6'd29: xpb[19] = 1024'd34234846618170307399110183927526316998531887860884287630083647603218911878688263862137906502875344967224749979676801637227593675850712551837016740288598775187909217429768022638533437472629065331375235546950008687062230474529381758525704092834077257290860094020302127408927400431743541257903749392825351542421;
            6'd30: xpb[19] = 1024'd18302710889952077806141717524363164792315963011158134220344207166781371552117633111175065869918263854447237991740485357879708790074361904030684886503194451444914269814301924476051109221131142657104009516377631076772740373620616057376248569182393100746845627825951572074048134505399713988573714568215798908114;
            6'd31: xpb[19] = 1024'd2370575161733848213173251121200012586100038161431980810604766730343831225547002360212225236961182741669726003804169078531823904298011256224353032717790127701919322198835826313568780969633219982832783485805253466483250272711850356226793045530708944202831161631601016739168868579055886719243679743606246273807;
            6'd32: xpb[19] = 1024'd110505135117640360019003712122851293124582540437441511528997181358883186236285510519264455818661775938335363423325346233763002859362880942973181303948716844892615049152940945488716691909652503029871755063620115702558121022023981428042316091562254236925636598851367519434396130726640692467032334745622288123831;
            6'd33: xpb[19] = 1024'd94572999389422130426035245719688140918366615587715358119257740922445645909714879768301615185704694825557851435389029954415117973586530295166849450163312521149620101537474847326234363658154580355600529033047738092268630921115215726892860567910570080381622132657016964099516864800296865197702299921012735489524;
            6'd34: xpb[19] = 1024'd78640863661203900833066779316524988712150690737989204709518300486008105583144249017338774552747613712780339447452713675067233087810179647360517596377908197406625153922008749163752035406656657681329303002475360481979140820206450025743405044258885923837607666462666408764637598873953037928372265096403182855217;
            6'd35: xpb[19] = 1024'd62708727932985671240098312913361836505934765888263051299778860049570565256573618266375933919790532600002827459516397395719348202033828999554185742592503873663630206306542651001269707155158735007058076971902982871689650719297684324593949520607201767293593200268315853429758332947609210659042230271793630220910;
            6'd36: xpb[19] = 1024'd46776592204767441647129846510198684299718841038536897890039419613133024930002987515413093286833451487225315471580081116371463316257478351747853888807099549920635258691076552838787378903660812332786850941330605261400160618388918623444493996955517610749578734073965298094879067021265383389712195447184077586603;
            6'd37: xpb[19] = 1024'd30844456476549212054161380107035532093502916188810744480299979176695484603432356764450252653876370374447803483643764837023578430481127703941522035021695226177640311075610454676305050652162889658515624910758227651110670517480152922295038473303833454205564267879614742759999801094921556120382160622574524952296;
            6'd38: xpb[19] = 1024'd14912320748330982461192913703872379887286991339084591070560538740257944276861726013487412020919289261670291495707448557675693544704777056135190181236290902434645363460144356513822722400664966984244398880185850040821180416571387221145582949652149297661549801685264187425120535168577728851052125797964972317989;
            6'd39: xpb[19] = 1024'd123046880704237494267023374705523660425769493615094121788952953368797299287600234172539642602619882458335928915228625712906872499769646742884018452467217619625341090414249475688970633340684250031283370458000712276896051165883518292961105995683694590384355238905030690120347797316162534598840780799981014168013;
            6'd40: xpb[19] = 1024'd107114744976019264674054908302360508219553568765367968379213512932359758961029603421576801969662801345558416927292309433558987613993296095077686598681813295882346142798783377526488305089186327357012144427428334666606561064974752591811650472032010433840340772710680134785468531389818707329510745975371461533706;
            6'd41: xpb[19] = 1024'd91182609247801035081086441899197356013337643915641814969474072495922218634458972670613961336705720232780904939355993154211102728216945447271354744896408972139351195183317279364005976837688404682740918396855957056317070964065986890662194948380326277296326306516329579450589265463474880060180711150761908899399;
            6'd42: xpb[19] = 1024'd75250473519582805488117975496034203807121719065915661559734632059484678307888341919651120703748639120003392951419676874863217842440594799465022891111004648396356247567851181201523648586190482008469692366283579446027580863157221189512739424728642120752311840321979024115709999537131052790850676326152356265092;
            6'd43: xpb[19] = 1024'd59318337791364575895149509092871051600905794216189508149995191623047137981317711168688280070791558007225880963483360595515332956664244151658691037325600324653361299952385083039041320334692559334198466335711201835738090762248455488363283901076957964208297374127628468780830733610787225521520641501542803630785;
            6'd44: xpb[19] = 1024'd43386202063146346302181042689707899394689869366463354740255751186609597654747080417725439437834476894448368975547044316167448070887893503852359183540196000910366352336918984876558992083194636659927240305138824225448600661339689787213828377425273807664282907933277913445951467684443398252190606676933250996478;
            6'd45: xpb[19] = 1024'd27454066334928116709212576286544747188473944516737201330516310750172057328176449666762598804877395781670856987610728036819563185111542856046027329754791677167371404721452886714076663831696713985656014274566446615159110560430924086064372853773589651120268441738927358111072201758099570982860571852323698362171;
            6'd46: xpb[19] = 1024'd11521930606709887116244109883381594982258019667011047920776870313734517001605818915799758171920314668893344999674411757471678299335192208239695475969387353424376457105986788551594335580198791311384788243994069004869620459522158384914917330121905494576253975544576802776192935831755743713530537027714145727864;
            6'd47: xpb[19] = 1024'd119656490562616398922074570885032875520740521943020578639169284942273872012344327074851988753620907865558982419195588912702857254400061894988523747200314070615072184060091907726742246520218074358423759821808931240944491208834289456730440376153450787299059412764343305471420197979340549461319192029730187577888;
            6'd48: xpb[19] = 1024'd103724354834398169329106104481869723314524597093294425229429844505836331685773696323889148120663826752781470431259272633354972368623711247182191893414909746872077236444625809564259918268720151684152533791236553630655001107925523755580984852501766630755044946569992750136540932052996722191989157205120634943581;
            6'd49: xpb[19] = 1024'd87792219106179939736137638078706571108308672243568271819690404069398791359203065572926307487706745640003958443322956354007087482847360599375860039629505423129082288829159711401777590017222229009881307760664176020365511007016758054431529328850082474211030480375642194801661666126652894922659122380511082309274;
            6'd50: xpb[19] = 1024'd71860083377961710143169171675543418902092747393842118409950963632961251032632434821963466854749664527226446455386640074659202597071009951569528185844101099386087341213693613239295261765724306335610081730091798410076020906107992353282073805198398317667016014181291639466782400200309067653329087555901529674967;
            6'd51: xpb[19] = 1024'd55927947649743480550200705272380266695876822544115965000211523196523710706061804071000626221792583414448934467450323795311317711294659303763196332058696775643092393598227515076812933514226383661338855699519420799786530805199226652132618281546714161123001547986941084131903134273965240383999052731291977040660;
            6'd52: xpb[19] = 1024'd39995811921525250957232238869217114489660897694389811590472082760086170379491173320037785588835502301671422479514007515963432825518308655956864478273292451900097445982761416914330605262728460987067629668947043189497040704290460950983162757895030004578987081792590528797023868347621413114669017906682424406353;
            6'd53: xpb[19] = 1024'd24063676193307021364263772466053962283444972844663658180732642323648630052920542569074944955878421188893910491577691236615547939741958008150532624487888128157102498367295318751848277011230538312796403638374665579207550603381695249833707234243345848034972615598239973462144602421277585845338983082072871772046;
            6'd54: xpb[19] = 1024'd8131540465088791771295306062890810077229047994937504770993201887211089726349911818112104322921340076116398503641374957267663053965607360344200770702483804414107550751829220589365948759732615638525177607802287968918060502472929548684251710591661691490958149403889418127265336494933758576008948257463319137739;
            6'd55: xpb[19] = 1024'd116266100420995303577125767064542090615711550270947035489385616515750444737088419977164334904621933272782035923162552112498842009030477047093029041933410521604803277705934339764513859699751898685564149185617150204992931251785060620499774756623206984213763586623655920822492598642518564323797603259479360987763;
            6'd56: xpb[19] = 1024'd100333964692777073984157300661378938409495625421220882079646176079312904410517789226201494271664852160004523935226235833150957123254126399286697188148006197861808330090468241602031531448253976011292923155044772594703441150876294919350319232971522827669749120429305365487613332716174737054467568434869808353456;
            6'd57: xpb[19] = 1024'd84401828964558844391188834258215786203279700571494728669906735642875364083947158475238653638707771047227011947289919553803072237477775751480365334362601874118813382475002143439549203196756053337021697124472394984413951049967529218200863709319838671125734654234954810152734066789830909785137533610260255719149;
            6'd58: xpb[19] = 1024'd68469693236340614798220367855052633997063775721768575260167295206437823757376527724275813005750689934449499959353603274455187351701425103674033480577197550375818434859536045277066874945258130662750471093900017374124460949058763517051408185668154514581720188040604254817854800863487082515807498785650703084842;
            6'd59: xpb[19] = 1024'd52537557508122385205251901451889481790847850872042421850427854770000283430805896973312972372793608821671987971417286995107302465925074455867701626791793226632823487244069947114584546693760207988479245063327639763834970848149997815901952662016470358037705721846253699482975534937143255246477463961041150450535;
            6'd60: xpb[19] = 1024'd36605421779904155612283435048726329584631926022316268440688414333562743104235266222350131739836527708894475983480970715759417580148723808061369773006388902889828539628603848952102218442262285314208019032755262153545480747241232114752497138364786201493691255651903144148096269010799427977147429136431597816228;
            6'd61: xpb[19] = 1024'd20673286051685926019314968645563177378416001172590115030948973897125202777664635471387291106879446596116963995544654436411532694372373160255037919220984579146833592013137750789619890190764362639936793002182884543255990646332466413603041614713102044949676789457552588813217003084455600707817394311822045181921;
            6'd62: xpb[19] = 1024'd4741150323467696426346502242400025172200076322863961621209533460687662451094004720424450473922365483339452007608338157063647808596022512448706065435580255403838644397671652627137561939266439965665566971610506932966500545423700712453586091061417888405662323263202033478337737158111773438487359487212492547614;
            6'd63: xpb[19] = 1024'd112875710279374208232176963244051305710682578598873492339601948089227017461832512879476681055622958680005089427129515312294826763660892199197534336666506972594534371351776771802285472879285723012704538549425369169041371294735831784269109137092963181128467760482968536173564999305696579186276014489228534397638;
        endcase
    end

    always_comb begin
        case(flag[6][16:12])
            5'd0: xpb[20] = 1024'd0;
            5'd1: xpb[20] = 1024'd96943574551155978639208496840888153504466653749147338929862507652789477135261882128513840422665877567227577439193199032946941877884541551391202482881102648851539423736310673639803144627787800338433312518852991558751881193827066083119653613441279024584453294288617980838685733379352751916945979664618981763331;
            5'd2: xpb[20] = 1024'd69820453418187215879618066276961874264234880372558993731593160240602058933214625347012609630674080825012005470928904631314819914927862768227244840745874256769388172903050129941976050064058394955556427429318743271139401537433235393274328657199328599902086685163118903647264938684776870816773269502612369042331;
            5'd3: xpb[20] = 1024'd42697332285218453120027635713035595024003106995970648533323812828414640731167368565511378838682284082796433502664610229682697951971183985063287198610645864687236922069789586244148955500328989572679542339784494983526921881039404703429003700957378175219720076037619826455844143990200989716600559340605756321331;
            5'd4: xpb[20] = 1024'd15574211152249690360437205149109315783771333619382303335054465416227222529120111784010148046690487340580861534400315828050575989014505201899329556475417472605085671236529042546321860936599584189802657250250246695914442224645574013583678744715427750537353466912120749264423349295625108616427849178599143600331;
            5'd5: xpb[20] = 1024'd112517785703405668999645701989997469288237987368529642264916973069016699664381993912523988469356364907808438973593514860997517866899046753290532039356520121456625094972839716186125005564387384528235969769103238254666323418472640096703332358156706775121806761200738730103109082674977860533373828843218125363662;
            5'd6: xpb[20] = 1024'd85394664570436906240055271426071190048006213991941297066647625656829281462334737131022757677364568165592867005329220459365395903942367970126574397221291729374473844139579172488297911000657979145359084679568989967053843762078809406858007401914756350439440152075239652911688287980401979433201118681211512642662;
            5'd7: xpb[20] = 1024'd58271543437468143480464840862144910807774440615352951868378278244641863260287480349521526885372771423377295037064926057733273940985689186962616755086063337292322593306318628790470816436928573762482199590034741679441364105684978717012682445672805925757073542949740575720267493285826098333028408519204899921662;
            5'd8: xpb[20] = 1024'd31148422304499380720874410298218631567542667238764606670108930832454445058240223568020296093380974681161723068800631656101151978029010403798659112950834945210171342473058085092643721873199168379605314500500493391828884449291148027167357489430855501074706933824241498528846698591250217232855698357198287200662;
            5'd9: xpb[20] = 1024'd4025301171530617961283979734292352327310893862176261471839583420267026856192966786519065301389177938946151100536337254469030015072331620634701470815606553128020091639797541394816627309469762996728429410966245104216404792897317337322032533188905076392340324698742421337425903896674336132682988195191674479662;
            5'd10: xpb[20] = 1024'd100968875722686596600492476575180505831777547611323600401702091073056503991454848915032905724055055506173728539729536287415971892956873172025903953696709201979559515376108215034619771937257563335161741929819236662968285986724383420441686146630184100976793618987360402176111637276027088049628967859810656242993;
            5'd11: xpb[20] = 1024'd73845754589717833840902046011254226591545774234735255203432743660869085789407592133531674932063258763958156571465241885783849930000194388861946311561480809897408264542847671336792677373528157952284856840284988375355806330330552730596361190388233676294427009861861324984690842581451206949456257697804043521993;
            5'd12: xpb[20] = 1024'd46722633456749071081311615447327947351314000858146910005163396248681667587360335352030444140071462021742584603200947484151727967043515605697988669426252417815257013709587127638965582809798752569407971750750740087743326673936722040751036234146283251612060400736362247793270047886875325849283547535797430800993;
            5'd13: xpb[20] = 1024'd19599512323780308321721184883401668111082227481558564806894048836494249385313078570529213348079665279527012634936653082519606004086836822534031027291024025733105762876326583941138488246069347186531086661216491800130847017542891350905711277904332826929693791610863170601849253192299444749110837373790818079993;
            5'd14: xpb[20] = 1024'd116543086874936286960929681724289821615548881230705903736756556489283726520574960699043053770745542846754590074129852115466547881971378373925233510172126674584645186612637257580941632873857147524964399180069483358882728211369957434025364891345611851514147085899481151440534986571652196666056817038409799843324;
            5'd15: xpb[20] = 1024'd89419965741967524201339251160363542375317107854117558538487209077096308318527703917541822978753746104539018105865557713834425919014699590761275868036898282502493935779376713883114538310127742142087514090535235071270248554976126744180039935103661426831780476773982074249114191877076315565884106876403187122324;
            5'd16: xpb[20] = 1024'd62296844608998761441748820596437263135085334477529213340217861664908890116480447136040592186761949362323446137601263312202303956058020807597318225901669890420342684946116170185287443746398336759210629001000986783657768898582296054334714978861711002149413867648482997057693397182500434465711396714396574401324;
            5'd17: xpb[20] = 1024'd35173723476029998682158390032510983894853561100940868141948514252721471914433190354539361394770152620107874169336968910570181993101342024433360583766441498338191434112855626487460349182668931376333743911466738496045289242188465364489390022619760577467047258522983919866272602487924553365538686552389961680324;
            5'd18: xpb[20] = 1024'd8050602343061235922567959468584704654621787724352522943679166840534053712385933573038130602778355877892302201072674508938060030144663241269402941631213106256040183279595082789633254618939525993456858821932490208432809585794634674644065066377810152784680649397484842674851807793348672265365976390383348959324;
            5'd19: xpb[20] = 1024'd104994176894217214561776456309472858159088441473499861873541674493323530847647815701551971025444233445119879640265873541885001908029204792660605424512315755107579607015905756429436399246727326331890171340785481767184690779621700757763718679819089177369133943686102823513537541172701424182311956055002330722655;
            5'd20: xpb[20] = 1024'd77871055761248451802186025745546578918856668096911516675272327081136112645600558920050740233452436702904307672001579140252879945072526009496647782377087363025428356182645212731609304682997920949013286251251233479572211123227870067918393723577138752686767334560603746322116746478125543082139245892995718001655;
            5'd21: xpb[20] = 1024'd50747934628279689042595595181620299678624894720323171477002979668948694443553302138549509441460639960688735703737284738620757982115847226332690140241858970943277105349384669033782210119268515566136401161716985191959731466834039378073068767335188328004400725435104669130695951783549661981966535730989105280655;
            5'd22: xpb[20] = 1024'd23624813495310926283005164617694020438393121343734826278733632256761276241506045357048278649468843218473163735472990336988636019159168443168732498106630578861125854516124125335955115555539110183259516072182736904347251810440208688227743811093237903322034116309605591939275157088973780881793825568982492559655;
            5'd23: xpb[20] = 1024'd120568388046466904922213661458582173942859775092882165208596139909550753376767927485562119072134720785700741174666189369935577897043709994559934980987733227712665278252434798975758260183326910521692828591035728463099133004267274771347397424534516927906487410598223572777960890468326532798739805233601474322986;
            5'd24: xpb[20] = 1024'd93445266913498142162623230894655894702628001716293820010326792497363335174720670704060888280142924043485169206401894968303455934087031211395977338852504835630514027419174255277931165619597505138815943501501480175486653347873444081502072468292566503224120801472724495586540095773750651698567095071594861601986;
            5'd25: xpb[20] = 1024'd66322145780529379403032800330729615462396228339705474812057445085175916972673413922559657488151127301269597238137600566671333971130352428232019696717276443548362776585913711580104071055868099755939058411967231887874173691479613391656747512050616078541754192347225418395119301079174770598394384909588248880986;
            5'd26: xpb[20] = 1024'd39199024647560616643442369766803336222164454963117129613788097672988498770626157141058426696159330559054025269873306165039212008173673645068062054582048051466211525752653167882276976492138694373062173322432983600261694035085782701811422555808665653859387583221726341203698506384598889498221674747581636159986;
            5'd27: xpb[20] = 1024'd12075903514591853883851939202877056981932681586528784415518750260801080568578900359557195904167533816838453301609011763407090045216994861904104412446819659384060274919392624184449881928409288990185288232898735312649214378691952011966097599566715229177020974096227264012277711690023008398048964585575023438986;
            5'd28: xpb[20] = 1024'd109019478065747832523060436043765210486399335335676123345381257913590557703840782488071036326833411384066030740802210796354031923101536413295306895327922308235599698655703297824253026556197089328618600751751726871401095572519018095085751213007994253761474268384845244850963445069375760314994944250194005202317;
            5'd29: xpb[20] = 1024'd81896356932779069763470005479838931246167561959087778147111910501403139501793525706569805534841614641850458772537916394721909960144857630131349253192693916153448447822442754126425931992467683945741715662217478583788615916125187405240426256766043829079107659259346167659542650374799879214822234088187392481317;
            5'd30: xpb[20] = 1024'd54773235799810307003879574915912652005935788582499432948842563089215721299746268925068574742849817899634886804273621993089787997188178846967391611057465524071297196989182210428598837428738278562864830572683230296176136259731356715395101300524093404396741050133847090468121855680223998114649523926180779760317;
            5'd31: xpb[20] = 1024'd27650114666841544244289144351986372765704015205911087750573215677028303097699012143567343950858021157419314836009327591457666034231500063803433968922237131989145946155921666730771742865008873179987945483148982008563656603337526025549776344282142979714374441008348013276701060985648117014476813764174167039317;
        endcase
    end

    always_comb begin
        case(flag[7][5:0])
            6'd0: xpb[21] = 1024'd0;
            6'd1: xpb[21] = 1024'd62296844608998761441748820596437263135085334477529213340217861664908890116480447136040592186761949362323446137601263312202303956058020807597318225901669890420342684946116170185287443746398336759210629001000986783657768898582296054334714978861711002149413867648482997057693397182500434465711396714396574401324;
            6'd2: xpb[21] = 1024'd526993533872781484698713788060093525472241829322742552303868264840884895651755362066113158866224415203742867745033189825544071274821280639476326787008739906994695322661123032944648301279467797111060393614733720951176946943695335704451388040192555032007831882848936085280266291072235914304103602167554318317;
            6'd3: xpb[21] = 1024'd62823838142871542926447534384497356660557576306851955892521729929749775012132202498106705345628173777527189005346296502027848027332842088236794552688678630327337380268777293218232092047677804556321689394615720504608945845525991390039166366901903557181421699531331933142973663473572670380015500316564128719641;
            6'd4: xpb[21] = 1024'd1053987067745562969397427576120187050944483658645485104607736529681769791303510724132226317732448830407485735490066379651088142549642561278952653574017479813989390645322246065889296602558935594222120787229467441902353893887390671408902776080385110064015663765697872170560532582144471828608207204335108636634;
            6'd5: xpb[21] = 1024'd63350831676744324411146248172557450186029818136174698444825598194590659907783957860172818504494398192730931873091329691853392098607663368876270879475687370234332075591438416251176740348957272353432749788230454225560122792469686725743617754942096112213429531414180869228253929764644906294319603918731683037958;
            6'd6: xpb[21] = 1024'd1580980601618344454096141364180280576416725487968227656911604794522654686955266086198339476598673245611228603235099569476632213824463841918428980361026219720984085967983369098833944903838403391333181180844201162853530840831086007113354164120577665096023495648546808255840798873216707742912310806502662954951;
            6'd7: xpb[21] = 1024'd63877825210617105895844961960617543711502059965497440997129466459431544803435713222238931663360622607934674740836362881678936169882484649515747206262696110141326770914099539284121388650236740150543810181845187946511299739413382061448069142982288667245437363297029805313534196055717142208623707520899237356275;
            6'd8: xpb[21] = 1024'd2107974135491125938794855152240374101888967317290970209215473059363539582607021448264452635464897660814971470980132759302176285099285122557905307148034959627978781290644492131778593205117871188444241574458934883804707787774781342817805552160770220128031327531395744341121065164288943657216414408670217273268;
            6'd9: xpb[21] = 1024'd64404818744489887380543675748677637236974301794820183549433334724272429699087468584305044822226847023138417608581396071504480241157305930155223533049704850048321466236760662317066036951516207947654870575459921667462476686357077397152520531022481222277445195179878741398814462346789378122927811123066791674592;
            6'd10: xpb[21] = 1024'd2634967669363907423493568940300467627361209146613712761519341324204424478258776810330565794331122076018714338725165949127720356374106403197381633935043699534973476613305615164723241506397338985555301968073668604755884734718476678522256940200962775160039159414244680426401331455361179571520518010837771591585;
            6'd11: xpb[21] = 1024'd64931812278362668865242389536737730762446543624142926101737202989113314594739223946371157981093071438342160476326429261330024312432127210794699859836713589955316161559421785350010685252795675744765930969074655388413653633300772732856971919062673777309453027062727677484094728637861614037231914725234345992909;
            6'd12: xpb[21] = 1024'd3161961203236688908192282728360561152833450975936455313823209589045309373910532172396678953197346491222457206470199138953264427648927683836857960722052439441968171935966738197667889807676806782666362361688402325707061681662172014226708328241155330192046991297093616511681597746433415485824621613005325909902;
            6'd13: xpb[21] = 1024'd65458805812235450349941103324797824287918785453465668654041071253954199490390979308437271139959295853545903344071462451155568383706948491434176186623722329862310856882082908382955333554075143541876991362689389109364830580244468068561423307102866332341460858945576613569374994928933849951536018327401900311226;
            6'd14: xpb[21] = 1024'd3688954737109470392890996516420654678305692805259197866127077853886194269562287534462792112063570906426200074215232328778808498923748964476334287509061179348962867258627861230612538108956274579777422755303136046658238628605867349931159716281347885224054823179942552596961864037505651400128725215172880228219;
            6'd15: xpb[21] = 1024'd65985799346108231834639817112857917813391027282788411206344939518795084386042734670503384298825520268749646211816495640981112454981769772073652513410731069769305552204744031415899981855354611338988051756304122830316007527188163404265874695143058887373468690828425549654655261220006085865840121929569454629543;
            6'd16: xpb[21] = 1024'd4215948270982251877589710304480748203777934634581940418430946118727079165214042896528905270929795321629942941960265518604352570198570245115810614296069919255957562581288984263557186410235742376888483148917869767609415575549562685635611104321540440256062655062791488682242130328577887314432828817340434546536;
            6'd17: xpb[21] = 1024'd66512792879981013319338530900918011338863269112111153758648807783635969281694490032569497457691744683953389079561528830806656526256591052713128840197739809676300247527405154448844630156634079136099112149918856551267184474131858739970326083183251442405476522711274485739935527511078321780144225531737008947860;
            6'd18: xpb[21] = 1024'd4742941804855033362288424092540841729250176463904682970734814383567964060865798258595018429796019736833685809705298708429896641473391525755286941083078659162952257903950107296501834711515210173999543542532603488560592522493258021340062492361732995288070486945640424767522396619650123228736932419507988864853;
            6'd19: xpb[21] = 1024'd67039786413853794804037244688978104864335510941433896310952676048476854177346245394635610616557969099157131947306562020632200597531412333352605166984748549583294942850066277481789278457913546933210172543533590272218361421075554075674777471223443997437484354594123421825215793802150557694448329133904563266177;
            6'd20: xpb[21] = 1024'd5269935338727814846987137880600935254722418293227425523038682648408848956517553620661131588662244152037428677450331898255440712748212806394763267870087399069946953226611230329446483012794677971110603936147337209511769469436953357044513880401925550320078318828489360852802662910722359143041036021675543183170;
            6'd21: xpb[21] = 1024'd67566779947726576288735958477038198389807752770756638863256544313317739072998000756701723775424193514360874815051595210457744668806233613992081493771757289490289638172727400514733926759193014730321232937148323993169538368019249411379228859263636552469492186476972357910496060093222793608752432736072117584494;
            6'd22: xpb[21] = 1024'd5796928872600596331685851668661028780194660122550168075342550913249733852169308982727244747528468567241171545195365088080984784023034087034239594657096138976941648549272353362391131314074145768221664329762070930462946416380648692748965268442118105352086150711338296938082929201794595057345139623843097501487;
            6'd23: xpb[21] = 1024'd68093773481599357773434672265098291915279994600079381415560412578158623968649756118767836934290417929564617682796628400283288740081054894631557820558766029397284333495388523547678575060472482527432293330763057714120715314962944747083680247303829107501500018359821293995776326384295029523056536338239671902811;
            6'd24: xpb[21] = 1024'd6323922406473377816384565456721122305666901951872910627646419178090618747821064344793357906394692982444914412940398277906528855297855367673715921444104878883936343871933476395335779615353613565332724723376804651414123363324344028453416656482310660384093982594187233023363195492866830971649243226010651819804;
            6'd25: xpb[21] = 1024'd68620767015472139258133386053158385440752236429402123967864280842999508864301511480833950093156642344768360550541661590108832811355876175271034147345774769304279028818049646580623223361751950324543353724377791435071892261906640082788131635344021662533507850242670230081056592675367265437360639940407226221128;
            6'd26: xpb[21] = 1024'd6850915940346159301083279244781215831139143781195653179950287442931503643472819706859471065260917397648657280685431467732072926572676648313192248231113618790931039194594599428280427916633081362443785116991538372365300310268039364157868044522503215416101814477036169108643461783939066885953346828178206138121;
            6'd27: xpb[21] = 1024'd69147760549344920742832099841218478966224478258724866520168149107840393759953266842900063252022866759972103418286694779934376882630697455910510474132783509211273724140710769613567871663031418121654414117992525156023069208850335418492583023384214217565515682125519166166336858966439501351664743542574780539445;
            6'd28: xpb[21] = 1024'd7377909474218940785781993032841309356611385610518395732254155707772388539124575068925584224127141812852400148430464657557616997847497928952668575018122358697925734517255722461225076217912549159554845510606272093316477257211734699862319432562695770448109646359885105193923728075011302800257450430345760456438;
            6'd29: xpb[21] = 1024'd69674754083217702227530813629278572491696720088047609072472017372681278655605022204966176410889091175175846286031727969759920953905518736549986800919792249118268419463371892646512519964310885918765474511607258876974246155794030754197034411424406772597523514008368102251617125257511737265968847144742334857762;
            6'd30: xpb[21] = 1024'd7904903008091722270480706820901402882083627439841138284558023972613273434776330430991697382993366228056143016175497847383161069122319209592144901805131098604920429839916845494169724519192016956665905904221005814267654204155430035566770820602888325480117478242734041279203994366083538714561554032513314774755;
            6'd31: xpb[21] = 1024'd70201747617090483712229527417338666017168961917370351624775885637522163551256777567032289569755315590379589153776761159585465025180340017189463127706800989025263114786033015679457168265590353715876534905221992597925423102737726089901485799464599327629531345891217038336897391548583973180272950746909889176079;
            6'd32: xpb[21] = 1024'd8431896541964503755179420608961496407555869269163880836861892237454158330428085793057810541859590643259885883920531037208705140397140490231621228592139838511915125162577968527114372820471484753776966297835739535218831151099125371271222208643080880512125310125582977364484260657155774628865657634680869093072;
            6'd33: xpb[21] = 1024'd70728741150963265196928241205398759542641203746693094177079753902363048446908532929098402728621540005583332021521794349411009096455161297828939454493809728932257810108694138712401816566869821512987595298836726318876600049681421425605937187504791882661539177774065974422177657839656209094577054349077443494396;
            6'd34: xpb[21] = 1024'd8958890075837285239878134397021589933028111098486623389165760502295043226079841155123923700725815058463628751665564227034249211671961770871097555379148578418909820485239091560059021121750952550888026691450473256170008098042820706975673596683273435544133142008431913449764526948228010543169761236848423411389;
            6'd35: xpb[21] = 1024'd71255734684836046681626954993458853068113445576015836729383622167203933342560288291164515887487764420787074889266827539236553167729982578468415781280818468839252505431355261745346464868149289310098655692451460039827776996625116761310388575544984437693547009656914910507457924130728445008881157951244997812713;
            6'd36: xpb[21] = 1024'd9485883609710066724576848185081683458500352927809365941469628767135928121731596517190036859592039473667371619410597416859793282946783051510573882166157318325904515807900214593003669423030420347999087085065206977121185044986516042680124984723465990576140973891280849535044793239300246457473864839015977729706;
            6'd37: xpb[21] = 1024'd71782728218708828166325668781518946593585687405338579281687490432044818238212043653230629046353988835990817757011860729062097239004803859107892108067827208746247200754016384778291113169428757107209716086066193760778953943568812097014839963585176992725554841539763846592738190421800680923185261553412552131030;
            6'd38: xpb[21] = 1024'd10012877143582848209275561973141776983972594757132108493773497031976813017383351879256150018458263888871114487155630606685337354221604332150050208953166058232899211130561337625948317724309888145110147478679940698072361991930211378384576372763658545608148805774129785620325059530372482371777968441183532048023;
            6'd39: xpb[21] = 1024'd72309721752581609651024382569579040119057929234661321833991358696885703133863799015296742205220213251194560624756893918887641310279625139747368434854835948653241896076677507811235761470708224904320776479680927481730130890512507432719291351625369547757562673422612782678018456712872916837489365155580106449347;
            6'd40: xpb[21] = 1024'd10539870677455629693974275761201870509444836586454851046077365296817697913035107241322263177324488304074857354900663796510881425496425612789526535740174798139893906453222460658892966025589355942221207872294674419023538938873906714089027760803851100640156637656978721705605325821444718286082072043351086366340;
            6'd41: xpb[21] = 1024'd72836715286454391135723096357639133644530171063984064386295226961726588029515554377362855364086437666398303492501927108713185381554446420386844761641844688560236591399338630844180409771987692701431836873295661202681307837456202768423742739665562102789570505305461718763298723003945152751793468757747660767664;
            6'd42: xpb[21] = 1024'd11066864211328411178672989549261964034917078415777593598381233561658582808686862603388376336190712719278600222645696986336425496771246893429002862527183538046888601775883583691837614326868823739332268265909408139974715885817602049793479148844043655672164469539827657790885592112516954200386175645518640684657;
            6'd43: xpb[21] = 1024'd73363708820327172620421810145699227170002412893306806938599095226567472925167309739428968522952662081602046360246960298538729452829267701026321088428853428467231286721999753877125058073267160498542897266910394923632484784399898104128194127705754657821578337188310654848578989295017388666097572359915215085981;
            6'd44: xpb[21] = 1024'd11593857745201192663371703337322057560389320245100336150685101826499467704338617965454489495056937134482343090390730176161969568046068174068479189314192277953883297098544706724782262628148291536443328659524141860925892832761297385497930536884236210704172301422676593876165858403589190114690279247686195002974;
            6'd45: xpb[21] = 1024'd73890702354199954105120523933759320695474654722629549490902963491408357820819065101495081681818886496805789227991993488364273524104088981665797415215862168374225982044660876910069706374546628295653957660525128644583661731343593439832645515745947212853586169071159590933859255586089624580401675962082769404298;
            6'd46: xpb[21] = 1024'd12120851279073974148070417125382151085861562074423078702988970091340352599990373327520602653923161549686085958135763365987513639320889454707955516101201017860877992421205829757726910929427759333554389053138875581877069779704992721202381924924428765736180133305525529961446124694661426028994382849853749321291;
            6'd47: xpb[21] = 1024'd74417695888072735589819237721819414220946896551952292043206831756249242716470820463561194840685110912009532095737026678189817595378910262305273742002870908281220677367321999943014354675826096092765018054139862365534838678287288775537096903786139767885594000954008527019139521877161860494705779564250323722615;
            6'd48: xpb[21] = 1024'd12647844812946755632769130913442244611333803903745821255292838356181237495642128689586715812789385964889828825880796555813057710595710735347431842888209757767872687743866952790671559230707227130665449446753609302828246726648688056906833312964621320768187965188374466046726390985733661943298486452021303639608;
            6'd49: xpb[21] = 1024'd74944689421945517074517951509879507746419138381275034595510700021090127612122575825627307999551335327213274963482059868015361666653731542944750068789879648188215372689983122975959002977105563889876078447754596086486015625230984111241548291826332322917601832836857463104419788168234096409009883166417878040932;
            6'd50: xpb[21] = 1024'd13174838346819537117467844701502338136806045733068563807596706621022122391293884051652828971655610380093571693625829745638601781870532015986908169675218497674867383066528075823616207531986694927776509840368343023779423673592383392611284701004813875800195797071223402132006657276805897857602590054188857957925;
            6'd51: xpb[21] = 1024'd75471682955818298559216665297939601271891380210597777147814568285931012507774331187693421158417559742417017831227093057840905737928552823584226395576888388095210068012644246008903651278385031686987138841369329807437192572174679446945999679866524877949609664719706399189700054459306332323313986768585432359249;
            6'd52: xpb[21] = 1024'd13701831880692318602166558489562431662278287562391306359900574885863007286945639413718942130521834795297314561370862935464145853145353296626384496462227237581862078389189198856560855833266162724887570233983076744730600620536078728315736089045006430832203628954072338217286923567878133771906693656356412276242;
            6'd53: xpb[21] = 1024'd75998676489691080043915379085999694797363622039920519700118436550771897403426086549759534317283784157620760698972126247666449809203374104223702722363897128002204763335305369041848299579664499484098199234984063528388369519118374782650451067906717432981617496602555335274980320750378568237618090370752986677566;
            6'd54: xpb[21] = 1024'd14228825414565100086865272277622525187750529391714048912204443150703892182597394775785055289388059210501057429115896125289689924420174577265860823249235977488856773711850321889505504134545630521998630627597810465681777567479774064020187477085198985864211460836921274302567189858950369686210797258523966594559;
            6'd55: xpb[21] = 1024'd76525670023563861528614092874059788322835863869243262252422304815612782299077841911825647476150008572824503566717159437491993880478195384863179049150905867909199458657966492074792947880943967281209259628598797249339546466062070118354902455946909988013625328485404271360260587041450804151922193972920540995883;
            6'd56: xpb[21] = 1024'd14755818948437881571563986065682618713222771221036791464508311415544777078249150137851168448254283625704800296860929315115233995694995857905337150036244717395851469034511444922450152435825098319109691021212544186632954514423469399724638865125391540896219292719770210387847456150022605600514900860691520912876;
            6'd57: xpb[21] = 1024'd77052663557436643013312806662119881848308105698566004804726173080453667194729597273891760635016232988028246434462192627317537951753016665502655375937914607816194153980627615107737596182223435078320320022213530970290723413005765454059353843987102543045633160368253207445540853332523040066226297575088095314200;
            6'd58: xpb[21] = 1024'd15282812482310663056262699853742712238695013050359534016812179680385661973900905499917281607120508040908543164605962504940778066969817138544813476823253457302846164357172567955394800737104566116220751414827277907584131461367164735429090253165584095928227124602619146473127722441094841514819004462859075231193;
            6'd59: xpb[21] = 1024'd77579657091309424498011520450179975373780347527888747357030041345294552090381352635957873793882457403231989302207225817143082023027837946142131702724923347723188849303288738140682244483502902875431380415828264691241900359949460789763805232027295098077640992251102143530821119623595275980530401177255649632517;
            6'd60: xpb[21] = 1024'd15809806016183444540961413641802805764167254879682276569116047945226546869552660861983394765986732456112286032350995694766322138244638419184289803610262197209840859679833690988339449038384033913331811808442011628535308408310860071133541641205776650960234956485468082558407988732167077429123108065026629549510;
            6'd61: xpb[21] = 1024'd78106650625182205982710234238240068899252589357211489909333909610135436986033107998023986952748681818435732169952259006968626094302659226781608029511932087630183544625949861173626892784782370672542440809442998412193077306893156125468256620067487653109648824133951079616101385914667511894834504779423203950834;
            6'd62: xpb[21] = 1024'd16336799550056226025660127429862899289639496709005019121419916210067431765204416224049507924852956871316028900096028884591866209519459699823766130397270937116835555002494814021284097339663501710442872202056745349486485355254555406837993029245969205992242788368317018643688255023239313343427211667194183867827;
            6'd63: xpb[21] = 1024'd78633644159054987467408948026300162424724831186534232461637777874976321881684863360090100111614906233639475037697292196794170165577480507421084356298940827537178239948610984206571541086061838469653501203057732133144254253836851461172708008107680208141656656016800015701381652205739747809138608381590758269151;
        endcase
    end

    always_comb begin
        case(flag[7][11:6])
            6'd0: xpb[22] = 1024'd0;
            6'd1: xpb[22] = 1024'd16863793083929007510358841217922992815111738538327761673723784474908316660856171586115621083719181286519771767841062074417410280794280980463242457184279677023830250325155937054228745640942969507553932595671479070437662302198250742542444417286161761024250620251165954728968521314311549257731315269361738186144;
            6'd2: xpb[22] = 1024'd33727586167858015020717682435845985630223477076655523347447568949816633321712343172231242167438362573039543535682124148834820561588561960926484914368559354047660500650311874108457491281885939015107865191342958140875324604396501485084888834572323522048501240502331909457937042628623098515462630538723476372288;
            6'd3: xpb[22] = 1024'd50591379251787022531076523653768978445335215614983285021171353424724949982568514758346863251157543859559315303523186223252230842382842941389727371552839031071490750975467811162686236922828908522661797787014437211312986906594752227627333251858485283072751860753497864186905563942934647773193945808085214558432;
            6'd4: xpb[22] = 1024'd67455172335716030041435364871691971260446954153311046694895137899633266643424686344462484334876725146079087071364248297669641123177123921852969828737118708095321001300623748216914982563771878030215730382685916281750649208793002970169777669144647044097002481004663818915874085257246197030925261077446952744576;
            6'd5: xpb[22] = 1024'd84318965419645037551794206089614964075558692691638808368618922374541583304280857930578105418595906432598858839205310372087051403971404902316212285921398385119151251625779685271143728204714847537769662978357395352188311510991253712712222086430808805121253101255829773644842606571557746288656576346808690930720;
            6'd6: xpb[22] = 1024'd101182758503574045062153047307537956890670431229966570042342706849449899965137029516693726502315087719118630607046372446504461684765685882779454743105678062142981501950935622325372473845657817045323595574028874422625973813189504455254666503716970566145503721506995728373811127885869295546387891616170429116864;
            6'd7: xpb[22] = 1024'd118046551587503052572511888525460949705782169768294331716066491324358216625993201102809347586034269005638402374887434520921871965559966863242697200289957739166811752276091559379601219486600786552877528169700353493063636115387755197797110921003132327169754341758161683102779649200180844804119206885532167303008;
            6'd8: xpb[22] = 1024'd10843648987307318684071802338569509776195481180886409261658420734289637949540233778909897455095775982715024735271003160760218405513027509150779532457906375256951328031676279096199725936026550339121263156984592717136937567365109167374576768606064638927185058595210579801641642440563761044731832328268311004821;
            6'd9: xpb[22] = 1024'd27707442071236326194430643556492502591307219719214170935382205209197954610396405365025518538814957269234796503112065235177628686307308489614021989642186052280781578356832216150428471576969519846675195752656071787574599869563359909917021185892226399951435678846376534530610163754875310302463147597630049190965;
            6'd10: xpb[22] = 1024'd44571235155165333704789484774415495406418958257541932609105989684106271271252576951141139622534138555754568270953127309595038967101589470077264446826465729304611828681988153204657217217912489354229128348327550858012262171761610652459465603178388160975686299097542489259578685069186859560194462866991787377109;
            6'd11: xpb[22] = 1024'd61435028239094341215148325992338488221530696795869694282829774159014587932108748537256760706253319842274340038794189384012449247895870450540506904010745406328442079007144090258885962858855458861783060943999029928449924473959861395001910020464549921999936919348708443988547206383498408817925778136353525563253;
            6'd12: xpb[22] = 1024'd78298821323023348725507167210261481036642435334197455956553558633922904592964920123372381789972501128794111806635251458429859528690151431003749361195025083352272329332300027313114708499798428369336993539670508998887586776158112137544354437750711683024187539599874398717515727697809958075657093405715263749397;
            6'd13: xpb[22] = 1024'd95162614406952356235866008428184473851754173872525217630277343108831221253821091709488002873691682415313883574476313532847269809484432411466991818379304760376102579657455964367343454140741397876890926135341988069325249078356362880086798855036873444048438159851040353446484249012121507333388408675077001935541;
            6'd14: xpb[22] = 1024'd112026407490881363746224849646107466666865912410852979304001127583739537914677263295603623957410863701833655342317375607264680090278713391930234275563584437399932829982611901421572199781684367384444858731013467139762911380554613622629243272323035205072688780102206308175452770326433056591119723944438740121685;
            6'd15: xpb[22] = 1024'd4823504890685629857784763459216026737279223823445056849593056993670959238224295971704173826472370678910277702700944247103026530231774037838316607731533073490072405738196621138170706231110131170688593718297706363836212832531967592206709119925967516830119496939255204874314763566815972831732349387174883823498;
            6'd16: xpb[22] = 1024'd21687297974614637368143604677139019552390962361772818523316841468579275899080467557819794910191551965430049470542006321520436811026055018301559064915812750513902656063352558192399451872053100678242526313969185434273875134730218334749153537212129277854370117190421159603283284881127522089463664656536622009642;
            6'd17: xpb[22] = 1024'd38551091058543644878502445895062012367502700900100580197040625943487592559936639143935415993910733251949821238383068395937847091820335998764801522100092427537732906388508495246628197512996070185796458909640664504711537436928469077291597954498291038878620737441587114332251806195439071347194979925898360195786;
            6'd18: xpb[22] = 1024'd55414884142472652388861287112985005182614439438428341870764410418395909220792810730051037077629914538469593006224130470355257372614616979228043979284372104561563156713664432300856943153939039693350391505312143575149199739126719819834042371784452799902871357692753069061220327509750620604926295195260098381930;
            6'd19: xpb[22] = 1024'd72278677226401659899220128330907997997726177976756103544488194893304225881648982316166658161349095824989364774065192544772667653408897959691286436468651781585393407038820369355085688794882009200904324100983622645586862041324970562376486789070614560927121977943919023790188848824062169862657610464621836568074;
            6'd20: xpb[22] = 1024'd89142470310330667409578969548830990812837916515083865218211979368212542542505153902282279245068277111509136541906254619190077934203178940154528893652931458609223657363976306409314434435824978708458256696655101716024524343523221304918931206356776321951372598195084978519157370138373719120388925733983574754218;
            6'd21: xpb[22] = 1024'd106006263394259674919937810766753983627949655053411626891935763843120859203361325488397900328787458398028908309747316693607488214997459920617771350837211135633053907689132243463543180076767948216012189292326580786462186645721472047461375623642938082975623218446250933248125891452685268378120241003345312940362;
            6'd22: xpb[22] = 1024'd122870056478188682430296651984676976443061393591739388565659548318029175864217497074513521412506639684548680077588378768024898495791740901081013808021490812656884158014288180517771925717710917723566121887998059856899848947919722790003820040929099843999873838697416887977094412766996817635851556272707051126506;
            6'd23: xpb[22] = 1024'd15667153877992948541856565797785536513474705004331466111251477727960597187764529750614071281568146661625302437971947407863244935744801546989096140189439448747023733769872900234370432167136681509809856875282299080973150399897076759581285888532032155757304555534465784675956406007379733876464181715443194828319;
            6'd24: xpb[22] = 1024'd32530946961921956052215407015708529328586443542659227784975262202868913848620701336729692365287327948145074205813009482280655216539082527452338597373719125770853984095028837288599177808079651017363789470953778151410812702095327502123730305818193916781555175785631739404924927321691283134195496984804933014463;
            6'd25: xpb[22] = 1024'd49394740045850963562574248233631522143698182080986989458699046677777230509476872922845313449006509234664845973654071556698065497333363507915581054557998802794684234420184774342827923449022620524917722066625257221848475004293578244666174723104355677805805796036797694133893448636002832391926812254166671200607;
            6'd26: xpb[22] = 1024'd66258533129779971072933089451554514958809920619314751132422831152685547170333044508960934532725690521184617741495133631115475778127644488378823511742278479818514484745340711397056669089965590032471654662296736292286137306491828987208619140390517438830056416287963648862861969950314381649658127523528409386751;
            6'd27: xpb[22] = 1024'd83122326213708978583291930669477507773921659157642512806146615627593863831189216095076555616444871807704389509336195705532886058921925468842065968926558156842344735070496648451285414730908559540025587257968215362723799608690079729751063557676679199854307036539129603591830491264625930907389442792890147572895;
            6'd28: xpb[22] = 1024'd99986119297637986093650771887400500589033397695970274479870400102502180492045387681192176700164053094224161277177257779950296339716206449305308426110837833866174985395652585505514160371851529047579519853639694433161461910888330472293507974962840960878557656790295558320799012578937480165120758062251885759039;
            6'd29: xpb[22] = 1024'd116849912381566993604009613105323493404145136234298036153594184577410497152901559267307797783883234380743933045018319854367706620510487429768550883295117510890005235720808522559742906012794498555133452449311173503599124213086581214835952392249002721902808277041461513049767533893249029422852073331613623945183;
            6'd30: xpb[22] = 1024'd9647009781371259715569526918432053474558447646890113699186113987341918476448591943408347652944741357820555405401888494206053060463548075676633215463066146980144811476393242276341412462220262341377187436595412727672425665063935184413418239851935033660238993878510409748629527133631945663464698774349767646996;
            6'd31: xpb[22] = 1024'd26510802865300267225928368136355046289670186185217875372909898462250235137304763529523968736663922644340327173242950568623463341257829056139875672647345824003975061801549179330570158103163231848931120032266891798110087967262185926955862657138096794684489614129676364477598048447943494921196014043711505833140;
            6'd32: xpb[22] = 1024'd43374595949229274736287209354278039104781924723545637046633682937158551798160935115639589820383103930860098941084012643040873622052110036603118129831625501027805312126705116384798903744106201356485052627938370868547750269460436669498307074424258555708740234380842319206566569762255044178927329313073244019284;
            6'd33: xpb[22] = 1024'd60238389033158282246646050572201031919893663261873398720357467412066868459017106701755210904102285217379870708925074717458283902846391017066360587015905178051635562451861053439027649385049170864038985223609849938985412571658687412040751491710420316732990854632008273935535091076566593436658644582434982205428;
            6'd34: xpb[22] = 1024'd77102182117087289757004891790124024735005401800201160394081251886975185119873278287870831987821466503899642476766136791875694183640671997529603044200184855075465812777016990493256395025992140371592917819281329009423074873856938154583195908996582077757241474883174228664503612390878142694389959851796720391572;
            6'd35: xpb[22] = 1024'd93965975201016297267363733008047017550117140338528922067805036361883501780729449873986453071540647790419414244607198866293104464434952977992845501384464532099296063102172927547485140666935109879146850414952808079860737176055188897125640326282743838781492095134340183393472133705189691952121275121158458577716;
            6'd36: xpb[22] = 1024'd110829768284945304777722574225970010365228878876856683741528820836791818441585621460102074155259829076939186012448260940710514745229233958456087958568744209123126313427328864601713886307878079386700783010624287150298399478253439639668084743568905599805742715385506138122440655019501241209852590390520196763860;
            6'd37: xpb[22] = 1024'd3626865684749570889282488039078570435642190289448761287120750246723239765132654136202624024321336054015808372831829580548861185182294604364170290736692845213265889182913584318312392757303843172944517997908526374371700930230793609245550591171837911563173432222555034821302648259884157450465215833256340465673;
            6'd38: xpb[22] = 1024'd20490658768678578399641329257001563250753928827776522960844534721631556425988825722318245108040517340535580140672891654966271465976575584827412747920972522237096139508069521372541138398246812680498450593580005444809363232429044351787995008457999672587424052473720989550271169574195706708196531102618078651817;
            6'd39: xpb[22] = 1024'd37354451852607585910000170474924556065865667366104284634568319196539873086844997308433866191759698627055351908513953729383681746770856565290655205105252199260926389833225458426769884039189782188052383189251484515247025534627295094330439425744161433611674672724886944279239690888507255965927846371979816837961;
            6'd40: xpb[22] = 1024'd54218244936536593420359011692847548880977405904432046308292103671448189747701168894549487275478879913575123676355015803801092027565137545753897662289531876284756640158381395480998629680132751695606315784922963585684687836825545836872883843030323194635925292976052899008208212202818805223659161641341555024105;
            6'd41: xpb[22] = 1024'd71082038020465600930717852910770541696089144442759807982015888146356506408557340480665108359198061200094895444196077878218502308359418526217140119473811553308586890483537332535227375321075721203160248380594442656122350139023796579415328260316484955660175913227218853737176733517130354481390476910703293210249;
            6'd42: xpb[22] = 1024'd87945831104394608441076694128693534511200882981087569655739672621264823069413512066780729442917242486614667212037139952635912589153699506680382576658091230332417140808693269589456120962018690710714180976265921726560012441222047321957772677602646716684426533478384808466145254831441903739121792180065031396393;
            6'd43: xpb[22] = 1024'd104809624188323615951435535346616527326312621519415331329463457096173139730269683652896350526636423773134438979878202027053322869947980487143625033842370907356247391133849206643684866602961660218268113571937400796997674743420298064500217094888808477708677153729550763195113776145753452996853107449426769582537;
            6'd44: xpb[22] = 1024'd121673417272252623461794376564539520141424360057743093003187241571081456391125855239011971610355605059654210747719264101470733150742261467606867491026650584380077641459005143697913612243904629725822046167608879867435337045618548807042661512174970238732927773980716717924082297460065002254584422718788507768681;
            6'd45: xpb[22] = 1024'd14470514672056889573354290377648080211837671470335170548779170981012877714672887915112521479417112036730833108102832741309079590695322113514949823194599220470217217214589863414512118693330393512065781154893119091508638497595902776620127359777902550490358490817765614622944290700447918495197048161524651470494;
            6'd46: xpb[22] = 1024'd31334307755985897083713131595571073026949410008662932222502955455921194375529059501228142563136293323250604875943894815726489871489603093978192280378878897494047467539745800468740864334273363019619713750564598161946300799794153519162571777064064311514609111068931569351912812014759467752928363430886389656638;
            6'd47: xpb[22] = 1024'd48198100839914904594071972813494065842061148546990693896226739930829511036385231087343763646855474609770376643784956890143900152283884074441434737563158574517877717864901737522969609975216332527173646346236077232383963101992404261705016194350226072538859731320097524080881333329071017010659678700248127842782;
            6'd48: xpb[22] = 1024'd65061893923843912104430814031417058657172887085318455569950524405737827697241402673459384730574655896290148411626018964561310433078165054904677194747438251541707968190057674577198355616159302034727578941907556302821625404190655004247460611636387833563110351571263478809849854643382566268390993969609866028926;
            6'd49: xpb[22] = 1024'd81925687007772919614789655249340051472284625623646217243674308880646144358097574259575005814293837182809920179467081038978720713872446035367919651931717928565538218515213611631427101257102271542281511537579035373259287706388905746789905028922549594587360971822429433538818375957694115526122309238971604215070;
            6'd50: xpb[22] = 1024'd98789480091701927125148496467263044287396364161973978917398093355554461018953745845690626898013018469329691947308143113396130994666727015831162109115997605589368468840369548685655846898045241049835444133250514443696950008587156489332349446208711355611611592073595388267786897272005664783853624508333342401214;
            6'd51: xpb[22] = 1024'd115653273175630934635507337685186037102508102700301740591121877830462777679809917431806247981732199755849463715149205187813541275461007996294404566300277282613198719165525485739884592538988210557389376728921993514134612310785407231874793863494873116635862212324761342996755418586317214041584939777695080587358;
            6'd52: xpb[22] = 1024'd8450370575435200747067251498294597172921414112893818136713807240394199003356950107906797850793706732926086075532773827651887715414068642202486898468225918703338294921110205456483098988413974343633111716206232738207913762762761201452259711097805428393292929161810239695617411826700130282197565220431224289171;
            6'd53: xpb[22] = 1024'd25314163659364208257426092716217589988033152651221579810437591715302515664213121694022418934512888019445857843373835902069297996208349622665729355652505595727168545246266142510711844629356943851187044311877711808645576064961011943994704128383967189417543549412976194424585933141011679539928880489792962475315;
            6'd54: xpb[22] = 1024'd42177956743293215767784933934140582803144891189549341484161376190210832325069293280138040018232069305965629611214897976486708277002630603128971812836785272750998795571422079564940590270299913358740976907549190879083238367159262686537148545670128950441794169664142149153554454455323228797660195759154700661459;
            6'd55: xpb[22] = 1024'd59041749827222223278143775152063575618256629727877103157885160665119148985925464866253661101951250592485401379055960050904118557796911583592214270021064949774829045896578016619169335911242882866294909503220669949520900669357513429079592962956290711466044789915308103882522975769634778055391511028516438847603;
            6'd56: xpb[22] = 1024'd75905542911151230788502616369986568433368368266204864831608945140027465646781636452369282185670431879005173146897022125321528838591192564055456727205344626798659296221733953673398081552185852373848842098892149019958562971555764171622037380242452472490295410166474058611491497083946327313122826297878177033747;
            6'd57: xpb[22] = 1024'd92769335995080238298861457587909561248480106804532626505332729614935782307637808038484903269389613165524944914738084199738939119385473544518699184389624303822489546546889890727626827193128821881402774694563628090396225273754014914164481797528614233514546030417640013340460018398257876570854141567239915219891;
            6'd58: xpb[22] = 1024'd109633129079009245809220298805832554063591845342860388179056514089844098968493979624600524353108794452044716682579146274156349400179754524981941641573903980846319796872045827781855572834071791388956707290235107160833887575952265656706926214814775994538796650668805968069428539712569425828585456836601653406035;
            6'd59: xpb[22] = 1024'd2430226478813511920780212618941114134005156755452465724648443499775520292041012300701074222170301429121339042962714913994695840132815170890023973741852616936459372627630547498454079283497555175200442277519346384907189027929619626284392062417708306296227367505854864768290532952952342069198082279337797107848;
            6'd60: xpb[22] = 1024'd19294019562742519431139053836864106949116895293780227398372227974683836952897183886816695305889482715641110810803776988412106120927096151353266430926132293960289622952786484552682824924440524682754374873190825455344851330127870368826836479703870067320477987757020819497259054267263891326929397548699535293992;
            6'd61: xpb[22] = 1024'd36157812646671526941497895054787099764228633832107989072096012449592153613753355472932316389608664002160882578644839062829516401721377131816508888110411970984119873277942421606911570565383494190308307468862304525782513632326121111369280896990031828344728608008186774226227575581575440584660712818061273480136;
            6'd62: xpb[22] = 1024'd53021605730600534451856736272710092579340372370435750745819796924500470274609527059047937473327845288680654346485901137246926682515658112279751345294691648007950123603098358661140316206326463697862240064533783596220175934524371853911725314276193589368979228259352728955196096895886989842392028087423011666280;
            6'd63: xpb[22] = 1024'd69885398814529541962215577490633085394452110908763512419543581399408786935465698645163558557047026575200426114326963211664336963309939092742993802478971325031780373928254295715369061847269433205416172660205262666657838236722622596454169731562355350393229848510518683684164618210198539100123343356784749852424;
        endcase
    end

    always_comb begin
        case(flag[7][16:12])
            5'd0: xpb[23] = 1024'd0;
            5'd1: xpb[23] = 1024'd86749191898458549472574418708556078209563849447091274093267365874317103596321870231279179640766207861720197882168025286081747244104220073206236259663251002055610624253410232769597807488212402712970105255876741737095500538920873338996614148848517111417480468761684638413133139524510088357854658626146488038568;
            5'd2: xpb[23] = 1024'd49431688112792357546349910012297723674429271768446864058402876683657311855334601552543288066874741413997246356878557137584430647367219811857312394310170963177530573937249248201565375784907599704630012903366243627826640227620849905028249728013804773568141034109252218796159750975091543698590627425667381592805;
            5'd3: xpb[23] = 1024'd12114184327126165620125401316039369139294694089802454023538387492997520114347332873807396492983274966274294831589088989087114050630219550508388528957090924299450523621088263633532944081602796696289920550855745518557779916320826471059885307179092435718801599456819799179186362425672999039326596225188275147042;
            5'd4: xpb[23] = 1024'd98863376225584715092699820024595447348858543536893728116805753367314623710669203105086576133749482827994492713757114275168861294734439623714624788620341926355061147874498496403130751569815199409260025806732487255653280455241699810056499456027609547136282068218504437592319501950183087397181254851334763185610;
            5'd5: xpb[23] = 1024'd61545872439918523166475311328337092813723965858249318081941264176654831969681934426350684559858016380271541188467646126671544697997439362365700923267261887476981097558337511835098319866510396400919933454221989146384420143941676376088135035192897209286942633566072017975346113400764542737917223650855656739847;
            5'd6: xpb[23] = 1024'd24228368654252331240250802632078738278589388179604908047076774985995040228694665747614792985966549932548589663178177978174228101260439101016777057914181848598901047242176527267065888163205593392579841101711491037115559832641652942119770614358184871437603198913639598358372724851345998078653192450376550294084;
            5'd7: xpb[23] = 1024'd110977560552710880712825221340634816488153237626696182140344140860312143825016535978893972626732757794268787545346203264255975345364659174223013317577432850654511671495586760036663695651417996105549946357588232774211060371562526281116384763206701982855083667675324236771505864375856086436507851076523038332652;
            5'd8: xpb[23] = 1024'd73660056767044688786600712644376461953018659948051772105479651669652352084029267300158081052841291346545836020056735115758658748627658912874089452224352811776431621179425775468631263948113193097209854005077734664942200060262502847148020342371989645005744233022891817154532475826437541777243819876043931886889;
            5'd9: xpb[23] = 1024'd36342552981378496860376203948118107417884082269407362070615162478992560343041998621422189478949824898822884494767266967261342151890658651525165586871272772898351570863264790900598832244808390088869761652567236555673339748962479413179655921537277307156404798370459397537559087277018997117979788675564825441126;
            5'd10: xpb[23] = 1024'd123091744879837046332950622656674185627447931716498636163882528353309663939363868852701369119716032760543082376935292253343089395994878724731401846534523774953962195116675023670196639733020792801839866908443978292768840287883352752176270070385794418573885267132144035950692226801529085475834447301711313479694;
            5'd11: xpb[23] = 1024'd85774241094170854406726113960415831092313354037854226129018039162649872198376600173965477545824566312820130851645824104845772799257878463382477981181443736075882144800514039102164208029715989793499774555933480183499979976583329318207905649551082080724545832479711616333718838252110540816570416101232207033931;
            5'd12: xpb[23] = 1024'd48456737308504662480501605264157476557178776359209816094153549971990080457389331495229585971933099865097179326356355956348456202520878202033554115828363697197802094484353054534131776326411186785159682203422982074231119665283305884239541228716369742875206397827279196716745449702691996157306384900753100588168;
            5'd13: xpb[23] = 1024'd11139233522838470554277096567899122022044198680565406059289060781330288716402062816493694398041633417374227801066887807851139605783877940684630250475283658319722044168192069966099344623106383776819589850912483964962259353983282450271176807881657405025866963174846777099772061153273451498042353700273994142405;
            5'd14: xpb[23] = 1024'd97888425421297020026851515276455200231608048127656680152556426655647392312723933047772874038807841279094425683234913093932886849888098013890866510138534660375332668421602302735697152111318786489789695106789225702057759892904155789267790956730174516443347431936531415512905200677783539855897012326420482180973;
            5'd15: xpb[23] = 1024'd60570921635630828100627006580196845696473470449012270117691937464987600571736664369036982464916374831371474157945444945435570253151097752541942644785454621497252618105441318167664720408013983481449602754278727592788899581604132355299426535895462178594007997284098995895931812128364995196632981125941375735210;
            5'd16: xpb[23] = 1024'd23253417849964636174402497883938491161338892770367860082827448274327808830749395690301090891024908383648522632655976796938253656414097491193018779432374582619172567789280333599632288704709180473109510401768229483520039270304108921331062115060749840744668562631666576278958423578946450537368949925462269289447;
            5'd17: xpb[23] = 1024'd110002609748423185646976916592494569370902742217459134176094814148644912427071265921580270531791116245368720514824002083020000900518317564399255039095625584674783192042690566369230096192921583186079615657644971220615539809224982260327676263909266952162149031393351214692091563103456538895223608551608757328015;
            5'd18: xpb[23] = 1024'd72685105962756993720752407896236214835768164538814724141230324957985120686083997242844378957899649797645768989534533934522684303781317303050331173742545545796703141726529581801197664489616780177739523305134473111346679497924958826359311843074554614312809596740918795075118174554037994235959577351129650882252;
            5'd19: xpb[23] = 1024'd35367602177090801794527899199977860300633586860170314106365835767325328945096728564108487384008183349922817464245065786025367707044317041701407308389465506918623091410368597233165232786311977169399430952623975002077819186624935392390947422239842276463470162088486375458144786004619449576695546150650544436489;
            5'd20: xpb[23] = 1024'd122116794075549351267102317908533938510197436307261588199633201641642432541418598795387667024774391211643015346413091072107114951148537114907643568052716508974233715663778830002763040274524379882369536208500716739173319725545808731387561571088359387880950630850171013871277925529129537934550204776797032475057;
            5'd21: xpb[23] = 1024'd84799290289883159340877809212275583975062858628617178164768712450982640800431330116651775450882924763920063821123622923609798354411536853558719702699636470096153665347617845434730608571219576874029443855990218629904459414245785297419197150253647050031611196197738594254304536979710993275286173576317926029294;
            5'd22: xpb[23] = 1024'd47481786504216967414653300516017229439928280949972768129904223260322849059444061437915883876991458316197112295834154775112481757674536592209795837346556431218073615031456860866698176867914773865689351503479720520635599102945761863450832729418934712182271761545306174637331148430292448616022142375838819583531;
            5'd23: xpb[23] = 1024'd10164282718550775488428791819758874904793703271328358095039734069663057318456792759179992303099991868474160770544686626615165160937536330860871971993476392339993564715295876298665745164609970857349259150969222411366738791645738429482468308584222374332932326892873755020357759880873903956758111175359713137768;
            5'd24: xpb[23] = 1024'd96913474617009324961003210528314953114357552718419632188307099943980160914778662990459171943866199730194358652712711912696912405041756404067108231656727394395604188968706109068263552652822373570319364406845964148462239330566611768479082457432739485750412795654558393433490899405383992314612769801506201176336;
            5'd25: xpb[23] = 1024'd59595970831343133034778701832056598579222975039775222153442610753320369173791394311723280369974733282471407127423243764199595808304756142718184366303647355517524138652545124500231120949517570561979272054335466039193379019266588334510718036598027147901073361002125973816517510855965447655348738601027094730573;
            5'd26: xpb[23] = 1024'd22278467045676941108554193135798244044088397361130812118578121562660577432804125632987388796083266834748455602133775615702279211567755881369260500950567316639444088336384139932198689246212767553639179701824967929924518707966564900542353615763314810051733926349693554199544122306546902996084707400547988284810;
            5'd27: xpb[23] = 1024'd109027658944135490581128611844354322253652246808222086211845487436977681029125995864266568436849474696468653484301800901784026455671975954575496760613818318695054712589794372701796496734425170266609284957701709667020019246887438239538967764611831921469214395111378192612677261831056991353939366026694476323378;
            5'd28: xpb[23] = 1024'd71710155158469298654904103148095967718517669129577676176980998246317889288138727185530676862958008248745701959012332753286709858934975693226572895260738279816974662273633388133764065031120367258269192605191211557751158935587414805570603343777119583619874960458945772995703873281638446694675334826215369877615;
            5'd29: xpb[23] = 1024'd34392651372803106728679594451837613183383091450933266142116509055658097547151458506794785289066541801022750433722864604789393262197975431877649029907658240938894611957472403565731633327815564249929100252680713448482298624287391371602238922942407245770535525806513353378730484732219902035411303625736263431852;
            5'd30: xpb[23] = 1024'd121141843271261656201254013160393691392946940898024540235383874929975201143473328738073964929832749662742948315890889890871140506302195505083885289570909242994505236210882636335329440816027966962899205508557455185577799163208264710598853071790924357188015994568197991791863624256729990393265962251882751470420;
            5'd31: xpb[23] = 1024'd83824339485595464275029504464135336857812363219380130200519385739315409402486060059338073355941283215019996790601421742373823909565195243734961424217829204116425185894721651767297009112723163954559113156046957076308938851908241276630488650956212019338676559915765572174890235707311445734001931051403645024657;
        endcase
    end

    always_comb begin
        case(flag[8][5:0])
            6'd0: xpb[24] = 1024'd0;
            6'd1: xpb[24] = 1024'd23253417849964636174402497883938491161338892770367860082827448274327808830749395690301090891024908383648522632655976796938253656414097491193018779432374582619172567789280333599632288704709180473109510401768229483520039270304108921331062115060749840744668562631666576278958423578946450537368949925462269289447;
            6'd2: xpb[24] = 1024'd46506835699929272348804995767876982322677785540735720165654896548655617661498791380602181782049816767297045265311953593876507312828194982386037558864749165238345135578560667199264577409418360946219020803536458967040078540608217842662124230121499681489337125263333152557916847157892901074737899850924538578894;
            6'd3: xpb[24] = 1024'd69760253549893908523207493651815473484016678311103580248482344822983426492248187070903272673074725150945567897967930390814760969242292473579056338297123747857517703367841000798896866114127541419328531205304688450560117810912326763993186345182249522234005687894999728836875270736839351612106849776386807868341;
            6'd4: xpb[24] = 1024'd93013671399858544697609991535753964645355571081471440331309793097311235322997582761204363564099633534594090530623907187753014625656389964772075117729498330476690271157121334398529154818836721892438041607072917934080157081216435685324248460242999362978674250526666305115833694315785802149475799701849077157788;
            6'd5: xpb[24] = 1024'd116267089249823180872012489419692455806694463851839300414137241371639044153746978451505454455124541918242613163279883984691268282070487455965093897161872913095862838946401667998161443523545902365547552008841147417600196351520544606655310575303749203723342813158332881394792117894732252686844749627311346447235;
            6'd6: xpb[24] = 1024'd15453811415663075647616059898816514223334929496471476368832834580989957647187235231791474131491775992447986388478367347050458097643364612602952551577916454781344732166110784260163493036737877117346864802222137054755874771603756755021394120681269595201191472375882399643644013399750070207095009726148021252351;
            6'd7: xpb[24] = 1024'd38707229265627711822018557782755005384673822266839336451660282855317766477936630922092565022516684376096509021134344143988711754057462103795971331010291037400517299955391117859795781741447057590456375203990366538275914041907865676352456235742019435945860035007548975922602436978696520744463959651610290541798;
            6'd8: xpb[24] = 1024'd61960647115592347996421055666693496546012715037207196534487731129645575308686026612393655913541592759745031653790320940926965410471559594988990110442665620019689867744671451459428070446156238063565885605758596021795953312211974597683518350802769276690528597639215552201560860557642971281832909577072559831245;
            6'd9: xpb[24] = 1024'd85214064965556984170823553550631987707351607807575056617315179403973384139435422302694746804566501143393554286446297737865219066885657086182008889875040202638862435533951785059060359150865418536675396007526825505315992582516083519014580465863519117435197160270882128480519284136589421819201859502534829120692;
            6'd10: xpb[24] = 1024'd108467482815521620345226051434570478868690500577942916700142627678301192970184817992995837695591409527042076919102274534803472723299754577375027669307414785258035003323232118658692647855574599009784906409295054988836031852820192440345642580924268958179865722902548704759477707715535872356570809427997098410139;
            6'd11: xpb[24] = 1024'd7654204981361515120829621913694537285330966222575092654838220887652106463625074773281857371958643601247450144300757897162662538872631734012886323723458326943516896542941234920694697368766573761584219202676044625991710272903404588711726126301789349657714382120098223008329603220553689876821069526833773215255;
            6'd12: xpb[24] = 1024'd30907622831326151295232119797633028446669858992942952737665669161979915294374470463582948262983551984895972776956734694100916195286729225205905103155832909562689464332221568520326986073475754234693729604444274109511749543207513510042788241362539190402382944751764799287288026799500140414190019452296042504702;
            6'd13: xpb[24] = 1024'd54161040681290787469634617681571519608008751763310812820493117436307724125123866153884039154008460368544495409612711491039169851700826716398923882588207492181862032121501902119959274778184934707803240006212503593031788813511622431373850356423289031147051507383431375566246450378446590951558969377758311794149;
            6'd14: xpb[24] = 1024'd77414458531255423644037115565510010769347644533678672903320565710635532955873261844185130045033368752193018042268688287977423508114924207591942662020582074801034599910782235719591563482894115180912750407980733076551828083815731352704912471484038871891720070015097951845204873957393041488927919303220581083596;
            6'd15: xpb[24] = 1024'd100667876381220059818439613449448501930686537304046532986148013984963341786622657534486220936058277135841540674924665084915677164529021698784961441452956657420207167700062569319223852187603295654022260809748962560071867354119840274035974586544788712636388632646764528124163297536339492026296869228682850373043;
            6'd16: xpb[24] = 1024'd123921294231184695992842111333386993092025430074414393068975462259291150617372053224787311827083185519490063307580641881853930820943119189977980220885331240039379735489342902918856140892312476127131771211517192043591906624423949195367036701605538553381057195278431104403121721115285942563665819154145119662490;
            6'd17: xpb[24] = 1024'd23108016397024590768445681812511051508665895719046569023671055468642064110812310005073331503450419593695436532779125244213120636515996346615838875301374781724861628709052019180858190405504450878931084004898181680747585044507161343733120246983058944858905854495980622651973616620303760083916079252981794467606;
            6'd18: xpb[24] = 1024'd46361434246989226942848179696449542670004788489414429106498503742969872941561705695374422394475327977343959165435102041151374292930093837808857654733749364344034196498332352780490479110213631352040594406666411164267624314811270265064182362043808785603574417127647198930932040199250210621285029178444063757053;
            6'd19: xpb[24] = 1024'd69614852096953863117250677580388033831343681259782289189325952017297681772311101385675513285500236360992481798091078838089627949344191329001876434166123946963206764287612686380122767814922811825150104808434640647787663585115379186395244477104558626348242979759313775209890463778196661158653979103906333046500;
            6'd20: xpb[24] = 1024'd92868269946918499291653175464326524992682574030150149272153400291625490603060497075976604176525144744641004430747055635027881605758288820194895213598498529582379332076893019979755056519631992298259615210202870131307702855419488107726306592165308467092911542390980351488848887357143111696022929029368602335947;
            6'd21: xpb[24] = 1024'd116121687796883135466055673348265016154021466800518009354980848565953299433809892766277695067550053128289527063403032431966135262172386311387913993030873112201551899866173353579387345224341172771369125611971099614827742125723597029057368707226058307837580105022646927767807310936089562233391878954830871625394;
            6'd22: xpb[24] = 1024'd15308409962723030241659243827389074570661932445150185309676441775304212927250149546563714743917287202494900288601515794325325077745263468025772647446916653887033793085882469841389394737533147523168438405352089251983420545806809177423452252603578699315428764240196446016659206441107379753642139053667546430510;
            6'd23: xpb[24] = 1024'd38561827812687666416061741711327565732000825215518045392503890049632021757999545236864805634942195586143422921257492591263578734159360959218791426879291236506206360875162803441021683442242327996277948807120318735503459816110918098754514367664328540060097326871863022295617630020053830291011088979129815719957;
            6'd24: xpb[24] = 1024'd61815245662652302590464239595266056893339717985885905475331338323959830588748940927165896525967103969791945553913469388201832390573458450411810206311665819125378928664443137040653972146951508469387459208888548219023499086415027020085576482725078380804765889503529598574576053599000280828380038904592085009404;
            6'd25: xpb[24] = 1024'd85068663512616938764866737479204548054678610756253765558158786598287639419498336617466987416992012353440468186569446185140086046987555941604828985744040401744551496453723470640286260851660688942496969610656777702543538356719135941416638597785828221549434452135196174853534477177946731365748988830054354298851;
            6'd26: xpb[24] = 1024'd108322081362581574939269235363143039216017503526621625640986234872615448250247732307768078308016920737088990819225422982078339703401653432797847765176414984363724064243003804239918549556369869415606480012425007186063577627023244862747700712846578062294103014766862751132492900756893181903117938755516623588298;
            6'd27: xpb[24] = 1024'd7508803528421469714872805842267097632657969171253801595681828081966361743687989088054097984384154811294364044423906344437529518974530589435706419592458526049205957462712920501920599069561844167405792805805996823219256047106457011113784258224098453771951673984412269381344796261910999423368198854353298393414;
            6'd28: xpb[24] = 1024'd30762221378386105889275303726205588793996861941621661678509276356294170574437384778355188875409063194942886677079883141375783175388628080628725199024833108668378525251993254101552887774271024640515303207574226306739295317410565932444846373284848294516620236616078845660303219840857449960737148779815567682861;
            6'd29: xpb[24] = 1024'd54015639228350742063677801610144079955335754711989521761336724630621979405186780468656279766433971578591409309735859938314036831802725571821743978457207691287551093041273587701185176478980205113624813609342455790259334587714674853775908488345598135261288799247745421939261643419803900498106098705277836972308;
            6'd30: xpb[24] = 1024'd77269057078315378238080299494082571116674647482357381844164172904949788235936176158957370657458879962239931942391836735252290488216823063014762757889582273906723660830553921300817465183689385586734324011110685273779373858018783775106970603406347976005957361879411998218220066998750351035475048630740106261755;
            6'd31: xpb[24] = 1024'd100522474928280014412482797378021062278013540252725241926991621179277597066685571849258461548483788345888454575047813532190544144630920554207781537321956856525896228619834254900449753888398566059843834412878914757299413128322892696438032718467097816750625924511078574497178490577696801572843998556202375551202;
            6'd32: xpb[24] = 1024'd123775892778244650586885295261959553439352433023093102009819069453605405897434967539559552439508696729536977207703790329128797801045018045400800316754331439145068796409114588500082042593107746532953344814647144240819452398627001617769094833527847657495294487142745150776136914156643252110212948481664644840649;
            6'd33: xpb[24] = 1024'd22962614944084545362488865741083611855992898667725277964514662662956319390875224319845572115875930803742350432902273691487987616617895202038658971170374980830550689628823704762084092106299721284752657608028133877975130818710213766135178378905368048973143146360294669024988809661661069630463208580501319645765;
            6'd34: xpb[24] = 1024'd46216032794049181536891363625022103017331791438093138047342110937284128221624620010146663006900839187390873065558250488426241273031992693231677750602749563449723257418104038361716380811008901757862168009796363361495170089014322687466240493966117889717811708991961245303947233240607520167832158505963588935212;
            6'd35: xpb[24] = 1024'd69469450644013817711293861508960594178670684208460998130169559211611937052374015700447753897925747571039395698214227285364494929446090184424696530035124146068895825207384371961348669515718082230971678411564592845015209359318431608797302609026867730462480271623627821582905656819553970705201108431425858224659;
            6'd36: xpb[24] = 1024'd92722868493978453885696359392899085340009576978828858212997007485939745883123411390748844788950655954687918330870204082302748585860187675617715309467498728688068392996664705560980958220427262704081188813332822328535248629622540530128364724087617571207148834255294397861864080398500421242570058356888127514106;
            6'd37: xpb[24] = 1024'd115976286343943090060098857276837576501348469749196718295824455760267554713872807081049935679975564338336440963526180879241002242274285166810734088899873311307240960785945039160613246925136443177190699215101051812055287899926649451459426839148367411951817396886960974140822503977446871779939008282350396803553;
            6'd38: xpb[24] = 1024'd15163008509782984835702427755961634917988935393828894250520048969618468207313063861335955356342798412541814188724664241600192057847162323448592743315916852992722854005654155422615296438328417928990012008482041449210966320009861599825510384525887803429666056104510492389674399482464689300189268381187071608669;
            6'd39: xpb[24] = 1024'd38416426359747621010104925639900126079327828164196754333347497243946277038062459551637046247367706796190336821380641038538445714261259814641611522748291435611895421794934489022247585143037598402099522410250270932731005590313970521156572499586637644174334618736177068668632823061411139837558218306649340898116;
            6'd40: xpb[24] = 1024'd61669844209712257184507423523838617240666720934564614416174945518274085868811855241938137138392615179838859454036617835476699370675357305834630302180666018231067989584214822621879873847746778875209032812018500416251044860618079442487634614647387484919003181367843644947591246640357590374927168232111610187563;
            6'd41: xpb[24] = 1024'd84923262059676893358909921407777108402005613704932474499002393792601894699561250932239228029417523563487382086692594632414953027089454797027649081613040600850240557373495156221512162552455959348318543213786729899771084130922188363818696729708137325663671743999510221226549670219304040912296118157573879477010;
            6'd42: xpb[24] = 1024'd108176679909641529533312419291715599563344506475300334581829842066929703530310646622540318920442431947135904719348571429353206683503552288220667861045415183469413125162775489821144451257165139821428053615554959383291123401226297285149758844768887166408340306631176797505508093798250491449665068083036148766457;
            6'd43: xpb[24] = 1024'd7363402075481424308915989770839657979984972119932510536525435276280617023750903402826338596809666021341277944547054791712396499076429444858526515461458725154895018382484606083146500770357114573227366408935949020446801821309509433515842390146407557886188965848726315754359989303268308969915328181872823571573;
            6'd44: xpb[24] = 1024'd30616819925446060483318487654778149141323864890300370619352883550608425854500299093127429487834574404989800577203031588650650155490526936051545294893833307774067586171764939682778789475066295046336876810704178503966841091613618354846904505207157398630857528480392892033318412882214759507284278107335092861020;
            6'd45: xpb[24] = 1024'd53870237775410696657720985538716640302662757660668230702180331824936234685249694783428520378859482788638323209859008385588903811904624427244564074326207890393240153961045273282411078179775475519446387212472407987486880361917727276177966620267907239375526091112059468312276836461161210044653228032797362150467;
            6'd46: xpb[24] = 1024'd77123655625375332832123483422655131464001650431036090785007780099264043515999090473729611269884391172286845842514985182527157468318721918437582853758582473012412721750325606882043366884484655992555897614240637471006919632221836197509028735328657080120194653743726044591235260040107660582022177958259631439914;
            6'd47: xpb[24] = 1024'd100377073475339969006525981306593622625340543201403950867835228373591852346748486164030702160909299555935368475170961979465411124732819409630601633190957055631585289539605940481675655589193836465665408016008866954526958902525945118840090850389406920864863216375392620870193683619054111119391127883721900729361;
            6'd48: xpb[24] = 1024'd123630491325304605180928479190532113786679435971771810950662676647919661177497881854331793051934207939583891107826938776403664781146916900823620412623331638250757857328886274081307944293903016938774918417777096438046998172830054040171152965450156761609531779007059197149152107198000561656760077809184170018808;
            6'd49: xpb[24] = 1024'd22817213491144499956532049669656172203319901616403986905358269857270574670938138634617812728301442013789264333025422138762854596719794057461479067039375179936239750548595390343309993807094991690574231211158086075202676592913266188537236510827677153087380438224608715398004002703018379177010337908020844823924;
            6'd50: xpb[24] = 1024'd46070631341109136130934547553594663364658794386771846988185718131598383501687534324918903619326350397437786965681398935701108253133891548654497846471749762555412318337875723942942282511804172163683741612926315558722715863217375109868298625888426993832049000856275291676962426281964829714379287833483114113371;
            6'd51: xpb[24] = 1024'd69324049191073772305337045437533154525997687157139707071013166405926192332436930015219994510351258781086309598337375732639361909547989039847516625904124345174584886127156057542574571216513352636793252014694545042242755133521484031199360740949176834576717563487941867955920849860911280251748237758945383402818;
            6'd52: xpb[24] = 1024'd92577467041038408479739543321471645687336579927507567153840614680254001163186325705521085401376167164734832230993352529577615565962086531040535405336498927793757453916436391142206859921222533109902762416462774525762794403825592952530422856009926675321386126119608444234879273439857730789117187684407652692265;
            6'd53: xpb[24] = 1024'd115830884891003044654142041205410136848675472697875427236668062954581809993935721395822176292401075548383354863649329326515869222376184022233554184768873510412930021705716724741839148625931713583012272818231004009282833674129701873861484971070676516066054688751275020513837697018804181326486137609869921981712;
            6'd54: xpb[24] = 1024'd15017607056842939429745611684534195265315938342507603191363656163932723487375978176108195968768309622588728088847812688875059037949061178871412839184917052098411914925425841003841198139123688334811585611611993646438512094212914022227568516448196907543903347968824538762689592523821998846736397708706596786828;
            6'd55: xpb[24] = 1024'd38271024906807575604148109568472686426654831112875463274191104438260532318125373866409286859793218006237250721503789485813312694363158670064431618617291634717584482714706174603473486843832868807921096013380223129958551364517022943558630631508946748288571910600491115041648016102768449384105347634168866076275;
            6'd56: xpb[24] = 1024'd61524442756772211778550607452411177587993723883243323357018552712588341148874769556710377750818126389885773354159766282751566350777256161257450398049666217336757050503986508203105775548542049281030606415148452613478590634821131864889692746569696589033240473232157691320606439681714899921474297559631135365722;
            6'd57: xpb[24] = 1024'd84777860606736847952953105336349668749332616653611183439846000986916149979624165247011468641843034773534295986815743079689820007191353652450469177482040799955929618293266841802738064253251229754140116816916682096998629905125240786220754861630446429777909035863824267599564863260661350458843247485093404655169;
            6'd58: xpb[24] = 1024'd108031278456701484127355603220288159910671509423979043522673449261243958810373560937312559532867943157182818619471719876628073663605451143643487956914415382575102186082547175402370352957960410227249627218684911580518669175429349707551816976691196270522577598495490843878523286839607800996212197410555673944616;
            6'd59: xpb[24] = 1024'd7218000622541378902959173699412218327311975068611219477369042470594872303813817717598579209235177231388191844670203238987263479178328300281346611330458924260584079302256291664372402471152384979048940012065901217674347595512561855917900522068716662000426257713040362127375182344625618516462457509392348749732;
            6'd60: xpb[24] = 1024'd30471418472506015077361671583350709488650867838979079560196490744922681134563213407899670100260085615036714477326180035925517135592425791474365390762833506879756647091536625264004691175861565452158450413834130701194386865816670777248962637129466502745094820344706938406333605923572069053831407434854618039179;
            6'd61: xpb[24] = 1024'd53724836322470651251764169467289200649989760609346939643023939019250489965312609098200760991284993998685237109982156832863770792006523282667384170195208089498929214880816958863636979880570745925267960815602360184714426136120779698580024752190216343489763382976373514685292029502518519591200357360316887328626;
            6'd62: xpb[24] = 1024'd76978254172435287426166667351227691811328653379714799725851387293578298796062004788501851882309902382333759742638133629802024448420620773860402949627582672118101782670097292463269268585279926398377471217370589668234465406424888619911086867250966184234431945608040090964250453081464970128569307285779156618073;
            6'd63: xpb[24] = 1024'd100231672022399923600569165235166182972667546150082659808678835567906107626811400478802942773334810765982282375294110426740278104834718265053421729059957254737274350459377626062901557289989106871486981619138819151754504676728997541242148982311716024979100508239706667243208876660411420665938257211241425907520;
        endcase
    end

    always_comb begin
        case(flag[8][11:6])
            6'd0: xpb[25] = 1024'd0;
            6'd1: xpb[25] = 1024'd123485089872364559774971663119104674134006438920450519891506283842233916457560796169104033664359719149630805007950087223678531761248815756246440508492331837356446918248657959662533845994698287344596492020907048635274543947033106462573211097372465865723769070871373243522167300239357871203307207136703695196967;
            6'd2: xpb[25] = 1024'd122903484060604378151144398833394915523314450715165355654880712619490937577812453428192996114061763989818460608442681012777999681656411177937720891968332633779203161927744701987437452797879368967882786433426857424184727043845316152181443625061702282180718238328629429014228072404787109389495724446781795909603;
            6'd3: xpb[25] = 1024'd122321878248844196527317134547685156912622462509880191418255141396747958698064110687281958563763808830006116208935274801877467602064006599629001275444333430201959405606831444312341059601060450591169080845946666213094910140657525841789676152750938698637667405785885614506288844570216347575684241756859896622239;
            6'd4: xpb[25] = 1024'd121740272437084014903489870261975398301930474304595027181629570174004979818315767946370921013465853670193771809427868590976935522471602021320281658920334226624715649285918186637244666404241532214455375258466475002005093237469735531397908680440175115094616573243141799998349616735645585761872759066937997334875;
            6'd5: xpb[25] = 1024'd121158666625323833279662605976265639691238486099309862945003998951262000938567425205459883463167898510381427409920462380076403442879197443011562042396335023047471892965004928962148273207422613837741669670986283790915276334281945221006141208129411531551565740700397985490410388901074823948061276377016098047511;
            6'd6: xpb[25] = 1024'd120577060813563651655835341690555881080546497894024698708378427728519022058819082464548845912869943350569083010413056169175871363286792864702842425872335819470228136644091671287051880010603695461027964083506092579825459431094154910614373735818647948008514908157654170982471161066504062134249793687094198760147;
            6'd7: xpb[25] = 1024'd119995455001803470032008077404846122469854509688739534471752856505776043179070739723637808362571988190756738610905649958275339283694388286394122809348336615892984380323178413611955486813784777084314258496025901368735642527906364600222606263507884364465464075614910356474531933231933300320438310997172299472783;
            6'd8: xpb[25] = 1024'd119413849190043288408180813119136363859162521483454370235127285283033064299322396982726770812274033030944394211398243747374807204101983708085403192824337412315740624002265155936859093616965858707600552908545710157645825624718574289830838791197120780922413243072166541966592705397362538506626828307250400185419;
            6'd9: xpb[25] = 1024'd118832243378283106784353548833426605248470533278169205998501714060290085419574054241815733261976077871132049811890837536474275124509579129776683576300338208738496867681351898261762700420146940330886847321065518946556008721530783979439071318886357197379362410529422727458653477562791776692815345617328500898055;
            6'd10: xpb[25] = 1024'd118250637566522925160526284547716846637778545072884041761876142837547106539825711500904695711678122711319705412383431325573743044917174551467963959776339005161253111360438640586666307223328021954173141733585327735466191818342993669047303846575593613836311577986678912950714249728221014879003862927406601610691;
            6'd11: xpb[25] = 1024'd117669031754762743536699020262007088027086556867598877525250571614804127660077368759993658161380167551507361012876025114673210965324769973159244343252339801584009355039525382911569914026509103577459436146105136524376374915155203358655536374264830030293260745443935098442775021893650253065192380237484702323327;
            6'd12: xpb[25] = 1024'd117087425943002561912871755976297329416394568662313713288625000392061148780329026019082620611082212391695016613368618903772678885732365394850524726728340598006765598718612125236473520829690185200745730558624945313286558011967413048263768901954066446750209912901191283934835794059079491251380897547562803035963;
            6'd13: xpb[25] = 1024'd116505820131242380289044491690587570805702580457028549051999429169318169900580683278171583060784257231882672213861212692872146806139960816541805110204341394429521842397698867561377127632871266824032024971144754102196741108779622737872001429643302863207159080358447469426896566224508729437569414857640903748599;
            6'd14: xpb[25] = 1024'd115924214319482198665217227404877812195010592251743384815373857946575191020832340537260545510486302072070327814353806481971614726547556238233085493680342190852278086076785609886280734436052348447318319383664562891106924205591832427480233957332539279664108247815703654918957338389937967623757932167719004461235;
            6'd15: xpb[25] = 1024'd115342608507722017041389963119168053584318604046458220578748286723832212141083997796349507960188346912257983414846400271071082646955151659924365877156342987275034329755872352211184341239233430070604613796184371680017107302404042117088466485021775696121057415272959840411018110555367205809946449477797105173871;
            6'd16: xpb[25] = 1024'd114761002695961835417562698833458294973626615841173056342122715501089233261335655055438470409890391752445639015338994060170550567362747081615646260632343783697790573434959094536087948042414511693890908208704180468927290399216251806696699012711012112578006582730216025903078882720796443996134966787875205886507;
            6'd17: xpb[25] = 1024'd114179396884201653793735434547748536362934627635887892105497144278346254381587312314527432859592436592633294615831587849270018487770342503306926644108344580120546817114045836860991554845595593317177202621223989257837473496028461496304931540400248529034955750187472211395139654886225682182323484097953306599143;
            6'd18: xpb[25] = 1024'd113597791072441472169908170262038777752242639430602727868871573055603275501838969573616395309294481432820950216324181638369486408177937924998207027584345376543303060793132579185895161648776674940463497033743798046747656592840671185913164068089484945491904917644728396887200427051654920368512001408031407311779;
            6'd19: xpb[25] = 1024'd113016185260681290546080905976329019141550651225317563632246001832860296622090626832705357758996526273008605816816775427468954328585533346689487411060346172966059304472219321510798768451957756563749791446263606835657839689652880875521396595778721361948854085101984582379261199217084158554700518718109508024415;
            6'd20: xpb[25] = 1024'd112434579448921108922253641690619260530858663020032399395620430610117317742342284091794320208698571113196261417309369216568422248993128768380767794536346969388815548151306063835702375255138838187036085858783415624568022786465090565129629123467957778405803252559240767871321971382513396740889036028187608737051;
            6'd21: xpb[25] = 1024'd111852973637160927298426377404909501920166674814747235158994859387374338862593941350883282658400615953383917017801963005667890169400724190072048178012347765811571791830392806160605982058319919810322380271303224413478205883277300254737861651157194194862752420016496953363382743547942634927077553338265709449687;
            6'd22: xpb[25] = 1024'd111271367825400745674599113119199743309474686609462070922369288164631359982845598609972245108102660793571572618294556794767358089808319611763328561488348562234328035509479548485509588861501001433608674683823033202388388980089509944346094178846430611319701587473753138855443515713371873113266070648343810162323;
            6'd23: xpb[25] = 1024'd110689762013640564050771848833489984698782698404176906685743716941888381103097255869061207557804705633759228218787150583866826010215915033454608944964349358657084279188566290810413195664682083056894969096342841991298572076901719633954326706535667027776650754931009324347504287878801111299454587958421910874959;
            6'd24: xpb[25] = 1024'd110108156201880382426944584547780226088090710198891742449118145719145402223348913128150170007506750473946883819279744372966293930623510455145889328440350155079840522867653033135316802467863164680181263508862650780208755173713929323562559234224903444233599922388265509839565060044230349485643105268500011587595;
            6'd25: xpb[25] = 1024'd109526550390120200803117320262070467477398721993606578212492574496402423343600570387239132457208795314134539419772338162065761851031105876837169711916350951502596766546739775460220409271044246303467557921382459569118938270526139013170791761914139860690549089845521695331625832209659587671831622578578112300231;
            6'd26: xpb[25] = 1024'd108944944578360019179290055976360708866706733788321413975867003273659444463852227646328094906910840154322195020264931951165229771438701298528450095392351747925353010225826517785124016074225327926753852333902268358029121367338348702779024289603376277147498257302777880823686604375088825858020139888656213012867;
            6'd27: xpb[25] = 1024'd108363338766599837555462791690650950256014745583036249739241432050916465584103884905417057356612884994509850620757525740264697691846296720219730478868352544348109253904913260110027622877406409550040146746422077146939304464150558392387256817292612693604447424760034066315747376540518064044208657198734313725503;
            6'd28: xpb[25] = 1024'd107781732954839655931635527404941191645322757377751085502615860828173486704355542164506019806314929834697506221250119529364165612253892141911010862344353340770865497584000002434931229680587491173326441158941885935849487560962768081995489344981849110061396592217290251807808148705947302230397174508812414438139;
            6'd29: xpb[25] = 1024'd107200127143079474307808263119231433034630769172465921265990289605430507824607199423594982256016974674885161821742713318463633532661487563602291245820354137193621741263086744759834836483768572796612735571461694724759670657774977771603721872671085526518345759674546437299868920871376540416585691818890515150775;
            6'd30: xpb[25] = 1024'd106618521331319292683980998833521674423938780967180757029364718382687528944858856682683944705719019515072817422235307107563101453069082985293571629296354933616377984942173487084738443286949654419899029983981503513669853754587187461211954400360321942975294927131802622791929693036805778602774209128968615863411;
            6'd31: xpb[25] = 1024'd106036915519559111060153734547811915813246792761895592792739147159944550065110513941772907155421064355260473022727900896662569373476678406984852012772355730039134228621260229409642050090130736043185324396501312302580036851399397150820186928049558359432244094589058808283990465202235016788962726439046716576047;
            6'd32: xpb[25] = 1024'd105455309707798929436326470262102157202554804556610428556113575937201571185362171200861869605123109195448128623220494685762037293884273828676132396248356526461890472300346971734545656893311817666471618809021121091490219948211606840428419455738794775889193262046314993776051237367664254975151243749124817288683;
            6'd33: xpb[25] = 1024'd104873703896038747812499205976392398591862816351325264319488004714458592305613828459950832054825154035635784223713088474861505214291869250367412779724357322884646715979433714059449263696492899289757913221540929880400403045023816530036651983428031192346142429503571179268112009533093493161339761059202918001319;
            6'd34: xpb[25] = 1024'd104292098084278566188671941690682639981170828146040100082862433491715613425865485719039794504527198875823439824205682263960973134699464672058693163200358119307402959658520456384352870499673980913044207634060738669310586141836026219644884511117267608803091596960827364760172781698522731347528278369281018713955;
            6'd35: xpb[25] = 1024'd103710492272518384564844677404972881370478839940754935846236862268972634546117142978128756954229243716011095424698276053060441055107060093749973546676358915730159203337607198709256477302855062536330502046580547458220769238648235909253117038806504025260040764418083550252233553863951969533716795679359119426591;
            6'd36: xpb[25] = 1024'd103128886460758202941017413119263122759786851735469771609611291046229655666368800237217719403931288556198751025190869842159908975514655515441253930152359712152915447016693941034160084106036144159616796459100356247130952335460445598861349566495740441716989931875339735744294326029381207719905312989437220139227;
            6'd37: xpb[25] = 1024'd102547280648998021317190148833553364149094863530184607372985719823486676786620457496306681853633333396386406625683463631259376895922250937132534313628360508575671690695780683359063690909217225782903090871620165036041135432272655288469582094184976858173939099332595921236355098194810445906093830299515320851863;
            6'd38: xpb[25] = 1024'd101965674837237839693362884547843605538402875324899443136360148600743697906872114755395644303335378236574062226176057420358844816329846358823814697104361304998427934374867425683967297712398307406189385284139973824951318529084864978077814621874213274630888266789852106728415870360239684092282347609593421564499;
            6'd39: xpb[25] = 1024'd101384069025477658069535620262133846927710887119614278899734577378000719027123772014484606753037423076761717826668651209458312736737441780515095080580362101421184178053954168008870904515579389029475679696659782613861501625897074667686047149563449691087837434247108292220476642525668922278470864919671522277135;
            6'd40: xpb[25] = 1024'd100802463213717476445708355976424088317018898914329114663109006155257740147375429273573569202739467916949373427161244998557780657145037202206375464056362897843940421733040910333774511318760470652761974109179591402771684722709284357294279677252686107544786601704364477712537414691098160464659382229749622989771;
            6'd41: xpb[25] = 1024'd100220857401957294821881091690714329706326910709043950426483434932514761267627086532662531652441512757137029027653838787657248577552632623897655847532363694266696665412127652658678118121941552276048268521699400191681867819521494046902512204941922524001735769161620663204598186856527398650847899539827723702407;
            6'd42: xpb[25] = 1024'd99639251590197113198053827405004571095634922503758786189857863709771782387878743791751494102143557597324684628146432576756716497960228045588936231008364490689452909091214394983581724925122633899334562934219208980592050916333703736510744732631158940458684936618876848696658959021956636837036416849905824415043;
            6'd43: xpb[25] = 1024'd99057645778436931574226563119294812484942934298473621953232292487028803508130401050840456551845602437512340228639026365856184418367823467280216614484365287112209152770301137308485331728303715522620857346739017769502234013145913426118977260320395356915634104076133034188719731187385875023224934159983925127679;
            6'd44: xpb[25] = 1024'd98476039966676749950399298833585053874250946093188457716606721264285824628382058309929419001547647277699995829131620154955652338775418888971496997960366083534965396449387879633388938531484797145907151759258826558412417109958123115727209788009631773372583271533389219680780503352815113209413451470062025840315;
            6'd45: xpb[25] = 1024'd97894434154916568326572034547875295263558957887903293479981150041542845748633715569018381451249692117887651429624213944055120259183014310662777381436366879957721640128474621958292545334665878769193446171778635347322600206770332805335442315698868189829532438990645405172841275518244351395601968780140126552951;
            6'd46: xpb[25] = 1024'd97312828343156386702744770262165536652866969682618129243355578818799866868885372828107343900951736958075307030116807733154588179590609732354057764912367676380477883807561364283196152137846960392479740584298444136232783303582542494943674843388104606286481606447901590664902047683673589581790486090218227265587;
            6'd47: xpb[25] = 1024'd96731222531396205078917505976455778042174981477332965006730007596056887989137030087196306350653781798262962630609401522254056099998205154045338148388368472803234127486648106608099758941028042015766034996818252925142966400394752184551907371077341022743430773905157776156962819849102827767979003400296327978223;
            6'd48: xpb[25] = 1024'd96149616719636023455090241690746019431482993272047800770104436373313909109388687346285268800355826638450618231101995311353524020405800575736618531864369269225990371165734848933003365744209123639052329409338061714053149497206961874160139898766577439200379941362413961649023592014532065954167520710374428690859;
            6'd49: xpb[25] = 1024'd95568010907875841831262977405036260820791005066762636533478865150570930229640344605374231250057871478638273831594589100452991940813395997427898915340370065648746614844821591257906972547390205262338623821857870502963332594019171563768372426455813855657329108819670147141084364179961304140356038020452529403495;
            6'd50: xpb[25] = 1024'd94986405096115660207435713119326502210099016861477472296853293927827951349892001864463193699759916318825929432087182889552459861220991419119179298816370862071502858523908333582810579350571286885624918234377679291873515690831381253376604954145050272114278276276926332633145136345390542326544555330530630116131;
            6'd51: xpb[25] = 1024'd94404799284355478583608448833616743599407028656192308060227722705084972470143659123552156149461961159013585032579776678651927781628586840810459682292371658494259102202995075907714186153752368508911212646897488080783698787643590942984837481834286688571227443734182518125205908510819780512733072640608730828767;
            6'd52: xpb[25] = 1024'd93823193472595296959781184547906984988715040450907143823602151482341993590395316382641118599164005999201240633072370467751395702036182262501740065768372454917015345882081818232617792956933450132197507059417296869693881884455800632593070009523523105028176611191438703617266680676249018698921589950686831541403;
            6'd53: xpb[25] = 1024'd93241587660835115335953920262197226378023052245621979586976580259599014710646973641730081048866050839388896233564964256850863622443777684193020449244373251339771589561168560557521399760114531755483801471937105658604064981268010322201302537212759521485125778648694889109327452841678256885110107260764932254039;
            6'd54: xpb[25] = 1024'd92659981849074933712126655976487467767331064040336815350351009036856035830898630900819043498568095679576551834057558045950331542851373105884300832720374047762527833240255302882425006563295613378770095884456914447514248078080220011809535064901995937942074946105951074601388225007107495071298624570843032966675;
            6'd55: xpb[25] = 1024'd92078376037314752088299391690777709156639075835051651113725437814113056951150288159908005948270140519764207434550151835049799463258968527575581216196374844185284076919342045207328613366476695002056390296976723236424431174892429701417767592591232354399024113563207260093448997172536733257487141880921133679311;
            6'd56: xpb[25] = 1024'd91496770225554570464472127405067950545947087629766486877099866591370078071401945418996968397972185359951863035042745624149267383666563949266861599672375640608040320598428787532232220169657776625342684709496532025334614271704639391026000120280468770855973281020463445585509769337965971443675659190999234391947;
            6'd57: xpb[25] = 1024'd90915164413794388840644863119358191935255099424481322640474295368627099191653602678085930847674230200139518635535339413248735304074159370958141983148376437030796564277515529857135826972838858248628979122016340814244797368516849080634232647969705187312922448477719631077570541503395209629864176501077335104583;
            6'd58: xpb[25] = 1024'd90333558602034207216817598833648433324563111219196158403848724145884120311905259937174893297376275040327174236027933202348203224481754792649422366624377233453552807956602272182039433776019939871915273534536149603154980465329058770242465175658941603769871615934975816569631313668824447816052693811155435817219;
            6'd59: xpb[25] = 1024'd89751952790274025592990334547938674713871123013910994167223152923141141432156917196263855747078319880514829836520526991447671144889350214340702750100378029876309051635689014506943040579201021495201567947055958392065163562141268459850697703348178020226820783392232002061692085834253686002241211121233536529855;
            6'd60: xpb[25] = 1024'd89170346978513843969163070262228916103179134808625829930597581700398162552408574455352818196780364720702485437013120780547139065296945636031983133576378826299065295314775756831846647382382103118487862359575767180975346658953478149458930231037414436683769950849488187553752857999682924188429728431311637242491;
            6'd61: xpb[25] = 1024'd88588741166753662345335805976519157492487146603340665693972010477655183672660231714441780646482409560890141037505714569646606985704541057723263517052379622721821538993862499156750254185563184741774156772095575969885529755765687839067162758726650853140719118306744373045813630165112162374618245741389737955127;
            6'd62: xpb[25] = 1024'd88007135354993480721508541690809398881795158398055501457346439254912204792911888973530743096184454401077796637998308358746074906112136479414543900528380419144577782672949241481653860988744266365060451184615384758795712852577897528675395286415887269597668285764000558537874402330541400560806763051467838667763;
            6'd63: xpb[25] = 1024'd87425529543233299097681277405099640271103170192770337220720868032169225913163546232619705545886499241265452238490902147845542826519731901105824284004381215567334026352035983806557467791925347988346745597135193547705895949390107218283627814105123686054617453221256744029935174495970638746995280361545939380399;
        endcase
    end

    always_comb begin
        case(flag[8][16:12])
            5'd0: xpb[26] = 1024'd0;
            5'd1: xpb[26] = 1024'd86843923731473117473854013119389881660411181987485172984095296809426247033415203491708667995588544081453107838983495936945010746927327322797104667480382011990090270031122726131461074595106429611633040009655002336616079046202316907891860341794360102511566620678512929521995946661399876933183797671624040093035;
            5'd2: xpb[26] = 1024'd49621151778821493548909098833965330576123936849234661840058738553875598729521268073402264776519413853463066270509498439310957653013434311039049209944432983046489865492674234925291909998695653501955882410922764826867797242183737042818742113905490755756313337942908801013885365248871120849248905516622485701739;
            5'd3: xpb[26] = 1024'd12398379826169869623964184548540779491836691710984150696022180298324950425627332655095861557450283625473024702035500941676904559099541299280993752408483954102889460954225743719122745402284877392278724812190527317119515438165157177745623886016621409001060055207304672505774783836342364765314013361620931310443;
            5'd4: xpb[26] = 1024'd99242303557642987097818197667930661152247873698469323680117477107751197459042536146804529553038827706926132541018996878621915306026868622078098419888865966092979730985348469850583819997391307003911764821845529653735594484367474085637484227810981511512626675885817602027770730497742241698497811033244971403478;
            5'd5: xpb[26] = 1024'd62019531604991363172873283382506110067960628560218812536080918852200549155148600728498126333969697478936090972544999380987862212112975610320042962352916937149379326446899978644414655400980530894234607223113292143987312680348894220564365999922112164757373393150213473519660149085213485614562918878243417012182;
            5'd6: xpb[26] = 1024'd24796759652339739247928369097081558983673383421968301392044360596649900851254665310191723114900567250946049404071001883353809118199082598561987504816967908205778921908451487438245490804569754784557449624381054634239030876330314355491247772033242818002120110414609345011549567672684729530628026723241862620886;
            5'd7: xpb[26] = 1024'd111640683383812856721782382216471440644084565409453474376139657406076147884669868801900391110489111332399157243054497820298819865126409921359092172297349920195869191939574213569706565399676184396190489634036056970855109922532631263383108113827602920513686731093122274533545514334084606463811824394865902713921;
            5'd8: xpb[26] = 1024'd74417911431161232796837467931046889559797320271202963232103099150525499580775933383593987891419981104409115674580500322664766771212516909601036714761400891252268787401125722363537400803265408286513332035303819461106828118514051398309989885938733573758433448357518146025434932921555850379876932239864348322625;
            5'd9: xpb[26] = 1024'd37195139478509608871892553645622338475510075132952452088066540894974851276881997965287584672350850876419074106106502825030713677298623897842981257225451862308668382862677231157368236206854632176836174436571581951358546314495471533236871658049864227003180165621914017517324351509027094295942040084862793931329;
            5'd10: xpb[26] = 1024'd124039063209982726345746566765012220135921257120437625072161837704401098310297201456996252667939394957872181945089998761975724424225951220640085924705833874298758652893799957288829310801961061788469214446226584287974625360697788441128731999844224329514746786300426947039320298170426971229125837756486834024364;
            5'd11: xpb[26] = 1024'd86816291257331102420801652479587669051634011982187113928125279448850450006403266038689849448870264729882140376616001264341671330312058208882030467169884845355158248355351466082660146205550285678792056847494346778226343556679208576055613771955354982759493503564822818531209716757898215145190945601485279633068;
            5'd12: xpb[26] = 1024'd49593519304679478495856738194163117967346766843936602784088721193299801702509330620383446229801134501892098808142003766707618236398165197123975009633935816411557843816902974876490981609139509569114899248762109268478061752660628710982495544066485636004240220829218690023099135345369459061256053446483725241772;
            5'd13: xpb[26] = 1024'd12370747352027854570911823908738566883059521705686091640052162937749153398615395202077043010732004273902057239668006269073565142484272185365919552097986787467957439278454483670321817012728733459437741650029871758729779948642048845909377316177616289248986938093614561514988553932840702977321161291482170850476;
            5'd14: xpb[26] = 1024'd99214671083500972044765837028128448543470703693171264624147459747175400432030598693785711006320548355355165078651502206018575889411599508163024219578368799458047709309577209801782891607835163071070781659684874095345858994844365753801237657971976391760553558772127491036984500594240579910504958963106210943511;
            5'd15: xpb[26] = 1024'd61991899130849348119820922742703897459183458554920753480110901491624752128136663275479307787251418127365123510177504708384522795497706496404968762042419770514447304771128718595613727011424386961393624060952636585597577190825785888728119430083107045005300276036523362528873919181711823826570066808104656552215;
            5'd16: xpb[26] = 1024'd24769127178197724194876008457279346374896213416670242336074343236074103824242727857172904568182287899375081941703507210750469701583813484646913304506470741570846900232680227389444562415013610851716466462220399075849295386807206023655001202194237698250046993300919234020763337769183067742635174653103102160919;
            5'd17: xpb[26] = 1024'd111613050909670841668730021576669228035307395404155415320169640045500350857657931348881572563770831980828189780687003147695480448511140807444017971986852753560937170263802953520905637010120040463349506471875401412465374433009522931546861543988597800761613613979432163542759284430582944675818972324727142253954;
            5'd18: xpb[26] = 1024'd74390278957019217743785107291244676951020150265904904176133081789949702553763995930575169344701701752838148212213005650061427354597247795685962514450903724617336765725354462314736472413709264353672348873143163902717092628990943066473743316099728454006360331243828035034648703018054188591884080169725587862658;
            5'd19: xpb[26] = 1024'd37167507004367593818840193005820125866732905127654393032096523534399054249870060512268766125632571524848106643739008152427374260683354783927907056914954695673736361186905971108567307817298488243995191274410926392968810824972363201400625088210859107251107048508223906526538121605525432507949188014724033471362;
            5'd20: xpb[26] = 1024'd124011430735840711292694206125210007527144087115139566016191820343825301283285264003977434121221115606301214482722504089372385007610682106725011724395336707663826631218028697240028382412404917855628231284065928729584889871174680109292485430005219209762673669186736836048534068266925309441132985686348073564397;
            5'd21: xpb[26] = 1024'd86788658783189087367749291839785456442856841976889054872155262088274652979391328585671030902151985378311172914248506591738331913696789094966956266859387678720226226679580206033859217815994141745951073685333691219836608067156100244219367202116349863007420386451132707540423486854396553357198093531346519173101;
            5'd22: xpb[26] = 1024'd49565886830537463442804377554360905358569596838638543728118703832724004675497393167364627683082855150321131345774509094104278819782896083208900809323438649776625822141131714827690053219583365636273916086601453710088326263137520379146248974227480516252167103715528579032312905441867797273263201376344964781805;
            5'd23: xpb[26] = 1024'd12343114877885839517859463268936354274282351700388032584082145577173356371603457749058224464013724922331089777300511596470225725869003071450845351787489620833025417602683223621520888623172589526596758487869216200340044459118940514073130746338611169496913820979924450524202324029339041189328309221343410390509;
            5'd24: xpb[26] = 1024'd99187038609358956991713476388326235934693533687873205568177442386599603405018661240766892459602269003784197616284007533415236472796330394247950019267871632823115687633805949752981963218279019138229798497524218536956123505321257421964991088132971272008480441658437380046198270690738918122512106892967450483544;
            5'd25: xpb[26] = 1024'd61964266656707333066768562102901684850406288549622694424140884131048955101124725822460489240533138775794156047810010035781183378882437382489894561731922603879515283095357458546812798621868243028552640898791981027207841701302677556891872860244101925253227158922833251538087689278210162038577214737965896092248;
            5'd26: xpb[26] = 1024'd24741494704055709141823647817477133766119043411372183280104325875498306797230790404154086021464008547804114479336012538147130284968544370731839104195973574935914878556908967340643634025457466918875483300059743517459559897284097691818754632355232578497973876187229123029977107865681405954642322582964341700952;
            5'd27: xpb[26] = 1024'd111585418435528826615677660936867015426530225398857356264199622684924553830645993895862754017052552629257222318319508475092141031895871693528943771676355586926005148588031693472104708620563896530508523309714745854075638943486414599710614974149592681009540496865742052551973054527081282887826120254588381793987;
            5'd28: xpb[26] = 1024'd74362646482877202690732746651442464342242980260606845120163064429373905526752058477556350797983422401267180749845510977458087937981978681770888314140406557982404744049583202265935544024153120420831365710982508344327357139467834734637496746260723334254287214130137924043862473114552526803891228099586827402691;
            5'd29: xpb[26] = 1024'd37139874530225578765787832366017913257955735122356333976126506173823257222858123059249947578914292173277139181371513479824034844068085670012832856604457529038804339511134711059766379427742344311154208112250270834579075335449254869564378518371853987499033931394533795535751891702023770719956335944585273011395;
            5'd30: xpb[26] = 1024'd123983798261698696239641845485407794918366917109841506960221802983249504256273326550958615574502836254730247020355009416769045590995412992809937524084839541028894609542257437191227454022848773922787248121905273171195154381651571777456238860166214090010600552073046725057747838363423647653140133616209313104430;
            5'd31: xpb[26] = 1024'd86761026309047072314696931199983243834079671971590995816185244727698855952379391132652212355433706026740205451881011919134992497081519981051882066548890512085294205003808945985058289426437997813110090523173035661446872577632991912383120632277344743255347269337442596549637256950894891569205241461207758713134;
        endcase
    end

endmodule





module xpb_lut_final
(
    input logic [16:0] flag[2],
    output logic [1023:0] xpb[6]
);
        
        
    always_comb begin
        case(flag[0][5:0])
            6'd0: xpb[0] = 1024'd0;
            6'd1: xpb[0] = 1024'd55702617802106849374131591674088040617099270768494973145298226092755780468191824222693406107749861711676964472413899923079725927973196287937687305623143083444077218855294267938671980409728888398142885343697765922473789832121566108508934540857597787896530607270469240209840717864551083287716666502998629652885;
            6'd2: xpb[0] = 1024'd111405235604213698748263183348176081234198541536989946290596452185511560936383648445386812215499723423353928944827799846159451855946392575875374611246286166888154437710588535877343960819457776796285770687395531844947579664243132217017869081715195575793061214540938480419681435729102166575433333005997259305770;
            6'd3: xpb[0] = 1024'd43041157722195806723595847617449689106599385179749235307762823213290446067266333758065147108591910825587744009784206334660113943078368529257901791853098209398540981996311586478385702037669459473118458422706057921057008646143801552561825052889563914422771918397290662599415625519724616846031309682370294474324;
            6'd4: xpb[0] = 1024'd98743775524302656097727439291537729723698655948244208453061049306046226535458157980758553216341772537264708482198106257739839871051564817195589097476241292842618200851605854417057682447398347871261343766403823843530798478265367661070759593747161702319302525667759902809256343384275700133747976185368924127209;
            6'd5: xpb[0] = 1024'd30379697642284764073060103560811337596099499591003497470227420333825111666340843293436888109433959939498523547154512746240501958183540770578116278083053335353004745137328905018099423665610030548094031501714349919640227460166036996614715564921530040949013229524112084988990533174898150404345952861741959295763;
            6'd6: xpb[0] = 1024'd86082315444391613447191695234899378213198770359498470615525646426580892134532667516130294217183821651175488019568412669320227886156737058515803583706196418797081963992623172956771404075338918946236916845412115842114017292287603105123650105779127828845543836794581325198831251039449233692062619364740588948648;
            6'd7: xpb[0] = 1024'd17718237562373721422524359504172986085599614002257759632692017454359777265415352828808629110276009053409303084524819157820889973288713011898330764313008461307468508278346223557813145293550601623069604580722641918223446274188272440667606076953496167475254540650933507378565440830071683962660596041113624117202;
            6'd8: xpb[0] = 1024'd73420855364480570796655951178261026702698884770752732777990243547115557733607177051502035218025870765086267556938719080900615901261909299836018069936151544751545727133640491496485125703279490021212489924420407840697236106309838549176540617811093955371785147921402747588406158694622767250377262544112253770087;
            6'd9: xpb[0] = 1024'd5056777482462678771988615447534634575099728413512021795156614574894442864489862364180370111118058167320082621895125569401277988393885253218545250542963587261932271419363542097526866921491172698045177659730933916806665088210507884720496588985462294001495851777754929768140348485245217520975239220485288938641;
            6'd10: xpb[0] = 1024'd60759395284569528146120207121622675192198999182006994940454840667650223332681686586873776218867919878997047094309025492481003916367081541156232556166106670706009490274657810036198847331220061096188063003428699839280454920332073993229431129843060081898026459048224169977981066349796300808691905723483918591526;
            6'd11: xpb[0] = 1024'd116462013086676377520251798795710715809298269950501968085753066760406003800873510809567182326617781590674011566722925415560729844340277829093919861789249754150086709129952077974870827740948949494330948347126465761754244752453640101738365670700657869794557066318693410187821784214347384096408572226482548244411;
            6'd12: xpb[0] = 1024'd48097935204658485495584463064984323681699113593261257102919437788184888931756196122245517219709968992907826631679331904061391931472253782476447042396061796660473253415675128575912568959160632171163636082436991837863673734354309437282321641875026208424267770175045592367555974004969834367006548902855583412965;
            6'd13: xpb[0] = 1024'd103800553006765334869716054739072364298798384361756230248217663880940669399948020344938923327459830704584791104093231827141117859445450070414134348019204880104550472270969396514584549368889520569306521426134757760337463566475875545791256182732623996320798377445514832577396691869520917654723215405854213065850;
            6'd14: xpb[0] = 1024'd35436475124747442845048719008345972171199228004515519265384034908719554530830705657617258220552018106818606169049638315641779946577426023796661528626016922614937016556692447115626290587101203246139209161445283836446892548376544881335212153906992334950509081301867014757130881660143367925321192082227248234404;
            6'd15: xpb[0] = 1024'd91139092926854292219180310682434012788298498773010492410682261001475334999022529880310664328301879818495570641463538238721505874550622311734348834249160006059014235411986715054298270996830091644282094505143049758920682380498110989844146694764590122847039688572336254966971599524694451213037858585225877887289;
            6'd16: xpb[0] = 1024'd22775015044836400194512974951707620660699342415769781427848632029254220129905215192988999221394067220729385706419944727222167961682598265116876014855972048569400779697709765655340012215041774321114782240453575835030111362398780325388102665938958461476750392428688437146705789315316901483635835261598913055843;
            6'd17: xpb[0] = 1024'd78477632846943249568644566625795661277798613184264754573146858122010000598097039415682405329143928932406350178833844650301893889655794553054563320479115132013477998553004033594011992624770662719257667584151341757503901194520346433897037206796556249373280999699157677356546507179867984771352501764597542708728;
            6'd18: xpb[0] = 1024'd10113554964925357543977230895069269150199456827024043590313229149788885728979724728360740222236116334640165243790251138802555976787770506437090501085927174523864542838727084195053733842982345396090355319461867833613330176421015769440993177970924588002991703555509859536280696970490435041950478440970577877282;
            6'd19: xpb[0] = 1024'd65816172767032206918108822569157309767298727595519016735611455242544666197171548951054146329985978046317129716204151061882281904760966794374777806709070257967941761694021352133725714252711233794233240663159633756087120008542581877949927718828522375899522310825979099746121414835041518329667144943969207530167;
            6'd20: xpb[0] = 1024'd121518790569139056292240414243245350384397998364013989880909681335300446665363373173747552437735839757994094188618050984962007832734163082312465112332213341412018980549315620072397694662440122192376126006857399678560909840664147986458862259686120163796052918096448339955962132699592601617383811446967837183052;
            6'd21: xpb[0] = 1024'd53154712687121164267573078512518958256798842006773278898076052363079331796246058486425887330828027160227909253574457473462669919866139035694992292939025383922405524835038670673439435880651804869208813742167925754670338822564817322002818230860488502425763621952800522135696322490215051887981788123340872351606;
            6'd22: xpb[0] = 1024'd108857330489228013641704670186606998873898112775268252043374278455835112264437882709119293438577888871904873725988357396542395847839335323632679598562168467366482743690332938612111416290380693267351699085865691677144128654686383430511752771718086290322294229223269762345537040354766135175698454626339502004491;
            6'd23: xpb[0] = 1024'd40493252607210121617037334455880606746298956418027541060540649483613997395320568021797628331670076274138688790944763885043057934971311277015206779168980509876869287976055989213153157508592375944184386821176217753253557636587052766055708742892454628952004933079621944525271230145388585446296431302712537173045;
            6'd24: xpb[0] = 1024'd96195870409316970991168926129968647363398227186522514205838875576369777863512392244491034439419937985815653263358663808122783862944507564952894084792123593320946506831350257151825137918321264342327272164873983675727347468708618874564643283750052416848535540350091184735111948009939668734013097805711166825930;
            6'd25: xpb[0] = 1024'd27831792527299078966501590399242255235799070829281803223005246604148662994395077557169369332512125388049468328315070296623445950076483518335421265398935635831333051117073307752866879136532947019159959900184509751836776450609288210108599254924420755478246244206443366914846137800562119004611074482084201994484;
            6'd26: xpb[0] = 1024'd83534410329405928340633182073330295852898341597776776368303472696904443462586901779862775440261987099726432800728970219703171878049679806273108571022078719275410269972367575691538859546261835417302845243882275674310566282730854318617533795782018543374776851476912607124686855665113202292327740985082831647369;
            6'd27: xpb[0] = 1024'd15170332447388036315965846342603903725299185240536065385469843724683328593469587092541110333354174501960247865685376708203833965181655759655635751628890761785796814258090626292580600764473518094135532979192801750419995264631523654161489766956386882004487555333264789304421045455735652562925717661455866815923;
            6'd28: xpb[0] = 1024'd70872950249494885690097438016691944342398456009031038530768069817439109061661411315234516441104036213637212338099276631283559893154852047593323057252033845229874033113384894231252581174202406492278418322890567672893785096753089762670424307813984669901018162603734029514261763320286735850642384164454496468808;
            6'd29: xpb[0] = 1024'd2508872367476993665430102285965552214799299651790327547934440845217994192544096627912851334196223615871027403055683119784221980286828000975850237858845887740260577399107944832294322392414089169111106058201093749003214078653759098214380278988353008530728866460086211693995953110909186121240360840827531637362;
            6'd30: xpb[0] = 1024'd58211490169583843039561693960053592831898570420285300693232666937973774660735920850606257441946085327547991875469583042863947908260024288913537543481988971184337796254402212770966302802142977567253991401898859671477003910775325206723314819845950796427259473730555451903836670975460269408957027343826161290247;
            6'd31: xpb[0] = 1024'd113914107971690692413693285634141633448997841188780273838530893030729555128927745073299663549695947039224956347883482965943673836233220576851224849105132054628415015109696480709638283211871865965396876745596625593950793742896891315232249360703548584323790081001024692113677388840011352696673693846824790943132;
            6'd32: xpb[0] = 1024'd45550030089672800389025949903415241321398684831539562855697264058508440259810430385977998442788134441458771412839889454444335923365196530233752029711944097138801559395419531310680024430083548642229564480907151670060222724797560650776205331877916922953500784857376874293411578630633802967271670523197826111686;
            6'd33: xpb[0] = 1024'd101252647891779649763157541577503281938497955600034536000995490151264220728002254608671404550537996153135735885253789377524061851338392818171439335335087180582878778250713799249352004839812437040372449824604917592534012556919126759285139872735514710850031392127846114503252296495184886254988337026196455764571;
            6'd34: xpb[0] = 1024'd32888570009761757738490205846776889810898799242793825018161861179043105858884939921349739443630183555369550950210195866024723938470368771553966515941899223093265322536436849850393746058024119717205137559915443668643441538819796094829095843909883049479742095984198296682986486285807336525586313702569490933125;
            6'd35: xpb[0] = 1024'd88591187811868607112621797520864930427998070011288798163460087271798886327076764144043145551380045267046515422624095789104449866443565059491653821565042306537342541391731117789065726467753008115348022903613209591117231370941362203338030384767480837376272703254667536892827204150358419813302980205568120586010;
            6'd36: xpb[0] = 1024'd20227109929850715087954461790138538300398913654048087180626458299577771457959449456721480444472232669280330487580502277605111953575541012874181002171854349047729085677454168390107467685964690792180710638923735667226660352842031538881986355941849176005983407111019719072561393940980870083900956881941155754564;
            6'd37: xpb[0] = 1024'd75929727731957564462086053464226578917498184422543060325924684392333551926151273679414886552222094380957294959994402200684837881548737300811868307794997432491806304532748436328779448095693579190323595982621501589700450184963597647390920896799446963902514014381488959282402111805531953371617623384939785407449;
            6'd38: xpb[0] = 1024'd7565649849939672437418717733500186789899028065302349343091055420112437057033958992093221445314281783191110024950808689185499968680713254194395488401809475002192848818471486929821189313905261867156283717932027665809879166864266982934876867973815302532224718237841141462136301596154403642215600061312820576003;
            6'd39: xpb[0] = 1024'd63268267652046521811550309407588227406998298833797322488389281512868217525225783214786627553064143494868074497364708612265225896653909542132082794024952558446270067673765754868493169723634150265299169061629793588283668998985833091443811408831413090428755325508310381671977019460705486929932266564311450228888;
            6'd40: xpb[0] = 1024'd118970885454153371185681901081676268024097569602292295633687507605623997993417607437480033660814005206545038969778608535344951824627105830069770099648095641890347286529060022807165150133363038663442054405327559510757458831107399199952745949689010878325285932778779621881817737325256570217648933067310079881773;
            6'd41: xpb[0] = 1024'd50606807572135479161014565350949875896498413245051584650853878633402883124300292750158368553906192608778854034735015023845613911759081783452297280254907684400733830814783073408206891351574721340274742140638085586866887813008068535496701920863379216954996636635131804061551927115879020488246909743683115050327;
            6'd42: xpb[0] = 1024'd106309425374242328535146157025037916513597684013546557796152104726158663592492116972851774661656054320455818507148914946925339839732278071389984585878050767844811049670077341346878871761303609738417627484335851509340677645129634644005636461720977004851527243905601044271392644980430103775963576246681744703212;
            6'd43: xpb[0] = 1024'd37945347492224436510478821294311524385998527656305846813318475753937548723374802285530109554748241722689633572105321435426001926864254024772511766484862810355197593955800391947920612979515292415250315219646377585450106627030303979549592432895345343481237947761953226451126834771052554046561552923054779871766;
            6'd44: xpb[0] = 1024'd93647965294331285884610412968399565003097798424800819958616701846693329191566626508223515662498103434366598044519221358505727854837450312710199072108005893799274812811094659886592593389244180813393200563344143507923896459151870088058526973752943131377768555032422466660967552635603637334278219426053409524651;
            6'd45: xpb[0] = 1024'd25283887412313393859943077237673172875498642067560108975783072874472214322449311820901850555590290836600413109475627847006389941969426266092726252714817936309661357096817710487634334607455863490225888298654669584033325441052539423602482944927311470007479258888774648840701742426226087604876196102426444693205;
            6'd46: xpb[0] = 1024'd80986505214420243234074668911761213492597912836055082121081298967227994790641136043595256663340152548277377581889527770086115869942622554030413558337961019753738575952111978426306315017184751888368773642352435506507115273174105532111417485784909257904009866159243889050542460290777170892592862605425074346090;
            6'd47: xpb[0] = 1024'd12622427332402351209407333181034821364998756478814371138247669995006879921523821356273591556432339950511192646845934258586777957074598507412940738944773062264125120237835029027348056235396434565201461377662961582616544255074774867655373456959277596533720570015596071230276650081399621163190839281798109514644;
            6'd48: xpb[0] = 1024'd68325045134509200583538924855122861982098027247309344283545896087762660389715645578966997664182201662188157119259834181666503885047794795350628044567916145708202339093129296966020036645125322963344346721360727505090334087196340976164307997816875384430251177286065311440117367945950704450907505784796739167529;
            6'd49: xpb[0] = 1024'd124027662936616049957670516529210902599197298015804317428844122180518440857907469801660403771932063373865121591673734104746229813020991083288315350191059229152279557948423564904692017054854211361487232065058493427564123919317907084673242538674473172326781784556534551649958085810501787738624172287795368820414;
            6'd50: xpb[0] = 1024'd55663585054598157933003180798484510471598141658563606446010493208297325988790155114338738665024250776098936656630140593246891900152967036670842530797871271662666102234146615505733758273065894038319919800369019503673552901218576420217198509848841510956492488412886733829692275601124238009222148964168403988968;
            6'd51: xpb[0] = 1024'd111366202856705007307134772472572551088697412427058579591308719301053106456981979337032144772774112487775901129044040516326617828126163324608529836421014355106743321089440883444405738682794782436462805144066785426147342733340142528726133050706439298853023095683355974039532993465675321296938815467167033641853;
            6'd52: xpb[0] = 1024'd43002124974687115282467436741846158961098256069817868608475090328831991587864664649710479665866299890009716194000447004827279915258139277991057017027826397617129865375163934045447479901006465113295492879377311502256771715240811864270089021880807637482733799539708156219267183256297771567536792143540068810407;
            6'd53: xpb[0] = 1024'd98704742776793964656599028415934199578197526838312841753773316421587772056056488872403885773616161601686680666414346927907005843231335565928744322650969481061207084230458201984119460310735353511438378223075077424730561547362377972779023562738405425379264406810177396429107901120848854855253458646538698463292;
            6'd54: xpb[0] = 1024'd30340664894776072631931692685207807450598370481072130770939687449366657186939174185082220666708349003920495731370753416407667930363311519311271503257781523571593628516181252585161201528947036188271065958385603500839990529263047308322979533912773764008975110666529578608842090911471305125851435322911733631846;
            6'd55: xpb[0] = 1024'd86043282696882922006063284359295848067697641249567103916237913542122437655130998407775626774458210715597460203784653339487393858336507807248958808880924607015670847371475520523833181938675924586413951302083369423313780361384613416831914074770371551905505717936998818818682808776022388413568101825910363284731;
            6'd56: xpb[0] = 1024'd17679204814865029981395948628569455940098484892326392933404284569901322786013683720453961667550398117831275268741059827988055945468483760631485989487736649526057391657198571124874923156887607263246639037393895499423209343285282752375870045944739890535216421793351000998416998566644838684166078502283398453285;
            6'd57: xpb[0] = 1024'd73381822616971879355527540302657496557197755660821366078702510662657103254205507943147367775300259829508239741154959751067781873441680048569173295110879732970134610512492839063546903566616495661389524381091661421896999175406848860884804586802337678431747029063820241208257716431195921971882745005282028106170;
            6'd58: xpb[0] = 1024'd5017744734953987330860204571931104429598599303580655095868881690435988385088193255825702668392447231742054806111366239568443960573656001951700475717691775480521154798215889664588644784828178338222212116402187498006428157307518196428760557976706017061457732920172423387991906221818372242480721681655063274724;
            6'd59: xpb[0] = 1024'd60720362537060836704991796246019145046697870072075628241167107783191768853280017478519108776142308943419019278525266162648169888546852289889387781340834858924598373653510157603260625194557066736365097460099953420480217989429084304937695098834303804957988340190641663597832624086369455530197388184653692927609;
            6'd60: xpb[0] = 1024'd116422980339167686079123387920107185663797140840570601386465333875947549321471841701212514883892170655095983750939166085727895816520048577827075086963977942368675592508804425541932605604285955134507982803797719342954007821550650413446629639691901592854518947461110903807673341950920538817914054687652322580494;
            6'd61: xpb[0] = 1024'd48058902457149794054456052189380793536197984483329890403631704903726434452354527013890849776984358057329798815895572574228557903652024531209602267570789984879062136794527476142974346822497637811340670539108245419063436803451319748990585610866269931484229651317463085987407531741542989088512031364025357749048;
            6'd62: xpb[0] = 1024'd103761520259256643428587643863468834153297255251824863548929930996482214920546351236584255884734219769006763288309472497308283831625220819147289573193933068323139355649821744081646327232226526209483555882806011341537226635572885857499520151723867719380760258587932326197248249606094072376228697867023987401933;
            6'd63: xpb[0] = 1024'd35397442377238751403920308132742442025698098894584152566096302024261100051429036549262590777826407171240578353265878985808945918757196772529816753800745110833525899935544794682688068450438208886316243618116537417646655617473555193043476122898236058010470962444284508376982439396716522646826674543397022570487;
        endcase
    end

    always_comb begin
        case(flag[0][11:6])
            6'd0: xpb[1] = 1024'd0;
            6'd1: xpb[1] = 1024'd91100060179345600778051899806830482642797369663079125711394528117016880519620860771955996885576268882917542825679778908888671846730393060467504059423888194277603118790839062621360048860167097284459128961814303340120445449595121301552410663755833845907001569714753748586823157261267605934543341046395652223372;
            6'd2: xpb[1] = 1024'd58133424674566460157304872208846532540896312200422567294657201169056865701932582633896922556494863456391936243902064383198279852619565786379847993831445347621515563012106907905089858528816988847608060315241366833876530048969345830139842757828438242547183236015390439143539786448606578851967992266165709962413;
            6'd3: xpb[1] = 1024'd25166789169787319536557844610862582438995254737766008877919874221096850884244304495837848227413458029866329662124349857507887858508738512292191928239002500965428007233374753188819668197466880410756991668668430327632614648343570358727274851901042639187364902316027129700256415635945551769392643485935767701454;
            6'd4: xpb[1] = 1024'd116266849349132920314609744417693065081792624400845134589314402338113731403865165267793845112989726912783872487804128766396559705239131572759695987662890695243031126024213815810179717057633977695216120630482733667753060097938691660279685515656876485094366472030780878287079572897213157703935984532331419924826;
            6'd5: xpb[1] = 1024'd83300213844353779693862716819709114979891566938188576172577075390153716586176887129734770783908321486258265906026414240706167711128304298672039922070447848586943570245481661093909526726283869258365051983909797161509144697312916188867117609729480881734548138331417568843796202084552130621360635752101477663867;
            6'd6: xpb[1] = 1024'd50333578339574639073115689221725164877990509475532017755839748442193701768488608991675696454826916059732659324248699715015775717017477024584383856478005001930856014466749506377639336394933760821513983337336860655265229296687140717454549703802085278374729804632054259400512831271891103538785286971871535402908;
            6'd7: xpb[1] = 1024'd17366942834795498452368661623741214776089452012875459339102421494233686950800330853616622125745510633207052742470985189325383722906649750496727790885562155274768458688017351661369146063583652384662914690763924149021313896061365246041981797874689675014911470932690949957229460459230076456209938191641593141949;
            6'd8: xpb[1] = 1024'd108467003014141099230420561430571697418886821675954585050496949611250567470421191625572619011321779516124595568150764098214055569637042810964231850309450349552371577478856414282729194923750749669122043652578227489141759345656486547594392461630523520921913040647444698544052617720497682390753279238037245365321;
            6'd9: xpb[1] = 1024'd75500367509361958609673533832587747316985764213298026633759622663290552652732913487513544682240374089598988986373049572523663575526215536876575784717007502896284021700124259566459004592400641232270975006005290982897843945030711076181824555703127917562094706948081389100769246907836655308177930457807303104362;
            6'd10: xpb[1] = 1024'd42533732004582817988926506234603797215084706750641468217022295715330537835044635349454470353158968663073382404595335046833271581415388262788919719124564656240196465921392104850188814261050532795419906359432354476653928544404935604769256649775732314202276373248718079657485876095175628225602581677577360843403;
            6'd11: xpb[1] = 1024'd9567096499803677368179478636619847113183649287984909800284968767370523017356357211395396024077563236547775822817620521142879587304560988701263653532121809584108910142659950133918623929700424358568837712859417970410013143779160133356688743848336710842458039549354770214202505282514601143027232897347418582444;
            6'd12: xpb[1] = 1024'd100667156679149278146231378443450329755981018951064035511679496884387403536977217983351392909653832119465318648497399430031551434034954049168767712956010003861712028933499012755278672789867521643027966674673721310530458593374281434909099407604170556749459609264108518801025662543782207077570573943743070805816;
            6'd13: xpb[1] = 1024'd67700521174370137525484350845466379654079961488407477094942169936427388719288939845292318580572426692939712066719684904341159439924126775081111647363567157205624473154766858039008482458517413206176898028100784804286543192748505963496531501676774953389641275564745209357742291731121179994995225163513128544857;
            6'd14: xpb[1] = 1024'd34733885669590996904737323247482429552178904025750918678204842988467373901600661707233244251491021266414105484941970378650767445813299500993455581771124310549536917376034703322738292127167304769325829381527848298042627792122730492083963595749379350029822941865381899914458920918460152912419876383283186283898;
            6'd15: xpb[1] = 1024'd1767250164811856283990295649498479450277846563094360261467516040507359083912383569174169922409615839888498903164255852960375451702472226905799516178681463893449361597302548606468101795817196332474760734954911791798712391496955020671395689821983746670004608166018590471175550105799125829844527603053244022939;
            6'd16: xpb[1] = 1024'd92867310344157457062042195456328962093075216226173485972862044157524239603533244341130166807985884722806041728844034761849047298432865287373303575602569658171052480388141611227828150655984293616933889696769215131919157841092076322223806353577817592577006177880772339057998707367066731764387868649448896246311;
            6'd17: xpb[1] = 1024'd59900674839378316441295167858345011991174158763516927556124717209564224785844966203071092478904479296280435147066320236158655304322038013285647510010126811514964924609409456511557960324634185180082821050196278625675242440466300850811238447650421989217187844181409029614715336554405704681812519869218953985352;
            6'd18: xpb[1] = 1024'd26934039334599175820548140260361061889273101300860369139387390261604209968156688065012018149823073869754828565288605710468263310211210739197991444417683964858877368830677301795287769993284076743231752403623342119431327039840525379398670541723026385857369510482045720171431965741744677599237171088989011724393;
            6'd19: xpb[1] = 1024'd118034099513944776598600040067191544532070470963939494850781918378621090487777548836968015035399342752672371390968384619356935156941603799665495503841572159136480487621516364416647818853451174027690881365437645459551772489435646680951081205478860231764371080196799468758255123003012283533780512135384663947765;
            6'd20: xpb[1] = 1024'd85067464009165635977853012469207594430169413501282936434044591430661075670089270698908940706317937326146764809190670093666543162830776525577839438249129312480392931842784209700377628522101065590839812718864708953307857088809871209538513299551464628404552746497436159314971752190351256451205163355154721686806;
            6'd21: xpb[1] = 1024'd52100828504386495357105984871223644328268356038626378017307264482701060852400992560849866377236531899621158227412955567976151168719949251490183372656686465824305376064052054984107438190750957153988744072291772447063941688184095738125945393624069025044734412798072849871688381377690229368629814574924779425847;
            6'd22: xpb[1] = 1024'd19134192999607354736358957273239694226367298575969819600569937534741046034712714422790792048155126473095551645635241042285759174609121977402527307064243619168217820285319900267837247859400848717137675425718835940820026287558320266713377487696673421684916079098709540428405010565029202286054465794694837164888;
            6'd23: xpb[1] = 1024'd110234253178952955514410857080070176869164668239048945311964465651757926554333575194746788933731395356013094471315019951174431021339515037870031366488131813445820939076158962889197296719567946001596804387533139280940471737153441568265788151452507267591917648813463289015228167826296808220597806841090489388260;
            6'd24: xpb[1] = 1024'd77267617674173814893663829482086226767263610776392386895227138703797911736645297056687714604649989929487487889537305425484039027228687763782375300895688966789733383297426808172927106388217837564745735740960202774696556336527666096853220245525111664232099315114099979571944797013635781138022458060860547127301;
            6'd25: xpb[1] = 1024'd44300982169394674272916801884102276665362553313735828478489811755837896918957018918628640275568584502961881307759590899793647033117860489694719235303246120133645827518694653456656916056867729127894667094387266268452640935901890625440652339597716060872280981414736670128661426200974754055447109280630604866342;
            6'd26: xpb[1] = 1024'd11334346664615533652169774286118326563461495851079270061752484807877882101268740780569565946487179076436274725981876374103255039007033215607063169710803273477558271739962498740386725725517620691043598447814329762208725535276115154028084433670320457512462647715373360685378055388313726972871760500400662605383;
            6'd27: xpb[1] = 1024'd102434406843961134430221674092948809206258865514158395773147012924894762620889601552525562832063447959353817551661655282991926885737426276074567229134691467755161390530801561361746774585684717975502727409628633102329170984871236455580495097426154303419464217430127109272201212649581332907415101546796314828755;
            6'd28: xpb[1] = 1024'd69467771339181993809474646494964859104357808051501837356409685976934747803201323414466488502982042532828210969883940757301534891626599001986911163542248621099073834752069406645476584254334609538651658763055696596085255584245460984167927191498758700059645883730763799828917841836920305824839752766566372567796;
            6'd29: xpb[1] = 1024'd36501135834402853188727618896980909002456750588845278939672359028974732985513045276407414173900637106302604388106226231611142897515771727899255097949805774442986278973337251929206393922984501101800590116482760089841340183619685512755359285571363096699827550031400490385634471024259278742264403986336430306837;
            6'd30: xpb[1] = 1024'd3534500329623712567980591298996958900555693126188720522935032081014718167824767138348339844819231679776997806328511705920750903404944453811599032357362927786898723194605097212936203591634392664949521469909823583597424782993910041342791379643967493340009216332037180942351100211598251659689055206106488045878;
            6'd31: xpb[1] = 1024'd94634560508969313346032491105827441543353062789267846234329560198031598687445627910304336730395500562694540632008290614809422750135337514279103091781251122064501841985444159834296252451801489949408650431724126923717870232589031342895202043399801339247010786046790929529174257472865857594232396252502140269250;
            6'd32: xpb[1] = 1024'd61667925004190172725285463507843491441452005326611287817592233250071583869757349772245262401314095136168934050230576089119030756024510240191447026188808275408414286206712005118026062120451381512557581785151190417473954831963255871482634137472405735887192452347427620085890886660204830511657047472272198008291;
            6'd33: xpb[1] = 1024'd28701289499411032104538435909859541339550947863954729400854906302111569052069071634186188072232689709643327468452861563428638761913682966103790960596365428752326730427979850401755871789101273075706513138578253911230039431337480400070066231545010132527374118648064310642607515847543803429081698692042255747332;
            6'd34: xpb[1] = 1024'd119801349678756632882590335716690023982348317527033855112249434419128449571689932406142184957808958592560870294132640472317310608644076026571295020020253623029929849218818913023115920649268370360165642100392557251350484880932601701622476895300843978434375688362818059229430673108811409363625039738437907970704;
            6'd35: xpb[1] = 1024'd86834714173977492261843308118706073880447260064377296695512107471168434754001654268083110628727553166035263712354925946626918614533248752483638954427810776373842293440086758306845730317918261923314573453819620745106569480306826230209908989373448375074557354663454749786147302296150382281049690958207965709745;
            6'd36: xpb[1] = 1024'd53868078669198351641096280520722123778546202601720738278774780523208419936313376130024036299646147739509657130577211420936526620422421478395982888835367929717754737661354603590575539986568153486463504807246684238862654079681050758797341083446052771714739020964091440342863931483489355198474342177978023448786;
            6'd37: xpb[1] = 1024'd20901443164419211020349252922738173676645145139064179862037453575248405118625097991964961970564742312984050548799496895246134626311594204308326823242925083061667181882622448874305349655218045049612436160673747732618738679055275287384773177518657168354920687264728130899580560670828328115898993397748081187827;
            6'd38: xpb[1] = 1024'd112001503343764811798401152729568656319442514802143305573431981692265285638245958763920958856141011195901593374479275804134806473041987264775830882666813277339270300673461511495665398515385142334071565122488051072739184128650396588937183841274491014261922256979481879486403717932095934050442334444143733411199;
            6'd39: xpb[1] = 1024'd79034867838985671177654125131584706217541457339486747156694654744305270820557680625861884527059605769375986792701561278444414478931159990688174817074370430683182744894729356779395208184035033897220496475915114566495268728024621117524615935347095410902103923280118570043120347119434906967866985663913791150240;
            6'd40: xpb[1] = 1024'd46068232334206530556907097533600756115640399876830188739957327796345256002869402487802810197978200342850380210923846752754022484820332716600518751481927584027095189115997202063125017852684925460369427829342178060251353327398845646112048029419699807542285589580755260599836976306773879885291636883683848889281;
            6'd41: xpb[1] = 1024'd13101596829427389936160069935616806013739342414173630323220000848385241185181124349743735868896794916324773629146132227063630490709505442512862685889484737371007633337265047346854827521334817023518359182769241554007437926773070174699480123492304204182467255881391951156553605494112852802716288103453906628322;
            6'd42: xpb[1] = 1024'd104201657008772990714211969742447288656536712077252756034614528965402121704801985121699732754473063799242316454825911135952302337439898502980366745313372931648610752128104109968214876381501914307977488144583544894127883376368191476251890787248138050089468825596145699743376762755380458737259629149849558851694;
            6'd43: xpb[1] = 1024'd71235021503993850093464942144463338554635654614596197617877202017442106887113706983640658425391658372716709873048196610261910343329071228892710679720930084992523196349371955251944686050151805871126419498010608387883967975742416004839322881320742446729650491896782390300093391942719431654684280369619616590735;
            6'd44: xpb[1] = 1024'd38268385999214709472717914546479388452734597151939639201139875069482092069425428845581584096310252946191103291270482084571518349218243954805054614128487238336435640570639800535674495718801697434275350851437671881640052575116640533426754975393346843369832158197419080856810021130058404572108931589389674329776;
            6'd45: xpb[1] = 1024'd5301750494435568851970886948495438350833539689283080784402548121522077251737150707522509767228847519665496709492767558881126355107416680717398548536044391680348084791907645819404305387451588997424282204864735375396137174490865062014187069465951240010013824498055771413526650317397377489533582809159732068817;
            6'd46: xpb[1] = 1024'd96401810673781169630022786755325920993630909352362206495797076238538957771358011479478506652805116402583039535172546467769798201837809741184902607959932585957951203582746708440764354247618686281883411166679038715516582624085986363566597733221785085917015394212809520000349807578664983424076923855555384292189;
            6'd47: xpb[1] = 1024'd63435175169002029009275759157341970891729851889705648079059749290578942953669733341419432323723710976057432953394831942079406207726982467097246542367489739301863647804014553724494163916268577845032342520106102209272667223460210892154029827294389482557197060513446210557066436766003956341501575075325442031230;
            6'd48: xpb[1] = 1024'd30468539664222888388528731559358020789828794427049089662322422342618928135981455203360357994642305549531826371617117416389014213616155193009590476775046892645776092025282399008223973584918469408181273873533165703028751822834435420741461921366993879197378726814082901113783065953342929258926226295095499770271;
            6'd49: xpb[1] = 1024'd121568599843568489166580631366188503432626164090128215373716950459635808655602315975316354880218574432449369197296896325277686060346548253477094536198935086923379210816121461629584022445085566692640402835347469043149197272429556722293872585122827725104380296528836649700606223214610535193469567341491151993643;
            6'd50: xpb[1] = 1024'd88601964338789348545833603768204553330725106627471656956979623511675793837914037837257280551137169005923762615519181799587294066235720979389438470606492240267291655037389306913313832113735458255789334188774532536905281871803781250881304679195432121744561962829473340257322852401949508110894218561261209732684;
            6'd51: xpb[1] = 1024'd55635328834010207925086576170220603228824049164815098540242296563715779020225759699198206222055763579398156033741467273896902072124893705301782405014049393611204099258657152197043641782385349818938265542201596030661366471178005779468736773268036518384743629130110030814039481589288481028318869781031267471725;
            6'd52: xpb[1] = 1024'd22668693329231067304339548572236653126922991702158540123504969615755764202537481561139131892974358152872549451963752748206510078014066431214126339421606546955116543479924997480773451451035241382087196895628659524417451070552230308056168867340640915024925295430746721370756110776627453945743521000801325210766;
            6'd53: xpb[1] = 1024'd113768753508576668082391448379067135769720361365237665834899497732772644722158342333095128778550627035790092277643531657095181924744459491681630398845494741232719662270764060102133500311202338666546325857442962864537896520147351609608579531096474760931926865145500469957579268037895059880286862047196977434138;
            6'd54: xpb[1] = 1024'd80802118003797527461644420781083185667819303902581107418162170784812629904470064195036054449469221609264485695865817131404789930633632217593974333253051894576632106492031905385863309979852230229695257210870026358293981119521576138196011625169079157572108531446137160514295897225234032797711513266967035173179;
            6'd55: xpb[1] = 1024'd47835482499018386840897393183099235565918246439924549001424843836852615086781786056976980120387816182738879114088102605714397936522804943506318267660609047920544550713299750669593119648502121792844188564297089852050065718895800666783443719241683554212290197746773851071012526412573005715136164486737092912220;
            6'd56: xpb[1] = 1024'd14868846994239246220150365585115285464017188977267990584687516888892600269093507918917905791306410756213272532310388080024005942411977669418662202068166201264456994934567595953322929317152013355993119917724153345806150318270025195370875813314287950852471864047410541627729155599911978632560815706507150651261;
            6'd57: xpb[1] = 1024'd105968907173584846998202265391945768106814558640347116296082045005909480788714368690873902676882679639130815357990166988912677789142370729886166261492054395542060113725406658574682978177319110640452248879538456685926595767865146496923286477070121796759473433762164290214552312861179584567104156752902802874633;
            6'd58: xpb[1] = 1024'd73002271668805706377455237793961818004913501177690557879344718057949465971026090552814828347801274212605208776212452463222285795031543455798510195899611548885972557946674503858412787845969002203601180232965520179682680367239371025510718571142726193399655100062800980771268942048518557484528807972672860613674;
            6'd59: xpb[1] = 1024'd40035636164026565756708210195977867903012443715033999462607391109989451153337812414755754018719868786079602194434737937531893800920716181710854130307168702229885002167942349142142597514618893766750111586392583673438764966613595554098150665215330590039836766363437671327985571235857530401953459192442918352715;
            6'd60: xpb[1] = 1024'd7069000659247425135961182597993917801111386252377441045870064162029436335649534276696679689638463359553995612657023411841501806809888907623198064714725855573797446389210194425872407183268785329899042939819647167194849565987820082685582759287934986680018432664074361884702200423196503319378110412212976091756;
            6'd61: xpb[1] = 1024'd98169060838593025914013082404824400443908755915456566757264592279046316855270395048652676575214732242471538438336802320730173653540281968090702124138614049851400565180049257047232456043435882614358171901633950507315295015582941384237993423043768832587020002378828110471525357684464109253921451458608628315128;
            6'd62: xpb[1] = 1024'd65202425333813885293266054806840450342007698452800008340527265331086302037582116910593602246133326815945931856559087795039781659429454694003046058546171203195313009401317102330962265712085774177507103255061014001071379614957165912825425517116373229227201668679464801028241986871803082171346102678378686054169;
            6'd63: xpb[1] = 1024'd32235789829034744672519027208856500240106640990143449923789938383126287219893838772534527917051921389420325274781373269349389665318627419915389992953728356539225453622584947614692075380735665740656034608488077494827464214331390441412857611188977625867383334980101491584958616059142055088770753898148743793210;
        endcase
    end

    always_comb begin
        case(flag[0][16:12])
            5'd0: xpb[2] = 1024'd0;
            5'd1: xpb[2] = 1024'd123335850008380345450570927015686982882904010653222575635184466500143167739514699544490524802628190272337868100461152178238061512049020480382894052377616550816828572413424010236052124240902763025115163570302380834947909663926511742965268274944811471774384904694855240171781773320409661023314094944544396016582;
            5'd2: xpb[2] = 1024'd122605004332635949502342926626559533021109594180709467142237077935309440141720260178965978390598706235232586793464810921897059183256820626210627979738902060699966470257276803134474009290288320328920129532217521823531458477632126712965557980206393494281949905975593422313457018566890689029509500062463197548833;
            5'd3: xpb[2] = 1024'd121874158656891553554114926237432083159315177708196358649289689370475712543925820813441431978569222198127305486468469665556056854464620772038361907100187570583104368101129596032895894339673877632725095494132662812115007291337741682965847685467975516789514907256331604455132263813371717035704905180381999081084;
            5'd4: xpb[2] = 1024'd121143312981147157605886925848304633297520761235683250156342300805641984946131381447916885566539738161022024179472128409215054525672420917866095834461473080466242265944982388931317779389059434936530061456047803800698556105043356652966137390729557539297079908537069786596807509059852745041900310298300800613335;
            5'd5: xpb[2] = 1024'd120412467305402761657658925459177183435726344763170141663394912240808257348336942082392339154510254123916742872475787152874052196880221063693829761822758590349380163788835181829739664438444992240335027417962944789282104918748971622966427095991139561804644909817807968738482754306333773048095715416219602145586;
            5'd6: xpb[2] = 1024'd119681621629658365709430925070049733573931928290657033170447523675974529750542502716867792742480770086811461565479445896533049868088021209521563689184044100232518061632687974728161549487830549544139993379878085777865653732454586592966716801252721584312209911098546150880157999552814801054291120534138403677837;
            5'd7: xpb[2] = 1024'd118950775953913969761202924680922283712137511818143924677500135111140802152748063351343246330451286049706180258483104640192047539295821355349297616545329610115655959476540767626583434537216106847944959341793226766449202546160201562967006506514303606819774912379284333021833244799295829060486525652057205210088;
            5'd8: xpb[2] = 1024'd118219930278169573812974924291794833850343095345630816184552746546307074554953623985818699918421802012600898951486763383851045210503621501177031543906615119998793857320393560525005319586601664151749925303708367755032751359865816532967296211775885629327339913660022515163508490045776857066681930769976006742339;
            5'd9: xpb[2] = 1024'd117489084602425177864746923902667383988548678873117707691605357981473346957159184620294153506392317975495617644490422127510042881711421647004765471267900629881931755164246353423427204635987221455554891265623508743616300173571431502967585917037467651834904914940760697305183735292257885072877335887894808274590;
            5'd10: xpb[2] = 1024'd116758238926680781916518923513539934126754262400604599198657969416639619359364745254769607094362833938390336337494080871169040552919221792832499398629186139765069653008099146321849089685372778759359857227538649732199848987277046472967875622299049674342469916221498879446858980538738913079072741005813609806841;
            5'd11: xpb[2] = 1024'd116027393250936385968290923124412484264959845928091490705710580851805891761570305889245060682333349901285055030497739614828038224127021938660233325990471649648207550851951939220270974734758336063164823189453790720783397800982661442968165327560631696850034917502237061588534225785219941085268146123732411339092;
            5'd12: xpb[2] = 1024'd115296547575191990020062922735285034403165429455578382212763192286972164163775866523720514270303865864179773723501398358487035895334822084487967253351757159531345448695804732118692859784143893366969789151368931709366946614688276412968455032822213719357599918782975243730209471031700969091463551241651212871343;
            5'd13: xpb[2] = 1024'd114565701899447594071834922346157584541371012983065273719815803722138436565981427158195967858274381827074492416505057102146033566542622230315701180713042669414483346539657525017114744833529450670774755113284072697950495428393891382968744738083795741865164920063713425871884716278181997097658956359570014403594;
            5'd14: xpb[2] = 1024'd113834856223703198123606921957030134679576596510552165226868415157304708968186987792671421446244897789969211109508715845805031237750422376143435108074328179297621244383510317915536629882915007974579721075199213686534044242099506352969034443345377764372729921344451608013559961524663025103854361477488815935845;
            5'd15: xpb[2] = 1024'd113104010547958802175378921567902684817782180038039056733921026592470981370392548427146875034215413752863929802512374589464028908958222521971169035435613689180759142227363110813958514932300565278384687037114354675117593055805121322969324148606959786880294922625189790155235206771144053110049766595407617468096;
            5'd16: xpb[2] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            5'd17: xpb[2] = 1024'd111642319196470010278922920789647785094193347093012839748026249462803526174803669696097782210156445678653367188519692076782024251373822813626636890158184708947034937915068696610802285031071679885994618960944636652284690683216351262969903559130123831895424925186666154438585697264106109122440576831245220532598;
            5'd18: xpb[2] = 1024'd110911473520725614330694920400520335232398930620499731255078860897969798577009230330573235798126961641548085881523350820441021922581622959454370817519470218830172835758921489509224170080457237189799584922859777640868239496921966232970193264391705854402989926467404336580260942510587137128635981949164022064849;
            5'd19: xpb[2] = 1024'd110180627844981218382466920011392885370604514147986622762131472333136070979214790965048689386097477604442804574527009564100019593789423105282104744880755728713310733602774282407646055129842794493604550884774918629451788310627581202970482969653287876910554927748142518721936187757068165134831387067082823597100;
            5'd20: xpb[2] = 1024'd109449782169236822434238919622265435508810097675473514269184083768302343381420351599524142974067993567337523267530668307759017264997223251109838672242041238596448631446627075306067940179228351797409516846690059618035337124333196172970772674914869899418119929028880700863611433003549193141026792185001625129351;
            5'd21: xpb[2] = 1024'd108718936493492426486010919233137985647015681202960405776236695203468615783625912233999596562038509530232241960534327051418014936205023396937572599603326748479586529290479868204489825228613909101214482808605200606618885938038811142971062380176451921925684930309618883005286678250030221147222197302920426661602;
            5'd22: xpb[2] = 1024'd107988090817748030537782918844010535785221264730447297283289306638634888185831472868475050150009025493126960653537985795077012607412823542765306526964612258362724427134332661102911710277999466405019448770520341595202434751744426112971352085438033944433249931590357065146961923496511249153417602420839228193853;
            5'd23: xpb[2] = 1024'd107257245142003634589554918454883085923426848257934188790341918073801160588037033502950503737979541456021679346541644538736010278620623688593040454325897768245862324978185454001333595327385023708824414732435482583785983565450041082971641790699615966940814932871095247288637168742992277159613007538758029726104;
            5'd24: xpb[2] = 1024'd106526399466259238641326918065755636061632431785421080297394529508967432990242594137425957325950057418916398039545303282395007949828423834420774381687183278129000222822038246899755480376770581012629380694350623572369532379155656052971931495961197989448379934151833429430312413989473305165808412656676831258355;
            5'd25: xpb[2] = 1024'd105795553790514842693098917676628186199838015312907971804447140944133705392448154771901410913920573381811116732548962026054005621036223980248508309048468788012138120665891039798177365426156138316434346656265764560953081192861271022972221201222780011955944935432571611571987659235954333172003817774595632790606;
            5'd26: xpb[2] = 1024'd105064708114770446744870917287500736338043598840394863311499752379299977794653715406376864501891089344705835425552620769713003292244024126076242236409754297895276018509743832696599250475541695620239312618180905549536630006566885992972510906484362034463509936713309793713662904482435361178199222892514434322857;
            5'd27: xpb[2] = 1024'd104333862439026050796642916898373286476249182367881754818552363814466250196859276040852318089861605307600554118556279513372000963451824271903976163771039807778413916353596625595021135524927252924044278580096046538120178820272500962972800611745944056971074937994047975855338149728916389184394628010433235855108;
            5'd28: xpb[2] = 1024'd103603016763281654848414916509245836614454765895368646325604975249632522599064836675327771677832121270495272811559938257030998634659624417731710091132325317661551814197449418493443020574312810227849244542011187526703727633978115932973090317007526079478639939274786157997013394975397417190590033128352037387359;
            5'd29: xpb[2] = 1024'd102872171087537258900186916120118386752660349422855537832657586684798795001270397309803225265802637233389991504563597000689996305867424563559444018493610827544689712041302211391864905623698367531654210503926328515287276447683730902973380022269108101986204940555524340138688640221878445196785438246270838919610;
            5'd30: xpb[2] = 1024'd102141325411792862951958915730990936890865932950342429339710198119965067403475957944278678853773153196284710197567255744348993977075224709387177945854896337427827609885155004290286790673083924835459176465841469503870825261389345872973669727530690124493769941836262522280363885468359473202980843364189640451861;
            5'd31: xpb[2] = 1024'd101410479736048467003730915341863487029071516477829320846762809555131339805681518578754132441743669159179428890570914488007991648283024855214911873216181847310965507729007797188708675722469482139264142427756610492454374075094960842973959432792272147001334943117000704422039130714840501209176248482108441984112;
        endcase
    end

    always_comb begin
        case(flag[1][5:0])
            6'd0: xpb[3] = 1024'd0;
            6'd1: xpb[3] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            6'd2: xpb[3] = 1024'd100679634060304071055502914952736037167277100005316212353815420990297612207887079213229586029714185122074147583574573231666989319490825001042645800577467357194103405572860590087130560771855039443069108389671751481037922888800575812974249138053854169508899944397738886563714375961321529215371653600027243516363;
            6'd3: xpb[3] = 1024'd88986103248393735883854908726696839378566436445106476466657203952957970643176049364836843437242440528389646671633113130210952058815627334286388638358035515324309771074505276461880721562023956303948563780314007298374703908090415332978884422239166529629939964889549800830518299905017977314498135486728068032379;
            6'd4: xpb[3] = 1024'd77292572436483400712206902500657641589855772884896740579498986915618329078465019516444100844770695934705145759691653028754914798140429667530131476138603673454516136576149962836630882352192873164828019170956263115711484927380254852983519706424478889750979985381360715097322223848714425413624617373428892548395;
            6'd5: xpb[3] = 1024'd65599041624573065540558896274618443801145109324687004692340769878278687513753989668051358252298951341020644847750192927298877537465232000773874313919171831584722502077794649211381043142361790025707474561598518933048265946670094372988154990609791249872020005873171629364126147792410873512751099260129717064411;
            6'd6: xpb[3] = 1024'd53905510812662730368910890048579246012434445764477268805182552840939045949042959819658615659827206747336143935808732825842840276790034334017617151699739989714928867579439335586131203932530706886586929952240774750385046965959933892992790274795103609993060026364982543630930071736107321611877581146830541580427;
            6'd7: xpb[3] = 1024'd42211980000752395197262883822540048223723782204267532918024335803599404384331929971265873067355462153651643023867272724386803016114836667261359989480308147845135233081084021960881364722699623747466385342883030567721827985249773412997425558980415970114100046856793457897733995679803769711004063033531366096443;
            6'd8: xpb[3] = 1024'd30518449188842060025614877596500850435013118644057797030866118766259762819620900122873130474883717559967142111925812622930765755439639000505102827260876305975341598582728708335631525512868540608345840733525286385058609004539612933002060843165728330235140067348604372164537919623500217810130544920232190612459;
            6'd9: xpb[3] = 1024'd18824918376931724853966871370461652646302455083848061143707901728920121254909870274480387882411972966282641199984352521474728494764441333748845665041444464105547964084373394710381686303037457469225296124167542202395390023829452453006696127351040690356180087840415286431341843567196665909257026806933015128475;
            6'd10: xpb[3] = 1024'd7131387565021389682318865144422454857591791523638325256549684691580479690198840426087645289940228372598140288042892420018691234089243666992588502822012622235754329586018081085131847093206374330104751514809798019732171043119291973011331411536353050477220108332226200698145767510893114008383508693633839644491;
            6'd11: xpb[3] = 1024'd119504552437235795909469786323197689813579555089164273497523322719217733462796949487709973912126158088356788783558925753141717814255266334791491465618911821299651369657233984797512247074892496912294404513839293683433312912630028265980945265404894859865080032238154172995056219528518195124628680406960258644838;
            6'd12: xpb[3] = 1024'd107811021625325460737821780097158492024868891528954537610365105681878091898085919639317231319654413494672287871617465651685680553580068668035234303399479979429857735158878671172262407865061413773173859904481549500770093931919867785985580549590207219986120052729965087261860143472214643223755162293661083160854;
            6'd13: xpb[3] = 1024'd96117490813415125566173773871119294236158227968744801723206888644538450333374889790924488727182668900987786959676005550229643292904871001278977141180048137560064100660523357547012568655230330634053315295123805318106874951209707305990215833775519580107160073221776001528664067415911091322881644180361907676870;
            6'd14: xpb[3] = 1024'd84423960001504790394525767645080096447447564408535065836048671607198808768663859942531746134710924307303286047734545448773606032229673334522719978960616295690270466162168043921762729445399247494932770685766061135443655970499546825994851117960831940228200093713586915795467991359607539422008126067062732192886;
            6'd15: xpb[3] = 1024'd72730429189594455222877761419040898658736900848325329948890454569859167203952830094139003542239179713618785135793085347317568771554475667766462816741184453820476831663812730296512890235568164355812226076408316952780436989789386345999486402146144300349240114205397830062271915303303987521134607953763556708902;
            6'd16: xpb[3] = 1024'd61036898377684120051229755193001700870026237288115594061732237532519525639241800245746260949767435119934284223851625245861531510879278001010205654521752611950683197165457416671263051025737081216691681467050572770117218009079225866004121686331456660470280134697208744329075839247000435620261089840464381224918;
            6'd17: xpb[3] = 1024'd49343367565773784879581748966962503081315573727905858174574020495179884074530770397353518357295690526249783311910165144405494250204080334253948492302320770080889562667102103046013211815905998077571136857692828587453999028369065386008756970516769020591320155189019658595879763190696883719387571727165205740934;
            6'd18: xpb[3] = 1024'd37649836753863449707933742740923305292604910167696122287415803457840242509819740548960775764823945932565282399968705042949456989528882667497691330082888928211095928168746789420763372606074914938450592248335084404790780047658904906013392254702081380712360175680830572862683687134393331818514053613866030256950;
            6'd19: xpb[3] = 1024'd25956305941953114536285736514884107503894246607486386400257586420500600945108710700568033172352201338880781488027244941493419728853685000741434167863457086341302293670391475795513533396243831799330047638977340222127561066948744426018027538887393740833400196172641487129487611078089779917640535500566854772966;
            6'd20: xpb[3] = 1024'd14262775130042779364637730288844909715183583047276650513099369383160959380397680852175290579880456745196280576085784840037382468178487333985177005644025244471508659172036162170263694186412748660209503029619596039464342086238583946022662823072706100954440216664452401396291535021786228016767017387267679288982;
            6'd21: xpb[3] = 1024'd2569244318132444192989724062805711926472919487066914625941152345821317815686651003782547987408712151511779664144324738581345207503289667228919843424593402601715024673680848545013854976581665521088958420261851856801123105528423466027298107258018461075480237156263315663095458965482676115893499273968503804998;
            6'd22: xpb[3] = 1024'd114942409190346850420140645241580946882460683052592862866914790373458571588284760065404876609594641867270428159660358071704371787669312335027822806221492601665612064744896752257394254958267788103278611419291347520502264975039159758996911961126560270463340161062191287960005910983107757232138670987294922805345;
            6'd23: xpb[3] = 1024'd103248878378436515248492639015541749093750019492383126979756573336118930023573730217012134017122897273585927247718897970248334526994114668271565644002060759795818430246541438632144415748436704964158066809933603337839045994328999279001547245311872630584380181554002202226809834926804205331265152873995747321361;
            6'd24: xpb[3] = 1024'd91555347566526180076844632789502551305039355932173391092598356298779288458862700368619391424651152679901426335777437868792297266318917001515308481782628917926024795748186125006894576538605621825037522200575859155175827013618838799006182529497184990705420202045813116493613758870500653430391634760696571837377;
            6'd25: xpb[3] = 1024'd79861816754615844905196626563463353516328692371963655205440139261439646894151670520226648832179408086216925423835977767336260005643719334759051319563197076056231161249830811381644737328774538685916977591218114972512608032908678319010817813682497350826460222537624030760417682814197101529518116647397396353393;
            6'd26: xpb[3] = 1024'd68168285942705509733548620337424155727618028811753919318281922224100005329440640671833906239707663492532424511894517665880222744968521668002794157343765234186437526751475497756394898118943455546796432981860370789849389052198517839015453097867809710947500243029434945027221606757893549628644598534098220869409;
            6'd27: xpb[3] = 1024'd56474755130795174561900614111384957938907365251544183431123705186760363764729610823441163647235918898847923599953057564424185484293324001246536995124333392316643892253120184131145058909112372407675888372502626607186170071488357359020088382053122071068540263521245859294025530701589997727771080420799045385425;
            6'd28: xpb[3] = 1024'd44781224318884839390252607885345760150196701691334447543965488149420722200018580975048421054764174305163422688011597462968148223618126334490279832904901550446850257754764870505895219699281289268555343763144882424522951090778196879024723666238434431189580284013056773560829454645286445826897562307499869901441;
            6'd29: xpb[3] = 1024'd33087693506974504218604601659306562361486038131124711656807271112081080635307551126655678462292429711478921776070137361512110962942928667734022670685469708577056623256409556880645380489450206129434799153787138241859732110068036399029358950423746791310620304504867687827633378588982893926024044194200694417457;
            6'd30: xpb[3] = 1024'd21394162695064169046956595433267364572775374570914975769649054074741439070596521278262935869820685117794420864128677260056073702267731000977765508466037866707262988758054243255395541279619122990314254544429394059196513129357875919033994234609059151431660324996678602094437302532679342025150526080901518933473;
            6'd31: xpb[3] = 1024'd9700631883153833875308589207228166784064711010705239882490837037401797505885491429870193277348940524109919952187217158600036441592533334221508346246606024837469354259698929630145702069788039851193709935071649876533294148647715439038629518794371511552700345488489516361241226476375790124277007967602343449489;
            6'd32: xpb[3] = 1024'd122073796755368240102459510386003401740052474576231188123464475065039051278483600491492521899534870239868568447703250491723063021758556002020411309043505223901366394330914833342526102051474162433383362934101145540234436018158451732008243372662913320940560269394417488658151678494000871240522179680928762449836;
            6'd33: xpb[3] = 1024'd110380265943457904930811504159964203951341811016021452236306258027699409713772570643099779307063125646184067535761790390267025761083358335264154146824073382031572759832559519717276262841643079294262818324743401357571217037448291252012878656848225681061600289886228402924955602437697319339648661567629586965852;
            6'd34: xpb[3] = 1024'd98686735131547569759163497933925006162631147455811716349148040990359768149061540794707036714591381052499566623820330288810988500408160668507896984604641540161779125334204206092026423631811996155142273715385657174907998056738130772017513941033538041182640310378039317191759526381393767438775143454330411481868;
            6'd35: xpb[3] = 1024'd86993204319637234587515491707885808373920483895601980461989823953020126584350510946314294122119636458815065711878870187354951239732963001751639822385209698291985490835848892466776584421980913016021729106027912992244779076027970292022149225218850401303680330869850231458563450325090215537901625341031235997884;
            6'd36: xpb[3] = 1024'd75299673507726899415867485481846610585209820335392244574831606915680485019639481097921551529647891865130564799937410085898913979057765334995382660165777856422191856337493578841526745212149829876901184496670168809581560095317809812026784509404162761424720351361661145725367374268786663637028107227732060513900;
            6'd37: xpb[3] = 1024'd63606142695816564244219479255807412796499156775182508687673389878340843454928451249528808937176147271446063887995949984442876718382567668239125497946346014552398221839138265216276906002318746737780639887312424626918341114607649332031419793589475121545760371853472059992171298212483111736154589114432885029916;
            6'd38: xpb[3] = 1024'd51912611883906229072571473029768215007788493214972772800515172841001201890217421401136066344704402677761562976054489882986839457707370001482868335726914172682604587340782951591027066792487663598660095277954680444255122133897488852036055077774787481666800392345282974258975222156179559835281071001133709545932;
            6'd39: xpb[3] = 1024'd40219081071995893900923466803729017219077829654763036913356955803661560325506391552743323752232658084077062064113029781530802197032172334726611173507482330812810952842427637965777227582656580459539550668596936261591903153187328372040690361960099841787840412837093888525779146099876007934407552887834534061948;
            6'd40: xpb[3] = 1024'd28525550260085558729275460577689819430367166094553301026198738766321918760795361704350581159760913490392561152171569680074764936356974667970354011288050488943017318344072324340527388372825497320419006059239192078928684172477167892045325646145412201908880433328904802792583070043572456033534034774535358577964;
            6'd41: xpb[3] = 1024'd16832019448175223557627454351650621641656502534343565139040521728982277196084331855957838567289168896708060240230109578618727675681777001214096849068618647073223683845717010715277549162994414181298461449881447896265465191767007412049960930330724562029920453820715717059386993987268904132660516661236183093980;
            6'd42: xpb[3] = 1024'd5138488636264888385979448125611423852945838974133829251882304691642635631373302007565095974817424303023559328288649477162690415006579334457839686849186805203430049347361697090027709953163331042177916840523703713602246211056846932054596214516036922150960474312526631326190917930965352231786998547937007609996;
            6'd43: xpb[3] = 1024'd117511653508479294613130369304386658808933602539659777492855942719279889403971411069187424597003354018782207823804682810285716995172602002256742649646086004267327089418577600802408109934849453624367569839553199377303388080567583225024210068384578731538820398218454603623101369948590433348032170261263426610343;
            6'd44: xpb[3] = 1024'd105818122696568959441482363078347461020222938979450041605697725681940247839260381220794682004531609425097706911863222708829679734497404335500485487426654162397533454920222287177158270725018370485247025230195455194640169099857422745028845352569891091659860418710265517889905293892286881447158652147964251126359;
            6'd45: xpb[3] = 1024'd94124591884658624269834356852308263231512275419240305718539508644600606274549351372401939412059864831413205999921762607373642473822206668744228325207222320527739820421866973551908431515187287346126480620837711011976950119147262265033480636755203451780900439202076432156709217835983329546285134034665075642375;
            6'd46: xpb[3] = 1024'd82431061072748289098186350626269065442801611859030569831381291607260964709838321524009196819588120237728705087980302505917605213147009001987971162987790478657946185923511659926658592305356204207005936011479966829313731138437101785038115920940515811901940459693887346423513141779679777645411615921365900158391;
            6'd47: xpb[3] = 1024'd70737530260837953926538344400229867654090948298820833944223074569921323145127291675616454227116375644044204176038842404461567952471811335231714000768358636788152551425156346301408753095525121067885391402122222646650512157726941305042751205125828172022980480185698260690317065723376225744538097808066724674407;
            6'd48: xpb[3] = 1024'd59043999448927618754890338174190669865380284738611098057064857532581681580416261827223711634644631050359703264097382303005530691796613668475456838548926794918358916926801032676158913885694037928764846792764478463987293177016780825047386489311140532144020500677509174957120989667072673843664579694767549190423;
            6'd49: xpb[3] = 1024'd47350468637017283583242331948151472076669621178401362169906640495242040015705231978830969042172886456675202352155922201549493431121416001719199676329494953048565282428445719050909074675862954789644302183406734281324074196306620345052021773496452892265060521169320089223924913610769121942791061581468373706439;
            6'd50: xpb[3] = 1024'd35656937825106948411594325722112274287958957618191626282748423457902398450994202130438226449701141862990701440214462100093456170446218334962942514110063111178771647930090405425659235466031871650523757574048990098660855215596459865056657057681765252386100541661131003490728837554465570041917543468169198222455;
            6'd51: xpb[3] = 1024'd23963407013196613239946319496073076499248294057981890395590206420562756886283172282045483857229397269306200528273001998637418909771020668206685351890631269308978013431735091800409396256200788511403212964691245915997636234886299385061292341867077612507140562152941917757532761498162018141044025354870022738471;
            6'd52: xpb[3] = 1024'd12269876201286278068298313270033878710537630497772154508431989383223115321572142433652741264757652675621699616331541897181381649095823001450428189671199427439184378933379778175159557046369705372282668355333501733334417254176138905065927626052389972628180582644752832024336685441858466240170507241570847254487;
            6'd53: xpb[3] = 1024'd576345389375942896650307043994680921826966937562418621273772345883473756861112585259998672285908081937198704390081795725344388420625334694171027451767585569390744435024464549909717836538622233162123745975757550671198273465978425070562910237702332749220603136563746291140609385554914339296989128271671770503;
            6'd54: xpb[3] = 1024'd112949510261590349123801228222769915877814730503088366862247410373520727529459221646882327294471837797695847199906115128848370968586648002493073990248666784633287784506240368262290117818224744815351776745005253214372340142976714718040176764106244142137080527042491718588051061403179995455542160841598090770850;
            6'd55: xpb[3] = 1024'd101255979449680013952153221996730718089104066942878630975089193336181085964748191798489584702000093204011346287964655027392333707911450335736816828029234942763494150007885054637040278608393661676231232135647509031709121162266554238044812048291556502258120547534302632854854985346876443554668642728298915286866;
            6'd56: xpb[3] = 1024'd89562448637769678780505215770691520300393403382668895087930976298841444400037161950096842109528348610326845376023194925936296447236252668980559665809803100893700515509529741011790439398562578537110687526289764849045902181556393758049447332476868862379160568026113547121658909290572891653795124614999739802882;
            6'd57: xpb[3] = 1024'd77868917825859343608857209544652322511682739822459159200772759261501802835326132101704099517056604016642344464081734824480259186561055002224302503590371259023906881011174427386540600188731495397990142916932020666382683200846233278054082616662181222500200588517924461388462833234269339752921606501700564318898;
            6'd58: xpb[3] = 1024'd66175387013949008437209203318613124722972076262249423313614542224162161270615102253311356924584859422957843552140274723024221925885857335468045341370939417154113246512819113761290760978900412258869598307574276483719464220136072798058717900847493582621240609009735375655266757177965787852048088388401388834914;
            6'd59: xpb[3] = 1024'd54481856202038673265561197092573926934261412702039687426456325186822519705904072404918614332113114829273342640198814621568184665210659668711788179151507575284319612014463800136040921769069329119749053698216532301056245239425912318063353185032805942742280629501546289922070681121662235951174570275102213350930;
            6'd60: xpb[3] = 1024'd42788325390128338093913190866534729145550749141829951539298108149482878141193042556525871739641370235588841728257354520112147404535462001955531016932075733414525977516108486510791082559238245980628509088858788118393026258715751838067988469218118302863320649993357204188874605065358684050301052161803037866946;
            6'd61: xpb[3] = 1024'd31094794578218002922265184640495531356840085581620215652139891112143236576482012708133129147169625641904340816315894418656110143860264335199273854712643891544732343017753172885541243349407162841507964479501043935729807278005591358072623753403430662984360670485168118455678529009055132149427534048503862382962;
            6'd62: xpb[3] = 1024'd19401263766307667750617178414456333568129422021410479764981674074803595011770982859740386554697881048219839904374434317200072883185066668443016692493212049674938708519397859260291404139576079702387419870143299753066588297295430878077259037588743023105400690976979032722482452952751580248554015935204686898978;
            6'd63: xpb[3] = 1024'd7707732954397332578969172188417135779418758461200743877823457037463953447059953011347643962226136454535338992432974215744035622509869001686759530273780207805145074021042545635041564929744996563266875260785555570403369316585270398081894321774055383226440711468789946989286376896448028347680497821905511414994;
        endcase
    end

    always_comb begin
        case(flag[1][11:6])
            6'd0: xpb[4] = 1024'd0;
            6'd1: xpb[4] = 1024'd120080897826611738806120093367192370735406522026726692118797095065101207219658062072969972584412066170293987487949007548867062202675891669485662493070679406869042114092258449347421964911431119145456528259815051234104511186096006691051508175642597192614300635374717919286196828914073109463925669535231930415341;
            6'd2: xpb[4] = 1024'd116095099969098736213441259329570308726114616927717700109462335065225519102006985235924873954166458031144825568440521663155060564510563004416164861125027772804393553614945681357213690631345032569602858911242862621844661521971116609138037781601964935961781367335318780542287129754217585910732649243838266346351;
            6'd3: xpb[4] = 1024'd112109302111585733620762425291948246716822711828708708100127575065349830984355908398879775323920849891995663648932035777443058926345234339346667229179376138739744993137632913367005416351258945993749189562670674009584811857846226527224567387561332679309262099295919641798377430594362062357539628952444602277361;
            6'd4: xpb[4] = 1024'd108123504254072731028083591254326184707530806729699716090792815065474142866704831561834676693675241752846501729423549891731057288179905674277169597233724504675096432660320145376797142071172859417895520214098485397324962193721336445311096993520700422656742831256520503054467731434506538804346608661050938208371;
            6'd5: xpb[4] = 1024'd104137706396559728435404757216704122698238901630690724081458055065598454749053754724789578063429633613697339809915064006019055650014577009207671965288072870610447872183007377386588867791086772842041850865526296785065112529596446363397626599480068166004223563217121364310558032274651015251153588369657274139381;
            6'd6: xpb[4] = 1024'd100151908539046725842725923179082060688946996531681732072123295065722766631402677887744479433184025474548177890406578120307054011849248344138174333342421236545799311705694609396380593511000686266188181516954108172805262865471556281484156205439435909351704295177722225566648333114795491697960568078263610070391;
            6'd7: xpb[4] = 1024'd96166110681533723250047089141459998679655091432672740062788535065847078513751601050699380802938417335399015970898092234595052373683919679068676701396769602481150751228381841406172319230914599690334512168381919560545413201346666199570685811398803652699185027138323086822738633954939968144767547786869946001401;
            6'd8: xpb[4] = 1024'd92180312824020720657368255103837936670363186333663748053453775065971390396100524213654282172692809196249854051389606348883050735518591013999179069451117968416502190751069073415964044950828513114480842819809730948285563537221776117657215417358171396046665759098923948078828934795084444591574527495476281932411;
            6'd9: xpb[4] = 1024'd88194514966507718064689421066215874661071281234654756044119015066095702278449447376609183542447201057100692131881120463171049097353262348929681437505466334351853630273756305425755770670742426538627173471237542336025713873096886035743745023317539139394146491059524809334919235635228921038381507204082617863421;
            6'd10: xpb[4] = 1024'd84208717108994715472010587028593812651779376135645764034784255066220014160798370539564084912201592917951530212372634577459047459187933683860183805559814700287205069796443537435547496390656339962773504122665353723765864208971995953830274629276906882741627223020125670591009536475373397485188486912688953794431;
            6'd11: xpb[4] = 1024'd80222919251481712879331752990971750642487471036636772025449495066344326043147293702518986281955984778802368292864148691747045821022605018790686173614163066222556509319130769445339222110570253386919834774093165111506014544847105871916804235236274626089107954980726531847099837315517873931995466621295289725441;
            6'd12: xpb[4] = 1024'd76237121393968710286652918953349688633195565937627780016114735066468637925496216865473887651710376639653206373355662806035044182857276353721188541668511432157907948841818001455130947830484166811066165425520976499246164880722215790003333841195642369436588686941327393103190138155662350378802446329901625656451;
            6'd13: xpb[4] = 1024'd72251323536455707693974084915727626623903660838618788006779975066592949807845140028428789021464768500504044453847176920323042544691947688651690909722859798093259388364505233464922673550398080235212496076948787886986315216597325708089863447155010112784069418901928254359280438995806826825609426038507961587461;
            6'd14: xpb[4] = 1024'd68265525678942705101295250878105564614611755739609795997445215066717261690194063191383690391219160361354882534338691034611040906526619023582193277777208164028610827887192465474714399270311993659358826728376599274726465552472435626176393053114377856131550150862529115615370739835951303272416405747114297518471;
            6'd15: xpb[4] = 1024'd64279727821429702508616416840483502605319850640600803988110455066841573572542986354338591760973552222205720614830205148899039268361290358512695645831556529963962267409879697484506124990225907083505157379804410662466615888347545544262922659073745599479030882823129976871461040676095779719223385455720633449481;
            6'd16: xpb[4] = 1024'd60293929963916699915937582802861440596027945541591811978775695066965885454891909517293493130727944083056558695321719263187037630195961693443198013885904895899313706932566929494297850710139820507651488031232222050206766224222655462349452265033113342826511614783730838127551341516240256166030365164326969380491;
            6'd17: xpb[4] = 1024'd56308132106403697323258748765239378586736040442582819969440935067090197337240832680248394500482335943907396775813233377475035992030633028373700381940253261834665146455254161504089576430053733931797818682660033437946916560097765380435981870992481086173992346744331699383641642356384732612837344872933305311501;
            6'd18: xpb[4] = 1024'd52322334248890694730579914727617316577444135343573827960106175067214509219589755843203295870236727804758234856304747491763034353865304363304202749994601627770016585977941393513881302149967647355944149334087844825687066895972875298522511476951848829521473078704932560639731943196529209059644324581539641242511;
            6'd19: xpb[4] = 1024'd48336536391377692137901080689995254568152230244564835950771415067338821101938679006158197239991119665609072936796261606051032715699975698234705118048949993705368025500628625523673027869881560780090479985515656213427217231847985216609041082911216572868953810665533421895822244036673685506451304290145977173521;
            6'd20: xpb[4] = 1024'd44350738533864689545222246652373192558860325145555843941436655067463132984287602169113098609745511526459911017287775720339031077534647033165207486103298359640719465023315857533464753589795474204236810636943467601167367567723095134695570688870584316216434542626134283151912544876818161953258283998752313104531;
            6'd21: xpb[4] = 1024'd40364940676351686952543412614751130549568420046546851932101895067587444866636525332067999979499903387310749097779289834627029439369318368095709854157646725576070904546003089543256479309709387628383141288371278988907517903598205052782100294829952059563915274586735144408002845716962638400065263707358649035541;
            6'd22: xpb[4] = 1024'd36379142818838684359864578577129068540276514947537859922767135067711756748985448495022901349254295248161587178270803948915027801203989703026212222211995091511422344068690321553048205029623301052529471939799090376647668239473314970868629900789319802911396006547336005664093146557107114846872243415964984966551;
            6'd23: xpb[4] = 1024'd32393344961325681767185744539507006530984609848528867913432375067836068631334371657977802719008687109012425258762318063203026163038661037956714590266343457446773783591377553562839930749537214476675802591226901764387818575348424888955159506748687546258876738507936866920183447397251591293679223124571320897561;
            6'd24: xpb[4] = 1024'd28407547103812679174506910501884944521692704749519875904097615067960380513683294820932704088763078969863263339253832177491024524873332372887216958320691823382125223114064785572631656469451127900822133242654713152127968911223534807041689112708055289606357470468537728176273748237396067740486202833177656828571;
            6'd25: xpb[4] = 1024'd24421749246299676581828076464262882512400799650510883894762855068084692396032217983887605458517470830714101419745346291779022886708003707817719326375040189317476662636752017582423382189365041324968463894082524539868119247098644725128218718667423032953838202429138589432364049077540544187293182541783992759581;
            6'd26: xpb[4] = 1024'd20435951388786673989149242426640820503108894551501891885428095068209004278381141146842506828271862691564939500236860406067021248542675042748221694429388555252828102159439249592215107909278954749114794545510335927608269582973754643214748324626790776301318934389739450688454349917685020634100162250390328690591;
            6'd27: xpb[4] = 1024'd16450153531273671396470408389018758493816989452492899876093335068333316160730064309797408198026254552415777580728374520355019610377346377678724062483736921188179541682126481602006833629192868173261125196938147315348419918848864561301277930586158519648799666350340311944544650757829497080907141958996664621601;
            6'd28: xpb[4] = 1024'd12464355673760668803791574351396696484525084353483907866758575068457628043078987472752309567780646413266615661219888634643017972212017712609226430538085287123530981204813713611798559349106781597407455848365958703088570254723974479387807536545526262996280398310941173200634951597973973527714121667603000552611;
            6'd29: xpb[4] = 1024'd8478557816247666211112740313774634475233179254474915857423815068581939925427910635707210937535038274117453741711402748931016334046689047539728798592433653058882420727500945621590285069020695021553786499793770090828720590599084397474337142504894006343761130271542034456725252438118449974521101376209336483621;
            6'd30: xpb[4] = 1024'd4492759958734663618433906276152572465941274155465923848089055068706251807776833798662112307289430134968291822202916863219014695881360382470231166646782018994233860250188177631382010788934608445700117151221581478568870926474194315560866748464261749691241862232142895712815553278262926421328081084815672414631;
            6'd31: xpb[4] = 1024'd506962101221661025755072238530510456649369056456931838754295068830563690125756961617013677043821995819129902694430977507013057716031717400733534701130384929585299772875409641173736508848521869846447802649392866309021262349304233647396354423629493038722594192743756968905854118407402868135060793422008345641;
            6'd32: xpb[4] = 1024'd120587859927833399831875165605722881192055891083183623957551390133931770909783819034586986261455888166113117390643438526374075260391923386886396027771809791798627413865133858988595701420279641015302976062464444100413532448445310924698904530066226685653023229567461676255102683032480512332060730328653938760982;
            6'd33: xpb[4] = 1024'd116602062070320397239196331568100819182763985984174631948216630134056082792132742197541887631210280026963955471134952640662073622226594721816898395826158157733978853387821090998387427140193554439449306713892255488153682784320420842785434136025594429000503961528062537511192983872624988778867710037260274691992;
            6'd34: xpb[4] = 1024'd112616264212807394646517497530478757173472080885165639938881870134180394674481665360496789000964671887814793551626466754950071984061266056747400763880506523669330292910508323008179152860107467863595637365320066875893833120195530760871963741984962172347984693488663398767283284712769465225674689745866610623002;
            6'd35: xpb[4] = 1024'd108630466355294392053838663492856695164180175786156647929547110134304706556830588523451690370719063748665631632117980869238070345895937391677903131934854889604681732433195555017970878580021381287741968016747878263633983456070640678958493347944329915695465425449264260023373585552913941672481669454472946554012;
            6'd36: xpb[4] = 1024'd104644668497781389461159829455234633154888270687147655920212350134429018439179511686406591740473455609516469712609494983526068707730608726608405499989203255540033171955882787027762604299935294711888298668175689651374133791945750597045022953903697659042946157409865121279463886393058418119288649163079282485022;
            6'd37: xpb[4] = 1024'd100658870640268386868480995417612571145596365588138663910877590134553330321528434849361493110227847470367307793101009097814067069565280061538907868043551621475384611478570019037554330019849208136034629319603501039114284127820860515131552559863065402390426889370465982535554187233202894566095628871685618416032;
            6'd38: xpb[4] = 1024'd96673072782755384275802161379990509136304460489129671901542830134677642203877358012316394479982239331218145873592523212102065431399951396469410236097899987410736051001257251047346055739763121560180959971031312426854434463695970433218082165822433145737907621331066843791644488073347371012902608580291954347042;
            6'd39: xpb[4] = 1024'd92687274925242381683123327342368447127012555390120679892208070134801954086226281175271295849736631192068983954084037326390063793234622731399912604152248353346087490523944483057137781459677034984327290622459123814594584799571080351304611771781800889085388353291667705047734788913491847459709588288898290278052;
            6'd40: xpb[4] = 1024'd88701477067729379090444493304746385117720650291111687882873310134926265968575204338226197219491023052919822034575551440678062155069294066330414972206596719281438930046631715066929507179590948408473621273886935202334735135446190269391141377741168632432869085252268566303825089753636323906516567997504626209062;
            6'd41: xpb[4] = 1024'd84715679210216376497765659267124323108428745192102695873538550135050577850924127501181098589245414913770660115067065554966060516903965401260917340260945085216790369569318947076721232899504861832619951925314746590074885471321300187477670983700536375780349817212869427559915390593780800353323547706110962140072;
            6'd42: xpb[4] = 1024'd80729881352703373905086825229502261099136840093093703864203790135174889733273050664135999958999806774621498195558579669254058878738636736191419708315293451152141809092006179086512958619418775256766282576742557977815035807196410105564200589659904119127830549173470288816005691433925276800130527414717298071082;
            6'd43: xpb[4] = 1024'd76744083495190371312407991191880199089844934994084711854869030135299201615621973827090901328754198635472336276050093783542057240573308071121922076369641817087493248614693411096304684339332688680912613228170369365555186143071520023650730195619271862475311281134071150072095992274069753246937507123323634002092;
            6'd44: xpb[4] = 1024'd72758285637677368719729157154258137080553029895075719845534270135423513497970896990045802698508590496323174356541607897830055602407979406052424444423990183022844688137380643106096410059246602105058943879598180753295336478946629941737259801578639605822792013094672011328186293114214229693744486831929969933102;
            6'd45: xpb[4] = 1024'd68772487780164366127050323116636075071261124796066727836199510135547825380319820153000704068262982357174012437033122012118053964242650740982926812478338548958196127660067875115888135779160515529205274531025992141035486814821739859823789407538007349170272745055272872584276593954358706140551466540536305864112;
            6'd46: xpb[4] = 1024'd64786689922651363534371489079014013061969219697057735826864750135672137262668743315955605438017374218024850517524636126406052326077322075913429180532686914893547567182755107125679861499074428953351605182453803528775637150696849777910319013497375092517753477015873733840366894794503182587358446249142641795122;
            6'd47: xpb[4] = 1024'd60800892065138360941692655041391951052677314598048743817529990135796449145017666478910506807771766078875688598016150240694050687911993410843931548587035280828899006705442339135471587218988342377497935833881614916515787486571959695996848619456742835865234208976474595096457195634647659034165425957748977726132;
            6'd48: xpb[4] = 1024'd56815094207625358349013821003769889043385409499039751808195230135920761027366589641865408177526157939726526678507664354982049049746664745774433916641383646764250446228129571145263312938902255801644266485309426304255937822447069614083378225416110579212714940937075456352547496474792135480972405666355313657142;
            6'd49: xpb[4] = 1024'd52829296350112355756334986966147827034093504400030759798860470136045072909715512804820309547280549800577364758999178469270047411581336080704936284695732012699601885750816803155055038658816169225790597136737237691996088158322179532169907831375478322560195672897676317608637797314936611927779385374961649588152;
            6'd50: xpb[4] = 1024'd48843498492599353163656152928525765024801599301021767789525710136169384792064435967775210917034941661428202839490692583558045773416007415635438652750080378634953325273504035164846764378730082649936927788165049079736238494197289450256437437334846065907676404858277178864728098155081088374586365083567985519162;
            6'd51: xpb[4] = 1024'd44857700635086350570977318890903703015509694202012775780190950136293696674413359130730112286789333522279040919982206697846044135250678750565941020804428744570304764796191267174638490098643996074083258439592860467476388830072399368342967043294213809255157136818878040120818398995225564821393344792174321450172;
            6'd52: xpb[4] = 1024'd40871902777573347978298484853281641006217789103003783770856190136418008556762282293685013656543725383129879000473720812134042497085350085496443388858777110505656204318878499184430215818557909498229589091020671855216539165947509286429496649253581552602637868779478901376908699835370041268200324500780657381182;
            6'd53: xpb[4] = 1024'd36886104920060345385619650815659578996925884003994791761521430136542320439111205456639915026298117243980717080965234926422040858920021420426945756913125476441007643841565731194221941538471822922375919742448483242956689501822619204516026255212949295950118600740079762632999000675514517715007304209386993312192;
            6'd54: xpb[4] = 1024'd32900307062547342792940816778037516987633978904985799752186670136666632321460128619594816396052509104831555161456749040710039220754692755357448124967473842376359083364252963204013667258385736346522250393876294630696839837697729122602555861172317039297599332700680623889089301515658994161814283917993329243202;
            6'd55: xpb[4] = 1024'd28914509205034340200261982740415454978342073805976807742851910136790944203809051782549717765806900965682393241948263154998037582589364090287950493021822208311710522886940195213805392978299649770668581045304106018436990173572839040689085467131684782645080064661281485145179602355803470608621263626599665174212;
            6'd56: xpb[4] = 1024'd24928711347521337607583148702793392969050168706967815733517150136915256086157974945504619135561292826533231322439777269286035944424035425218452861076170574247061962409627427223597118698213563194814911696731917406177140509447948958775615073091052525992560796621882346401269903195947947055428243335206001105222;
            6'd57: xpb[4] = 1024'd20942913490008335014904314665171330959758263607958823724182390137039567968506898108459520505315684687384069402931291383574034306258706760148955229130518940182413401932314659233388844418127476618961242348159728793917290845323058876862144679050420269340041528582483207657360204036092423502235223043812337036232;
            6'd58: xpb[4] = 1024'd16957115632495332422225480627549268950466358508949831714847630137163879850855821271414421875070076548234907483422805497862032668093378095079457597184867306117764841455001891243180570138041390043107572999587540181657441181198168794948674285009788012687522260543084068913450504876236899949042202752418672967242;
            6'd59: xpb[4] = 1024'd12971317774982329829546646589927206941174453409940839705512870137288191733204744434369323244824468409085745563914319612150031029928049430009959965239215672053116280977689123252972295857955303467253903651015351569397591517073278713035203890969155756035002992503684930169540805716381376395849182461025008898252;
            6'd60: xpb[4] = 1024'd8985519917469327236867812552305144931882548310931847696178110137412503615553667597324224614578860269936583644405833726438029391762720764940462333293564037988467720500376355262764021577869216891400234302443162957137741852948388631121733496928523499382483724464285791425631106556525852842656162169631344829262;
            6'd61: xpb[4] = 1024'd4999722059956324644188978514683082922590643211922855686843350137536815497902590760279125984333252130787421724897347840726027753597392099870964701347912403923819160023063587272555747297783130315546564953870974344877892188823498549208263102887891242729964456424886652681721407396670329289463141878237680760272;
            6'd62: xpb[4] = 1024'd1013924202443322051510144477061020913298738112913863677508590137661127380251513923234027354087643991638259805388861955014026115432063434801467069402260769859170599545750819282347473017697043739692895605298785732618042524698608467294792708847258986077445188385487513937811708236814805736270121586844016691282;
            6'd63: xpb[4] = 1024'd121094822029055060857630237844253391648705260139640555796305685202762334599909575996203999938499710161932247293337869503881088318107955104287129562472940176728212713638009268629769437929128162885149423865113836966722553710794615158346300884489856178691745823760205433224008537150887915200195791122075947106623;
        endcase
    end

    always_comb begin
        case(flag[1][16:12])
            5'd0: xpb[5] = 1024'd0;
            5'd1: xpb[5] = 1024'd117109024171542058264951403806631329639413355040631563786970925202886646482258499159158901308254102022783085373829383618169086679942626439217631930527288542663564153160696500639561163649042076309295754516541648354462704046669725076432830490449223922039226555720806294480098837991032391647002770830682283037633;
            5'd2: xpb[5] = 1024'd110151352658959375131103880208448226534128282955527443445809995340796397627207859408302731401850529736123021340201273801759109519044032543880103736038246044393437631751821783941492088106566946897281311424696056862561047243118553379900682411215218394811633208027495530930091147908136150276886851834738971590935;
            5'd3: xpb[5] = 1024'd103193681146376691997256356610265123428843210870423323104649065478706148772157219657446561495446957449462957306573163985349132358145438648542575541549203546123311110342947067243423012564091817485266868332850465370659390439567381683368534331981212867584039860334184767380083457825239908906770932838795660144237;
            5'd4: xpb[5] = 1024'd96236009633794008863408833012082020323558138785319202763488135616615899917106579906590391589043385162802893272945054168939155197246844753205047347060161047853184588934072350545353937021616688073252425241004873878757733636016209986836386252747207340356446512640874003830075767742343667536655013842852348697539;
            5'd5: xpb[5] = 1024'd89278338121211325729561309413898917218273066700215082422327205754525651062055940155734221682639812876142829239316944352529178036348250857867519152571118549583058067525197633847284861479141558661237982149159282386856076832465038290304238173513201813128853164947563240280068077659447426166539094846909037250841;
            5'd6: xpb[5] = 1024'd82320666608628642595713785815715814112987994615110962081166275892435402207005300404878051776236240589482765205688834536119200875449656962529990958082076051312931546116322917149215785936666429249223539057313690894954420028913866593772090094279196285901259817254252476730060387576551184796423175850965725804143;
            5'd7: xpb[5] = 1024'd75362995096045959461866262217532711007702922530006841740005346030345153351954660654021881869832668302822701172060724719709223714551063067192462763593033553042805024707448200451146710394191299837209095965468099403052763225362694897239942015045190758673666469560941713180052697493654943426307256855022414357445;
            5'd8: xpb[5] = 1024'd68405323583463276328018738619349607902417850444902721398844416168254904496904020903165711963429096016162637138432614903299246553652469171854934569103991054772678503298573483753077634851716170425194652873622507911151106421811523200707793935811185231446073121867630949630045007410758702056191337859079102910747;
            5'd9: xpb[5] = 1024'd61447652070880593194171215021166504797132778359798601057683486306164655641853381152309542057025523729502573104804505086889269392753875276517406374614948556502551981889698767055008559309241041013180209781776916419249449618260351504175645856577179704218479774174320186080037317327862460686075418863135791464049;
            5'd10: xpb[5] = 1024'd54489980558297910060323691422983401691847706274694480716522556444074406786802741401453372150621951442842509071176395270479292231855281381179878180125906058232425460480824050356939483766765911601165766689931324927347792814709179807643497777343174176990886426481009422530029627244966219315959499867192480017351;
            5'd11: xpb[5] = 1024'd47532309045715226926476167824800298586562634189590360375361626581984157931752101650597202244218379156182445037548285454069315070956687485842349985636863559962298939071949333658870408224290782189151323598085733435446136011158008111111349698109168649763293078787698658980021937162069977945843580871249168570653;
            5'd12: xpb[5] = 1024'd40574637533132543792628644226617195481277562104486240034200696719893909076701461899741032337814806869522381003920175637659337910058093590504821791147821061692172417663074616960801332681815652777136880506240141943544479207606836414579201618875163122535699731094387895430014247079173736575727661875305857123955;
            5'd13: xpb[5] = 1024'd33616966020549860658781120628434092375992490019382119693039766857803660221650822148884862431411234582862316970292065821249360749159499695167293596658778563422045896254199900262732257139340523365122437414394550451642822404055664718047053539641157595308106383401077131880006556996277495205611742879362545677257;
            5'd14: xpb[5] = 1024'd26659294507967177524933597030250989270707417934277999351878836995713411366600182398028692525007662296202252936663956004839383588260905799829765402169736065151919374845325183564663181596865393953107994322548958959741165600504493021514905460407152068080513035707766368329998866913381253835495823883419234230559;
            5'd15: xpb[5] = 1024'd19701622995384494391086073432067886165422345849173879010717907133623162511549542647172522618604090009542188903035846188429406427362311904492237207680693566881792853436450466866594106054390264541093551230703367467839508796953321324982757381173146540852919688014455604779991176830485012465379904887475922783861;
            5'd16: xpb[5] = 1024'd12743951482801811257238549833884783060137273764069758669556977271532913656498902896316352712200517722882124869407736372019429266463718009154709013191651068611666332027575750168525030511915135129079108138857775975937851993402149628450609301939141013625326340321144841229983486747588771095263985891532611337163;
            5'd17: xpb[5] = 1024'd5786279970219128123391026235701679954852201678965638328396047409442664801448263145460182805796945436222060835779626555609452105565124113817180818702608570341539810618701033470455954969440005717064665047012184484036195189850977931918461222705135486397732992627834077679975796664692529725148066895589299890465;
            5'd18: xpb[5] = 1024'd122895304141761186388342430042333009594265556719597202115366972612329311283706762304619084114051047459005146209609010173778538785507750553034812749229897113005103963779397534110017118618482082026360419563553832838498899236520703008351291713154359408436959548348640372160074634655724921372150837726271582928098;
            5'd19: xpb[5] = 1024'd115937632629178503254494906444149906488980484634493081774206042750239062428656122553762914207647475172345082175980900357368561624609156657697284554740854614734977442370522817411948043076006952614345976471708241346597242432969531311819143633920353881209366200655329608610066944572828680002034918730328271481400;
            5'd20: xpb[5] = 1024'd108979961116595820120647382845966803383695412549388961433045112888148813573605482802906744301243902885685018142352790540958584463710562762359756360251812116464850920961648100713878967533531823202331533379862649854695585629418359615286995554686348353981772852962018845060059254489932438631918999734384960034702;
            5'd21: xpb[5] = 1024'd102022289604013136986799859247783700278410340464284841091884183026058564718554843052050574394840330599024954108724680724548607302811968867022228165762769618194724399552773384015809891991056693790317090288017058362793928825867187918754847475452342826754179505268708081510051564407036197261803080738441648588004;
            5'd22: xpb[5] = 1024'd95064618091430453852952335649600597173125268379180720750723253163968315863504203301194404488436758312364890075096570908138630141913374971684699971273727119924597878143898667317740816448581564378302647196171466870892272022316016222222699396218337299526586157575397317960043874324139955891687161742498337141306;
            5'd23: xpb[5] = 1024'd88106946578847770719104812051417494067840196294076600409562323301878067008453563550338234582033186025704826041468461091728652981014781076347171776784684621654471356735023950619671740906106434966288204104325875378990615218764844525690551316984331772298992809882086554410036184241243714521571242746555025694608;
            5'd24: xpb[5] = 1024'd81149275066265087585257288453234390962555124208972480068401393439787818153402923799482064675629613739044762007840351275318675820116187181009643582295642123384344835326149233921602665363631305554273761012480283887088958415213672829158403237750326245071399462188775790860028494158347473151455323750611714247910;
            5'd25: xpb[5] = 1024'd74191603553682404451409764855051287857270052123868359727240463577697569298352284048625894769226041452384697974212241458908698659217593285672115387806599625114218313917274517223533589821156176142259317920634692395187301611662501132626255158516320717843806114495465027310020804075451231781339404754668402801212;
            5'd26: xpb[5] = 1024'd67233932041099721317562241256868184751984980038764239386079533715607320443301644297769724862822469165724633940584131642498721498318999390334587193317557126844091792508399800525464514278681046730244874828789100903285644808111329436094107079282315190616212766802154263760013113992554990411223485758725091354514;
            5'd27: xpb[5] = 1024'd60276260528517038183714717658685081646699907953660119044918603853517071588251004546913554956418896879064569906956021826088744337420405494997058998828514628573965271099525083827395438736205917318230431736943509411383988004560157739561959000048309663388619419108843500210005423909658749041107566762781779907816;
            5'd28: xpb[5] = 1024'd53318589015934355049867194060501978541414835868555998703757673991426822733200364796057385050015324592404505873327912009678767176521811599659530804339472130303838749690650367129326363193730787906215988645097917919482331201008986043029810920814304136161026071415532736659997733826762507670991647766838468461118;
            5'd29: xpb[5] = 1024'd46360917503351671916019670462318875436129763783451878362596744129336573878149725045201215143611752305744441839699802193268790015623217704322002609850429632033712228281775650431257287651255658494201545553252326427580674397457814346497662841580298608933432723722221973109990043743866266300875728770895157014420;
            5'd30: xpb[5] = 1024'd39403245990768988782172146864135772330844691698347758021435814267246325023099085294345045237208180019084377806071692376858812854724623808984474415361387133763585706872900933733188212108780529082187102461406734935679017593906642649965514762346293081705839376028911209559982353660970024930759809774951845567722;
            5'd31: xpb[5] = 1024'd32445574478186305648324623265952669225559619613243637680274884405156076168048445543488875330804607732424313772443582560448835693826029913646946220872344635493459185464026217035119136566305399670172659369561143443777360790355470953433366683112287554478246028335600446009974663578073783560643890779008534121024;
        endcase
    end



endmodule
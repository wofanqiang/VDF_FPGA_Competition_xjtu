module xpb_4_260
(
    input [4:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    4'b0000 : xpb = 1024'h0;
    4'b0001 : xpb = 1024'h9dadfaf9f421c3b5ee4049696b8d0127cde11ab194c9d5c9152eb87c40dccd135360bc17fff418f6e2d569833bf50bed4012f5e6d4753736f2f8b93b74e90b958eb03679d20808e3540c18b5dd1e90d185aee0031ea4b50d6474e2dae3d9818369de5b3c7c6f85062f64e24bfd6cf71263ed7b46bbbcd46d6f7dc53125434e55;
    4'b0010 : xpb = 1024'h8aaeb09e265552a3117b1afbc6bfbafe2a4c3232541c0b1aac80b7a2ceb6ed1ea378fab735c1b35f264c93bf948c07101c0bc3e786379e2235523318aeffa279a9113844f47f1481957e2ec921615d721758c66db0c33d0a135d33bb0d886074a4b5244f4816117ed809ddb90309c7fb790117ab272e4baa988c0f5dc1a4363f;
    4'b0011 : xpb = 1024'h77af66425888e19034b5ec8e21f274d486b749b3136e406c43d2b6c95c910d29f39139566b8f4dc769c3bdfbed230232f80491e837fa050d77abacf5e916395dc3723a1016f6201fd6f044dc65a42a12a902acd842e1c506c245849b37373f65df8bed6213bc9df780aed92608a698e48e14b40f929fc2e7c19a598a5e051e29;
    4'b0100 : xpb = 1024'h64b01be68abc707d57f0be207d252eaae3226133d2c075bddb24b5efea6b2d3543a977f5a15ce82fad3ae83845b9fd55d3fd5fe8e9bc6bf8ba0526d3232cd041ddd33bdb396d2bbe18625aefa9e6f6b33aac9342d5004d03712dd57b60e61e571a62b674df632a702953d4930e4369cda3285073fe113a24eaa8a3b6fa660613;
    4'b0101 : xpb = 1024'h51b0d18abcefff6a7b2b8fb2d857e8813f8d78b49212ab0f7276b51678454d4093c1b694d72a8297f0b212749e50f878aff62de99b7ed2e3fc5ea0b05d436725f8343da65be4375c59d47102ee29c353cc5679ad671ed5002016265b8a94fd4855397f87ab09b6e8d1f8d00013e03ab6b83becd86982b16213b6ede396c6edfd;
    4'b0110 : xpb = 1024'h3eb1872eef238e579e666145338aa2579bf890355164e06109c8b43d061f6d4be3d9f5340cf81d0034293cb0f6e7f39b8beefbea4d4139cf3eb81a8d9759fe0a12953f717e5b42fa9b468716326c8ff45e006017f93d5cfccefe773bb443dc399010489a76b043617a9dcb6d197d0b9fcd4f893cd4f4289f3cc538103327d5e7;
    4'b0111 : xpb = 1024'h2bb23cd321571d44c1a132d78ebd5c2df863a7b610b715b2a11ab36393f98d5733f233d342c5b76877a066ed4f7eeebe67e7c9eaff03a0ba8111946ad17094ee2cf6413ca0d24e98dcb89d2976af5c94efaa46828b5be4f97de6c81bddf2bb2acae711ad4256cfda2342c6da1f19dc88e26325a140659fdc65d3823ccf88bdd1;
    4'b1000 : xpb = 1024'h18b2f277538aac31e4dc0469e9f0160454cebf36d0094b04386cb28a21d3ad62840a7272789351d0bb179129a815e9e143e097ebb0c607a5c36b0e480b872bd247574307c3495a371e2ab33cbaf2293581542ced1d7a6cf62ccf18fc07a19a1c05bddac00dfd5c52cbe7c24724b6ad71f776c205abd717198ee1cc696be9a5bb;
    4'b1001 : xpb = 1024'h5b3a81b85be3b1f0816d5fc4522cfdab139d6b78f5b8055cfbeb1b0afadcd6dd422b111ae60ec38fe8ebb6600ace5041fd965ec62886e9105c48825459dc2b661b844d2e5c065d55f9cc94fff34f5d612fe1357af98f4f2dbb769dc3150790d4094a3d2d9a3e8cb748cbdb42a537e5b0c8a5e6a17488e56b7f01696084a8da5;
    4'b1010 : xpb = 1024'ha361a31579dffed4f6571f65b0afd1027f1af1692425561ee4ed6a2cf08a9a8127836d29ae55052fe16424e93ca1f0f15fec5bd336fda5c7f8bd4160ba86ce4bf0687b4cb7c86eb8b3a8e205dc5386a798acf35ace3daa00402c4cb71529fa90aa72ff0f56136dd1a3f1a00027c0756d7077d9b0d30562c4276ddbc72d8ddbfa;
    4'b1011 : xpb = 1024'h906258b9ac138dc21991f0f80be28ad8db8608e9e3778b707c3f69537e64ba8c779babc8e4229f9824db4f259538ec143be529d3e8c00cb33b16bb3df49d65300ac97d17da3f7a56f51af819209653482a56d9c5605c31fcef149d973ed8d981e549c82221b9fa4a4c969b6d2d5d4656858b76153e76da01507c25f3c9eec3e4;
    4'b1100 : xpb = 1024'h7d630e5dde471caf3cccc28a671544af37f1206aa2c9c0c21391687a0c3eda97c7b3ea6819f03a0068527961edcfe73717ddf7d49a82739e7d70351b2eb3fc14252a7ee2fcb685f5368d0e2c64d91fe8bc00c02ff27ab9f99dfcee776887b87320209134ed6086c2f53b96da32fa173f9a9f1279a9e8513e798a7020664fabce;
    4'b1101 : xpb = 1024'h6a63c402107aab9c6007941cc247fe85945c37eb621bf613aae367a09a18faa317cc29074fbdd468abc9a39e4666e259f3d6c5d54c44da89bfc9aef868ca92f83f8b80ae1f2d919377ff243fa91bec894daaa69a849941f64ce53f57923697645af75a47b907133b9de092473896e828afb2aede1559c87ba298ba4d02b093b8;
    4'b1110 : xpb = 1024'h576479a642ae3a89834265af1d7ab85bf0c74f6c216e2b65423566c727f31aae67e467a6858b6ed0ef40cdda9efddd7ccfcf93d5fe074175022328d5a2e129dc59ec827941a49d31b9713a52ed5eb929df548d0516b7c9f2fbcd9037bbe5765595ce235a84ad9fb446858db43e33b911c4c64b4280cb3fb8cba704799f117ba2;
    4'b1111 : xpb = 1024'h44652f4a74e1c976a67d374178ad72324d3266ece0c060b6d98765edb5cd3ab9b7fca645bb59093932b7f816f794d89fabc861d6afc9a860447ca2b2dcf7c0c0744d8444641ba8cffae3506631a185ca70fe736fa8d651efaab5e117e5945546d0a4ec6d50542c2cef2a892143d089fad9d9e7a6ec3cb6f5f4b54ea63b72638c;
    endcase
end

endmodule

module xpb_5_245
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h44adf529557f81a3fbe6129f995c0e86b88bdcebb6bcd3615dec701fb2b771ff917d5a16e5b38a659dfc25ff5ef34e2ce35772dc2e166e457a2b2c5111102bd1f942cef8bb8ddda2650ba952691a56b5b0dce26a7dd57cd9c2cc56bfdd06ce381972a31b0f02770bfd0702853ba7514f489d13afaa8762c8a69bc02ac39f5b1a;
    5'b00010 : xpb = 1024'h895bea52aaff0347f7cc253f32b81d0d7117b9d76d79a6c2bbd8e03f656ee3ff22fab42dcb6714cb3bf84bfebde69c59c6aee5b85c2cdc8af45658a2222057a3f2859df1771bbb44ca1752a4d234ad6b61b9c4d4fbaaf9b38598ad7fba0d9c7032e546361e04ee17fa0e050a774ea29e913a275f550ec5914d378055873eb634;
    5'b00011 : xpb = 1024'h1d5c9a263e90502328acc007bbb9e442b82d93924ebed9ac9be897096523a8f6b12f90cbe6f420a23a9632b7397bd9bc45ec30ae67907a84bde24594f85e0ec47779383b83189ba21c88f954a2733ff01e91ada6ecfa497c92d87244dce9c8161d5057277c3e6c96705520b0bb25cdc48afd5c2caf4acb29ad63c57bc1fbaae3;
    5'b00100 : xpb = 1024'h620a8f4f940fd1c72492d2a75515f2c970b9707e057bad0df9d5072917db1af642aceae2cca7ab07d89258b6986f27e92943a38a95a6e8ca380d71e6096e3a9670bc07343ea679448194a2a70b8d96a5cf6e90116acfc65655a4c904b9f0964e36c2fa428b40e3a26d5c2335f6cd1f13d39a6fdc59d22df253ff85a6859b05fd;
    5'b00101 : xpb = 1024'ha6b88478e98f536b2078e546ee72015029454d69bc38806f57c17748ca928cf5d42a44f9b25b356d768e7eb5f76276160c9b1666c3bd570fb2389e371a7e666869fed62cfa3456e6e6a04bf974a7ed5b804b727be8a5433018711fc496f7648650359d5d9a435aae6a6325bb327470631c37838c045990bafa9b45d1493a6117;
    5'b00110 : xpb = 1024'h3ab9344c7d20a0465159800f7773c885705b27249d7db35937d12e12ca4751ed625f2197cde84144752c656e72f7b3788bd8615ccf20f5097bc48b29f0bc1d88eef27077063137443911f2a944e67fe03d235b4dd9f492f925b0e489b9d3902c3aa0ae4ef87cd92ce0aa4161764b9b8915fab8595e9596535ac78af783f755c6;
    5'b00111 : xpb = 1024'h7f672975d2a021ea4d3f92af10cfd70c28e70410543a86ba95bd9e327cfec3ecf3dc7baeb39bcbaa13288b6dd1eb01a56f2fd438fd37634ef5efb77b01cc495ae8353f6fc1bf14e69e1d9bfbae00d695ee003db857ca0fd2e87d3b4996da5e645413516a077f5038ddb143e6b1f2ecd85e97cc09091cf91c01634b224796b0e0;
    5'b01000 : xpb = 1024'h1367d94966316ec57e202d7799d19e416ffcddcb357fb9a475cd54fc7cb388e48211584ccf28d78111c672264d803f07ee6d1f2f089b0148bf7ba46dd80a007b6d28d9b9cdbbf543f08f42ab7e3f691aaad8268a49195f9bf5bd000eb9b68a0a3e7e625b65b8ceb753f85f8cf5ca17fe585b00d66358feb4618f90488253a58f;
    5'b01001 : xpb = 1024'h5815ce72bbb0f0697a064017332dacc82888bab6ec3c8d05d3b9c51c2f6afae4138eb263b4dc61e6afc29825ac738d34d1c4920b36b16f8e39a6d0bee91a2c4d666ba8b28949d2e6559aebfde759bfd05bb508f4c6eedc75b88956ce96bd584257f1057674bb45c350ff62123171694da0f814860de0617d082b507345f300a9;
    5'b01010 : xpb = 1024'h9cc3c39c1130720d75ec52b6cc89bb4ee11497a2a2f9606731a6353be2226ce3a50c0c7a9a8fec4c4dbebe250b66db61b51c04e764c7ddd3b3d1fd0ffa2a581f5fae77ab44d7b088baa69550507416860c91eb5f44c4594f7b55ad8e73c4267a7163a89183bdbccf4e0664976d18ba9ce9952835b867c445aec7109e09925bc3;
    5'b01011 : xpb = 1024'h30c4736fa4c1bee8a6cced7f558b8284282a715d843e935111b5ec05e1d731db3340e918b61cf8234c5ca4dd86fc18c434594fdd702b7bcd7d5dea02d0680f3fe4a211f550d490e60d183c0020b2a90ac969d4313613a9188895725396a052205bceb982e1f73b4dc44d803db0efe5c2e3585d0312a3c9de0ef355c4444f5072;
    5'b01100 : xpb = 1024'h75726898fa41408ca2b3001eeee7910ae0b64e493afb66b26fa25c25948ea3dac4be432f9bd08288ea58cadce5ef66f117b0c2b99e41ea12f7891653e1783b11dde4e0ee0c626e887223e55289ccffc07a46b69bb3e925f24b61c91373a7205875415c9df0f9b259c15482c2ec9737122bf570b2bd2b2ca6b58f15ef07eeab8c;
    5'b01101 : xpb = 1024'h973186c8dd28d67d3939ae777e9584027cc28041c40999c4fb212ef944368d252f31fcdb75d8e5fe8f6b1956184a45396ee0dafa9a5880cc1150346b7b5f23262d87b38185f4ee5c4958c025a0b9245371e9f6da53875bb58a18dd896834bfe5fac6d8f4f3330d8379b9e69306e623825b8a5801767323f15bb5b1542aba03b;
    5'b01110 : xpb = 1024'h4e210d95e3520f0bcf79ad87114566c6e05804efd2fd6cfdad9e830f46fadad1e47079e49d1118c586f2d794c077f2807a45808bd7bbf6523b402f97c8c61e045c1b4a30d3ed2c8829a13554c325e8fae7fb81d8230df2951b6de498738a1a36791f10aa5e35a7e434a2a0ee6c15b3876e55b92fc1ee9507bc571b40064afb55;
    5'b01111 : xpb = 1024'h92cf02bf38d190afcb5fc026aaa1754d98e3e1db89ba405f0b8af32ef9b24cd175edd3fb82c4a32b24eefd941f6b40ad5d9cf36805d26497b56b5be8d9d649d6555e19298f7b0a2a8eacdea72c403fb098d86442a0e36f6ede3a3b585090e86e9291b3c56d381ef031a9a373a7bd04d6b6f2ccdf6c75f7d062f2db6ac9ea566f;
    5'b10000 : xpb = 1024'h26cfb292cc62dd8afc405aef33a33c82dff9bb966aff7348eb9aa9f8f96711c90422b0999e51af02238ce44c9b007e0fdcda3e5e113602917ef748dbb01400f6da51b3739b77ea87e11e8556fc7ed23555b04d149232bf37eb7a001d736d14147cfcc4b6cb719d6ea7f0bf19eb942ffcb0b601acc6b1fd68c31f209104a74b1e;
    5'b10001 : xpb = 1024'h6b7da7bc21e25f2ef8266d8eccff4b099885988221bc46aa49871a18ac1e83c895a00ab084053967c1890a4bf9f3cc3cc031b13a3f4c70d6f922752cc1242cc8d394826c5705c82a462a2ea9659928eb068d2f7f10083c11ae4656dd5073e24c966f67d1da74147aa4f7c19f273b814bf953155c7139603169bae0bbc846a638;
    5'b10010 : xpb = 1024'hb02b9ce57761e0d2f40c802e665b59905111756dd8791a0ba7738a385ed5f5c8271d64c769b8c3cd5f85304b58e71a69a38924166d62df1c734da17dd234589accd751651293a5ccab35d7fbceb37fa0b76a11e98dddb8eb7112ad9d2d7ab084afe20aece9768b86a1fec42462e2d29b41f0290c1bc0c2fa1056a0e68be60152;
    5'b10011 : xpb = 1024'h442c4cb90af32dae24ed1af6ef5d20c598274f28b9be4cf5878341025e8ababfb55241658545cfa45e231703d47c57cc22c66f0c78c67d163cd98e70a8720fbb51caebaf1e908629fda77eab9ef212257441fabb7f2d08b47e5272625056dc2a9a4d1bde47b00a051845dfcaa6b9fdc13bb35dd975fcc8927082e60cc6a2f601;
    5'b10100 : xpb = 1024'h88da41e26072af5220d32d9688b92f4c50b32c14707b2056e56fb12211422cbf46cf9b7c6af95a09fc1f3d03336fa5f9061de1e8a6dceb5bb704bac1b9823b8d4b0dbaa7da1e63cc62b327fe080c68db251edd25fd02858e411ec9222d5daa62b3bfbef956b28111154ce24fe2614f108450718920842b5b171ea6378a42511b;
    5'b10101 : xpb = 1024'h1cdaf1b5f403fc2d51b3c85f11baf68197c905cf51c05340c57f67ec10f6f1b6d504781a868665e0fabd23bbaf04e35b855b2cdeb24089558090a7b48fbff2add00154f1e61b4429b524ceadd84afb5fe1f6c5f7ee51d5574e5e8de75039d6089e2acfeab4ebff8f8b93fdf626387a367e13a6567ac030f3774aeb5dc4ff45ca;
    5'b10110 : xpb = 1024'h6188e6df49837dd14d99dafeab1705085054e2bb087d26a2236bd80bc3ae63b66681d2316c39f04698b949bb0df8318868b29fbae056f79afabbd405a0d01e7fc94423eaa1a921cc1a3078004165521592d3a8626c275231112ae4a72d40a440b79d7305c3ee769b889b007b61dfcb85c6b0ba06254793bc1de6ab88889ea0e4;
    5'b10111 : xpb = 1024'ha636dc089f02ff75497fed9e4473138f08e0bfa6bf39fa038158482b7665d5b5f7ff2c4851ed7aac36b56fba6ceb7fb54c0a12970e6d65e074e70056b1e04a51c286f2e35d36ff6e7f3c2152aa7fa8cb43b08acce9fccf0ad3f73b670a477278d1101620d2f0eda785a203009d871cd50f4dcdb5cfcef684c4826bb34c3dfbfe;
    5'b11000 : xpb = 1024'h3a378bdc32944c507a608866cd74dac44ff69961a07f2ced6167fef5761a9aad863408e66d7a868335535672e880bd17cb475d8d19d103da3e72ed49881e0172477a8d2d6933dfcbd1adc8027abe3b500088739edb4c1ed3e137002c2d239e1ebb7b2712312a6c25fbe91ea6e15e47fb091102832a0afc1d24aeb0d986faf0ad;
    5'b11001 : xpb = 1024'h7ee581058813cdf476469b0666d0e94b0882764d573c004ebf546f1528d20cad17b162fd532e10e8d34f7c7247740b44ae9ed06947e7721fb89e199a992e2d4440bd5c2624c1bd6e36b97154e3d89205b165560959219bada40356ec0a2a6c56d4edca2d402ce331f8f0212c1d05994a51ae1632d4925ee5cb4a71044a9a4bc7;
    5'b11010 : xpb = 1024'h12e630d91ba51acfa72735ceefd2b0804f985008388133389f6425df2886d1a4a5e63f9b6ebb1cbfd1ed632ac30948a72ddc1b5f534b1019822a068d6f6be464c5b0f67030be9dcb892b1804b417248a6e3d3edb4a70eb76b1431bb12d0697fcbf58db1e9e6661b06f373cd260dcc4704b714b002ece647e2b76b62a85574076;
    5'b11011 : xpb = 1024'h5794260271249c73a30d486e892ebf0708242cf3ef3e0699fd5095fedb3e43a4376399b2546ea7256fe9892a21fc96d411338e3b81617e5efc5532de807c1036bef3c568ec4c7b6dee36c1571d317b401f1a2145c8466850740f72710a0d6634d8cb7e39ad68d8bc6c3e3f579c8415bf940e5eafd955c746d212765548f69b90;
    5'b11100 : xpb = 1024'h9c421b2bc6a41e179ef35b0e228acd8dc0b009dfa5fad9fb5b3d061e8df5b5a3c8e0f3c93a22318b0de5af2980efe500f48b0117af77eca476805f2f918c3c08b8369461a7da591053426aa9864bd1f5cff703b0461be52a36dbc930e714346cf23e2154bc6b4fc8694541dcd82b670edcab725f83dd2a0f78ae36800c95f6aa;
    5'b11101 : xpb = 1024'h3042caff5a356af2cfd3f5d6ab8c94c307c5e39a87400ce53b4cbce88daa7a9b5715d06755af3d620c8395e1fc85226373c84c0dbadb8a9e400c4c2267c9f3293d2a2eabb3d7396da5b41159568a647a8cceec82376b34f3441b8df609f06012dca932461aa4ce46df8c5d831c029234d66ea72cde192fa7d8da7ba64752eb59;
    5'b11110 : xpb = 1024'h74f0c028afb4ec96cbba087644e8a349c051c0863dfce04699392d084061ec9ae8932a7e3b62c7c7aa7fbbe15b787090571fbee9e8f1f8e3ba37787378da1efb366cfda46f6517100abfbaabbfa4bb303dabceecb540b1cd06e7e4b5e6f72e4af61bd56129a74552dc93600857a9e3841f0bbadc88a092707f763bd10af24673;
    5'b11111 : xpb = 1024'h8f16ffc43463971fc9aa33ecdea6a7f07679a411f4213307948e3d24016b19276c8071c56efd39ea91da299d70dadf2d65d09dff45596dd83c365664f17d61bbb6097ee7b61f76d5d31615b8fe34db4fa83b7bea69001961427a97b09d359f0e086e65287e0c3d152da7bae9b810eaa18ceefa9e2dc9808dfa280f745af3b22;
    endcase
end

endmodule

module xpb_5_780
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h15ee98e055c3b100969a71dea06f6f0d795f549c70e736513e66c35d197b7c729f9aa21fc932ed2d5d6e8134a1b70c9096ca951e22bf752f1f5b2cff7d60b2b5135f3bb4d5a5709235939753fa3ecef048f7e973b3525043857d9eb65b2dbfec9b152d068933324774176560750fb8c7b14cfde9fd40b7e06724c4a52da62a3a;
    5'b00010 : xpb = 1024'h2bdd31c0ab8762012d34e3bd40dede1af2bea938e1ce6ca27ccd86ba32f6f8e53f35443f9265da5abadd0269436e19212d952a3c457eea5e3eb659fefac1656a26be7769ab4ae1246b272ea7f47d9de091efd2e766a4a0870afb3d6cb65b7fd9362a5a0d1266648ee82ecac0ea1f718f6299fbd3fa816fc0ce49894a5b4c5474;
    5'b00011 : xpb = 1024'h41cbcaa1014b1301c3cf559be14e4d286c1dfdd552b5a2f3bb344a174c727557decfe65f5b98c788184b839de52525b1c45fbf5a683e5f8d5e1186fe7822181f3a1db31e80f051b6a0bac5fbeebc6cd0dae7bc5b19f6f0ca9078dc2311893fc5d13f87139b9996d65c4630215f2f2a5713e6f9bdf7c227a1356e4def88f27eae;
    5'b00100 : xpb = 1024'h57ba6381570ec4025a69c77a81bdbc35e57d5271c39cd944f99b0d7465edf1ca7e6a887f24cbb4b575ba04d286dc32425b2a54788afdd4bc7d6cb3fdf582cad44d7ceed35695c248d64e5d4fe8fb3bc123dfa5cecd49410e15f67ad96cb6ffb26c54b41a24ccc91dd05d9581d43ee31ec533f7a7f502df819c931294b698a8e8;
    5'b00101 : xpb = 1024'h6da8fc61acd27502f1043959222d2b435edca70e34840f963801d0d17f696e3d1e052a9eedfea1e2d328860728933ed2f1f4e996adbd49eb9cc7e0fd72e37d8960dc2a882c3b32db0be1f4a3e33a0ab16cd78f42809b91519b74198fc7e4bf9f0769e120adfffb654474fae2494e9be67680f591f243976203b7d739e43ed322;
    5'b00110 : xpb = 1024'h8397954202962603879eab37c29c9a50d83bfbaaa56b45e77668942e98e4eaafbd9fccbeb7318f103097073bca4a4b6388bf7eb4d07cbf1abc230dfcf044303e743b663d01e0a36d41758bf7dd78d9a1b5cf78b633ede19520f1b84623127f8ba27f0e2737332dacb88c6042be5e54ae27cdf37bef844f426adc9bdf11e4fd5c;
    5'b00111 : xpb = 1024'h99862e225859d7041e391d16630c095e519b504716527c38b4cf578bb26067225d3a6ede80647c3d8e0588706c0157f41f8a13d2f33c3449db7e3afc6da4e2f3879aa1f1d78613ff7709234bd7b7a891fec76229e74031d8a66f56fc7e403f783d943b2dc0665ff42ca3c5a3336e0d75d91af165ecc50722d20160843f8b2796;
    5'b01000 : xpb = 1024'haf74c702ae1d8804b4d38ef5037b786bcafaa4e38739b289f3361ae8cbdbe394fcd510fe4997696aeb7409a50db86484b654a8f115fba978fad967fbeb0595a89af9dda6ad2b8491ac9cba9fd1f6778247bf4b9d9a92821c2becf5b2d96dff64d8a968344999923ba0bb2b03a87dc63d8a67ef4fea05bf03392625296d3151d0;
    5'b01001 : xpb = 1024'h14b61a8d41f3043c806888fc9390a027d2e3f64f22a94863b3c024f03254b2ff992735a548a3d809a9844b92cc11604ae905162916084e5c6995559d2d93d3ac3a09e4acd33ff7decf964f51335982419cb23b78c15ea54efbde026e7a711cbf44b703112203cbf58e12a98525bd58dbecdb0e5796fb19b359db6eca11f5159f;
    5'b01010 : xpb = 1024'h2aa4b36d97b6b53d1702fadb34000f354c434aeb93907eb4f226e84d4bd02f7238c1d7c511d6c53706f2ccc76dc86cdb7fcfab4738c7c38b88f0829caaf486614d692061a8e568710529e6a52d985131e5aa24ec74b0f592815ba124d59edcabdfcc3017ab36fe3d022a0ee59acd11a39e280c41943bd193c100336f3f9b3fd9;
    5'b01011 : xpb = 1024'h40934c4ded7a663dad9d6cb9d46f7e42c5a29f880477b506308dabaa654babe4d85c79e4db09b26464614dfc0f7f796c169a40655b8738baa84baf9c2855391660c85c167e8ad9033abd7df927d720222ea20e60280345d606d93fdb30cc9c987ae15d1e346a3084764174460fdcca6b4f750a2b917c89742824f8146d416a13;
    5'b01100 : xpb = 1024'h5681e52e433e173e4437de9874deed503f01f424755eeb576ef46f077ec7285777f71c04a43c9f91c1cfcf30b13685fcad64d5837e46ade9c7a6dc9ba5b5ebcb742797cb543049957051154d2215ef127799f7d3db5596198c56de918bfa5c8515f68a24bd9d62cbea58d9a684ec833300c208158ebd41548f49bcb99ae7944d;
    5'b01101 : xpb = 1024'h6c707e0e9901c83edad25077154e5c5db86148c0e64621a8ad5b32649842a4ca1791be246d6f8cbf1f3e506552ed928d442f6aa1a1062318e702099b23169e808786d38029d5ba27a5e4aca11c54be02c091e1478ea7e65d11d47d47e7281c71b10bb72b46d095135e703f06f9fc3bfab20f05ff8bfdf934f66e815ec88dbe87;
    5'b01110 : xpb = 1024'h825f16eeeec5793f716cc255b5bdcb6b31c09d5d572d57f9ebc1f5c1b1be213cb72c604436a279ec7cacd199f4a49f1ddaf9ffbfc3c59848065d369aa07751359ae60f34ff7b2ab9db7843f516938cf30989cabb41fa36a097521bfe4255dc5e4c20e431d003c75ad287a4676f0bf4c2635c03e9893eb1155d934603f633e8c1;
    5'b01111 : xpb = 1024'h984dafcf44892a4008073434562d3a78ab1ff1f9c8148e4b2a28b91ecb399daf56c70263ffd56719da1b52ce965babae71c494dde6850d7725b8639a1dd803eaae454ae9d5209b4c110bdb4910d25be35281b42ef54c86e41ccfbab49d839c4ae73611385936f9a2469f09c7e41bad8a14a901d3867f68f5c4b80aa923da12fb;
    5'b10000 : xpb = 1024'hae3c48af9a4cdb409ea1a612f69ca986247f469638fbc49c688f7c7be4b51a21f661a483c90854473789d4033812b83f088f29fc094482a6451390999b38b69fc1a4869eaac60bde469f729d0b112ad39b799da2a89ed727a24d596af8b15c37824b3e3ee26a2be9bab66f28592b6651c5f5ffbd83c020d62bdccf4e51803d35;
    5'b10001 : xpb = 1024'h137d9c3a2e2257786a36a01a86b1d1422c689801d46b5a76291986834b2de98c92b3c92ac814c2e5f59a15f0f66bb4053b3f973409512789b3cf7e3addc6f4a360b48da4d0da7f2b6999074e6c743592f06c8d7dcf6afa5a723e662699b47991ee58d91bbad465a3a80deda9d66af8f028691ec530b57b864c9218eef6440104;
    5'b10010 : xpb = 1024'h296c351a83e6087900d111f92721404fa5c7ec9e455290c7678049e064a965ff324e6b4a9147b013530897259822c095d20a2c522c109cb8d32aab3a5b27a7587413c959a67fefbd9f2c9ea266b30483396476f182bd4a9df7bc04dcf4e2397e896e0622440797eb1c25530a4b7ab1b7d9b61caf2df63366b3b6dd9423ea2b3e;
    5'b10011 : xpb = 1024'h3f5acdfad9a9b979976b83d7c790af5d1f27413ab639c718a5e70d3d7e24e271d1e90d6a5a7a9d40b077185a39d9cd2668d4c1704ed011e7f285d839d8885a0d8773050e7c25604fd4c035f660f1d373825c6065360f9ae17d39a393500ff96b24833328cd3aca32903cb86ac08a6a7f8b031a992b36eb471adba23951905578;
    5'b10100 : xpb = 1024'h554966db2f6d6a7a2e05f5b668001e6a988695d72720fd69e44dd09a97a05ee47183af8a23ad8a6e0de5998edb90d9b6ff9f568e718f871711e1053955e90cc29ad240c351cad0e20a53cd4a5b30a263cb5449d8e961eb2502b74249ab3db957bf98602f566dfc7a04541dcb359a23473c5018832877a327820066de7f367fb2;
    5'b10101 : xpb = 1024'h6b37ffbb85311b7ac4a06795086f8d7811e5ea73980833bb22b493f7b11bdb57111e51a9ece0779b6b541ac37d47e6479669ebac944efc46313c3238d349bf77ae317c78277041743fe7649e556f7154144c334c9cb43b688834e100066b79445aad8d35dfa12ec1786b832baaa9dc0eed9d166d25b85b07e9252b83acdca9ec;
    5'b10110 : xpb = 1024'h8126989bdaf4cc7b5b3ad973a8defc858b453f1008ef6a0c611b5754ca9757c9b0b8f3c9b61364c8c8c29bf81efef2d82d3480cab70e717550975f3850aa722cc190b82cfd15b206757afbf24fae40445d441cc050068bac0db27fb661993930f5c2ba3c68d46108ec82e88c1fb994d69eea145722f912e85049f028da82d426;
    5'b10111 : xpb = 1024'h9715317c30b87d7bf1d54b52494e6b9304a493ac79d6a05d9f821ab1e412d43c505395e97f4651f626311d2cc0b5ff68c3ff15e8d9cde6a46ff28c37ce0b24e1d4eff3e1d2bb2298ab0e934649ed0f34a63c06340358dbef93301e6cbcc6f91d90d7e742f2079350609a4dec94c94d9e503712412039cac8b76eb4ce0828fe60;
    5'b11000 : xpb = 1024'had03ca5c867c2e7c886fbd30e9bddaa07e03e848eabdd6aedde8de0efd8e50aeefee380948793f23839f9e61626d0bf95ac9ab06fc8d5bd38f4db9374b6bd796e84f2f96a860932ae0a22a9a442bde24ef33efa7b6ab2c3318adbd2317f4b90a2bed14497b3ac597d4b1b34d09d906660184102b1d7a82a91e93797335cf289a;
    5'b11001 : xpb = 1024'h12451de71a51aab45404b73879d3025c85ed39b4862d6c889e72e816640720198c405cb04785adc241afe04f20c607bf8d7a183efc9a00b6fe09a6d88dfa159a875f369cce750678039bbf4ba58ee8e44426df82dd774f65e89ec9deb8f7d66497faaf2653a4ff51c20931ce8718990463f72f32ca6fdd593f48c313da92ec69;
    5'b11010 : xpb = 1024'h2833b6c770155bb4ea9f29171a427169ff4c8e50f714a2d9dcd9ab737d829c8c2bdafed010b89aef9f1e6183c27d14502444ad5d1f5975e61d64d3d80b5ac84f9abe7251a41a770a392f569f9fcdb7d48d1ec8f690c99fa96e1c689514259651330fdc2cdcd831993620972efc2851cc15442d1cc7b09539a66d87b9083916a3;
    5'b11011 : xpb = 1024'h3e224fa7c5d90cb581399af5bab1e07778abe2ed67fbd92b1b406ed096fe18fecb75a0efd9eb881cfc8ce2b8643420e0bb0f427b4218eb153cc000d788bb7b04ae1dae0679bfe79c6ec2edf39a0c86c4d616b26a441befecf39a074b6f53563dce250933660b63e0aa37fc8f71380a93c6912b06c4f14d1a0d924c5e35df40dd;
    5'b11100 : xpb = 1024'h5410e8881b9cbdb617d40cd45b214f84f20b3789d8e30f7c59a7322db07995716b10430fa31e754a59fb63ed05eb2d7151d9d79964d860445c1b2dd7061c2db9c17ce9bb4f65582ea4568547944b55b51f0e9bddf76e40307917a601ca81162a693a3639ef3e96281e4f61efe647c35b77de28f0c23204fa74b7110363856b17;
    5'b11101 : xpb = 1024'h69ff816871606eb6ae6e7eb2fb90be926b6a8c2649ca45cd980df58ac9f511e40aaae52f6c516277b769e521a7a23a01e8a46cb78797d5737b765ad6837ce06ed4dc2570250ac8c0d9ea1c9b8e8a24a568068551aac09073fe9544b825aed617044f63407871c86f9266c7505b577c23292b26dabf72bcdadbdbd5a8912b9551;
    5'b11110 : xpb = 1024'h7fee1a48c7241fb74508f0919c002d9fe4c9e0c2bab17c1ed674b8e7e3708e56aa45874f35844fa514d86656495946927f6f01d5aa574aa29ad187d600dd9323e83b6124fab039530f7db3ef88c8f395b0fe6ec55e12e0b78412e36e80dc96039f64904701a4fab7067e2cb0d06734eada7824c4bcb374bb43009a4dbed1bf8b;
    5'b11111 : xpb = 1024'h95dcb3291ce7d0b7dba362703c6f9cad5e29355f2b98b27014db7c44fcec0ac949e0296efeb73cd27246e78aeb105323163996f3cd16bfd1ba2cb4d57e3e45d8fb9a9cd9d055a9e545114b438307c285f9f65839116530fb09908224dc0a55f03a79bd4d8ad82cfe7a9592114576edb28bc522aeb9f42c9baa255ef2ec77e9c5;
    endcase
end

endmodule

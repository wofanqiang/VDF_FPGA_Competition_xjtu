module xpb_5_475
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha2b024067d7790dc0506c6f5b325c2c8baee409f263bdf301a779c995fbe81c499e11ce2cbc5c36ca4abcd597184ad9fcd3f76393f226210ce69be010baf472c2894b1663c4a8d3e950369643ebd7f181a26ab36f5bbbef6978e20f702b7df397f8510dc7832667b4335999a7674c9c8f87206b3de947e0d3cf52163c516dd13;
    5'b00010 : xpb = 1024'h94b302b73900ecef3f08161455f13e4004667e0d77001de8b7127fdd0c7a56813079bc4ccd65084aa9f95b6bffab4a753664c48c5b91f3d5ec343ca3dc8c19a6dcda2e1dc9041d38176cd025e49f39ff40485cd55ef150dc798faff34b451be0d0028f8f3f9bd468ffab4c55f5196d68a20a2e856cdd9eea337ac7c3014b53bb;
    5'b00011 : xpb = 1024'h86b5e167f48a490279096532f8bcb9b74ddebb7bc7c45ca153ad6320b9362b3dc7125bb6cf044d28af46e97e8dd1e74a9f8a12df7801859b09febb46ad68ec21911faad555bdad3199d636e78a80f4e6666a0e73c826e2c25b913eef93d2588820800e4207054256bc20ff1173be11084ba25656fb26bfc72a006e223d7fca63;
    5'b00100 : xpb = 1024'h78b8c018b013a515b30ab4519b88352e9756f8ea18889b59f048466465f1fffa5daafb20d0a39206b49477911bf8842008af61329471176027c939e97e45be9c4565278ce2773d2b1c3f9da93062afcd8c8bc012315c74a83d92cdebdc5f952f70fd8cf4ce6eb0447896b1ccf262b4a7f53a7e28896fe0a42086148179b4410b;
    5'b00101 : xpb = 1024'h6abb9ec96b9d0128ed0c03703e53b0a5e0cf3658694cda128ce329a812add4b6f4439a8ad242d6e4b9e205a3aa1f20f571d4af85b0e0a9254593b88c4f229116f9aaa4446f30cd249ea9046ad6446ab4b2ad71b09a92068e1f945ce824ecd1d6c17b0ba795d81e32350c6488710758479ed2a5fa17b90181170bbae0b5e8b7b3;
    5'b00110 : xpb = 1024'h5cbe7d7a27265d3c270d528ee11f2c1d2a4773c6ba1118cb297e0cebbf69a9738adc39f4d3e21bc2bf2f93b63845bdcadaf9fdd8cd503aea635e372f1fff6391adf020fbfbea5d1e21126b2c7c26259bd8cf234f03c798740195ebe46d7a0e7e11f88a5a5d418c1ff1821743efabfbe7486acdcba602225e0d91613ff21d2e5b;
    5'b00111 : xpb = 1024'h4ec15c2ae2afb94f610ea1ad83eaa79473bfb1350ad55783c618f02f6c257e302174d95ed58160a0c47d21c8c66c5aa0441f4c2be9bfccaf8128b5d1f0dc360c62359db388a3ed17a37bd1ee2207e082fef0d4ed6cfd2a59e3977ae0b6074b256276090d24aafa0dadf7c9ff6e509f86f202f59d344b433b0417079f2e51a503;
    5'b01000 : xpb = 1024'h40c43adb9e3915629b0ff0cc26b6230bbd37eea35b99963c62b3d37318e152ecb80d78c8d720a57ec9caafdb5492f775ad449a7f062f5e749ef33474c1b90887167b1a6b155d7d1125e538afc7e99b6a2512868bd632bc3fc59909dcfe9487ccb2f387bfec1467fb6a6d7cbaecf543269b9b1d6ec2946417fa9cadfe6a861bab;
    5'b01001 : xpb = 1024'h32c7198c59c27175d5113feac9819e8306b02c11ac5dd4f4ff4eb6b6c59d27a94ea61832d8bfea5ccf183dede2b9944b1669e8d2229ef039bcbdb3179295db01cac09722a2170d0aa84e9f716dcb56514b34382a3f684e25a79a98d94721c47403710672b37dd5e926e32f766b99e6c64533454050dd84f4f122545da6ba9253;
    5'b01010 : xpb = 1024'h24c9f83d154bcd890f128f096c4d19fa5028697ffd2213ad9be999fa7258fc65e53eb79cda5f2f3ad465cc0070e031207f8f37253f0e81feda8831ba6372ad7c7f0613da2ed09d042ab8063313ad11387155e9c8a89de00b899c27d58faf011b53ee85257ae743d6e358e231ea3e8a65eecb6d11df26a5d1e7a7fabce2ef08fb;
    5'b01011 : xpb = 1024'h16ccd6edd0d5299c4913de280f18957199a0a6ee4de6526638847d3e1f14d1227bd75706dbfe7418d9b35a12ff06cdf5e8b485785b7e13c3f852b05d344f7ff7334b9091bb8a2cfdad216cf4b98ecc1f97779b6711d371f16b9db6d1d83c3dc2a46c03d84250b1c49fce94ed68e32e05986394e36d6fc6aede2da11c1f237fa3;
    5'b01100 : xpb = 1024'h8cfb59e8c5e85af83152d46b1e410e8e318e45c9eaa911ed51f6081cbd0a5df126ff670dd9db8f6df00e8258d2d6acb51d9d3cb77eda589161d2f00052c5271e7910d494843bcf72f8ad3b65f708706bd994d057b0903d74d9f45ce20c97a69f4e9828b09ba1fb25c4447a8e787d1a541fbbcb4fbb8e78bd4b3477b5b57f64b;
    5'b01101 : xpb = 1024'hab7fd9a509d6168b881bf43c6509d3b19e0724fbc4e6704eef96fd1b2b8f27a3ac511353a9637c6383acb57efeb2186b1f194a04b7100799e486ed0110db999e1025beaf848e4a35c48e3d1a9e2e061ed7bff83c70c4c2cde52d66c5238159a3746e936781ec862d9f79e1435dfc9b6e3a6dc368da4d659911a868df206ed35e;
    5'b01110 : xpb = 1024'h9d82b855c55f729ec21d435b07d54f28e77f626a15aaaf078c31e05ed84afc6042e9b2bdab02c14188fa43918cd8b540883e9857d37f995f02516ba3e1b86c18c46b3b671147da2f46f7a3dc440fc105fde1a9dad9fa54b3c72ef5c16c0e964ac4ec121a4955f41b5bef93fedca13f0de405eb3a68968676082e0f3e5ca34a06;
    5'b01111 : xpb = 1024'h8f85970680e8ceb1fc1e9279aaa0caa030f79fd8666eedc028ccc3a28506d11cd9825227aca2061f8e47d1a41aff5215f163e6aaefef2b24201bea46b2953e9378b0b81e9e016a28c9610a9de9f17bed24035b79432fe699a93084bdb49bd2f2156990cd10bf6209186546ba5b45e2ad8d9e130bf6dfa752feb3b59d98d7c0ae;
    5'b10000 : xpb = 1024'h818875b73c722ac5361fe1984d6c46177a6fdd46b7332c78c567a6e631c2a5d9701af191ae414afd93955fb6a925eeeb5a8934fe0c5ebce93de668e98372110e2cf634d62abafa224bca715f8fd336d44a250d17ac65787f8b3213b9fd290f9965e70f7fd828cff6d4daf975d9ea864d37363add8528c82ff5395bfcd50c3756;
    5'b10001 : xpb = 1024'h738b5467f7fb86d8702130b6f037c18ec3e81ab507f76b3162028a29de7e7a9606b390fbafe08fdb98e2edc9374c8bc0c3ae835128ce4eae5bb0e78c544ee388e13bb18db7748a1bce33d82135b4f1bb7046beb6159b0a656d33a2b645b64c40b6648e329f923de49150ac31588f29ece0ce62af1371e90cebbf025c1140adfe;
    5'b10010 : xpb = 1024'h658e3318b384e2ebaa227fd593033d060d60582358bba9e9fe9d6d6d8b3a4f529d4c3065b17fd4b99e307bdbc57328962cd3d1a4453de073797b662f252bb60395812e45442e1a15509d3ee2db96aca2966870547ed09c4b4f3531b28e4388e806e20ce566fbabd24dc65eecd733cd8c8a668a80a1bb09e9e244a8bb4d7524a6;
    5'b10011 : xpb = 1024'h579111c96f0e3efee423cef435ceb87d56d89591a97fe8a29b3850b137f6240f33e4cfcfb31f1997a37e09ee5399c56b95f91ff761ad72389745e4d1f608887e49c6aafcd0e7aa0ed306a5a481786789bc8a21f2e8062e313136c0aed6d0c58f575f8b982e6519c00a3c11a855d8712c33feb25230042ac6d8ca4f1a89a99b4e;
    5'b10100 : xpb = 1024'h4993f07a2a979b121e251e12d89a33f4a050d2fffa44275b37d333f4e4b1f8cbca7d6f39b4be5e75a8cb9800e1c06240ff1e6e4a7e1d03fdb5106374c6e55af8fe0c27b45da13a0855700c66275a2270e2abd391513bc01713384fab1f5e0236a7dd0a4af5ce87adc6b1c463d47d14cbdd96da23be4d4ba3cf4ff579c5de11f6;
    5'b10101 : xpb = 1024'h3b96cf2ae620f72558266d317b65af6be9c9106e4b086613d46e1738916dcd8861160ea3b65da353ae1926136fe6ff166843bc9d9a8c95c2d2dae21797c22d73b251a46bea5aca01d7d97327cd3bdd5808cd852fba7151fcf539dea767eb3eddf85a88fdbd37f59b8327771f5321b86b872f01f54c966c80c5d59bd90212889e;
    5'b10110 : xpb = 1024'h2d99addba1aa53389227bc501e312ae333414ddc9bcca4cc7108fa7c3e29a244f7aeae0db7fce831b366b425fe0d9bebd1690af0b6fc2787f0a560ba689effee66972123771459fb5a42d9e9731d983f2eef36ce23a6e3e2d73b6da3b0787b8548d807b084a163893f9d29dad1c65c0b30c729c6dadf8d5dbc5b42383e46ff46;
    5'b10111 : xpb = 1024'h1f9c8c8c5d33af4bcc290b6ec0fca65a7cb98b4aec90e3850da3ddbfeae577018e474d77b99c2d0fb8b442388c3438c13a8e5943d36bb94d0e6fdf5d397bd2691adc9ddb03cde9f4dcac40ab18ff53265510e86c8cdc75c8b93cfc9ff905b82c995586634c0ad176fc12dc96506affaada5f51986928ae3ab2e0e8977a7b75ee;
    5'b11000 : xpb = 1024'h119f6b3d18bd0b5f062a5a8d63c821d1c631c8b93d55223daa3ec10397a14bbe24dfece1bb3b71edbe01d04b1a5ad596a3b3a796efdb4b122c3a5e000a58a4e3cf221a92908779ee5f15a76cbee10e0d7b329a0af61207ae9b3e8b9c4192f4d3e9d3051613743f64b8888f51cf0fa34a83f77969f771cf17a9668ef6b6afec96;
    5'b11001 : xpb = 1024'h3a249edd4466772402ba9ac06939d490faa06278e1960f646d9a447445d207abb788c4bbcdab6cbc34f5e5da881726c0cd8f5ea0c4adcd74a04dca2db35775e8367974a1d4109e7e17f0e2e64c2c8f4a1544ba95f4799947d401a988a20317b3a5083c8daddad5274fe420d4db446ea2d8fa13b85baeff49fec3555f2e4633e;
    5'b11010 : xpb = 1024'ha6526df451bdf84e453270a1b9b96011ca9846c6b4554026615140e0a41ba23f5559a92e88a07a3867fb2bb71a06200bda186c234b6d3ee8186e9aa3e6e4be8aabfc48b0598b972676827792a380480cbb7af6e05503588b14ce3b8f8cd810b4b9d594a5531013cdb833dba7c42910b32601a7ef644f6e01dce156b9b7fb4051;
    5'b11011 : xpb = 1024'h98554ca50d4754617f33bfc05c84db891410843505197edefdec242450d776fbebf248988a3fbf166d48b9c9a82cbce1433dba7667dcd0ad36391946b7c191056041c567e645271ff8ebde54496202f3e19ca87ebe38ea70f6cfca8bd5654d5c0a5313581a7981bb74a98e6342cdb452cf99cfc0f2988eded366fd18f42fb6f9;
    5'b11100 : xpb = 1024'h8a582b55c8d0b074b9350edeff5057005d88c1a355ddbd979a870767fd934bb8828ae8028bdf03f4729647dc365359b6ac6308c9844c6272540397e9889e63801487421f72feb7197b554515ef43bddb07be5a1d276e7c56d8d159881df28a035ad0920ae1e2efa9311f411ec17257f27931f79280e1afbbc9eca37830642da1;
    5'b11101 : xpb = 1024'h7c5b0a06845a0c87f3365dfda21bd277a700ff11a6a1fc503721eaabaa4f20751923876c8d7e48d277e3d5eec479f68c1588571ca0bbf43771ce168c597b35fac8ccbed6ffb84712fdbeabd7952578c22de00bbb90a40e3cbad2e884667fc6aaab4e10bda94c5d96ed94f3da4016fb9222ca1f640f2ad098c07249d76c98a449;
    5'b11110 : xpb = 1024'h6e5de8b73fe3689b2d37ad1c44e74deef0793c7ff7663b08d3bccdef570af531afbc26d68f1d8db07d31640152a093617eada56fbd2b85fc8f98952f2a5808757d123b8e8c71d70c802812993b0733a95401bd59f9d9a0229cd47780af0d0351fbcb8f7070b5cb84aa0aa695bebb9f31cc6247359d73f175b6f7f036a8cd1af1;
    5'b11111 : xpb = 1024'h6060c767fb6cc4ae6738fc3ae7b2c96639f179ee482a79c17057b13303c6c9ee4654c64090bcd28e827ef213e0c73036e7d2f3c2d99b17c1ad6313d1fb34daf03157b846192b67060291795ae0e8ee907a236ef8630f32087ed6067cf79a3ff94c490e23381f3972668059513d6042d175fa6f072bbd1252ad7d9695e5019199;
    endcase
end

endmodule

module xpb_5_135
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hfb3a999adf61c967399c4eb54e2ed0a52e2575e9db1987fad14c1a17e5486bc7e1381a0993096e8dae6cfbaf6fbd0d25ee8d063ef5d9acdb777e7924360078b7aa427098ed50a5048e622b87bcfd255796478c6009e35ac3640cd30468864dab7305d3ca6e080fce5bdedb3a64dae8fecf940bd3bd3bbcbea199d3195e4400e;
    5'b00010 : xpb = 1024'h1f6753335bec392ce73389d6a9c5da14a5c4aebd3b6330ff5a298342fca90d78fc27034132612dd1b5cd9f75edf7a1a4bdd1a0c7debb359b6eefcf2486c00f16f5484e131daa14a091cc4570f79fa4aaf2c8f18c013c6b586c819a608d10c9b56e60ba794dc101f9cb7bdb674c9b5d1fd9f2817a77a77797d4333a632bc8801c;
    5'b00011 : xpb = 1024'h2f1afccd09e255c35acd4ec1fea8c71ef8a7061bd914c97f073e44e47afd94357a3a84e1cb91c4ba90b46f30e4f372771cba712bce18d0692667b6b6ca2016a26fec751cac7f1ef0dab26829736f77006c2d6a5201daa104a2c26790d3992e90259117b5f4a182f6b139c91af2e90bafc6ebc237b37b3363be4cd794c1acc02a;
    5'b00100 : xpb = 1024'h3ecea666b7d87259ce6713ad538bb4294b895d7a76c661feb4530685f9521af1f84e068264c25ba36b9b3eebdbef43497ba3418fbd766b36dddf9e490d801e2dea909c263b54294123988ae1ef3f4955e591e3180278d6b0d90334c11a21936adcc174f29b8203f396f7b6ce9936ba3fb3e502f4ef4eef2fa86674c657910038;
    5'b00101 : xpb = 1024'h4e82500065ce8ef04200d898a86ea1339e6bb4d91477fa7e6167c82777a6a1ae76618822fdf2f28c46820ea6d2eb141bda8c11f3acd40604955785db50e025b96534c32fca2933916c7ead9a6b0f1bab5ef65bde03170c5d0f4401f160a9f84593f1d22f426284f07cb5a4823f8468cfa0de43b22b22aafb928011f7ed754046;
    5'b00110 : xpb = 1024'h5e35f99a13c4ab86b59a9d83fd518e3df14e0c37b22992fe0e7c89c8f5fb286af47509c3972389752168de61c9e6e4ee3974e2579c31a0d24ccf6d6d94402d44dfd8ea3958fe3de1b564d052e6deee00d85ad4a403b542094584cf21a7325d204b222f6be94305ed62739235e5d2175f8dd7846f66f666c77c99af2983598054;
    5'b00111 : xpb = 1024'h6de9a333c1bac81d2934626f52347b48443063964fdb2b7dbb914b6a744faf2772888b643054205dfc4fae1cc0e2b5c0985db2bb8b8f3ba0044754ffd7a034d05a7d1142e7d34831fe4af30b62aec05651bf4d6a045377b57bc59c51edbac1fb02528ca8902386ea48317fe98c1fc5ef7ad0c52ca2ca229366b34c5b193dc062;
    5'b01000 : xpb = 1024'h7d9d4ccd6fb0e4b39cce275aa71768529712baf4ed8cc3fd68a60d0bf2a435e3f09c0d04c984b746d7367dd7b7de8692f746831f7aecd66dbbbf3c921b003c5bd521384c76a85282473115c3de7e92abcb23c63004f1ad61b2066982344326d5b982e9e5370407e72def6d9d326d747f67ca05e9de9dde5f50cce98caf220070;
    5'b01001 : xpb = 1024'h8d50f6671da7014a1067ec45fbfa555ce9f512538b3e5c7d15bacead70f8bca06eaf8ea562b54e2fb21d4d92aeda5765562f53836a4a713b733724245e6043e74fc55f56057d5cd29017387c5a4e650144883ef6058fe30de84736b27acb8bb070b34721dde488e413ad5b50d8bb230f54c346a71a719a2b3ae686be4506407e;
    5'b01010 : xpb = 1024'h9d04a000cb9d1de08401b13150dd42673cd769b228eff4fcc2cf904eef4d435cecc31045fbe5e5188d041d4da5d62837b51823e759a80c092aaf0bb6a1c04b72ca69865f94526722d8fd5b34d61e3756bdecb7bc062e18ba1e8803e2c153f08b27e3a45e84c509e0f96b49047f08d19f41bc8764564555f7250023efdaea808c;
    5'b01011 : xpb = 1024'hacb8499a79933a76f79b761ca5c02f718fb9c110c6a18d7c6fe451f06da1ca196ad691e695167c0167eaed089cd1f90a1400f44b4905a6d6e226f348e52052fe450dad692327717321e37ded51ee09ac3751308206cc4e6654c8d11307dc5565df14019b2ba58adddf2936b82556802f2eb5c821921911c30f19c12170cec09a;
    5'b01100 : xpb = 1024'hbbeadde659b2244a02fc330ea48d52a7126153e8edb85849f1c5a3c38f3a3cde5a1960e6420945ba3737d7cb06fb9120ecf9cc915b07158e8ff9b7cedade5d84b629fc4026b7e7e582f9e0334e217d0bcb0afaf7ae45701d57d0c48943a17ae673cccae21bd134d3e273d8cd3d40895ccd529fc7da1705eb2c3e34e7dd09a3d;
    5'b01101 : xpb = 1024'h1b72577813913edb13c9881c3f2bc234c4086c9d2c8d1e044c311bddb7482a8a63b517aefd512b447e5a4d37a76b89e46db86d2d050e0c26a077830f310ded63c606c6cd914088cea115c0bbb0b1ea26361528757b828cae0bbdd978dac27c891e6d29eac89d944a23e52b407a21b725b9ce6ab9b9752c2a9cdd808013b4da4b;
    5'b01110 : xpb = 1024'h2b260111c1875b7187634d07940eaf3f16eac3fbca3eb683f945dd7f359cb146e1c8994f9681c22d59411cf29e675ab6cca13d90f46ba6f457ef6aa1746df4ef40aaedd72015931ee9fbe3742c81bc7baf79a13b7c20c25a41fea6a9214ae163d59d87276f7e154709a318f4206f65b5a6c7ab76f548e7f686f71db1a9991a59;
    5'b01111 : xpb = 1024'h3ad9aaab6f7d7807fafd11f2e8f19c4969cd1b5a67f04f03a65a9f20b3f138035fdc1af02fb259163427ecad95632b892b8a0df4e3c941c20f675233b7cdfc7abb4f14e0aeea9d6f32e2062ca8518ed128de1a017cbef806783f73d967d3463e8ccde464165e9643ef6106a7c6bd144593c0ec34311ca3c27110bae33f7d5a67;
    5'b10000 : xpb = 1024'h4a8d54451d73949e6e96d6de3dd48953bcaf72b905a1e783536f60c23245bebfddef9c90c8e2efff0f0ebc688c5efc5b8a72de58d326dc8fc6df39c5fb2e040635f33bea3dbfa7bf7bc828e524216126a24292c77d5d2db2ae804109ae5bab1943fe41a0bd3f1740d51ef45b6d0ac2d580ba2cf16cf05f8e5b2a5814d5619a75;
    5'b10001 : xpb = 1024'h5a40fddecb69b134e2309bc992b7765e0f91ca17a353800300842263b09a457c5c031e31621386e7e9f58c23835acd2de95baebcc284775d7e5721583e8e0b91b09762f3cc94b20fc4ae4b9d9ff1337c1ba70b8d7dfb635ee4c10e39f4e40ff3fb2e9edd641f983dbadce20f135871656db36daea8c41b5a4543f5466b45da83;
    5'b10010 : xpb = 1024'h69f4a778795fcdcb55ca60b4e79a63686274217641051882ad98e4052eeecc38da169fd1fb441dd0c4dc5bde7a569e0048447f20b1e2122b35cf08ea81ee131d2b3b89fd5b69bc600d946e561bc105d1950b84537e99990b1b01db6a3b6c74ceb25efc1a0b00193aa09acfc2b9a61ff55aacae6be497d7262f5d9278012a1a91;
    5'b10011 : xpb = 1024'h79a851122755ea61c96425a03c7d5072b55678d4deb6b1025aada5a6ad4352f5582a21729474b4b99fc32b9971526ed2a72d4f84a13facf8ed46f07cc54e1aa8a5dfb106ea3ec6b0567a910e9790d8270e6ffd197f37ceb75142a89a81f4d9a9698f5956b1e09a378658bd765ff3ce8547a5ef29206b92f219772fa9970e5a9f;
    5'b10100 : xpb = 1024'h895bfaabd54c06f83cfdea8b91603d7d0838d0337c68498207c267482b97d9b1d63da3132da54ba27aa9fb54684e3fa506161fe8909d47c6a4bed80f08ae22342083d8107913d1009f60b3c71360aa7c87d475df7fd60463878375cac87d3e8420bfb69358c11b346c16ab2a06417d15349f2fe65c3f4ebe0390ccdb2cf29aad;
    5'b10101 : xpb = 1024'h990fa4458342238eb097af76e6432a875b1b27921a19e201b4d728e9a9ec606e545124b3c6d5e28b5590cb0f5f4a107764fef04c7ffae2945c36bfa14c0e29bf9b27ff1a07e8db50e846d67f8f307cd20138eea580743a0fbdc442fb0f05a35ed7f013cfffa19c3151d498ddac8f2ba5219870a398130a89edaa6a0cc2d6dabb;
    5'b10110 : xpb = 1024'ha8c34ddf31384025243174623b261791adfd7ef0b7cb7a8161ebea8b2840e72ad264a6546006797430779aca5645e149c3e7c0b06f587d6213aea7338f6e314b15cc262396bde5a1312cf9380b004f277a9d676b81126fbbf405102b558e08398f20710ca6821d2e3792869152dcda350e91b160d3e6c655d7c4073e58bb1ac9;
    5'b10111 : xpb = 1024'h7c9b2231d4027f2ccc5c1767faebd4a8f69d31e800572899123f2d6f392c0df4d2faa7c2f1091ce6c002b3e69e3a151beb6692e3c0347e41a874f6797fbc4251c21187e7601f2ac6779194dedf45d4bfffce698f52a785774b94b60e1ebca8217493c1f9c99a59d96908d66015a629bacb1133bbf6f24f17b6e296b65bcf46c;
    5'b11000 : xpb = 1024'h177d5bbccb364489405f8661d491aa54e24c2a7d1db70b093e38b47871e7479bcb432c1cc84128b746e6faf960df72241d9f39922b60e2b1d1ff36f9db5bcbb096c53f8804d6fcfcb05f3c0669c42fa179615f5ef5c8ae03aafa189128742f5cce79995c437a269a7c4e7b19a7a8112b99aa53f8fb42e0bd6587c69cfba1347a;
    5'b11001 : xpb = 1024'h27310556792c611fb3f94b4d2974975f352e81dbbb68a388eb4d7619f03bce584956adbd6171bfa021cdcab457db42f67c8809f61abe7d7f89771e8c1ebbd33c1169669193ac074cf9455ebee59401f6f2c5d824f666e3afe13ae5c16efc943785a9f698ea5aa797620c68cd4df5bfbb86a394b637169c894fa163ce91857488;
    5'b11010 : xpb = 1024'h36e4aef027227db6279310387e5784698810d93a591a3c08986237bb6e905514c76a2f5dfaa25688fcb49a6f4ed713c8db70da5a0a1c184d40ef061e621bdac78c0d8d9b2281119d422b81776163d44c6c2a50eaf705195c177bb2f1b584f9123cda53d5913b289447ca5680f4436e4b739cd57372ea585539bb01002769b496;
    5'b11011 : xpb = 1024'h46985889d5189a4c9b2cd523d33a7173daf33098f6cbd4884576f95cece4dbd1457db0fe93d2ed71d79b6a2a45d2e49b3a59aabdf979b31af866edb0a57be25306b1b4a4b1561bed8b11a42fdd33a6a1e58ec9b0f7a34f084dbc8021fc0d5decf40ab112381ba9912d8844349a911cdb60961630aebe142123d49e31bd4df4a4;
    5'b11100 : xpb = 1024'h564c0223830eb6e30ec69a0f281d5e7e2dd587f7947d6d07f28bbafe6b39628dc391329f2d03845ab28239e53cceb56d99427b21e8d74de8afded542e8dbe9de8155dbae402b263dd3f7c6e8590378f75ef34276f84184b483fd4d524295c2c7ab3b0e4edefc2a8e134631e840decb6b4d8f56edea91cfed0dee3b63533234b2;
    5'b11101 : xpb = 1024'h65ffabbd3104d37982605efa7d004b8880b7df56322f05879fa07c9fe98de94a41a4b43fc6341b438d6909a033ca863ff82b4b85d834e8b66756bcd52c3bf169fbfa02b7cf00308e1cdde9a0d4d34b4cd857bb3cf8dfba60ba3e1a82891e27a2626b6b8b85dcab8af9041f9be72c79fb3a8897ab26658bb8f807d894e91674c0;
    5'b11110 : xpb = 1024'h75b35556defaf00ff5fa23e5d1e33892d39a36b4cfe09e074cb53e4167e27006bfb835e05f64b22c684fd95b2ac6571257141be9c79283841ecea4676f9bf8f5769e29c15dd53ade65c40c5950a31da251bc3402f97df00cf07ee7b2cfa68c7d199bc8c82cbd2c87dec20d4f8d7a288b2781d86862394784e22175c67efab4ce;
    5'b11111 : xpb = 1024'h8566fef08cf10ca66993e8d126c6259d267c8e136d923686f9c9ffe2e636f6c33dcbb780f89549154336a91621c227e4b5fcec4db6f01e51d6468bf9b2fc0080f14250caecaa452eaeaa2f11cc72eff7cb20acc8fa1c25b926bfb4e3162ef157d0cc2604d39dad84c47ffb0333c7d71b147b19259e0d0350cc3b12f814def4dc;
    endcase
end

endmodule

module xpb_5_5
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h40dd8a97273283eb8504775b0fc72f5d9ccb6d39a4812a876256b299d584e88f68f9744bad15425f5d10a1432518fba2034cd4a5c3de926643629d116e2f081d19c4889c73f27d96a85386c88882bf34271b2696bfe3e6ff60bdc4f28c56c9bb8ca3bc823be35691c98483ef78992493d4d9f3559275415357f7e52f675198c6;
    5'b00010 : xpb = 1024'h81bb152e4e6507d70a08eeb61f8e5ebb3996da734902550ec4ad6533ab09d11ed1f2e8975a2a84beba2142864a31f7440699a94b87bd24cc86c53a22dc5e103a33891138e7e4fb2d50a70d9111057e684e364d2d7fc7cdfec17b89e518ad93771947790477c6ad23930907def1324927a9b3e6ab24ea82a6afefca5ecea3318c;
    5'b00011 : xpb = 1024'h11eb5a6fb3a956f9c407ee3a1efb46c764ec447c180bdf1ea9275e77cd8c0ca637a3df6a3d19488f77d3a4828bece21ba5cc560b28e8e6e7198897d60fbaa3a5d8fe6526ac467b7ee66091b700ac796b814c7a2bb32587ed6cacbcdcead9baa076e3a35d02e10b27d5cda4ef71fb47922fb3fb1e671466c9c1783489ad1263e7;
    5'b00100 : xpb = 1024'h52c8e506dadbdae5490c65952ec2762501b7b1b5bc8d09a60b7e1111a310f535a09d53b5ea2e8aeed4e445c5b105ddbda9192ab0ecc7794d5ceb34e77de9abc2f2c2edc32038f9158eb4187f892f389fa867a0c273096eeccd6a81cf7730845c03875fdf3ec461b99f5228deea946c26048dee73f989a81d197019b91463fcad;
    5'b00101 : xpb = 1024'h93a66f9e020e5ed0ce10dcf03e89a5829e831eef610e342d6dd4c3ab7895ddc50996c8019743cd4e31f4e708d61ed95fac65ff56b0a60bb3a04dd1f8ec18b3e00c87765f942b76ac37079f4811b1f7d3cf82c75932ed55ec2e2846c203874e17902b1c617aa7b84b68d6acce632d90b9d967e1c98bfee9707167fee87bb59573;
    5'b00110 : xpb = 1024'h23d6b4df6752adf3880fdc743df68d8ec9d888f83017be3d524ebcef9b18194c6f47bed47a32911eefa7490517d9c4374b98ac1651d1cdce33112fac1f75474bb1fcca4d588cf6fdccc1236e0158f2d70298f457664b0fdad95979b9d5b37540edc746ba05c2164fab9b49dee3f68f245f67f63cce28cd9382f069135a24c7ce;
    5'b00111 : xpb = 1024'h64b43f768e8531df0d1453cf4dbdbcec66a3f631d498e8c4b4a56f89709d01dbd84133202747d37e4cb7ea483cf2bfd94ee580bc15b060347673ccbd8da44f68cbc152e9cc7f74947514aa3689dbb20b29b41aee262ef6da3a173eac620a3efc7a6b033c41a56ce1751fcdce5c8fb3b83441e992609e0ee6dae84e42c1766094;
    5'b01000 : xpb = 1024'ha591ca0db5b7b5ca9218cb2a5d84ec4a036f636b791a134c16fc22234621ea6b413aa76bd45d15dda9c88b8b620bbb7b52325561d98ef29ab9d669cefbd35785e585db864071f22b1d6830ff125e713f50cf4184e612ddd99ad5039eee6108b8070ebfbe7d88c3733ea451bdd528d84c091bdce7f313503a32e0337228c7f95a;
    5'b01001 : xpb = 1024'h35c20f4f1afc04ed4c17caae5cf1d4562ec4cd7448239d5bfb761b6768a425f2a6eb9e3eb74bd9ae677aed87a3c6a652f16502217abab4b54c99c7822f2feaf18afb2f7404d3727cb321b52502056c4283e56e83197097c846063696c08d2fe164aaea1708a321778168eece55f1d6b68f1bf15b353d345d44689d9d07372bb5;
    5'b01010 : xpb = 1024'h769f99e6422e88d8d11c42096cb903b3cb903aadeca4c7e35dccce013e290e820fe5128a64611c0dc48b8ecac8dfa1f4f4b1d6c73e99471b8ffc64939d5ef30ea4bfb81078c5f0135b753bed8a882b76ab009519d9547ec7a6c3fb894ce3f99cf14ea699448678094aed72bdce8afb4a63f5e4b0c7b275b09c6082cc6e88c47b;
    5'b01011 : xpb = 1024'h6cfdf27a772d7fb8b1b418d6c25ebbff6e5a4b6bbae51f34246c74560ab4a097596095d474fdfde823df0c70a9a8ccc93e48386dfc5093622bfc246d0bb867a4a350bfe3d277064f12ec0137a2f2679de16c2180cb238b651f52e811f1020c64eead0f1cfa0d60d8db20fce4f53f9b4e9f5f92409dc59d3ade8ecf74cf7f6d6;
    5'b01100 : xpb = 1024'h47ad69becea55be7101fb8e87bed1b1d93b111f0602f7c7aa49d79df36303298de8f7da8f465223ddf4e920a2fb3886e9731582ca3a39b9c66225f583eea8e9763f9949ab119edfb998246dc02b1e5ae0531e8aecc961fb5b2b2f373ab66ea81db8e8d740b842c9f573693bdc7ed1e48becfec799c519b2705e0d226b4498f9c;
    5'b01101 : xpb = 1024'h888af455f5d7dfd2952430438bb44a7b307c7f2a04b0a70206f42c790bb51b284788f1f4a17a649d3c5f334d54cc84109a7e2cd267822e02a984fc69ad1996b47dbe1d37250c6b9241d5cda48b34a4e22c4d0f458c7a06b51370b86637bdb43d683249f64767833120bb17ad408642dc93a9dfcf2ec6dc7a5dd8b7561b9b2862;
    5'b01110 : xpb = 1024'h18bb39975b1c2ef54f232fc78b2132875bd1e932d3ba3111eb6e25bd2e3756afad39e8c78469286dfa11954996876ee839b0d99208adf01d3c485a1ce0762a2023337124e96debe3d78f51ca7adb9fe55f633c43bfd7c0a3bea1eb5e09e9db66c5ce744ed281e135637fb4bdc14f414719a9f44270f0c09d6f612180fa0a5abd;
    5'b01111 : xpb = 1024'h5998c42e824eb2e0d427a7229ae861e4f89d566c783b5b994dc4d85703bc3f3f16335d13317e6acd5722368cbba06a8a3cfdae37cc8c82837faaf72e4ea5323d3cf7f9c15d60697a7fe2d893035e5f19867e62da7fbba7a31f5fb0509640a522527230d10e6537c72d0438ad39e865daee83e798036601f0c75906b0615bf383;
    5'b10000 : xpb = 1024'h9a764ec5a98136cc592c1e7daaaf91429568c3a61cbc8620b01b8af0d94127ce7f2cd15ede93ad2cb432d7cfe0b9662c404a82dd906b14e9c30d943fbcd43a5a56bc825dd152e71128365f5b8be11e4dad9989713f9f8ea2801d754322976edddf15ed534a488e58f688bc9cb2818a6ec35ddaed95db43441f50ebdfc8ad8c49;
    5'b10001 : xpb = 1024'h2aa694070ec585ef132b1e01aa1c794ec0be2daeebc6103094958434fbc36355e4ddc831c18270fd71e539cc22745103df7d2f9d3196d70455d0f1f2f030cdc5fc31d64b95b46762bdefe3817b881950e0afb66f72fd48912b4ea83af4c396073cb217abd562ec5d394d59ad334a88d9495def60d805276730d9560aa71cbea4;
    5'b10010 : xpb = 1024'h6b841e9e35f809da982f955cb9e3a8ac5d899ae890473ab7f6ec36ced1484be54dd73c7d6e97b35ccef5db0f478d4ca5e2ca0442f575696a99338f045e5fd5e315f65ee809a6e4f966436a4a040ad88507cadd0632e12f908c0c6d2d811a5fc2c955d42e114642ef02d1dd9cabe3ad6d1e37e2b66a7a68ba88d13b3a0e6e576a;
    5'b10011 : xpb = 1024'hac61a9355d2a8dc61d340cb7c9aad809fa55082234c8653f5942e968a6cd3474b6d0b0c91bacf5bc2c067c526ca64847e616d8e8b953fbd0dc962c15cc8ede002fbae7847d9962900e96f1128c8d97b92ee6039cf2c5168fecca32200d71297e55f990b04d299980cc56618c247cd200f311d60bfcefaa0de0c9206975bff030;
    5'b10100 : xpb = 1024'h3c91ee76c26edce8d7330c3bc917c01625aa722b03d1ef4f3dbce2acc94f6ffc1c81a79bfe9bb98ce9b8de4eae61331f854985a85a7fbdeb6f5989c8ffeb716bd5303b7241fae2e1a45075387c3492bc61fc309b2622d07e97fb6517df9d50a7b395bb08d843f7850f1afe9ca545d06b7911ea7f3f198e30f2518a94542f228b;
    5'b10101 : xpb = 1024'h7d6f790de9a160d45c378396d8deef73c275df64a85319d6a01395469ed4588b857b1be7abb0fbec46c97f91d37a2ec188965a4e1e5e5051b2bc26da6e1a7988eef4c40eb5ed60784ca3fc0104b751f089175731e606b77df8b92a0a6bf41a634039778b14274e16d89f828c1ddef4ff4debddd4d18ecf844a496fc3bb80bb51;
    5'b10110 : xpb = 1024'hd9fbe4f4ee5aff71636831ad84bd77fedcb496d775ca3e6848d8e8ac1569412eb2c12ba8e9fbfbd047be18e1535199927c9070dbf8a126c457f848da1770cf4946a17fc7a4ee0c9e25d8026f45e4cf3bc2d84301964716ca3ea5d023e20418c9dd5a1e39f41ac1b1b641f9c9ea7f369d3ebf24813b8b3a75bd1d9ee99efedac;
    5'b10111 : xpb = 1024'h4e7d48e6761833e29b3afa75e81306dd8a96b6a71bddce6de6e4412496db7ca2542587063bb5021c618c82d13a4e153b2b15dbb38368a4d288e2219f0fa61511ae2ea098ee415e608ab106ef7ce10c27e348aac6d948586c04a821f4ca770b482a795e65db2502ace4e8a38c174117fda8c5e59da62df4fab3c9bf1e01418672;
    5'b11000 : xpb = 1024'h8f5ad37d9d4ab7ce203f71d0f7da363b276223e0c05ef8f5493af3be6c606531bd1efb51e8ca447bbe9d24145f6710dd2e62b05947473738cc44beb07dd51d2ec7f329356233dbf733048db80563cb5c0a63d15d992c3f6b6565e6e756cdd503b71d1ae81708593eae6d277b8fda3c917d9fd8f338a3364e0bc1a44d68931f38;
    5'b11001 : xpb = 1024'h1f8b18bf028f06f0da3e7154f7471e4752b78de98f6883052db4ed028ee2a0b922cff224cbb9084c7c4f8610a121fbb4cd955d18e872f9535f081c63b131b09a6d687d2326955c48c8be11ddf50ac65f3d79fe5bcc89f95a109719df28f9fc2d14b94540a222b742f131c48c10a33afc039fed667acd1a711d4a0e7847025193;
    5'b11010 : xpb = 1024'h6068a35629c18adc5f42e8b0070e4da4ef82fb2333e9ad8c900b9f9c646789488bc9667078ce4aabd9602753c63af756d0e231beac518bb9a26ab9751f60b8b7872d05bf9a87d9df711198a67d8d8593649524f28c6de0597154ded1b550c5e8a15d01c2de060dd4bab6487b893c5f8fd879e0bc0d425bc47541f3a7ae53ea59;
    5'b11011 : xpb = 1024'ha1462ded50f40ec7e447600b16d57d028c4e685cd86ad813f262523639ec71d7f4c2dabc25e38d0b3670c896eb53f2f8d42f066470301e1fe5cd56868d8fc0d4a0f18e5c0e7a577619651f6f061044c78bb04b894c51c758d212a3c441a78fa42e00be4519e96466843acc6b01d58423ad53d4119fb79d17cd39d8d715a5831f;
    5'b11100 : xpb = 1024'h3176732eb6385dea9e465f8f1642650eb7a3d265a7746223d6dc4b7a5c6ead5f5a73d18f08d250dbf4232a932d0eddd07361b324115be03a7890b439c0ec54404666e249d2dbd7c7af1ea394f5b73fcabec678877faf81477d43d6bc13d3b6cd8b9ce89da503c26ac6ff697b829e828e3353e884e1e1813adec24301f414b57a;
    5'b11101 : xpb = 1024'h7253fdc5dd6ae1d6234ad6ea2609946c546f3f9f4bf58cab3932fe1431f395eec36d45dab5e7933b5133cbd65227d97276ae87c9d53a72a0bbf3514b2f1b5c5d602b6ae646ce555e57722a5d7e39fefee5e19f1e3f936846de019baea02a80891840a51fe0e718fc9083ed6afb37a722082ddbda7456c28e36ba28315b664e40;
    5'b11110 : xpb = 1024'h284430742af30f8dd49d66e25767c787fc4a9a81aff16bb1dacf7585475d176291e3cad98d6570c0ee62dd293e2c44a15e13489766634bb4eb6aefe6277efc905a0bed40b2fd5afed2bae836de0fa0218f7cc1c72f122358932cea67256a7b275dccf786c017700d3488a7b7c00a58c8e2df04db680a6b14842925c39d5809b;
    5'b11111 : xpb = 1024'h4361cd9e69e1b4e4624e4dc9353dabd61c9016e1bf8041428003a9f229faba059217b0f945eb996b6bf6cf15b8fbbfec192e092f3a44c72192194c0fd0a6f7e61f6547707f225346957f354bf663b9364012f2b332d50934e9f09398fead716e02808bfaa7e4cd929ccd0e6af499ca206307e3a348f5e804a03a778ba1271961;
    endcase
end

endmodule

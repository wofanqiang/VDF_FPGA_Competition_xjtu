module xpb_5_445
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h57548b22dd8c9bede5bc71ace86e2fa3f070a2c6c61ed5f6ff6541f52a1b35f8609ca6e21df9de1cea93a639f317353a3f41b57fc03c1e0fe85645180ecc230b704f1a5c3535ff013353e56e9fdd95286b9ef6e2e2588871eb617cfab6f1a8195290ea60aef5c43323264cb1fb34a7885cdc5b44da17ee909c2a8254afaf56c9;
    5'b00010 : xpb = 1024'haea91645bb1937dbcb78e359d0dc5f47e0e1458d8c3dabedfeca83ea54366bf0c1394dc43bf3bc39d5274c73e62e6a747e836aff80783c1fd0ac8a301d984616e09e34b86a6bfe0266a7cadd3fbb2a50d73dedc5c4b110e3d6c2f9f56de35032a521d4c15deb8866464c9963f6694f10b9b8b689b42fdd21385504a95f5ead92;
    5'b00011 : xpb = 1024'h55505c12d6b79f00e62fdd2fa8f0479a5fdbe5237ce4e16d80530c89cb4ef4e11e8d772d8fc71bc8205cb366f5e78ee459aaf8991e0189e408638fe9f191f470dc9e1a65f010ffbe8761ada946bcfb484ed7eb101a836c450c97e4f56aaa55b9c8ab2cf85c18540be2b2ff36f9cdd06fc7bb32ec3dfc6e818e100bf9862b9df0;
    5'b00100 : xpb = 1024'haca4e735b4443aeecbec4edc915e773e504c87ea4303b7647fb84e7ef56a2ad97f2a1e0fadc0f9e50af059a0e8fec41e98ecae18de3da7f3f0b9d502005e177c4ced34c22546febfbab59317e69a9070ba76e1f2fcdbf4b6f7f961f0219bfdd31b3c17590b0e183f05d94be8f50277f824978e3118145d122a3a8e4e35daf4b9;
    5'b00101 : xpb = 1024'h534c2d02cfe2a213e6a348b269725f90cf47278033aaece40140d71e6c82b3c9dc7e4779019459735625c093f8b7e88e74143bb27bc6f5b82870dabbd457c5d648ed1a6faaec007bdb6f75e3ed9c61683210df3d52ae50182dce4cf01e63035a3ec56f90093ae3e4a23fb1bbf866f957329a0a93a1e0ee727ff5959e5ca7e517;
    5'b00110 : xpb = 1024'haaa0b825ad6f3e01cc5fba5f51e08f34bfb7ca46f9c9c2db00a61913969de9c23d1aee5b1f8e379040b966cdebcf1dc8b355f1323c0313c810c71fd3e323e8e1b93c34cbe021ff7d0ec35b528d79f6909dafd6203506d88a192fc9ead554ab73915659f0b830a817c565fe6df39ba0df8f7665d87bf8dd031c2017f30c573be0;
    5'b00111 : xpb = 1024'h5147fdf2c90da526e716b43529f477873eb269dcea70f85a822ea1b30db672b29a6f17c47361971e8beecdc0fb8842388e7d7ecbd98c618c487e258db71d973bb53c1a7965c701392f7d3e1e947bc7881549d36a8ad933eb4f04b4ead21bb0fab4dfb227b65d73bd61cc6440f700223e9d78e23b05c56e6371db1f4333242c3e;
    5'b01000 : xpb = 1024'ha89c8915a69a4114ccd325e21262a72b2f230ca3b08fce518193e3a837d1a8aafb0bbea6915b753b768273faee9f7772cdbf344b99c87f9c30d46aa5c5e9ba47258b34d59afd003a62d1238d34595cb080e8ca4d6d31bc5d3a6631e5890d591407709c88655337f084f2b0f2f234c9c6fa553d7fdfdd5cf40e05a197e2d38307;
    5'b01001 : xpb = 1024'h4f43cee2c238a839e78a1fb7ea768f7dae1dac39a13703d1031c6c47aeea319b585fe80fe52ed4c9c1b7daedfe589be2a8e6c1e53751cd60688b705f99e368a1218b1a8320a201f6838b06593b5b2da7f882c797c30417be703b1ce585d45e9b2af9f4bf63800396215916c5f5994b260857b9e269a9ee5463c0a8e809a07365;
    5'b01010 : xpb = 1024'ha6985a059fc54427cd469164d2e4bf219e8e4f006755d9c80281ae3cd9056793b8fc8ef20328b2e6ac4b8127f16fd11ce8287764f78deb7050e1b577a8af8bac91da34df55d800f7b6deebc7db38c2d06421be7aa55ca0305b9c99e03cc606b47d8adf201275c7c9447f6377f0cdf2ae6534152743c1dce4ffeb2b3cb94fca2e;
    5'b01011 : xpb = 1024'h4d3f9fd2bb63ab4ce7fd8b3aaaf8a7741d88ee9657fd0f47840a36dc501df0841650b85b56fc1274f780e81b0128f58cc35004fe951739348898bb317ca93a068dda1a8cdb7d02b3d798ce93e23a93c7dbbbbbc4fb2efb91917184e0398d0c3ba114375710a2936ee0e5c94af432740d73369189cd8e6e4555a6328ce01cba8c;
    5'b01100 : xpb = 1024'ha4942af598f0473acdb9fce79366d7180df9915d1e1be53e836f78d17a39267c76ed5f3d74f5f091e2148e54f4402ac70291ba7e5553574470ef00498b755d11fe2934e910b301b50aecb402821828f0475ab2a7dd8784037cd301daf07eb454f3a521b7bf9857a2040c15fcef671b95d012eccea7a65cd5f1d0b4e18fcc1155;
    5'b01101 : xpb = 1024'h4b3b70c2b48eae5fe870f6bd6b7abf6a8cf430f30ec31abe04f80170f151af6cd44188a6c8c950202d49f54803f94f36ddb94817f2dca508a8a606035f6f0b6bfa291a96965803712ba696ce8919f9e7bef4aff23359df64b2a7ecdaed45b9dc172e79eebdc52347a0727bcff2cb9cf4de1569313172ee36478bbc31b69901b3;
    5'b01110 : xpb = 1024'ha28ffbe5921b4a4dce2d686a53e8ef0e7d64d3b9d4e1f0b5045d43661b6ce56534de2f88e6c32e3d17dd9b81f71084711cfafd97b318c31890fc4b1b6e3b2e776a7834f2cb8e02725efa7c3d28f78f102a93a6d515b267d69e0969d5a43761f569bf644f6cbae77ac398c881ee00447d3af1c4760b8adcc6e3b63e866648587c;
    5'b01111 : xpb = 1024'h493741b2adb9b172e8e462402bfcd760fc5f734fc589263485e5cc0592856e55923258f23a968dcb6313027506c9a8e0f8228b3150a210dcc8b350d54234dcd166781aa05133042e7fb45f092ff96007a22da41f6b84c337d3de54d5a0fe677c8d48bc866ae7b3205fff2e54f164c5dc48f440d895576e27397145d68d1548da;
    5'b10000 : xpb = 1024'ha08bccd58b464d60cea0d3ed146b0704ecd016168ba7fc2b854b0dfabca0a44df2ceffd458906be84da6a8aef9e0de1b376440b110de2eecb10995ed5100ffdcd6c734fc8669032fb3084477cfd6f5300dcc9b024ddd4ba9bf3fd1d057f00f95dfd9a6e719dd775383257b06ec996d64a5d09c1d6f6f5cb7d59bc82b3cc49fa3;
    5'b10001 : xpb = 1024'h473312a2a6e4b485e957cdc2ec7eef576bcab5ac7c4f31ab06d3969a33b92d3e5023293dac63cb7698dc0fa2099a028b128bce4aae677cb0e8c09ba724faae36d2c71aaa0c0e04ebd3c22743d6d8c6278566984ca3afa70af514bcd054b7151d0362ff1e180a42f91f8be0d9effdeec3b3d3187ff93bee182b56cf7b63919001;
    5'b10010 : xpb = 1024'h9e879dc584715073cf143f6fd4ed1efb5c3b5873426e07a20638d88f5dd46336b0bfd01fca5da993836fb5dbfcb137c551cd83ca6ea39ac0d116e0bf33c6d14243163506414403ed07160cb276b65b4ff1058f2f86082f7ce07639cb0ba8bd3655f3e97ec700072c42b22d8beb32964c10af73c4d353dca8c78151d01340e6ca;
    5'b10011 : xpb = 1024'h452ee392a00fb798e9cb3945ad01074ddb35f80933153d2187c1612ed4ecec270e13f9891e310921cea51ccf0c6a5c352cf511640c2ce88508cde67907c07f9c3f161ab3c6e905a927cfef7e7db82c47689f8c79dbda8ade164b24cb086fc2bd797d41b5c52cd2d1df18935eee9717ab1eb1f0275d206e091d3c59203a0dd728;
    5'b10100 : xpb = 1024'h9c836eb57d9c5386cf87aaf2956f36f1cba69acff93413188726a323ff08221f6eb0a06b3c2ae73eb938c308ff81916f6c36c6e3cc690694f1242b91168ca2a7af65350ffc1f04aa5b23d4ed1d95c16fd43e835cbe33135001aca1c5bf616ad6cc0e2c1674229705023ee010e9cbbf337b8e4b6c37385c99b966db74e9bd2df1;
    5'b10101 : xpb = 1024'h432ab482993abaabea3ea4c86d831f444aa13a65e9db489808af2bc37620ab0fcc04c9d48ffe46cd046e29fc0f3ab5df475e547d69f2545928db314aea865101ab651abd81c406667bddb7b9249792674bd880a714056eb137818cc5bc28705def97844d724f62aa9ea545e3ed3040928990c7cec104edfa0f21e2c5108a1e4f;
    5'b10110 : xpb = 1024'h9a7f3fa576c75699cffb167555f14ee83b11dd2caffa1e8f08146db8a03be1082ca170b6adf824e9ef01d0360251eb1986a009fd2a2e726911317662f952740d1bb43519b6fa0567af319d27c475278fb7777789f65df72322e309c0731a187742286eae214526ddc1cb9295e864e81ae66d23139b1cdc8aab4c6519c0397518;
    5'b10111 : xpb = 1024'h412685729265bdbeeab2104b2e05373aba0c7cc2a0a1540e899cf658175469f889f59a2001cb84783a373729120b0f8961c79796c7b7c02d48e87c1ccd4c226717b41ac73c9f0723cfeb7ff3cb76f8872f1174d44c30528458b7f4c06fe11dfe65b1c6e51f71f2835e31f868ebc96979f46f9f7624e96deb01076c69e7066576;
    5'b11000 : xpb = 1024'h987b10956ff259acd06e81f8167366deaa7d1f8966c02a058902384d416f9ff0ea9241021fc5629524cadd63052244c3a1094d1687f3de3d313ec134dc1845728803352371d50625033f65626b548daf9ab06bb72e88daf6441971bb26d2c617b842b145ce67b6b68158451ae6fe1102514bfabaff015c7b9d31eebe96b5bc3f;
    5'b11001 : xpb = 1024'h3f2256628b90c0d1eb257bcdee874f312977bf1f57675f850a8ac0ecb88828e147e66a6b7398c2237000445614db69337c30dab0257d2c0168f5c6eeb011f3cc84031ad0f77a07e123f9482e72565ea7124a6901845b365779ee5cbb2399cb9edbcc097ccc94825c1dbeaaedea6292615f4e771d88cdeddbf2ecf60ebd82ac9d;
    5'b11010 : xpb = 1024'h9676e185691d5cbfd0e1ed7ad6f57ed519e861e61d86357c09f002e1e2a35ed9a883114d9192a0405a93ea9007f29e6dbb72902fe5b94a11514c0c06bede16d7f452352d2cb006e2574d2d9d1233f3cf7de95fe466b3bec9654fd9b5da8b73b82e5cf3dd7b8a468f40e4f79fe59739e9bc2ad26262e5dc6c8f1778636d320366;
    5'b11011 : xpb = 1024'h3d1e275284bbc3e4eb98e750af09672798e3017c0e2d6afb8b788b8159bbe7ca05d73ab6e565ffcea5c9518317abc2dd969a1dc9834297d5890311c092d7c531f0521adab255089e780710691935c4c6f5835d2ebc861a2a9b24c4b5d752793f51e64c1479b71234dd4b5d72e8fbbb48ca2d4ec4ecb26dcce4d27fb393fef3c4;
    5'b11100 : xpb = 1024'h9472b27562485fd2d15558fd977796cb8953a442d44c40f28addcd7683d71dc26673e199035fddeb905cf7bd0ac2f817d5dbd349437eb5e5715956d8a1a3e83d60a13536e78b079fab5af5d7b91359ef612254119edea29c868641b08e442158a477367528acd6680071aa24e43062d12709aa09c6ca5c5d80fd020843ae4a8d;
    5'b11101 : xpb = 1024'h3b19f8427de6c6f7ec0c52d36f8b7f1e084e43d8c4f376720c665615faefa6b2c3c80b0257333d79db925eb01a7c1c87b10360e2e10803a9a9105c92759d96975ca11ae46d30095bcc14d8a3c0152ae6d8bc515bf4b0fdfdbc5b2cb08b0b26dfc8008eac26d9a20d9cd80ff7e794e430350c266c5096edbdd6b809586a7b3aeb;
    5'b11110 : xpb = 1024'h926e83655b7362e5d1c8c48057f9aec1f8bee69f8b124c690bcb980b250adcab2464b1e4752d1b96c62604ea0d9351c1f0451662a14421b99166a1aa8469b9a2ccf03540a266085cff68be125ff2c00f445b483ed709866fa7bca9ab41fccef91a91790cd5cf6640bffe5ca9e2c98bb891e881b12aaedc4e72e28bad1a2a91b4;
    5'b11111 : xpb = 1024'h3915c9327711ca0aec7fbe56300d971477b986357bb981e88d5420aa9c23659b81b8db4dc9007b25115b6bdd1d4c7631cb6ca3fc3ecd6f7dc91da764586367fcc8f01aee280b0a192022a0de66f49106bbf545892cdbe1d0dd9194ab3ec3d4803e1ad143d3fc31e65c64c27ce62e0d179feafe13b47b6daec89d92fd40f78212;
    endcase
end

endmodule

module xpb_5_600
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h58bde9c9b0f8ee4243c72abefd15a315697b3e3cb9854f2ac81ccf3504006e729abeefea601f7c0a5c40932aac0b43e15a85ea0efe0c12b534c87ab6a506b4825ad050fd1f9753041ef2cd2be5c2e5de402324fc7a82fb025c5364f86d7df616fee625e546dbb49088ca6476576a211ff89659abac7b1782155578194a79ed31;
    5'b00010 : xpb = 1024'hce8e3da003a7bbbc88dda6e9d0fed9618079489d92fdde125ce51454fe2fdd3235625bf61879861922e70e74b876f850f1ac37d965551eb8f1b60f0f3af45341516d4b8f9da8c32b4b97b532aa078b8c415060687fc8f4031a37f620d1499bcec4b9a0dcee70938ad4e20db7041c16a252d47508aad1d3e43b752e0c1173f7;
    5'b00011 : xpb = 1024'h598c780750fc95fe00500865e6e6a1eecafbb78557184d08da79b44958fe9e4fccf452465637f59075637a3920c3bad9ab779646d77167d3edba30c5b441a8d59c21be48af34fbc74a3e64e1186ced69cc64755ce302c3f65f6d9cee8e4f3fb2cdaadf8623ca2524139f46840e6e3d369ae92e20b525e955f990ed47568b6128;
    5'b00100 : xpb = 1024'h19d1c7b40074f777911bb4dd3a1fdb2c300f2913b25fbbc24b9ca28a9fc5fba646ac4b7ec30f30c3245ce1ce970edf0a1e3586fb2caaa3d71e36c1e1e75e8a682a2da971f3b518656972f6a65540f171882a0c0d0ff91e806346fec41a293379d897341b9dce12715a9c41b6e08382d44a5a8ea1155a3a7c876ea5c1822e7ee;
    5'b00101 : xpb = 1024'h5a5b0644f1003db9bcd8e60cd0b7a0c82c7c30cdf4ab4ae6ecd6995dadfcce2cff29b4a24c506f168e866147957c31d1fc69427eb0d6bcf2a6abe6d4c37c9d28dd732b943ed2a48a7589fc964b16f4f558a5c5bd4b828cea6287d4e4af20894e9c6f992700b895b79e742891c572594d3d3c0295bdd0bb29ddcc6275629cd51f;
    5'b00110 : xpb = 1024'h26baab8e00af733359a98f4bd72fc8c24816bd9d8b8f99a3716af3cfefa8f9796a02713e2496c924b68b52b5e2964e8f2d504a78c2fff5c2ad5222d2db0dcf9c3f447e2aed8fa4981e2c71f97fe16a2a4c3f121397f5adc094ea7e26273dcd36c4e2ce296cb51baa07ea629250c5443e6f87d5f1a00757bacb25f8a24345be5;
    5'b00111 : xpb = 1024'h5b2994829103e5757961c3b3ba889fa18dfcaa16923e48c4ff337e7202fafe0a315f16fe4268e89ca7a948560a34a8ca4d5aeeb68a3c12115f9d9ce3d2b7917c1ec498dfce704d4da0d5944b7dc0fc80e4e7161db40255de65a20cdacff1d2ea6b3452c7dda7064b29490a9f7c767563df8ed70ac67b8cfdc207d7a36eae4916;
    5'b01000 : xpb = 1024'h33a38f6800e9eeef223769ba743fb658601e522764bf7784973945153f8bf74c8d5896fd861e618648b9c39d2e1dbe143c6b0df6595547ae3c6d83c3cebd14d0545b52e3e76a30cad2e5ed4caa81e2e31054181a1ff23d00c68dfd88345266f3b12e68373b9c24e2b538836dc10705a894b51d422ab474f90edd4b83045cfdc;
    5'b01001 : xpb = 1024'h5bf822c031078d3135eaa15aa4599e7aef7d235f2fd146a31190638657f92de76394795a38816222c0cc2f647eed1fc29e4c9aee63a16730188f52f2e1f285cf6016062b5e0df610cc212c00b06b040c7128667e1c821ed268bc44d0f0c31c8639f90c68ba9576deb41decad337a917a81e1ab7fcf265ed1a6434cd17abfbd0d;
    5'b01010 : xpb = 1024'h408c734201246aaaeac54429114fa3ee7825e6b13def5565bd07965a8f6ef51fb0aebcbce7a5f9e7dae8348479a52d994b85d173efaa9999cb88e4b4c26c5a046972279ce144bcfd879f689fd5225b9bd4691e20a7eecc40f8317cea416700b09d7a02450a832e1b6286a4493148c712b9e26492b561923752949e63c5743d3;
    5'b01011 : xpb = 1024'h5cc6b0fdd10b34ecf2737f018e2a9d5450fd9ca7cd64448123ed489aacf75dc495c9dbb62e99dba8d9ef1672f3a596baef3e47263d06bc4ed1810901f12d7a22a1677376edab9ed3f76cc3b5e3150b97fd69b6de8501e7c66bd67cc71194662208bdc6099783e7723ef2cebaea7ead9124347ff4d7d130a58a7ec1ff86d13104;
    5'b01100 : xpb = 1024'h4d75571c015ee666b3531e97ae5f9184902d7b3b171f3346e2d5e79fdf51f2f2d404e27c492d92496d16a56bc52c9d1e5aa094f185ffeb855aa445a5b61b9f387e88fc55db1f49303c58e3f2ffc2d454987e24272feb5b8129d4fc4c4e7b9a6d89c59c52d96a37540fd4c524a18a887cdf0fabe3400eaf75964bf144868b7ca;
    5'b01101 : xpb = 1024'h5d953f3b710edca8aefc5ca877fb9c2db27e15f06af7425f364a2daf01f58da1c7ff3e1224b2552ef311fd81685e0db3402ff35e166c116d8a72bf1100686e75e2b8e0c27d49479722b85b6b15bf132389ab073eed81b0ba6ef0b4bd3265afbdd7827faa74725805c9c7b0c8a182c9a7c6875469e07c02796eba372d92e2a4fb;
    5'b01110 : xpb = 1024'h5a5e3af6019962227be0f9064b6f7f1aa8350fc4f04f112808a438e52f34f0c5f75b083baab52aaaff45165310b40ca369bb586f1c553d70e9bfa696a9cae46c939fd10ed4f9d562f1125f462a634d0d5c932a2db7e7eac15b787bae5b90342a76113660a851408cbd22e60011cc49e7043cf333cabbccb3da03442547a2bc1;
    5'b01111 : xpb = 1024'h5e63cd79111284646b853a4f61cc9b0713fe8f39088a403d48a712c356f3bd7efa34a06e1acaceb50c34e48fdd1684ab91219f95efd1668c436475200fa362c9240a4e0e0ce6f05a4e03f32048691aaf15ec579f560179ae720aecb35336f959a647394b5160c899549c92d65886e5be68da28dee926d44d52f5ac5b9ef418f2;
    5'b10000 : xpb = 1024'h67471ed001d3ddde446ed374e87f6cb0c03ca44ec97eef092e728a2a7f17ee991ab12dfb0c3cc30c9173873a5c3b7c2878d61becb2aa8f5c78db07879d7a29a0a8b6a5c7ced46195a5cbda995503c5c620a830343fe47a018d1bfb1068a4cde7625cd06e773849c56a7106db820e0b51296a3a845568e9f21dba970608b9fb8;
    5'b10001 : xpb = 1024'h5f325bb6b1162c20280e17f64b9d99e0757f0881a61d3e1b5b03f7d7abf1ed5c2c6a02ca10e3483b2557cb9e51cefba3e2134bcdc936bbaafc562b2f1ede571c655bbb599c84991d794f8ad57b13223aa22da7ffbe8142a2752524a9740842f5750bf2ec2e4f392cdf7174e40f8b01d50b2cfd53f1d1a62137312189ab058ce9;
    5'b10010 : xpb = 1024'h743002aa020e599a0cfcade3858f5a46d84438d8a2aeccea5440db6fcefaec6c3e0753ba6dc45b6e23a1f821a7c2ebad87f0df6a48ffe14807f6687891296ed4bdcd7a80c8aeedc85a8555ec7fa43e7ee4bd363ac7e10941bebf7a7275b967a44ea86a7c461f52fe17bf27b6f24fccbb4e9781d4e01607306171e9e6c9d13af;
    5'b10011 : xpb = 1024'h6000e9f45119d3dbe496f59d356e98b9d6ff81ca43b03bf96d60dcec00f01d395e9f652606fbc1c13e7ab2acc687729c3304f805a29c10c9b547e13e2e194b6fa6ad28a52c2241e0a49b228aadbd29c62e6ef86027010b96783f5c9f94d98c9143d0ac8d0b3da9c06a4656f1c68f1debad7fd1c8fa7c77f51b6c96b7b71700e0;
    5'b10100 : xpb = 1024'h8118e6840248d555d58a8852229f47dcf04bcd627bdeaacb7a0f2cb51eddea3f615d7979cf4bf3cfb5d06908f34a5b32970ba2e7df5533339711c96984d8b408d2e44f39c28979fb0f3ed13faa44b737a8d23c414fdd9881f062f9d482ce01613af4048a15065c36c50d489262918e2573c4c9256ac3246ea5293cc78ae87a6;
    5'b10101 : xpb = 1024'h60cf7831f11d7b97a11fd3441f3f9793387ffb12e14339d77fbdc20055ee4d1690d4c781fd143b47579d99bb3b3fe99483f6a43d7c0165e86e39974d3d543fc2e7fe95f0bbbfeaa3cfe6ba3fe0673151bab048c08f80d48a7b599495b5aad62d1295662de82c1a53f51b38ff7d933a024fd2a63e032749c8ffa80be5c32874d7;
    5'b10110 : xpb = 1024'h8e01ca5e028351119e1862c0bfaf3573085361ec550e88ac9fdd7dfa6ec0e81284b39f3930d38c3147fed9f03ed1cab7a626666575aa851f262d2a5a7887f93ce7fb23f2bc64062dc3f84c92d4e52ff06ce74247d7da27c2220679368fe29b1e273f9e97e3ed656f725b696dd2d34f8f98f21075f57041ace8e08fa84bffb9d;
    5'b10111 : xpb = 1024'h619e066f912123535da8b0eb0910966c9a00745b7ed637b5921aa714aaec7cf3c30a29ddf32cb4cd70c080c9aff8608cd4e850755566bb07272b4d5c4c8f34162950033c4b5d9366fb3251f5131138dd46f19920f8009d7e7e73cc8bd67c1fc8e15a1fcec51a8ae77ff01b0d34975618f2257ab30bd21b9ce3e38113cf39e8ce;
    5'b11000 : xpb = 1024'h9aeaae3802bdcccd66a63d2f5cbf2309205af6762e3e668dc5abcf3fbea3e5e5a809c4f8925b2492da2d4ad78a593a3cb54129e30bffd70ab5488b4b6c373e70fd11f8abb63e926078b1c7e5ff85a8a930fc484e5fd6b70253a9f8989cf734db138b38a5b2d46ea81fa98a49431510f9be1f57c6801d5eeb2c97e2890d16f94;
    5'b11001 : xpb = 1024'h626c94ad3124cb0f1a318e91f2e19545fb80eda41c693593a4778c28ffeaacd0f53f8c39e9452e5389e367d824b0d78525d9fcad2ecc1025e01d036b5bca28696aa17087dafb3c2a267de9aa45bb4068d332e98160806672818e0481f74d6964b01ed96fa208fb7b0ac4fd1aeb9b722f94784f28147ced70c81ef641db4b5cc5;
    5'b11010 : xpb = 1024'ha7d3921202f848892f34179df9cf109f38628b00076e446eeb7a20850e86e3b8cb5feab7f3e2bcf46c5bbbbed5e0a9c1c45bed60a25528f64463ec3c5fe683a51228cd64b0191e932d6b43392a262161f5114e54e7d34642854d77faaa0bce97ffd6d2b381bb77e0ccf7ab24b356d263e34c9f170aca7c29704f3569ce2e38b;
    5'b11011 : xpb = 1024'h633b22ead12872cad6ba6c38dcb2941f5d0166ecb9fc3371b6d4713d54e8dcae2774ee95df5da7d9a3064ee699694e7d76cba8e508316544990eb97a6b051cbcabf2ddd36a98e4ed51c9815f786547f45f7439e1c9002f6684a83c78181eb3007ee393107ef76c0e9599df28a29f8e4636cb239d1d27bf44ac5a6b6fe75cd0bc;
    5'b11100 : xpb = 1024'hb4bc75ec0332c444f7c1f20c96defe35506a1f89e09e2250114871ca5e69e18beeb61077556a5555fe8a2ca621681946d376b0de38aa7ae1d37f4d2d5395c8d9273fa21da9f3aac5e224be8c54c69a1ab926545b6fcfd582b6f0f75cb7206854ec226cc150a281197a45cc00239893ce0879e66795779967b406884a8f45782;
    5'b11101 : xpb = 1024'h6409b128712c1a86934349dfc68392f8be81e035578f314fc9315651a9e70c8b59aa50f1d576215fbc2935f50e21c575c7bd551ce196ba6352006f897a40110fed444b1efa368db07d151914ab0f4f7febb58a42317ff85a87c2746e38effc9c4da84cb15be5dca2206ec13659a3aa5cd91df81225d291189095e09df36e44b3;
    5'b11110 : xpb = 1024'hc1a559c6036d4000c04fcc7b33eeebcb6871b413b9ce00313716c30fae4cdf5f120c3636b6f1edb790b89d8d6cef88cbe291745bceffcccd629aae1e47450e0d3c5676d6a3ce36f896de39df7f6712d37d3b5a61f7cc64c2e89476bec4350211d86e06cf1f898a522793ecdb93da55382da72db82024b6a5f7bddb2b505cb79;
    5'b11111 : xpb = 1024'h64d83f66112fc2424fcc2786b05491d22002597df5222f2ddb8e3b65fee53c688bdfb34dcb8e9ae5d54c1d0382da3c6e18af0154bafc0f820af22598897b05632e95b86a89d43673a860b0c9ddb9570b77f6daa299ffc14e8adcac6459c146381c6d065238d44d35ab43a34410a7c6737b70cc872e7d62ec74d155cbff7fb8aa;
    endcase
end

endmodule

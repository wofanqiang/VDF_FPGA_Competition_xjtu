module compressor_array_8_6_1288
(
    input  [7:0] col_in_0,
    input  [7:0] col_in_1,
    input  [7:0] col_in_2,
    input  [7:0] col_in_3,
    input  [7:0] col_in_4,
    input  [7:0] col_in_5,
    input  [7:0] col_in_6,
    input  [7:0] col_in_7,
    input  [7:0] col_in_8,
    input  [7:0] col_in_9,
    input  [7:0] col_in_10,
    input  [7:0] col_in_11,
    input  [7:0] col_in_12,
    input  [7:0] col_in_13,
    input  [7:0] col_in_14,
    input  [7:0] col_in_15,
    input  [7:0] col_in_16,
    input  [7:0] col_in_17,
    input  [7:0] col_in_18,
    input  [7:0] col_in_19,
    input  [7:0] col_in_20,
    input  [7:0] col_in_21,
    input  [7:0] col_in_22,
    input  [7:0] col_in_23,
    input  [7:0] col_in_24,
    input  [7:0] col_in_25,
    input  [7:0] col_in_26,
    input  [7:0] col_in_27,
    input  [7:0] col_in_28,
    input  [7:0] col_in_29,
    input  [7:0] col_in_30,
    input  [7:0] col_in_31,
    input  [7:0] col_in_32,
    input  [7:0] col_in_33,
    input  [7:0] col_in_34,
    input  [7:0] col_in_35,
    input  [7:0] col_in_36,
    input  [7:0] col_in_37,
    input  [7:0] col_in_38,
    input  [7:0] col_in_39,
    input  [7:0] col_in_40,
    input  [7:0] col_in_41,
    input  [7:0] col_in_42,
    input  [7:0] col_in_43,
    input  [7:0] col_in_44,
    input  [7:0] col_in_45,
    input  [7:0] col_in_46,
    input  [7:0] col_in_47,
    input  [7:0] col_in_48,
    input  [7:0] col_in_49,
    input  [7:0] col_in_50,
    input  [7:0] col_in_51,
    input  [7:0] col_in_52,
    input  [7:0] col_in_53,
    input  [7:0] col_in_54,
    input  [7:0] col_in_55,
    input  [7:0] col_in_56,
    input  [7:0] col_in_57,
    input  [7:0] col_in_58,
    input  [7:0] col_in_59,
    input  [7:0] col_in_60,
    input  [7:0] col_in_61,
    input  [7:0] col_in_62,
    input  [7:0] col_in_63,
    input  [7:0] col_in_64,
    input  [7:0] col_in_65,
    input  [7:0] col_in_66,
    input  [7:0] col_in_67,
    input  [7:0] col_in_68,
    input  [7:0] col_in_69,
    input  [7:0] col_in_70,
    input  [7:0] col_in_71,
    input  [7:0] col_in_72,
    input  [7:0] col_in_73,
    input  [7:0] col_in_74,
    input  [7:0] col_in_75,
    input  [7:0] col_in_76,
    input  [7:0] col_in_77,
    input  [7:0] col_in_78,
    input  [7:0] col_in_79,
    input  [7:0] col_in_80,
    input  [7:0] col_in_81,
    input  [7:0] col_in_82,
    input  [7:0] col_in_83,
    input  [7:0] col_in_84,
    input  [7:0] col_in_85,
    input  [7:0] col_in_86,
    input  [7:0] col_in_87,
    input  [7:0] col_in_88,
    input  [7:0] col_in_89,
    input  [7:0] col_in_90,
    input  [7:0] col_in_91,
    input  [7:0] col_in_92,
    input  [7:0] col_in_93,
    input  [7:0] col_in_94,
    input  [7:0] col_in_95,
    input  [7:0] col_in_96,
    input  [7:0] col_in_97,
    input  [7:0] col_in_98,
    input  [7:0] col_in_99,
    input  [7:0] col_in_100,
    input  [7:0] col_in_101,
    input  [7:0] col_in_102,
    input  [7:0] col_in_103,
    input  [7:0] col_in_104,
    input  [7:0] col_in_105,
    input  [7:0] col_in_106,
    input  [7:0] col_in_107,
    input  [7:0] col_in_108,
    input  [7:0] col_in_109,
    input  [7:0] col_in_110,
    input  [7:0] col_in_111,
    input  [7:0] col_in_112,
    input  [7:0] col_in_113,
    input  [7:0] col_in_114,
    input  [7:0] col_in_115,
    input  [7:0] col_in_116,
    input  [7:0] col_in_117,
    input  [7:0] col_in_118,
    input  [7:0] col_in_119,
    input  [7:0] col_in_120,
    input  [7:0] col_in_121,
    input  [7:0] col_in_122,
    input  [7:0] col_in_123,
    input  [7:0] col_in_124,
    input  [7:0] col_in_125,
    input  [7:0] col_in_126,
    input  [7:0] col_in_127,
    input  [7:0] col_in_128,
    input  [7:0] col_in_129,
    input  [7:0] col_in_130,
    input  [7:0] col_in_131,
    input  [7:0] col_in_132,
    input  [7:0] col_in_133,
    input  [7:0] col_in_134,
    input  [7:0] col_in_135,
    input  [7:0] col_in_136,
    input  [7:0] col_in_137,
    input  [7:0] col_in_138,
    input  [7:0] col_in_139,
    input  [7:0] col_in_140,
    input  [7:0] col_in_141,
    input  [7:0] col_in_142,
    input  [7:0] col_in_143,
    input  [7:0] col_in_144,
    input  [7:0] col_in_145,
    input  [7:0] col_in_146,
    input  [7:0] col_in_147,
    input  [7:0] col_in_148,
    input  [7:0] col_in_149,
    input  [7:0] col_in_150,
    input  [7:0] col_in_151,
    input  [7:0] col_in_152,
    input  [7:0] col_in_153,
    input  [7:0] col_in_154,
    input  [7:0] col_in_155,
    input  [7:0] col_in_156,
    input  [7:0] col_in_157,
    input  [7:0] col_in_158,
    input  [7:0] col_in_159,
    input  [7:0] col_in_160,
    input  [7:0] col_in_161,
    input  [7:0] col_in_162,
    input  [7:0] col_in_163,
    input  [7:0] col_in_164,
    input  [7:0] col_in_165,
    input  [7:0] col_in_166,
    input  [7:0] col_in_167,
    input  [7:0] col_in_168,
    input  [7:0] col_in_169,
    input  [7:0] col_in_170,
    input  [7:0] col_in_171,
    input  [7:0] col_in_172,
    input  [7:0] col_in_173,
    input  [7:0] col_in_174,
    input  [7:0] col_in_175,
    input  [7:0] col_in_176,
    input  [7:0] col_in_177,
    input  [7:0] col_in_178,
    input  [7:0] col_in_179,
    input  [7:0] col_in_180,
    input  [7:0] col_in_181,
    input  [7:0] col_in_182,
    input  [7:0] col_in_183,
    input  [7:0] col_in_184,
    input  [7:0] col_in_185,
    input  [7:0] col_in_186,
    input  [7:0] col_in_187,
    input  [7:0] col_in_188,
    input  [7:0] col_in_189,
    input  [7:0] col_in_190,
    input  [7:0] col_in_191,
    input  [7:0] col_in_192,
    input  [7:0] col_in_193,
    input  [7:0] col_in_194,
    input  [7:0] col_in_195,
    input  [7:0] col_in_196,
    input  [7:0] col_in_197,
    input  [7:0] col_in_198,
    input  [7:0] col_in_199,
    input  [7:0] col_in_200,
    input  [7:0] col_in_201,
    input  [7:0] col_in_202,
    input  [7:0] col_in_203,
    input  [7:0] col_in_204,
    input  [7:0] col_in_205,
    input  [7:0] col_in_206,
    input  [7:0] col_in_207,
    input  [7:0] col_in_208,
    input  [7:0] col_in_209,
    input  [7:0] col_in_210,
    input  [7:0] col_in_211,
    input  [7:0] col_in_212,
    input  [7:0] col_in_213,
    input  [7:0] col_in_214,
    input  [7:0] col_in_215,
    input  [7:0] col_in_216,
    input  [7:0] col_in_217,
    input  [7:0] col_in_218,
    input  [7:0] col_in_219,
    input  [7:0] col_in_220,
    input  [7:0] col_in_221,
    input  [7:0] col_in_222,
    input  [7:0] col_in_223,
    input  [7:0] col_in_224,
    input  [7:0] col_in_225,
    input  [7:0] col_in_226,
    input  [7:0] col_in_227,
    input  [7:0] col_in_228,
    input  [7:0] col_in_229,
    input  [7:0] col_in_230,
    input  [7:0] col_in_231,
    input  [7:0] col_in_232,
    input  [7:0] col_in_233,
    input  [7:0] col_in_234,
    input  [7:0] col_in_235,
    input  [7:0] col_in_236,
    input  [7:0] col_in_237,
    input  [7:0] col_in_238,
    input  [7:0] col_in_239,
    input  [7:0] col_in_240,
    input  [7:0] col_in_241,
    input  [7:0] col_in_242,
    input  [7:0] col_in_243,
    input  [7:0] col_in_244,
    input  [7:0] col_in_245,
    input  [7:0] col_in_246,
    input  [7:0] col_in_247,
    input  [7:0] col_in_248,
    input  [7:0] col_in_249,
    input  [7:0] col_in_250,
    input  [7:0] col_in_251,
    input  [7:0] col_in_252,
    input  [7:0] col_in_253,
    input  [7:0] col_in_254,
    input  [7:0] col_in_255,
    input  [7:0] col_in_256,
    input  [7:0] col_in_257,
    input  [7:0] col_in_258,
    input  [7:0] col_in_259,
    input  [7:0] col_in_260,
    input  [7:0] col_in_261,
    input  [7:0] col_in_262,
    input  [7:0] col_in_263,
    input  [7:0] col_in_264,
    input  [7:0] col_in_265,
    input  [7:0] col_in_266,
    input  [7:0] col_in_267,
    input  [7:0] col_in_268,
    input  [7:0] col_in_269,
    input  [7:0] col_in_270,
    input  [7:0] col_in_271,
    input  [7:0] col_in_272,
    input  [7:0] col_in_273,
    input  [7:0] col_in_274,
    input  [7:0] col_in_275,
    input  [7:0] col_in_276,
    input  [7:0] col_in_277,
    input  [7:0] col_in_278,
    input  [7:0] col_in_279,
    input  [7:0] col_in_280,
    input  [7:0] col_in_281,
    input  [7:0] col_in_282,
    input  [7:0] col_in_283,
    input  [7:0] col_in_284,
    input  [7:0] col_in_285,
    input  [7:0] col_in_286,
    input  [7:0] col_in_287,
    input  [7:0] col_in_288,
    input  [7:0] col_in_289,
    input  [7:0] col_in_290,
    input  [7:0] col_in_291,
    input  [7:0] col_in_292,
    input  [7:0] col_in_293,
    input  [7:0] col_in_294,
    input  [7:0] col_in_295,
    input  [7:0] col_in_296,
    input  [7:0] col_in_297,
    input  [7:0] col_in_298,
    input  [7:0] col_in_299,
    input  [7:0] col_in_300,
    input  [7:0] col_in_301,
    input  [7:0] col_in_302,
    input  [7:0] col_in_303,
    input  [7:0] col_in_304,
    input  [7:0] col_in_305,
    input  [7:0] col_in_306,
    input  [7:0] col_in_307,
    input  [7:0] col_in_308,
    input  [7:0] col_in_309,
    input  [7:0] col_in_310,
    input  [7:0] col_in_311,
    input  [7:0] col_in_312,
    input  [7:0] col_in_313,
    input  [7:0] col_in_314,
    input  [7:0] col_in_315,
    input  [7:0] col_in_316,
    input  [7:0] col_in_317,
    input  [7:0] col_in_318,
    input  [7:0] col_in_319,
    input  [7:0] col_in_320,
    input  [7:0] col_in_321,
    input  [7:0] col_in_322,
    input  [7:0] col_in_323,
    input  [7:0] col_in_324,
    input  [7:0] col_in_325,
    input  [7:0] col_in_326,
    input  [7:0] col_in_327,
    input  [7:0] col_in_328,
    input  [7:0] col_in_329,
    input  [7:0] col_in_330,
    input  [7:0] col_in_331,
    input  [7:0] col_in_332,
    input  [7:0] col_in_333,
    input  [7:0] col_in_334,
    input  [7:0] col_in_335,
    input  [7:0] col_in_336,
    input  [7:0] col_in_337,
    input  [7:0] col_in_338,
    input  [7:0] col_in_339,
    input  [7:0] col_in_340,
    input  [7:0] col_in_341,
    input  [7:0] col_in_342,
    input  [7:0] col_in_343,
    input  [7:0] col_in_344,
    input  [7:0] col_in_345,
    input  [7:0] col_in_346,
    input  [7:0] col_in_347,
    input  [7:0] col_in_348,
    input  [7:0] col_in_349,
    input  [7:0] col_in_350,
    input  [7:0] col_in_351,
    input  [7:0] col_in_352,
    input  [7:0] col_in_353,
    input  [7:0] col_in_354,
    input  [7:0] col_in_355,
    input  [7:0] col_in_356,
    input  [7:0] col_in_357,
    input  [7:0] col_in_358,
    input  [7:0] col_in_359,
    input  [7:0] col_in_360,
    input  [7:0] col_in_361,
    input  [7:0] col_in_362,
    input  [7:0] col_in_363,
    input  [7:0] col_in_364,
    input  [7:0] col_in_365,
    input  [7:0] col_in_366,
    input  [7:0] col_in_367,
    input  [7:0] col_in_368,
    input  [7:0] col_in_369,
    input  [7:0] col_in_370,
    input  [7:0] col_in_371,
    input  [7:0] col_in_372,
    input  [7:0] col_in_373,
    input  [7:0] col_in_374,
    input  [7:0] col_in_375,
    input  [7:0] col_in_376,
    input  [7:0] col_in_377,
    input  [7:0] col_in_378,
    input  [7:0] col_in_379,
    input  [7:0] col_in_380,
    input  [7:0] col_in_381,
    input  [7:0] col_in_382,
    input  [7:0] col_in_383,
    input  [7:0] col_in_384,
    input  [7:0] col_in_385,
    input  [7:0] col_in_386,
    input  [7:0] col_in_387,
    input  [7:0] col_in_388,
    input  [7:0] col_in_389,
    input  [7:0] col_in_390,
    input  [7:0] col_in_391,
    input  [7:0] col_in_392,
    input  [7:0] col_in_393,
    input  [7:0] col_in_394,
    input  [7:0] col_in_395,
    input  [7:0] col_in_396,
    input  [7:0] col_in_397,
    input  [7:0] col_in_398,
    input  [7:0] col_in_399,
    input  [7:0] col_in_400,
    input  [7:0] col_in_401,
    input  [7:0] col_in_402,
    input  [7:0] col_in_403,
    input  [7:0] col_in_404,
    input  [7:0] col_in_405,
    input  [7:0] col_in_406,
    input  [7:0] col_in_407,
    input  [7:0] col_in_408,
    input  [7:0] col_in_409,
    input  [7:0] col_in_410,
    input  [7:0] col_in_411,
    input  [7:0] col_in_412,
    input  [7:0] col_in_413,
    input  [7:0] col_in_414,
    input  [7:0] col_in_415,
    input  [7:0] col_in_416,
    input  [7:0] col_in_417,
    input  [7:0] col_in_418,
    input  [7:0] col_in_419,
    input  [7:0] col_in_420,
    input  [7:0] col_in_421,
    input  [7:0] col_in_422,
    input  [7:0] col_in_423,
    input  [7:0] col_in_424,
    input  [7:0] col_in_425,
    input  [7:0] col_in_426,
    input  [7:0] col_in_427,
    input  [7:0] col_in_428,
    input  [7:0] col_in_429,
    input  [7:0] col_in_430,
    input  [7:0] col_in_431,
    input  [7:0] col_in_432,
    input  [7:0] col_in_433,
    input  [7:0] col_in_434,
    input  [7:0] col_in_435,
    input  [7:0] col_in_436,
    input  [7:0] col_in_437,
    input  [7:0] col_in_438,
    input  [7:0] col_in_439,
    input  [7:0] col_in_440,
    input  [7:0] col_in_441,
    input  [7:0] col_in_442,
    input  [7:0] col_in_443,
    input  [7:0] col_in_444,
    input  [7:0] col_in_445,
    input  [7:0] col_in_446,
    input  [7:0] col_in_447,
    input  [7:0] col_in_448,
    input  [7:0] col_in_449,
    input  [7:0] col_in_450,
    input  [7:0] col_in_451,
    input  [7:0] col_in_452,
    input  [7:0] col_in_453,
    input  [7:0] col_in_454,
    input  [7:0] col_in_455,
    input  [7:0] col_in_456,
    input  [7:0] col_in_457,
    input  [7:0] col_in_458,
    input  [7:0] col_in_459,
    input  [7:0] col_in_460,
    input  [7:0] col_in_461,
    input  [7:0] col_in_462,
    input  [7:0] col_in_463,
    input  [7:0] col_in_464,
    input  [7:0] col_in_465,
    input  [7:0] col_in_466,
    input  [7:0] col_in_467,
    input  [7:0] col_in_468,
    input  [7:0] col_in_469,
    input  [7:0] col_in_470,
    input  [7:0] col_in_471,
    input  [7:0] col_in_472,
    input  [7:0] col_in_473,
    input  [7:0] col_in_474,
    input  [7:0] col_in_475,
    input  [7:0] col_in_476,
    input  [7:0] col_in_477,
    input  [7:0] col_in_478,
    input  [7:0] col_in_479,
    input  [7:0] col_in_480,
    input  [7:0] col_in_481,
    input  [7:0] col_in_482,
    input  [7:0] col_in_483,
    input  [7:0] col_in_484,
    input  [7:0] col_in_485,
    input  [7:0] col_in_486,
    input  [7:0] col_in_487,
    input  [7:0] col_in_488,
    input  [7:0] col_in_489,
    input  [7:0] col_in_490,
    input  [7:0] col_in_491,
    input  [7:0] col_in_492,
    input  [7:0] col_in_493,
    input  [7:0] col_in_494,
    input  [7:0] col_in_495,
    input  [7:0] col_in_496,
    input  [7:0] col_in_497,
    input  [7:0] col_in_498,
    input  [7:0] col_in_499,
    input  [7:0] col_in_500,
    input  [7:0] col_in_501,
    input  [7:0] col_in_502,
    input  [7:0] col_in_503,
    input  [7:0] col_in_504,
    input  [7:0] col_in_505,
    input  [7:0] col_in_506,
    input  [7:0] col_in_507,
    input  [7:0] col_in_508,
    input  [7:0] col_in_509,
    input  [7:0] col_in_510,
    input  [7:0] col_in_511,
    input  [7:0] col_in_512,
    input  [7:0] col_in_513,
    input  [7:0] col_in_514,
    input  [7:0] col_in_515,
    input  [7:0] col_in_516,
    input  [7:0] col_in_517,
    input  [7:0] col_in_518,
    input  [7:0] col_in_519,
    input  [7:0] col_in_520,
    input  [7:0] col_in_521,
    input  [7:0] col_in_522,
    input  [7:0] col_in_523,
    input  [7:0] col_in_524,
    input  [7:0] col_in_525,
    input  [7:0] col_in_526,
    input  [7:0] col_in_527,
    input  [7:0] col_in_528,
    input  [7:0] col_in_529,
    input  [7:0] col_in_530,
    input  [7:0] col_in_531,
    input  [7:0] col_in_532,
    input  [7:0] col_in_533,
    input  [7:0] col_in_534,
    input  [7:0] col_in_535,
    input  [7:0] col_in_536,
    input  [7:0] col_in_537,
    input  [7:0] col_in_538,
    input  [7:0] col_in_539,
    input  [7:0] col_in_540,
    input  [7:0] col_in_541,
    input  [7:0] col_in_542,
    input  [7:0] col_in_543,
    input  [7:0] col_in_544,
    input  [7:0] col_in_545,
    input  [7:0] col_in_546,
    input  [7:0] col_in_547,
    input  [7:0] col_in_548,
    input  [7:0] col_in_549,
    input  [7:0] col_in_550,
    input  [7:0] col_in_551,
    input  [7:0] col_in_552,
    input  [7:0] col_in_553,
    input  [7:0] col_in_554,
    input  [7:0] col_in_555,
    input  [7:0] col_in_556,
    input  [7:0] col_in_557,
    input  [7:0] col_in_558,
    input  [7:0] col_in_559,
    input  [7:0] col_in_560,
    input  [7:0] col_in_561,
    input  [7:0] col_in_562,
    input  [7:0] col_in_563,
    input  [7:0] col_in_564,
    input  [7:0] col_in_565,
    input  [7:0] col_in_566,
    input  [7:0] col_in_567,
    input  [7:0] col_in_568,
    input  [7:0] col_in_569,
    input  [7:0] col_in_570,
    input  [7:0] col_in_571,
    input  [7:0] col_in_572,
    input  [7:0] col_in_573,
    input  [7:0] col_in_574,
    input  [7:0] col_in_575,
    input  [7:0] col_in_576,
    input  [7:0] col_in_577,
    input  [7:0] col_in_578,
    input  [7:0] col_in_579,
    input  [7:0] col_in_580,
    input  [7:0] col_in_581,
    input  [7:0] col_in_582,
    input  [7:0] col_in_583,
    input  [7:0] col_in_584,
    input  [7:0] col_in_585,
    input  [7:0] col_in_586,
    input  [7:0] col_in_587,
    input  [7:0] col_in_588,
    input  [7:0] col_in_589,
    input  [7:0] col_in_590,
    input  [7:0] col_in_591,
    input  [7:0] col_in_592,
    input  [7:0] col_in_593,
    input  [7:0] col_in_594,
    input  [7:0] col_in_595,
    input  [7:0] col_in_596,
    input  [7:0] col_in_597,
    input  [7:0] col_in_598,
    input  [7:0] col_in_599,
    input  [7:0] col_in_600,
    input  [7:0] col_in_601,
    input  [7:0] col_in_602,
    input  [7:0] col_in_603,
    input  [7:0] col_in_604,
    input  [7:0] col_in_605,
    input  [7:0] col_in_606,
    input  [7:0] col_in_607,
    input  [7:0] col_in_608,
    input  [7:0] col_in_609,
    input  [7:0] col_in_610,
    input  [7:0] col_in_611,
    input  [7:0] col_in_612,
    input  [7:0] col_in_613,
    input  [7:0] col_in_614,
    input  [7:0] col_in_615,
    input  [7:0] col_in_616,
    input  [7:0] col_in_617,
    input  [7:0] col_in_618,
    input  [7:0] col_in_619,
    input  [7:0] col_in_620,
    input  [7:0] col_in_621,
    input  [7:0] col_in_622,
    input  [7:0] col_in_623,
    input  [7:0] col_in_624,
    input  [7:0] col_in_625,
    input  [7:0] col_in_626,
    input  [7:0] col_in_627,
    input  [7:0] col_in_628,
    input  [7:0] col_in_629,
    input  [7:0] col_in_630,
    input  [7:0] col_in_631,
    input  [7:0] col_in_632,
    input  [7:0] col_in_633,
    input  [7:0] col_in_634,
    input  [7:0] col_in_635,
    input  [7:0] col_in_636,
    input  [7:0] col_in_637,
    input  [7:0] col_in_638,
    input  [7:0] col_in_639,
    input  [7:0] col_in_640,
    input  [7:0] col_in_641,
    input  [7:0] col_in_642,
    input  [7:0] col_in_643,
    input  [7:0] col_in_644,
    input  [7:0] col_in_645,
    input  [7:0] col_in_646,
    input  [7:0] col_in_647,
    input  [7:0] col_in_648,
    input  [7:0] col_in_649,
    input  [7:0] col_in_650,
    input  [7:0] col_in_651,
    input  [7:0] col_in_652,
    input  [7:0] col_in_653,
    input  [7:0] col_in_654,
    input  [7:0] col_in_655,
    input  [7:0] col_in_656,
    input  [7:0] col_in_657,
    input  [7:0] col_in_658,
    input  [7:0] col_in_659,
    input  [7:0] col_in_660,
    input  [7:0] col_in_661,
    input  [7:0] col_in_662,
    input  [7:0] col_in_663,
    input  [7:0] col_in_664,
    input  [7:0] col_in_665,
    input  [7:0] col_in_666,
    input  [7:0] col_in_667,
    input  [7:0] col_in_668,
    input  [7:0] col_in_669,
    input  [7:0] col_in_670,
    input  [7:0] col_in_671,
    input  [7:0] col_in_672,
    input  [7:0] col_in_673,
    input  [7:0] col_in_674,
    input  [7:0] col_in_675,
    input  [7:0] col_in_676,
    input  [7:0] col_in_677,
    input  [7:0] col_in_678,
    input  [7:0] col_in_679,
    input  [7:0] col_in_680,
    input  [7:0] col_in_681,
    input  [7:0] col_in_682,
    input  [7:0] col_in_683,
    input  [7:0] col_in_684,
    input  [7:0] col_in_685,
    input  [7:0] col_in_686,
    input  [7:0] col_in_687,
    input  [7:0] col_in_688,
    input  [7:0] col_in_689,
    input  [7:0] col_in_690,
    input  [7:0] col_in_691,
    input  [7:0] col_in_692,
    input  [7:0] col_in_693,
    input  [7:0] col_in_694,
    input  [7:0] col_in_695,
    input  [7:0] col_in_696,
    input  [7:0] col_in_697,
    input  [7:0] col_in_698,
    input  [7:0] col_in_699,
    input  [7:0] col_in_700,
    input  [7:0] col_in_701,
    input  [7:0] col_in_702,
    input  [7:0] col_in_703,
    input  [7:0] col_in_704,
    input  [7:0] col_in_705,
    input  [7:0] col_in_706,
    input  [7:0] col_in_707,
    input  [7:0] col_in_708,
    input  [7:0] col_in_709,
    input  [7:0] col_in_710,
    input  [7:0] col_in_711,
    input  [7:0] col_in_712,
    input  [7:0] col_in_713,
    input  [7:0] col_in_714,
    input  [7:0] col_in_715,
    input  [7:0] col_in_716,
    input  [7:0] col_in_717,
    input  [7:0] col_in_718,
    input  [7:0] col_in_719,
    input  [7:0] col_in_720,
    input  [7:0] col_in_721,
    input  [7:0] col_in_722,
    input  [7:0] col_in_723,
    input  [7:0] col_in_724,
    input  [7:0] col_in_725,
    input  [7:0] col_in_726,
    input  [7:0] col_in_727,
    input  [7:0] col_in_728,
    input  [7:0] col_in_729,
    input  [7:0] col_in_730,
    input  [7:0] col_in_731,
    input  [7:0] col_in_732,
    input  [7:0] col_in_733,
    input  [7:0] col_in_734,
    input  [7:0] col_in_735,
    input  [7:0] col_in_736,
    input  [7:0] col_in_737,
    input  [7:0] col_in_738,
    input  [7:0] col_in_739,
    input  [7:0] col_in_740,
    input  [7:0] col_in_741,
    input  [7:0] col_in_742,
    input  [7:0] col_in_743,
    input  [7:0] col_in_744,
    input  [7:0] col_in_745,
    input  [7:0] col_in_746,
    input  [7:0] col_in_747,
    input  [7:0] col_in_748,
    input  [7:0] col_in_749,
    input  [7:0] col_in_750,
    input  [7:0] col_in_751,
    input  [7:0] col_in_752,
    input  [7:0] col_in_753,
    input  [7:0] col_in_754,
    input  [7:0] col_in_755,
    input  [7:0] col_in_756,
    input  [7:0] col_in_757,
    input  [7:0] col_in_758,
    input  [7:0] col_in_759,
    input  [7:0] col_in_760,
    input  [7:0] col_in_761,
    input  [7:0] col_in_762,
    input  [7:0] col_in_763,
    input  [7:0] col_in_764,
    input  [7:0] col_in_765,
    input  [7:0] col_in_766,
    input  [7:0] col_in_767,
    input  [7:0] col_in_768,
    input  [7:0] col_in_769,
    input  [7:0] col_in_770,
    input  [7:0] col_in_771,
    input  [7:0] col_in_772,
    input  [7:0] col_in_773,
    input  [7:0] col_in_774,
    input  [7:0] col_in_775,
    input  [7:0] col_in_776,
    input  [7:0] col_in_777,
    input  [7:0] col_in_778,
    input  [7:0] col_in_779,
    input  [7:0] col_in_780,
    input  [7:0] col_in_781,
    input  [7:0] col_in_782,
    input  [7:0] col_in_783,
    input  [7:0] col_in_784,
    input  [7:0] col_in_785,
    input  [7:0] col_in_786,
    input  [7:0] col_in_787,
    input  [7:0] col_in_788,
    input  [7:0] col_in_789,
    input  [7:0] col_in_790,
    input  [7:0] col_in_791,
    input  [7:0] col_in_792,
    input  [7:0] col_in_793,
    input  [7:0] col_in_794,
    input  [7:0] col_in_795,
    input  [7:0] col_in_796,
    input  [7:0] col_in_797,
    input  [7:0] col_in_798,
    input  [7:0] col_in_799,
    input  [7:0] col_in_800,
    input  [7:0] col_in_801,
    input  [7:0] col_in_802,
    input  [7:0] col_in_803,
    input  [7:0] col_in_804,
    input  [7:0] col_in_805,
    input  [7:0] col_in_806,
    input  [7:0] col_in_807,
    input  [7:0] col_in_808,
    input  [7:0] col_in_809,
    input  [7:0] col_in_810,
    input  [7:0] col_in_811,
    input  [7:0] col_in_812,
    input  [7:0] col_in_813,
    input  [7:0] col_in_814,
    input  [7:0] col_in_815,
    input  [7:0] col_in_816,
    input  [7:0] col_in_817,
    input  [7:0] col_in_818,
    input  [7:0] col_in_819,
    input  [7:0] col_in_820,
    input  [7:0] col_in_821,
    input  [7:0] col_in_822,
    input  [7:0] col_in_823,
    input  [7:0] col_in_824,
    input  [7:0] col_in_825,
    input  [7:0] col_in_826,
    input  [7:0] col_in_827,
    input  [7:0] col_in_828,
    input  [7:0] col_in_829,
    input  [7:0] col_in_830,
    input  [7:0] col_in_831,
    input  [7:0] col_in_832,
    input  [7:0] col_in_833,
    input  [7:0] col_in_834,
    input  [7:0] col_in_835,
    input  [7:0] col_in_836,
    input  [7:0] col_in_837,
    input  [7:0] col_in_838,
    input  [7:0] col_in_839,
    input  [7:0] col_in_840,
    input  [7:0] col_in_841,
    input  [7:0] col_in_842,
    input  [7:0] col_in_843,
    input  [7:0] col_in_844,
    input  [7:0] col_in_845,
    input  [7:0] col_in_846,
    input  [7:0] col_in_847,
    input  [7:0] col_in_848,
    input  [7:0] col_in_849,
    input  [7:0] col_in_850,
    input  [7:0] col_in_851,
    input  [7:0] col_in_852,
    input  [7:0] col_in_853,
    input  [7:0] col_in_854,
    input  [7:0] col_in_855,
    input  [7:0] col_in_856,
    input  [7:0] col_in_857,
    input  [7:0] col_in_858,
    input  [7:0] col_in_859,
    input  [7:0] col_in_860,
    input  [7:0] col_in_861,
    input  [7:0] col_in_862,
    input  [7:0] col_in_863,
    input  [7:0] col_in_864,
    input  [7:0] col_in_865,
    input  [7:0] col_in_866,
    input  [7:0] col_in_867,
    input  [7:0] col_in_868,
    input  [7:0] col_in_869,
    input  [7:0] col_in_870,
    input  [7:0] col_in_871,
    input  [7:0] col_in_872,
    input  [7:0] col_in_873,
    input  [7:0] col_in_874,
    input  [7:0] col_in_875,
    input  [7:0] col_in_876,
    input  [7:0] col_in_877,
    input  [7:0] col_in_878,
    input  [7:0] col_in_879,
    input  [7:0] col_in_880,
    input  [7:0] col_in_881,
    input  [7:0] col_in_882,
    input  [7:0] col_in_883,
    input  [7:0] col_in_884,
    input  [7:0] col_in_885,
    input  [7:0] col_in_886,
    input  [7:0] col_in_887,
    input  [7:0] col_in_888,
    input  [7:0] col_in_889,
    input  [7:0] col_in_890,
    input  [7:0] col_in_891,
    input  [7:0] col_in_892,
    input  [7:0] col_in_893,
    input  [7:0] col_in_894,
    input  [7:0] col_in_895,
    input  [7:0] col_in_896,
    input  [7:0] col_in_897,
    input  [7:0] col_in_898,
    input  [7:0] col_in_899,
    input  [7:0] col_in_900,
    input  [7:0] col_in_901,
    input  [7:0] col_in_902,
    input  [7:0] col_in_903,
    input  [7:0] col_in_904,
    input  [7:0] col_in_905,
    input  [7:0] col_in_906,
    input  [7:0] col_in_907,
    input  [7:0] col_in_908,
    input  [7:0] col_in_909,
    input  [7:0] col_in_910,
    input  [7:0] col_in_911,
    input  [7:0] col_in_912,
    input  [7:0] col_in_913,
    input  [7:0] col_in_914,
    input  [7:0] col_in_915,
    input  [7:0] col_in_916,
    input  [7:0] col_in_917,
    input  [7:0] col_in_918,
    input  [7:0] col_in_919,
    input  [7:0] col_in_920,
    input  [7:0] col_in_921,
    input  [7:0] col_in_922,
    input  [7:0] col_in_923,
    input  [7:0] col_in_924,
    input  [7:0] col_in_925,
    input  [7:0] col_in_926,
    input  [7:0] col_in_927,
    input  [7:0] col_in_928,
    input  [7:0] col_in_929,
    input  [7:0] col_in_930,
    input  [7:0] col_in_931,
    input  [7:0] col_in_932,
    input  [7:0] col_in_933,
    input  [7:0] col_in_934,
    input  [7:0] col_in_935,
    input  [7:0] col_in_936,
    input  [7:0] col_in_937,
    input  [7:0] col_in_938,
    input  [7:0] col_in_939,
    input  [7:0] col_in_940,
    input  [7:0] col_in_941,
    input  [7:0] col_in_942,
    input  [7:0] col_in_943,
    input  [7:0] col_in_944,
    input  [7:0] col_in_945,
    input  [7:0] col_in_946,
    input  [7:0] col_in_947,
    input  [7:0] col_in_948,
    input  [7:0] col_in_949,
    input  [7:0] col_in_950,
    input  [7:0] col_in_951,
    input  [7:0] col_in_952,
    input  [7:0] col_in_953,
    input  [7:0] col_in_954,
    input  [7:0] col_in_955,
    input  [7:0] col_in_956,
    input  [7:0] col_in_957,
    input  [7:0] col_in_958,
    input  [7:0] col_in_959,
    input  [7:0] col_in_960,
    input  [7:0] col_in_961,
    input  [7:0] col_in_962,
    input  [7:0] col_in_963,
    input  [7:0] col_in_964,
    input  [7:0] col_in_965,
    input  [7:0] col_in_966,
    input  [7:0] col_in_967,
    input  [7:0] col_in_968,
    input  [7:0] col_in_969,
    input  [7:0] col_in_970,
    input  [7:0] col_in_971,
    input  [7:0] col_in_972,
    input  [7:0] col_in_973,
    input  [7:0] col_in_974,
    input  [7:0] col_in_975,
    input  [7:0] col_in_976,
    input  [7:0] col_in_977,
    input  [7:0] col_in_978,
    input  [7:0] col_in_979,
    input  [7:0] col_in_980,
    input  [7:0] col_in_981,
    input  [7:0] col_in_982,
    input  [7:0] col_in_983,
    input  [7:0] col_in_984,
    input  [7:0] col_in_985,
    input  [7:0] col_in_986,
    input  [7:0] col_in_987,
    input  [7:0] col_in_988,
    input  [7:0] col_in_989,
    input  [7:0] col_in_990,
    input  [7:0] col_in_991,
    input  [7:0] col_in_992,
    input  [7:0] col_in_993,
    input  [7:0] col_in_994,
    input  [7:0] col_in_995,
    input  [7:0] col_in_996,
    input  [7:0] col_in_997,
    input  [7:0] col_in_998,
    input  [7:0] col_in_999,
    input  [7:0] col_in_1000,
    input  [7:0] col_in_1001,
    input  [7:0] col_in_1002,
    input  [7:0] col_in_1003,
    input  [7:0] col_in_1004,
    input  [7:0] col_in_1005,
    input  [7:0] col_in_1006,
    input  [7:0] col_in_1007,
    input  [7:0] col_in_1008,
    input  [7:0] col_in_1009,
    input  [7:0] col_in_1010,
    input  [7:0] col_in_1011,
    input  [7:0] col_in_1012,
    input  [7:0] col_in_1013,
    input  [7:0] col_in_1014,
    input  [7:0] col_in_1015,
    input  [7:0] col_in_1016,
    input  [7:0] col_in_1017,
    input  [7:0] col_in_1018,
    input  [7:0] col_in_1019,
    input  [7:0] col_in_1020,
    input  [7:0] col_in_1021,
    input  [7:0] col_in_1022,
    input  [7:0] col_in_1023,
    input  [7:0] col_in_1024,
    input  [7:0] col_in_1025,
    input  [7:0] col_in_1026,
    input  [7:0] col_in_1027,
    input  [7:0] col_in_1028,
    input  [7:0] col_in_1029,
    input  [7:0] col_in_1030,
    input  [7:0] col_in_1031,
    input  [7:0] col_in_1032,
    input  [7:0] col_in_1033,
    input  [7:0] col_in_1034,
    input  [7:0] col_in_1035,
    input  [7:0] col_in_1036,
    input  [7:0] col_in_1037,
    input  [7:0] col_in_1038,
    input  [7:0] col_in_1039,
    input  [7:0] col_in_1040,
    input  [7:0] col_in_1041,
    input  [7:0] col_in_1042,
    input  [7:0] col_in_1043,
    input  [7:0] col_in_1044,
    input  [7:0] col_in_1045,
    input  [7:0] col_in_1046,
    input  [7:0] col_in_1047,
    input  [7:0] col_in_1048,
    input  [7:0] col_in_1049,
    input  [7:0] col_in_1050,
    input  [7:0] col_in_1051,
    input  [7:0] col_in_1052,
    input  [7:0] col_in_1053,
    input  [7:0] col_in_1054,
    input  [7:0] col_in_1055,
    input  [7:0] col_in_1056,
    input  [7:0] col_in_1057,
    input  [7:0] col_in_1058,
    input  [7:0] col_in_1059,
    input  [7:0] col_in_1060,
    input  [7:0] col_in_1061,
    input  [7:0] col_in_1062,
    input  [7:0] col_in_1063,
    input  [7:0] col_in_1064,
    input  [7:0] col_in_1065,
    input  [7:0] col_in_1066,
    input  [7:0] col_in_1067,
    input  [7:0] col_in_1068,
    input  [7:0] col_in_1069,
    input  [7:0] col_in_1070,
    input  [7:0] col_in_1071,
    input  [7:0] col_in_1072,
    input  [7:0] col_in_1073,
    input  [7:0] col_in_1074,
    input  [7:0] col_in_1075,
    input  [7:0] col_in_1076,
    input  [7:0] col_in_1077,
    input  [7:0] col_in_1078,
    input  [7:0] col_in_1079,
    input  [7:0] col_in_1080,
    input  [7:0] col_in_1081,
    input  [7:0] col_in_1082,
    input  [7:0] col_in_1083,
    input  [7:0] col_in_1084,
    input  [7:0] col_in_1085,
    input  [7:0] col_in_1086,
    input  [7:0] col_in_1087,
    input  [7:0] col_in_1088,
    input  [7:0] col_in_1089,
    input  [7:0] col_in_1090,
    input  [7:0] col_in_1091,
    input  [7:0] col_in_1092,
    input  [7:0] col_in_1093,
    input  [7:0] col_in_1094,
    input  [7:0] col_in_1095,
    input  [7:0] col_in_1096,
    input  [7:0] col_in_1097,
    input  [7:0] col_in_1098,
    input  [7:0] col_in_1099,
    input  [7:0] col_in_1100,
    input  [7:0] col_in_1101,
    input  [7:0] col_in_1102,
    input  [7:0] col_in_1103,
    input  [7:0] col_in_1104,
    input  [7:0] col_in_1105,
    input  [7:0] col_in_1106,
    input  [7:0] col_in_1107,
    input  [7:0] col_in_1108,
    input  [7:0] col_in_1109,
    input  [7:0] col_in_1110,
    input  [7:0] col_in_1111,
    input  [7:0] col_in_1112,
    input  [7:0] col_in_1113,
    input  [7:0] col_in_1114,
    input  [7:0] col_in_1115,
    input  [7:0] col_in_1116,
    input  [7:0] col_in_1117,
    input  [7:0] col_in_1118,
    input  [7:0] col_in_1119,
    input  [7:0] col_in_1120,
    input  [7:0] col_in_1121,
    input  [7:0] col_in_1122,
    input  [7:0] col_in_1123,
    input  [7:0] col_in_1124,
    input  [7:0] col_in_1125,
    input  [7:0] col_in_1126,
    input  [7:0] col_in_1127,
    input  [7:0] col_in_1128,
    input  [7:0] col_in_1129,
    input  [7:0] col_in_1130,
    input  [7:0] col_in_1131,
    input  [7:0] col_in_1132,
    input  [7:0] col_in_1133,
    input  [7:0] col_in_1134,
    input  [7:0] col_in_1135,
    input  [7:0] col_in_1136,
    input  [7:0] col_in_1137,
    input  [7:0] col_in_1138,
    input  [7:0] col_in_1139,
    input  [7:0] col_in_1140,
    input  [7:0] col_in_1141,
    input  [7:0] col_in_1142,
    input  [7:0] col_in_1143,
    input  [7:0] col_in_1144,
    input  [7:0] col_in_1145,
    input  [7:0] col_in_1146,
    input  [7:0] col_in_1147,
    input  [7:0] col_in_1148,
    input  [7:0] col_in_1149,
    input  [7:0] col_in_1150,
    input  [7:0] col_in_1151,
    input  [7:0] col_in_1152,
    input  [7:0] col_in_1153,
    input  [7:0] col_in_1154,
    input  [7:0] col_in_1155,
    input  [7:0] col_in_1156,
    input  [7:0] col_in_1157,
    input  [7:0] col_in_1158,
    input  [7:0] col_in_1159,
    input  [7:0] col_in_1160,
    input  [7:0] col_in_1161,
    input  [7:0] col_in_1162,
    input  [7:0] col_in_1163,
    input  [7:0] col_in_1164,
    input  [7:0] col_in_1165,
    input  [7:0] col_in_1166,
    input  [7:0] col_in_1167,
    input  [7:0] col_in_1168,
    input  [7:0] col_in_1169,
    input  [7:0] col_in_1170,
    input  [7:0] col_in_1171,
    input  [7:0] col_in_1172,
    input  [7:0] col_in_1173,
    input  [7:0] col_in_1174,
    input  [7:0] col_in_1175,
    input  [7:0] col_in_1176,
    input  [7:0] col_in_1177,
    input  [7:0] col_in_1178,
    input  [7:0] col_in_1179,
    input  [7:0] col_in_1180,
    input  [7:0] col_in_1181,
    input  [7:0] col_in_1182,
    input  [7:0] col_in_1183,
    input  [7:0] col_in_1184,
    input  [7:0] col_in_1185,
    input  [7:0] col_in_1186,
    input  [7:0] col_in_1187,
    input  [7:0] col_in_1188,
    input  [7:0] col_in_1189,
    input  [7:0] col_in_1190,
    input  [7:0] col_in_1191,
    input  [7:0] col_in_1192,
    input  [7:0] col_in_1193,
    input  [7:0] col_in_1194,
    input  [7:0] col_in_1195,
    input  [7:0] col_in_1196,
    input  [7:0] col_in_1197,
    input  [7:0] col_in_1198,
    input  [7:0] col_in_1199,
    input  [7:0] col_in_1200,
    input  [7:0] col_in_1201,
    input  [7:0] col_in_1202,
    input  [7:0] col_in_1203,
    input  [7:0] col_in_1204,
    input  [7:0] col_in_1205,
    input  [7:0] col_in_1206,
    input  [7:0] col_in_1207,
    input  [7:0] col_in_1208,
    input  [7:0] col_in_1209,
    input  [7:0] col_in_1210,
    input  [7:0] col_in_1211,
    input  [7:0] col_in_1212,
    input  [7:0] col_in_1213,
    input  [7:0] col_in_1214,
    input  [7:0] col_in_1215,
    input  [7:0] col_in_1216,
    input  [7:0] col_in_1217,
    input  [7:0] col_in_1218,
    input  [7:0] col_in_1219,
    input  [7:0] col_in_1220,
    input  [7:0] col_in_1221,
    input  [7:0] col_in_1222,
    input  [7:0] col_in_1223,
    input  [7:0] col_in_1224,
    input  [7:0] col_in_1225,
    input  [7:0] col_in_1226,
    input  [7:0] col_in_1227,
    input  [7:0] col_in_1228,
    input  [7:0] col_in_1229,
    input  [7:0] col_in_1230,
    input  [7:0] col_in_1231,
    input  [7:0] col_in_1232,
    input  [7:0] col_in_1233,
    input  [7:0] col_in_1234,
    input  [7:0] col_in_1235,
    input  [7:0] col_in_1236,
    input  [7:0] col_in_1237,
    input  [7:0] col_in_1238,
    input  [7:0] col_in_1239,
    input  [7:0] col_in_1240,
    input  [7:0] col_in_1241,
    input  [7:0] col_in_1242,
    input  [7:0] col_in_1243,
    input  [7:0] col_in_1244,
    input  [7:0] col_in_1245,
    input  [7:0] col_in_1246,
    input  [7:0] col_in_1247,
    input  [7:0] col_in_1248,
    input  [7:0] col_in_1249,
    input  [7:0] col_in_1250,
    input  [7:0] col_in_1251,
    input  [7:0] col_in_1252,
    input  [7:0] col_in_1253,
    input  [7:0] col_in_1254,
    input  [7:0] col_in_1255,
    input  [7:0] col_in_1256,
    input  [7:0] col_in_1257,
    input  [7:0] col_in_1258,
    input  [7:0] col_in_1259,
    input  [7:0] col_in_1260,
    input  [7:0] col_in_1261,
    input  [7:0] col_in_1262,
    input  [7:0] col_in_1263,
    input  [7:0] col_in_1264,
    input  [7:0] col_in_1265,
    input  [7:0] col_in_1266,
    input  [7:0] col_in_1267,
    input  [7:0] col_in_1268,
    input  [7:0] col_in_1269,
    input  [7:0] col_in_1270,
    input  [7:0] col_in_1271,
    input  [7:0] col_in_1272,
    input  [7:0] col_in_1273,
    input  [7:0] col_in_1274,
    input  [7:0] col_in_1275,
    input  [7:0] col_in_1276,
    input  [7:0] col_in_1277,
    input  [7:0] col_in_1278,
    input  [7:0] col_in_1279,
    input  [7:0] col_in_1280,
    input  [7:0] col_in_1281,
    input  [7:0] col_in_1282,
    input  [7:0] col_in_1283,
    input  [7:0] col_in_1284,
    input  [7:0] col_in_1285,
    input  [7:0] col_in_1286,
    input  [7:0] col_in_1287,

    output [5:0] col_out_0,
    output [5:0] col_out_1,
    output [5:0] col_out_2,
    output [5:0] col_out_3,
    output [5:0] col_out_4,
    output [5:0] col_out_5,
    output [5:0] col_out_6,
    output [5:0] col_out_7,
    output [5:0] col_out_8,
    output [5:0] col_out_9,
    output [5:0] col_out_10,
    output [5:0] col_out_11,
    output [5:0] col_out_12,
    output [5:0] col_out_13,
    output [5:0] col_out_14,
    output [5:0] col_out_15,
    output [5:0] col_out_16,
    output [5:0] col_out_17,
    output [5:0] col_out_18,
    output [5:0] col_out_19,
    output [5:0] col_out_20,
    output [5:0] col_out_21,
    output [5:0] col_out_22,
    output [5:0] col_out_23,
    output [5:0] col_out_24,
    output [5:0] col_out_25,
    output [5:0] col_out_26,
    output [5:0] col_out_27,
    output [5:0] col_out_28,
    output [5:0] col_out_29,
    output [5:0] col_out_30,
    output [5:0] col_out_31,
    output [5:0] col_out_32,
    output [5:0] col_out_33,
    output [5:0] col_out_34,
    output [5:0] col_out_35,
    output [5:0] col_out_36,
    output [5:0] col_out_37,
    output [5:0] col_out_38,
    output [5:0] col_out_39,
    output [5:0] col_out_40,
    output [5:0] col_out_41,
    output [5:0] col_out_42,
    output [5:0] col_out_43,
    output [5:0] col_out_44,
    output [5:0] col_out_45,
    output [5:0] col_out_46,
    output [5:0] col_out_47,
    output [5:0] col_out_48,
    output [5:0] col_out_49,
    output [5:0] col_out_50,
    output [5:0] col_out_51,
    output [5:0] col_out_52,
    output [5:0] col_out_53,
    output [5:0] col_out_54,
    output [5:0] col_out_55,
    output [5:0] col_out_56,
    output [5:0] col_out_57,
    output [5:0] col_out_58,
    output [5:0] col_out_59,
    output [5:0] col_out_60,
    output [5:0] col_out_61,
    output [5:0] col_out_62,
    output [5:0] col_out_63,
    output [5:0] col_out_64,
    output [5:0] col_out_65,
    output [5:0] col_out_66,
    output [5:0] col_out_67,
    output [5:0] col_out_68,
    output [5:0] col_out_69,
    output [5:0] col_out_70,
    output [5:0] col_out_71,
    output [5:0] col_out_72,
    output [5:0] col_out_73,
    output [5:0] col_out_74,
    output [5:0] col_out_75,
    output [5:0] col_out_76,
    output [5:0] col_out_77,
    output [5:0] col_out_78,
    output [5:0] col_out_79,
    output [5:0] col_out_80,
    output [5:0] col_out_81,
    output [5:0] col_out_82,
    output [5:0] col_out_83,
    output [5:0] col_out_84,
    output [5:0] col_out_85,
    output [5:0] col_out_86,
    output [5:0] col_out_87,
    output [5:0] col_out_88,
    output [5:0] col_out_89,
    output [5:0] col_out_90,
    output [5:0] col_out_91,
    output [5:0] col_out_92,
    output [5:0] col_out_93,
    output [5:0] col_out_94,
    output [5:0] col_out_95,
    output [5:0] col_out_96,
    output [5:0] col_out_97,
    output [5:0] col_out_98,
    output [5:0] col_out_99,
    output [5:0] col_out_100,
    output [5:0] col_out_101,
    output [5:0] col_out_102,
    output [5:0] col_out_103,
    output [5:0] col_out_104,
    output [5:0] col_out_105,
    output [5:0] col_out_106,
    output [5:0] col_out_107,
    output [5:0] col_out_108,
    output [5:0] col_out_109,
    output [5:0] col_out_110,
    output [5:0] col_out_111,
    output [5:0] col_out_112,
    output [5:0] col_out_113,
    output [5:0] col_out_114,
    output [5:0] col_out_115,
    output [5:0] col_out_116,
    output [5:0] col_out_117,
    output [5:0] col_out_118,
    output [5:0] col_out_119,
    output [5:0] col_out_120,
    output [5:0] col_out_121,
    output [5:0] col_out_122,
    output [5:0] col_out_123,
    output [5:0] col_out_124,
    output [5:0] col_out_125,
    output [5:0] col_out_126,
    output [5:0] col_out_127,
    output [5:0] col_out_128,
    output [5:0] col_out_129,
    output [5:0] col_out_130,
    output [5:0] col_out_131,
    output [5:0] col_out_132,
    output [5:0] col_out_133,
    output [5:0] col_out_134,
    output [5:0] col_out_135,
    output [5:0] col_out_136,
    output [5:0] col_out_137,
    output [5:0] col_out_138,
    output [5:0] col_out_139,
    output [5:0] col_out_140,
    output [5:0] col_out_141,
    output [5:0] col_out_142,
    output [5:0] col_out_143,
    output [5:0] col_out_144,
    output [5:0] col_out_145,
    output [5:0] col_out_146,
    output [5:0] col_out_147,
    output [5:0] col_out_148,
    output [5:0] col_out_149,
    output [5:0] col_out_150,
    output [5:0] col_out_151,
    output [5:0] col_out_152,
    output [5:0] col_out_153,
    output [5:0] col_out_154,
    output [5:0] col_out_155,
    output [5:0] col_out_156,
    output [5:0] col_out_157,
    output [5:0] col_out_158,
    output [5:0] col_out_159,
    output [5:0] col_out_160,
    output [5:0] col_out_161,
    output [5:0] col_out_162,
    output [5:0] col_out_163,
    output [5:0] col_out_164,
    output [5:0] col_out_165,
    output [5:0] col_out_166,
    output [5:0] col_out_167,
    output [5:0] col_out_168,
    output [5:0] col_out_169,
    output [5:0] col_out_170,
    output [5:0] col_out_171,
    output [5:0] col_out_172,
    output [5:0] col_out_173,
    output [5:0] col_out_174,
    output [5:0] col_out_175,
    output [5:0] col_out_176,
    output [5:0] col_out_177,
    output [5:0] col_out_178,
    output [5:0] col_out_179,
    output [5:0] col_out_180,
    output [5:0] col_out_181,
    output [5:0] col_out_182,
    output [5:0] col_out_183,
    output [5:0] col_out_184,
    output [5:0] col_out_185,
    output [5:0] col_out_186,
    output [5:0] col_out_187,
    output [5:0] col_out_188,
    output [5:0] col_out_189,
    output [5:0] col_out_190,
    output [5:0] col_out_191,
    output [5:0] col_out_192,
    output [5:0] col_out_193,
    output [5:0] col_out_194,
    output [5:0] col_out_195,
    output [5:0] col_out_196,
    output [5:0] col_out_197,
    output [5:0] col_out_198,
    output [5:0] col_out_199,
    output [5:0] col_out_200,
    output [5:0] col_out_201,
    output [5:0] col_out_202,
    output [5:0] col_out_203,
    output [5:0] col_out_204,
    output [5:0] col_out_205,
    output [5:0] col_out_206,
    output [5:0] col_out_207,
    output [5:0] col_out_208,
    output [5:0] col_out_209,
    output [5:0] col_out_210,
    output [5:0] col_out_211,
    output [5:0] col_out_212,
    output [5:0] col_out_213,
    output [5:0] col_out_214,
    output [5:0] col_out_215,
    output [5:0] col_out_216,
    output [5:0] col_out_217,
    output [5:0] col_out_218,
    output [5:0] col_out_219,
    output [5:0] col_out_220,
    output [5:0] col_out_221,
    output [5:0] col_out_222,
    output [5:0] col_out_223,
    output [5:0] col_out_224,
    output [5:0] col_out_225,
    output [5:0] col_out_226,
    output [5:0] col_out_227,
    output [5:0] col_out_228,
    output [5:0] col_out_229,
    output [5:0] col_out_230,
    output [5:0] col_out_231,
    output [5:0] col_out_232,
    output [5:0] col_out_233,
    output [5:0] col_out_234,
    output [5:0] col_out_235,
    output [5:0] col_out_236,
    output [5:0] col_out_237,
    output [5:0] col_out_238,
    output [5:0] col_out_239,
    output [5:0] col_out_240,
    output [5:0] col_out_241,
    output [5:0] col_out_242,
    output [5:0] col_out_243,
    output [5:0] col_out_244,
    output [5:0] col_out_245,
    output [5:0] col_out_246,
    output [5:0] col_out_247,
    output [5:0] col_out_248,
    output [5:0] col_out_249,
    output [5:0] col_out_250,
    output [5:0] col_out_251,
    output [5:0] col_out_252,
    output [5:0] col_out_253,
    output [5:0] col_out_254,
    output [5:0] col_out_255,
    output [5:0] col_out_256,
    output [5:0] col_out_257,
    output [5:0] col_out_258,
    output [5:0] col_out_259,
    output [5:0] col_out_260,
    output [5:0] col_out_261,
    output [5:0] col_out_262,
    output [5:0] col_out_263,
    output [5:0] col_out_264,
    output [5:0] col_out_265,
    output [5:0] col_out_266,
    output [5:0] col_out_267,
    output [5:0] col_out_268,
    output [5:0] col_out_269,
    output [5:0] col_out_270,
    output [5:0] col_out_271,
    output [5:0] col_out_272,
    output [5:0] col_out_273,
    output [5:0] col_out_274,
    output [5:0] col_out_275,
    output [5:0] col_out_276,
    output [5:0] col_out_277,
    output [5:0] col_out_278,
    output [5:0] col_out_279,
    output [5:0] col_out_280,
    output [5:0] col_out_281,
    output [5:0] col_out_282,
    output [5:0] col_out_283,
    output [5:0] col_out_284,
    output [5:0] col_out_285,
    output [5:0] col_out_286,
    output [5:0] col_out_287,
    output [5:0] col_out_288,
    output [5:0] col_out_289,
    output [5:0] col_out_290,
    output [5:0] col_out_291,
    output [5:0] col_out_292,
    output [5:0] col_out_293,
    output [5:0] col_out_294,
    output [5:0] col_out_295,
    output [5:0] col_out_296,
    output [5:0] col_out_297,
    output [5:0] col_out_298,
    output [5:0] col_out_299,
    output [5:0] col_out_300,
    output [5:0] col_out_301,
    output [5:0] col_out_302,
    output [5:0] col_out_303,
    output [5:0] col_out_304,
    output [5:0] col_out_305,
    output [5:0] col_out_306,
    output [5:0] col_out_307,
    output [5:0] col_out_308,
    output [5:0] col_out_309,
    output [5:0] col_out_310,
    output [5:0] col_out_311,
    output [5:0] col_out_312,
    output [5:0] col_out_313,
    output [5:0] col_out_314,
    output [5:0] col_out_315,
    output [5:0] col_out_316,
    output [5:0] col_out_317,
    output [5:0] col_out_318,
    output [5:0] col_out_319,
    output [5:0] col_out_320,
    output [5:0] col_out_321,
    output [5:0] col_out_322,
    output [5:0] col_out_323,
    output [5:0] col_out_324,
    output [5:0] col_out_325,
    output [5:0] col_out_326,
    output [5:0] col_out_327,
    output [5:0] col_out_328,
    output [5:0] col_out_329,
    output [5:0] col_out_330,
    output [5:0] col_out_331,
    output [5:0] col_out_332,
    output [5:0] col_out_333,
    output [5:0] col_out_334,
    output [5:0] col_out_335,
    output [5:0] col_out_336,
    output [5:0] col_out_337,
    output [5:0] col_out_338,
    output [5:0] col_out_339,
    output [5:0] col_out_340,
    output [5:0] col_out_341,
    output [5:0] col_out_342,
    output [5:0] col_out_343,
    output [5:0] col_out_344,
    output [5:0] col_out_345,
    output [5:0] col_out_346,
    output [5:0] col_out_347,
    output [5:0] col_out_348,
    output [5:0] col_out_349,
    output [5:0] col_out_350,
    output [5:0] col_out_351,
    output [5:0] col_out_352,
    output [5:0] col_out_353,
    output [5:0] col_out_354,
    output [5:0] col_out_355,
    output [5:0] col_out_356,
    output [5:0] col_out_357,
    output [5:0] col_out_358,
    output [5:0] col_out_359,
    output [5:0] col_out_360,
    output [5:0] col_out_361,
    output [5:0] col_out_362,
    output [5:0] col_out_363,
    output [5:0] col_out_364,
    output [5:0] col_out_365,
    output [5:0] col_out_366,
    output [5:0] col_out_367,
    output [5:0] col_out_368,
    output [5:0] col_out_369,
    output [5:0] col_out_370,
    output [5:0] col_out_371,
    output [5:0] col_out_372,
    output [5:0] col_out_373,
    output [5:0] col_out_374,
    output [5:0] col_out_375,
    output [5:0] col_out_376,
    output [5:0] col_out_377,
    output [5:0] col_out_378,
    output [5:0] col_out_379,
    output [5:0] col_out_380,
    output [5:0] col_out_381,
    output [5:0] col_out_382,
    output [5:0] col_out_383,
    output [5:0] col_out_384,
    output [5:0] col_out_385,
    output [5:0] col_out_386,
    output [5:0] col_out_387,
    output [5:0] col_out_388,
    output [5:0] col_out_389,
    output [5:0] col_out_390,
    output [5:0] col_out_391,
    output [5:0] col_out_392,
    output [5:0] col_out_393,
    output [5:0] col_out_394,
    output [5:0] col_out_395,
    output [5:0] col_out_396,
    output [5:0] col_out_397,
    output [5:0] col_out_398,
    output [5:0] col_out_399,
    output [5:0] col_out_400,
    output [5:0] col_out_401,
    output [5:0] col_out_402,
    output [5:0] col_out_403,
    output [5:0] col_out_404,
    output [5:0] col_out_405,
    output [5:0] col_out_406,
    output [5:0] col_out_407,
    output [5:0] col_out_408,
    output [5:0] col_out_409,
    output [5:0] col_out_410,
    output [5:0] col_out_411,
    output [5:0] col_out_412,
    output [5:0] col_out_413,
    output [5:0] col_out_414,
    output [5:0] col_out_415,
    output [5:0] col_out_416,
    output [5:0] col_out_417,
    output [5:0] col_out_418,
    output [5:0] col_out_419,
    output [5:0] col_out_420,
    output [5:0] col_out_421,
    output [5:0] col_out_422,
    output [5:0] col_out_423,
    output [5:0] col_out_424,
    output [5:0] col_out_425,
    output [5:0] col_out_426,
    output [5:0] col_out_427,
    output [5:0] col_out_428,
    output [5:0] col_out_429,
    output [5:0] col_out_430,
    output [5:0] col_out_431,
    output [5:0] col_out_432,
    output [5:0] col_out_433,
    output [5:0] col_out_434,
    output [5:0] col_out_435,
    output [5:0] col_out_436,
    output [5:0] col_out_437,
    output [5:0] col_out_438,
    output [5:0] col_out_439,
    output [5:0] col_out_440,
    output [5:0] col_out_441,
    output [5:0] col_out_442,
    output [5:0] col_out_443,
    output [5:0] col_out_444,
    output [5:0] col_out_445,
    output [5:0] col_out_446,
    output [5:0] col_out_447,
    output [5:0] col_out_448,
    output [5:0] col_out_449,
    output [5:0] col_out_450,
    output [5:0] col_out_451,
    output [5:0] col_out_452,
    output [5:0] col_out_453,
    output [5:0] col_out_454,
    output [5:0] col_out_455,
    output [5:0] col_out_456,
    output [5:0] col_out_457,
    output [5:0] col_out_458,
    output [5:0] col_out_459,
    output [5:0] col_out_460,
    output [5:0] col_out_461,
    output [5:0] col_out_462,
    output [5:0] col_out_463,
    output [5:0] col_out_464,
    output [5:0] col_out_465,
    output [5:0] col_out_466,
    output [5:0] col_out_467,
    output [5:0] col_out_468,
    output [5:0] col_out_469,
    output [5:0] col_out_470,
    output [5:0] col_out_471,
    output [5:0] col_out_472,
    output [5:0] col_out_473,
    output [5:0] col_out_474,
    output [5:0] col_out_475,
    output [5:0] col_out_476,
    output [5:0] col_out_477,
    output [5:0] col_out_478,
    output [5:0] col_out_479,
    output [5:0] col_out_480,
    output [5:0] col_out_481,
    output [5:0] col_out_482,
    output [5:0] col_out_483,
    output [5:0] col_out_484,
    output [5:0] col_out_485,
    output [5:0] col_out_486,
    output [5:0] col_out_487,
    output [5:0] col_out_488,
    output [5:0] col_out_489,
    output [5:0] col_out_490,
    output [5:0] col_out_491,
    output [5:0] col_out_492,
    output [5:0] col_out_493,
    output [5:0] col_out_494,
    output [5:0] col_out_495,
    output [5:0] col_out_496,
    output [5:0] col_out_497,
    output [5:0] col_out_498,
    output [5:0] col_out_499,
    output [5:0] col_out_500,
    output [5:0] col_out_501,
    output [5:0] col_out_502,
    output [5:0] col_out_503,
    output [5:0] col_out_504,
    output [5:0] col_out_505,
    output [5:0] col_out_506,
    output [5:0] col_out_507,
    output [5:0] col_out_508,
    output [5:0] col_out_509,
    output [5:0] col_out_510,
    output [5:0] col_out_511,
    output [5:0] col_out_512,
    output [5:0] col_out_513,
    output [5:0] col_out_514,
    output [5:0] col_out_515,
    output [5:0] col_out_516,
    output [5:0] col_out_517,
    output [5:0] col_out_518,
    output [5:0] col_out_519,
    output [5:0] col_out_520,
    output [5:0] col_out_521,
    output [5:0] col_out_522,
    output [5:0] col_out_523,
    output [5:0] col_out_524,
    output [5:0] col_out_525,
    output [5:0] col_out_526,
    output [5:0] col_out_527,
    output [5:0] col_out_528,
    output [5:0] col_out_529,
    output [5:0] col_out_530,
    output [5:0] col_out_531,
    output [5:0] col_out_532,
    output [5:0] col_out_533,
    output [5:0] col_out_534,
    output [5:0] col_out_535,
    output [5:0] col_out_536,
    output [5:0] col_out_537,
    output [5:0] col_out_538,
    output [5:0] col_out_539,
    output [5:0] col_out_540,
    output [5:0] col_out_541,
    output [5:0] col_out_542,
    output [5:0] col_out_543,
    output [5:0] col_out_544,
    output [5:0] col_out_545,
    output [5:0] col_out_546,
    output [5:0] col_out_547,
    output [5:0] col_out_548,
    output [5:0] col_out_549,
    output [5:0] col_out_550,
    output [5:0] col_out_551,
    output [5:0] col_out_552,
    output [5:0] col_out_553,
    output [5:0] col_out_554,
    output [5:0] col_out_555,
    output [5:0] col_out_556,
    output [5:0] col_out_557,
    output [5:0] col_out_558,
    output [5:0] col_out_559,
    output [5:0] col_out_560,
    output [5:0] col_out_561,
    output [5:0] col_out_562,
    output [5:0] col_out_563,
    output [5:0] col_out_564,
    output [5:0] col_out_565,
    output [5:0] col_out_566,
    output [5:0] col_out_567,
    output [5:0] col_out_568,
    output [5:0] col_out_569,
    output [5:0] col_out_570,
    output [5:0] col_out_571,
    output [5:0] col_out_572,
    output [5:0] col_out_573,
    output [5:0] col_out_574,
    output [5:0] col_out_575,
    output [5:0] col_out_576,
    output [5:0] col_out_577,
    output [5:0] col_out_578,
    output [5:0] col_out_579,
    output [5:0] col_out_580,
    output [5:0] col_out_581,
    output [5:0] col_out_582,
    output [5:0] col_out_583,
    output [5:0] col_out_584,
    output [5:0] col_out_585,
    output [5:0] col_out_586,
    output [5:0] col_out_587,
    output [5:0] col_out_588,
    output [5:0] col_out_589,
    output [5:0] col_out_590,
    output [5:0] col_out_591,
    output [5:0] col_out_592,
    output [5:0] col_out_593,
    output [5:0] col_out_594,
    output [5:0] col_out_595,
    output [5:0] col_out_596,
    output [5:0] col_out_597,
    output [5:0] col_out_598,
    output [5:0] col_out_599,
    output [5:0] col_out_600,
    output [5:0] col_out_601,
    output [5:0] col_out_602,
    output [5:0] col_out_603,
    output [5:0] col_out_604,
    output [5:0] col_out_605,
    output [5:0] col_out_606,
    output [5:0] col_out_607,
    output [5:0] col_out_608,
    output [5:0] col_out_609,
    output [5:0] col_out_610,
    output [5:0] col_out_611,
    output [5:0] col_out_612,
    output [5:0] col_out_613,
    output [5:0] col_out_614,
    output [5:0] col_out_615,
    output [5:0] col_out_616,
    output [5:0] col_out_617,
    output [5:0] col_out_618,
    output [5:0] col_out_619,
    output [5:0] col_out_620,
    output [5:0] col_out_621,
    output [5:0] col_out_622,
    output [5:0] col_out_623,
    output [5:0] col_out_624,
    output [5:0] col_out_625,
    output [5:0] col_out_626,
    output [5:0] col_out_627,
    output [5:0] col_out_628,
    output [5:0] col_out_629,
    output [5:0] col_out_630,
    output [5:0] col_out_631,
    output [5:0] col_out_632,
    output [5:0] col_out_633,
    output [5:0] col_out_634,
    output [5:0] col_out_635,
    output [5:0] col_out_636,
    output [5:0] col_out_637,
    output [5:0] col_out_638,
    output [5:0] col_out_639,
    output [5:0] col_out_640,
    output [5:0] col_out_641,
    output [5:0] col_out_642,
    output [5:0] col_out_643,
    output [5:0] col_out_644,
    output [5:0] col_out_645,
    output [5:0] col_out_646,
    output [5:0] col_out_647,
    output [5:0] col_out_648,
    output [5:0] col_out_649,
    output [5:0] col_out_650,
    output [5:0] col_out_651,
    output [5:0] col_out_652,
    output [5:0] col_out_653,
    output [5:0] col_out_654,
    output [5:0] col_out_655,
    output [5:0] col_out_656,
    output [5:0] col_out_657,
    output [5:0] col_out_658,
    output [5:0] col_out_659,
    output [5:0] col_out_660,
    output [5:0] col_out_661,
    output [5:0] col_out_662,
    output [5:0] col_out_663,
    output [5:0] col_out_664,
    output [5:0] col_out_665,
    output [5:0] col_out_666,
    output [5:0] col_out_667,
    output [5:0] col_out_668,
    output [5:0] col_out_669,
    output [5:0] col_out_670,
    output [5:0] col_out_671,
    output [5:0] col_out_672,
    output [5:0] col_out_673,
    output [5:0] col_out_674,
    output [5:0] col_out_675,
    output [5:0] col_out_676,
    output [5:0] col_out_677,
    output [5:0] col_out_678,
    output [5:0] col_out_679,
    output [5:0] col_out_680,
    output [5:0] col_out_681,
    output [5:0] col_out_682,
    output [5:0] col_out_683,
    output [5:0] col_out_684,
    output [5:0] col_out_685,
    output [5:0] col_out_686,
    output [5:0] col_out_687,
    output [5:0] col_out_688,
    output [5:0] col_out_689,
    output [5:0] col_out_690,
    output [5:0] col_out_691,
    output [5:0] col_out_692,
    output [5:0] col_out_693,
    output [5:0] col_out_694,
    output [5:0] col_out_695,
    output [5:0] col_out_696,
    output [5:0] col_out_697,
    output [5:0] col_out_698,
    output [5:0] col_out_699,
    output [5:0] col_out_700,
    output [5:0] col_out_701,
    output [5:0] col_out_702,
    output [5:0] col_out_703,
    output [5:0] col_out_704,
    output [5:0] col_out_705,
    output [5:0] col_out_706,
    output [5:0] col_out_707,
    output [5:0] col_out_708,
    output [5:0] col_out_709,
    output [5:0] col_out_710,
    output [5:0] col_out_711,
    output [5:0] col_out_712,
    output [5:0] col_out_713,
    output [5:0] col_out_714,
    output [5:0] col_out_715,
    output [5:0] col_out_716,
    output [5:0] col_out_717,
    output [5:0] col_out_718,
    output [5:0] col_out_719,
    output [5:0] col_out_720,
    output [5:0] col_out_721,
    output [5:0] col_out_722,
    output [5:0] col_out_723,
    output [5:0] col_out_724,
    output [5:0] col_out_725,
    output [5:0] col_out_726,
    output [5:0] col_out_727,
    output [5:0] col_out_728,
    output [5:0] col_out_729,
    output [5:0] col_out_730,
    output [5:0] col_out_731,
    output [5:0] col_out_732,
    output [5:0] col_out_733,
    output [5:0] col_out_734,
    output [5:0] col_out_735,
    output [5:0] col_out_736,
    output [5:0] col_out_737,
    output [5:0] col_out_738,
    output [5:0] col_out_739,
    output [5:0] col_out_740,
    output [5:0] col_out_741,
    output [5:0] col_out_742,
    output [5:0] col_out_743,
    output [5:0] col_out_744,
    output [5:0] col_out_745,
    output [5:0] col_out_746,
    output [5:0] col_out_747,
    output [5:0] col_out_748,
    output [5:0] col_out_749,
    output [5:0] col_out_750,
    output [5:0] col_out_751,
    output [5:0] col_out_752,
    output [5:0] col_out_753,
    output [5:0] col_out_754,
    output [5:0] col_out_755,
    output [5:0] col_out_756,
    output [5:0] col_out_757,
    output [5:0] col_out_758,
    output [5:0] col_out_759,
    output [5:0] col_out_760,
    output [5:0] col_out_761,
    output [5:0] col_out_762,
    output [5:0] col_out_763,
    output [5:0] col_out_764,
    output [5:0] col_out_765,
    output [5:0] col_out_766,
    output [5:0] col_out_767,
    output [5:0] col_out_768,
    output [5:0] col_out_769,
    output [5:0] col_out_770,
    output [5:0] col_out_771,
    output [5:0] col_out_772,
    output [5:0] col_out_773,
    output [5:0] col_out_774,
    output [5:0] col_out_775,
    output [5:0] col_out_776,
    output [5:0] col_out_777,
    output [5:0] col_out_778,
    output [5:0] col_out_779,
    output [5:0] col_out_780,
    output [5:0] col_out_781,
    output [5:0] col_out_782,
    output [5:0] col_out_783,
    output [5:0] col_out_784,
    output [5:0] col_out_785,
    output [5:0] col_out_786,
    output [5:0] col_out_787,
    output [5:0] col_out_788,
    output [5:0] col_out_789,
    output [5:0] col_out_790,
    output [5:0] col_out_791,
    output [5:0] col_out_792,
    output [5:0] col_out_793,
    output [5:0] col_out_794,
    output [5:0] col_out_795,
    output [5:0] col_out_796,
    output [5:0] col_out_797,
    output [5:0] col_out_798,
    output [5:0] col_out_799,
    output [5:0] col_out_800,
    output [5:0] col_out_801,
    output [5:0] col_out_802,
    output [5:0] col_out_803,
    output [5:0] col_out_804,
    output [5:0] col_out_805,
    output [5:0] col_out_806,
    output [5:0] col_out_807,
    output [5:0] col_out_808,
    output [5:0] col_out_809,
    output [5:0] col_out_810,
    output [5:0] col_out_811,
    output [5:0] col_out_812,
    output [5:0] col_out_813,
    output [5:0] col_out_814,
    output [5:0] col_out_815,
    output [5:0] col_out_816,
    output [5:0] col_out_817,
    output [5:0] col_out_818,
    output [5:0] col_out_819,
    output [5:0] col_out_820,
    output [5:0] col_out_821,
    output [5:0] col_out_822,
    output [5:0] col_out_823,
    output [5:0] col_out_824,
    output [5:0] col_out_825,
    output [5:0] col_out_826,
    output [5:0] col_out_827,
    output [5:0] col_out_828,
    output [5:0] col_out_829,
    output [5:0] col_out_830,
    output [5:0] col_out_831,
    output [5:0] col_out_832,
    output [5:0] col_out_833,
    output [5:0] col_out_834,
    output [5:0] col_out_835,
    output [5:0] col_out_836,
    output [5:0] col_out_837,
    output [5:0] col_out_838,
    output [5:0] col_out_839,
    output [5:0] col_out_840,
    output [5:0] col_out_841,
    output [5:0] col_out_842,
    output [5:0] col_out_843,
    output [5:0] col_out_844,
    output [5:0] col_out_845,
    output [5:0] col_out_846,
    output [5:0] col_out_847,
    output [5:0] col_out_848,
    output [5:0] col_out_849,
    output [5:0] col_out_850,
    output [5:0] col_out_851,
    output [5:0] col_out_852,
    output [5:0] col_out_853,
    output [5:0] col_out_854,
    output [5:0] col_out_855,
    output [5:0] col_out_856,
    output [5:0] col_out_857,
    output [5:0] col_out_858,
    output [5:0] col_out_859,
    output [5:0] col_out_860,
    output [5:0] col_out_861,
    output [5:0] col_out_862,
    output [5:0] col_out_863,
    output [5:0] col_out_864,
    output [5:0] col_out_865,
    output [5:0] col_out_866,
    output [5:0] col_out_867,
    output [5:0] col_out_868,
    output [5:0] col_out_869,
    output [5:0] col_out_870,
    output [5:0] col_out_871,
    output [5:0] col_out_872,
    output [5:0] col_out_873,
    output [5:0] col_out_874,
    output [5:0] col_out_875,
    output [5:0] col_out_876,
    output [5:0] col_out_877,
    output [5:0] col_out_878,
    output [5:0] col_out_879,
    output [5:0] col_out_880,
    output [5:0] col_out_881,
    output [5:0] col_out_882,
    output [5:0] col_out_883,
    output [5:0] col_out_884,
    output [5:0] col_out_885,
    output [5:0] col_out_886,
    output [5:0] col_out_887,
    output [5:0] col_out_888,
    output [5:0] col_out_889,
    output [5:0] col_out_890,
    output [5:0] col_out_891,
    output [5:0] col_out_892,
    output [5:0] col_out_893,
    output [5:0] col_out_894,
    output [5:0] col_out_895,
    output [5:0] col_out_896,
    output [5:0] col_out_897,
    output [5:0] col_out_898,
    output [5:0] col_out_899,
    output [5:0] col_out_900,
    output [5:0] col_out_901,
    output [5:0] col_out_902,
    output [5:0] col_out_903,
    output [5:0] col_out_904,
    output [5:0] col_out_905,
    output [5:0] col_out_906,
    output [5:0] col_out_907,
    output [5:0] col_out_908,
    output [5:0] col_out_909,
    output [5:0] col_out_910,
    output [5:0] col_out_911,
    output [5:0] col_out_912,
    output [5:0] col_out_913,
    output [5:0] col_out_914,
    output [5:0] col_out_915,
    output [5:0] col_out_916,
    output [5:0] col_out_917,
    output [5:0] col_out_918,
    output [5:0] col_out_919,
    output [5:0] col_out_920,
    output [5:0] col_out_921,
    output [5:0] col_out_922,
    output [5:0] col_out_923,
    output [5:0] col_out_924,
    output [5:0] col_out_925,
    output [5:0] col_out_926,
    output [5:0] col_out_927,
    output [5:0] col_out_928,
    output [5:0] col_out_929,
    output [5:0] col_out_930,
    output [5:0] col_out_931,
    output [5:0] col_out_932,
    output [5:0] col_out_933,
    output [5:0] col_out_934,
    output [5:0] col_out_935,
    output [5:0] col_out_936,
    output [5:0] col_out_937,
    output [5:0] col_out_938,
    output [5:0] col_out_939,
    output [5:0] col_out_940,
    output [5:0] col_out_941,
    output [5:0] col_out_942,
    output [5:0] col_out_943,
    output [5:0] col_out_944,
    output [5:0] col_out_945,
    output [5:0] col_out_946,
    output [5:0] col_out_947,
    output [5:0] col_out_948,
    output [5:0] col_out_949,
    output [5:0] col_out_950,
    output [5:0] col_out_951,
    output [5:0] col_out_952,
    output [5:0] col_out_953,
    output [5:0] col_out_954,
    output [5:0] col_out_955,
    output [5:0] col_out_956,
    output [5:0] col_out_957,
    output [5:0] col_out_958,
    output [5:0] col_out_959,
    output [5:0] col_out_960,
    output [5:0] col_out_961,
    output [5:0] col_out_962,
    output [5:0] col_out_963,
    output [5:0] col_out_964,
    output [5:0] col_out_965,
    output [5:0] col_out_966,
    output [5:0] col_out_967,
    output [5:0] col_out_968,
    output [5:0] col_out_969,
    output [5:0] col_out_970,
    output [5:0] col_out_971,
    output [5:0] col_out_972,
    output [5:0] col_out_973,
    output [5:0] col_out_974,
    output [5:0] col_out_975,
    output [5:0] col_out_976,
    output [5:0] col_out_977,
    output [5:0] col_out_978,
    output [5:0] col_out_979,
    output [5:0] col_out_980,
    output [5:0] col_out_981,
    output [5:0] col_out_982,
    output [5:0] col_out_983,
    output [5:0] col_out_984,
    output [5:0] col_out_985,
    output [5:0] col_out_986,
    output [5:0] col_out_987,
    output [5:0] col_out_988,
    output [5:0] col_out_989,
    output [5:0] col_out_990,
    output [5:0] col_out_991,
    output [5:0] col_out_992,
    output [5:0] col_out_993,
    output [5:0] col_out_994,
    output [5:0] col_out_995,
    output [5:0] col_out_996,
    output [5:0] col_out_997,
    output [5:0] col_out_998,
    output [5:0] col_out_999,
    output [5:0] col_out_1000,
    output [5:0] col_out_1001,
    output [5:0] col_out_1002,
    output [5:0] col_out_1003,
    output [5:0] col_out_1004,
    output [5:0] col_out_1005,
    output [5:0] col_out_1006,
    output [5:0] col_out_1007,
    output [5:0] col_out_1008,
    output [5:0] col_out_1009,
    output [5:0] col_out_1010,
    output [5:0] col_out_1011,
    output [5:0] col_out_1012,
    output [5:0] col_out_1013,
    output [5:0] col_out_1014,
    output [5:0] col_out_1015,
    output [5:0] col_out_1016,
    output [5:0] col_out_1017,
    output [5:0] col_out_1018,
    output [5:0] col_out_1019,
    output [5:0] col_out_1020,
    output [5:0] col_out_1021,
    output [5:0] col_out_1022,
    output [5:0] col_out_1023,
    output [5:0] col_out_1024,
    output [5:0] col_out_1025,
    output [5:0] col_out_1026,
    output [5:0] col_out_1027,
    output [5:0] col_out_1028,
    output [5:0] col_out_1029,
    output [5:0] col_out_1030,
    output [5:0] col_out_1031,
    output [5:0] col_out_1032,
    output [5:0] col_out_1033,
    output [5:0] col_out_1034,
    output [5:0] col_out_1035,
    output [5:0] col_out_1036,
    output [5:0] col_out_1037,
    output [5:0] col_out_1038,
    output [5:0] col_out_1039,
    output [5:0] col_out_1040,
    output [5:0] col_out_1041,
    output [5:0] col_out_1042,
    output [5:0] col_out_1043,
    output [5:0] col_out_1044,
    output [5:0] col_out_1045,
    output [5:0] col_out_1046,
    output [5:0] col_out_1047,
    output [5:0] col_out_1048,
    output [5:0] col_out_1049,
    output [5:0] col_out_1050,
    output [5:0] col_out_1051,
    output [5:0] col_out_1052,
    output [5:0] col_out_1053,
    output [5:0] col_out_1054,
    output [5:0] col_out_1055,
    output [5:0] col_out_1056,
    output [5:0] col_out_1057,
    output [5:0] col_out_1058,
    output [5:0] col_out_1059,
    output [5:0] col_out_1060,
    output [5:0] col_out_1061,
    output [5:0] col_out_1062,
    output [5:0] col_out_1063,
    output [5:0] col_out_1064,
    output [5:0] col_out_1065,
    output [5:0] col_out_1066,
    output [5:0] col_out_1067,
    output [5:0] col_out_1068,
    output [5:0] col_out_1069,
    output [5:0] col_out_1070,
    output [5:0] col_out_1071,
    output [5:0] col_out_1072,
    output [5:0] col_out_1073,
    output [5:0] col_out_1074,
    output [5:0] col_out_1075,
    output [5:0] col_out_1076,
    output [5:0] col_out_1077,
    output [5:0] col_out_1078,
    output [5:0] col_out_1079,
    output [5:0] col_out_1080,
    output [5:0] col_out_1081,
    output [5:0] col_out_1082,
    output [5:0] col_out_1083,
    output [5:0] col_out_1084,
    output [5:0] col_out_1085,
    output [5:0] col_out_1086,
    output [5:0] col_out_1087,
    output [5:0] col_out_1088,
    output [5:0] col_out_1089,
    output [5:0] col_out_1090,
    output [5:0] col_out_1091,
    output [5:0] col_out_1092,
    output [5:0] col_out_1093,
    output [5:0] col_out_1094,
    output [5:0] col_out_1095,
    output [5:0] col_out_1096,
    output [5:0] col_out_1097,
    output [5:0] col_out_1098,
    output [5:0] col_out_1099,
    output [5:0] col_out_1100,
    output [5:0] col_out_1101,
    output [5:0] col_out_1102,
    output [5:0] col_out_1103,
    output [5:0] col_out_1104,
    output [5:0] col_out_1105,
    output [5:0] col_out_1106,
    output [5:0] col_out_1107,
    output [5:0] col_out_1108,
    output [5:0] col_out_1109,
    output [5:0] col_out_1110,
    output [5:0] col_out_1111,
    output [5:0] col_out_1112,
    output [5:0] col_out_1113,
    output [5:0] col_out_1114,
    output [5:0] col_out_1115,
    output [5:0] col_out_1116,
    output [5:0] col_out_1117,
    output [5:0] col_out_1118,
    output [5:0] col_out_1119,
    output [5:0] col_out_1120,
    output [5:0] col_out_1121,
    output [5:0] col_out_1122,
    output [5:0] col_out_1123,
    output [5:0] col_out_1124,
    output [5:0] col_out_1125,
    output [5:0] col_out_1126,
    output [5:0] col_out_1127,
    output [5:0] col_out_1128,
    output [5:0] col_out_1129,
    output [5:0] col_out_1130,
    output [5:0] col_out_1131,
    output [5:0] col_out_1132,
    output [5:0] col_out_1133,
    output [5:0] col_out_1134,
    output [5:0] col_out_1135,
    output [5:0] col_out_1136,
    output [5:0] col_out_1137,
    output [5:0] col_out_1138,
    output [5:0] col_out_1139,
    output [5:0] col_out_1140,
    output [5:0] col_out_1141,
    output [5:0] col_out_1142,
    output [5:0] col_out_1143,
    output [5:0] col_out_1144,
    output [5:0] col_out_1145,
    output [5:0] col_out_1146,
    output [5:0] col_out_1147,
    output [5:0] col_out_1148,
    output [5:0] col_out_1149,
    output [5:0] col_out_1150,
    output [5:0] col_out_1151,
    output [5:0] col_out_1152,
    output [5:0] col_out_1153,
    output [5:0] col_out_1154,
    output [5:0] col_out_1155,
    output [5:0] col_out_1156,
    output [5:0] col_out_1157,
    output [5:0] col_out_1158,
    output [5:0] col_out_1159,
    output [5:0] col_out_1160,
    output [5:0] col_out_1161,
    output [5:0] col_out_1162,
    output [5:0] col_out_1163,
    output [5:0] col_out_1164,
    output [5:0] col_out_1165,
    output [5:0] col_out_1166,
    output [5:0] col_out_1167,
    output [5:0] col_out_1168,
    output [5:0] col_out_1169,
    output [5:0] col_out_1170,
    output [5:0] col_out_1171,
    output [5:0] col_out_1172,
    output [5:0] col_out_1173,
    output [5:0] col_out_1174,
    output [5:0] col_out_1175,
    output [5:0] col_out_1176,
    output [5:0] col_out_1177,
    output [5:0] col_out_1178,
    output [5:0] col_out_1179,
    output [5:0] col_out_1180,
    output [5:0] col_out_1181,
    output [5:0] col_out_1182,
    output [5:0] col_out_1183,
    output [5:0] col_out_1184,
    output [5:0] col_out_1185,
    output [5:0] col_out_1186,
    output [5:0] col_out_1187,
    output [5:0] col_out_1188,
    output [5:0] col_out_1189,
    output [5:0] col_out_1190,
    output [5:0] col_out_1191,
    output [5:0] col_out_1192,
    output [5:0] col_out_1193,
    output [5:0] col_out_1194,
    output [5:0] col_out_1195,
    output [5:0] col_out_1196,
    output [5:0] col_out_1197,
    output [5:0] col_out_1198,
    output [5:0] col_out_1199,
    output [5:0] col_out_1200,
    output [5:0] col_out_1201,
    output [5:0] col_out_1202,
    output [5:0] col_out_1203,
    output [5:0] col_out_1204,
    output [5:0] col_out_1205,
    output [5:0] col_out_1206,
    output [5:0] col_out_1207,
    output [5:0] col_out_1208,
    output [5:0] col_out_1209,
    output [5:0] col_out_1210,
    output [5:0] col_out_1211,
    output [5:0] col_out_1212,
    output [5:0] col_out_1213,
    output [5:0] col_out_1214,
    output [5:0] col_out_1215,
    output [5:0] col_out_1216,
    output [5:0] col_out_1217,
    output [5:0] col_out_1218,
    output [5:0] col_out_1219,
    output [5:0] col_out_1220,
    output [5:0] col_out_1221,
    output [5:0] col_out_1222,
    output [5:0] col_out_1223,
    output [5:0] col_out_1224,
    output [5:0] col_out_1225,
    output [5:0] col_out_1226,
    output [5:0] col_out_1227,
    output [5:0] col_out_1228,
    output [5:0] col_out_1229,
    output [5:0] col_out_1230,
    output [5:0] col_out_1231,
    output [5:0] col_out_1232,
    output [5:0] col_out_1233,
    output [5:0] col_out_1234,
    output [5:0] col_out_1235,
    output [5:0] col_out_1236,
    output [5:0] col_out_1237,
    output [5:0] col_out_1238,
    output [5:0] col_out_1239,
    output [5:0] col_out_1240,
    output [5:0] col_out_1241,
    output [5:0] col_out_1242,
    output [5:0] col_out_1243,
    output [5:0] col_out_1244,
    output [5:0] col_out_1245,
    output [5:0] col_out_1246,
    output [5:0] col_out_1247,
    output [5:0] col_out_1248,
    output [5:0] col_out_1249,
    output [5:0] col_out_1250,
    output [5:0] col_out_1251,
    output [5:0] col_out_1252,
    output [5:0] col_out_1253,
    output [5:0] col_out_1254,
    output [5:0] col_out_1255,
    output [5:0] col_out_1256,
    output [5:0] col_out_1257,
    output [5:0] col_out_1258,
    output [5:0] col_out_1259,
    output [5:0] col_out_1260,
    output [5:0] col_out_1261,
    output [5:0] col_out_1262,
    output [5:0] col_out_1263,
    output [5:0] col_out_1264,
    output [5:0] col_out_1265,
    output [5:0] col_out_1266,
    output [5:0] col_out_1267,
    output [5:0] col_out_1268,
    output [5:0] col_out_1269,
    output [5:0] col_out_1270,
    output [5:0] col_out_1271,
    output [5:0] col_out_1272,
    output [5:0] col_out_1273,
    output [5:0] col_out_1274,
    output [5:0] col_out_1275,
    output [5:0] col_out_1276,
    output [5:0] col_out_1277,
    output [5:0] col_out_1278,
    output [5:0] col_out_1279,
    output [5:0] col_out_1280,
    output [5:0] col_out_1281,
    output [5:0] col_out_1282,
    output [5:0] col_out_1283,
    output [5:0] col_out_1284,
    output [5:0] col_out_1285,
    output [5:0] col_out_1286,
    output [5:0] col_out_1287,
    output [5:0] col_out_1288
);



//--compressor_array input and output----------------------

wire [8:0] u_ca_in_0;
wire [8:0] u_ca_in_1;
wire [8:0] u_ca_in_2;
wire [8:0] u_ca_in_3;
wire [8:0] u_ca_in_4;
wire [8:0] u_ca_in_5;
wire [8:0] u_ca_in_6;
wire [8:0] u_ca_in_7;
wire [8:0] u_ca_in_8;
wire [8:0] u_ca_in_9;
wire [8:0] u_ca_in_10;
wire [8:0] u_ca_in_11;
wire [8:0] u_ca_in_12;
wire [8:0] u_ca_in_13;
wire [8:0] u_ca_in_14;
wire [8:0] u_ca_in_15;
wire [8:0] u_ca_in_16;
wire [8:0] u_ca_in_17;
wire [8:0] u_ca_in_18;
wire [8:0] u_ca_in_19;
wire [8:0] u_ca_in_20;
wire [8:0] u_ca_in_21;
wire [8:0] u_ca_in_22;
wire [8:0] u_ca_in_23;
wire [8:0] u_ca_in_24;
wire [8:0] u_ca_in_25;
wire [8:0] u_ca_in_26;
wire [8:0] u_ca_in_27;
wire [8:0] u_ca_in_28;
wire [8:0] u_ca_in_29;
wire [8:0] u_ca_in_30;
wire [8:0] u_ca_in_31;
wire [8:0] u_ca_in_32;
wire [8:0] u_ca_in_33;
wire [8:0] u_ca_in_34;
wire [8:0] u_ca_in_35;
wire [8:0] u_ca_in_36;
wire [8:0] u_ca_in_37;
wire [8:0] u_ca_in_38;
wire [8:0] u_ca_in_39;
wire [8:0] u_ca_in_40;
wire [8:0] u_ca_in_41;
wire [8:0] u_ca_in_42;
wire [8:0] u_ca_in_43;
wire [8:0] u_ca_in_44;
wire [8:0] u_ca_in_45;
wire [8:0] u_ca_in_46;
wire [8:0] u_ca_in_47;
wire [8:0] u_ca_in_48;
wire [8:0] u_ca_in_49;
wire [8:0] u_ca_in_50;
wire [8:0] u_ca_in_51;
wire [8:0] u_ca_in_52;
wire [8:0] u_ca_in_53;
wire [8:0] u_ca_in_54;
wire [8:0] u_ca_in_55;
wire [8:0] u_ca_in_56;
wire [8:0] u_ca_in_57;
wire [8:0] u_ca_in_58;
wire [8:0] u_ca_in_59;
wire [8:0] u_ca_in_60;
wire [8:0] u_ca_in_61;
wire [8:0] u_ca_in_62;
wire [8:0] u_ca_in_63;
wire [8:0] u_ca_in_64;
wire [8:0] u_ca_in_65;
wire [8:0] u_ca_in_66;
wire [8:0] u_ca_in_67;
wire [8:0] u_ca_in_68;
wire [8:0] u_ca_in_69;
wire [8:0] u_ca_in_70;
wire [8:0] u_ca_in_71;
wire [8:0] u_ca_in_72;
wire [8:0] u_ca_in_73;
wire [8:0] u_ca_in_74;
wire [8:0] u_ca_in_75;
wire [8:0] u_ca_in_76;
wire [8:0] u_ca_in_77;
wire [8:0] u_ca_in_78;
wire [8:0] u_ca_in_79;
wire [8:0] u_ca_in_80;
wire [8:0] u_ca_in_81;
wire [8:0] u_ca_in_82;
wire [8:0] u_ca_in_83;
wire [8:0] u_ca_in_84;
wire [8:0] u_ca_in_85;
wire [8:0] u_ca_in_86;
wire [8:0] u_ca_in_87;
wire [8:0] u_ca_in_88;
wire [8:0] u_ca_in_89;
wire [8:0] u_ca_in_90;
wire [8:0] u_ca_in_91;
wire [8:0] u_ca_in_92;
wire [8:0] u_ca_in_93;
wire [8:0] u_ca_in_94;
wire [8:0] u_ca_in_95;
wire [8:0] u_ca_in_96;
wire [8:0] u_ca_in_97;
wire [8:0] u_ca_in_98;
wire [8:0] u_ca_in_99;
wire [8:0] u_ca_in_100;
wire [8:0] u_ca_in_101;
wire [8:0] u_ca_in_102;
wire [8:0] u_ca_in_103;
wire [8:0] u_ca_in_104;
wire [8:0] u_ca_in_105;
wire [8:0] u_ca_in_106;
wire [8:0] u_ca_in_107;
wire [8:0] u_ca_in_108;
wire [8:0] u_ca_in_109;
wire [8:0] u_ca_in_110;
wire [8:0] u_ca_in_111;
wire [8:0] u_ca_in_112;
wire [8:0] u_ca_in_113;
wire [8:0] u_ca_in_114;
wire [8:0] u_ca_in_115;
wire [8:0] u_ca_in_116;
wire [8:0] u_ca_in_117;
wire [8:0] u_ca_in_118;
wire [8:0] u_ca_in_119;
wire [8:0] u_ca_in_120;
wire [8:0] u_ca_in_121;
wire [8:0] u_ca_in_122;
wire [8:0] u_ca_in_123;
wire [8:0] u_ca_in_124;
wire [8:0] u_ca_in_125;
wire [8:0] u_ca_in_126;
wire [8:0] u_ca_in_127;
wire [8:0] u_ca_in_128;
wire [8:0] u_ca_in_129;
wire [8:0] u_ca_in_130;
wire [8:0] u_ca_in_131;
wire [8:0] u_ca_in_132;
wire [8:0] u_ca_in_133;
wire [8:0] u_ca_in_134;
wire [8:0] u_ca_in_135;
wire [8:0] u_ca_in_136;
wire [8:0] u_ca_in_137;
wire [8:0] u_ca_in_138;
wire [8:0] u_ca_in_139;
wire [8:0] u_ca_in_140;
wire [8:0] u_ca_in_141;
wire [8:0] u_ca_in_142;
wire [8:0] u_ca_in_143;
wire [8:0] u_ca_in_144;
wire [8:0] u_ca_in_145;
wire [8:0] u_ca_in_146;
wire [8:0] u_ca_in_147;
wire [8:0] u_ca_in_148;
wire [8:0] u_ca_in_149;
wire [8:0] u_ca_in_150;
wire [8:0] u_ca_in_151;
wire [8:0] u_ca_in_152;
wire [8:0] u_ca_in_153;
wire [8:0] u_ca_in_154;
wire [8:0] u_ca_in_155;
wire [8:0] u_ca_in_156;
wire [8:0] u_ca_in_157;
wire [8:0] u_ca_in_158;
wire [8:0] u_ca_in_159;
wire [8:0] u_ca_in_160;
wire [8:0] u_ca_in_161;
wire [8:0] u_ca_in_162;
wire [8:0] u_ca_in_163;
wire [8:0] u_ca_in_164;
wire [8:0] u_ca_in_165;
wire [8:0] u_ca_in_166;
wire [8:0] u_ca_in_167;
wire [8:0] u_ca_in_168;
wire [8:0] u_ca_in_169;
wire [8:0] u_ca_in_170;
wire [8:0] u_ca_in_171;
wire [8:0] u_ca_in_172;
wire [8:0] u_ca_in_173;
wire [8:0] u_ca_in_174;
wire [8:0] u_ca_in_175;
wire [8:0] u_ca_in_176;
wire [8:0] u_ca_in_177;
wire [8:0] u_ca_in_178;
wire [8:0] u_ca_in_179;
wire [8:0] u_ca_in_180;
wire [8:0] u_ca_in_181;
wire [8:0] u_ca_in_182;
wire [8:0] u_ca_in_183;
wire [8:0] u_ca_in_184;
wire [8:0] u_ca_in_185;
wire [8:0] u_ca_in_186;
wire [8:0] u_ca_in_187;
wire [8:0] u_ca_in_188;
wire [8:0] u_ca_in_189;
wire [8:0] u_ca_in_190;
wire [8:0] u_ca_in_191;
wire [8:0] u_ca_in_192;
wire [8:0] u_ca_in_193;
wire [8:0] u_ca_in_194;
wire [8:0] u_ca_in_195;
wire [8:0] u_ca_in_196;
wire [8:0] u_ca_in_197;
wire [8:0] u_ca_in_198;
wire [8:0] u_ca_in_199;
wire [8:0] u_ca_in_200;
wire [8:0] u_ca_in_201;
wire [8:0] u_ca_in_202;
wire [8:0] u_ca_in_203;
wire [8:0] u_ca_in_204;
wire [8:0] u_ca_in_205;
wire [8:0] u_ca_in_206;
wire [8:0] u_ca_in_207;
wire [8:0] u_ca_in_208;
wire [8:0] u_ca_in_209;
wire [8:0] u_ca_in_210;
wire [8:0] u_ca_in_211;
wire [8:0] u_ca_in_212;
wire [8:0] u_ca_in_213;
wire [8:0] u_ca_in_214;
wire [8:0] u_ca_in_215;
wire [8:0] u_ca_in_216;
wire [8:0] u_ca_in_217;
wire [8:0] u_ca_in_218;
wire [8:0] u_ca_in_219;
wire [8:0] u_ca_in_220;
wire [8:0] u_ca_in_221;
wire [8:0] u_ca_in_222;
wire [8:0] u_ca_in_223;
wire [8:0] u_ca_in_224;
wire [8:0] u_ca_in_225;
wire [8:0] u_ca_in_226;
wire [8:0] u_ca_in_227;
wire [8:0] u_ca_in_228;
wire [8:0] u_ca_in_229;
wire [8:0] u_ca_in_230;
wire [8:0] u_ca_in_231;
wire [8:0] u_ca_in_232;
wire [8:0] u_ca_in_233;
wire [8:0] u_ca_in_234;
wire [8:0] u_ca_in_235;
wire [8:0] u_ca_in_236;
wire [8:0] u_ca_in_237;
wire [8:0] u_ca_in_238;
wire [8:0] u_ca_in_239;
wire [8:0] u_ca_in_240;
wire [8:0] u_ca_in_241;
wire [8:0] u_ca_in_242;
wire [8:0] u_ca_in_243;
wire [8:0] u_ca_in_244;
wire [8:0] u_ca_in_245;
wire [8:0] u_ca_in_246;
wire [8:0] u_ca_in_247;
wire [8:0] u_ca_in_248;
wire [8:0] u_ca_in_249;
wire [8:0] u_ca_in_250;
wire [8:0] u_ca_in_251;
wire [8:0] u_ca_in_252;
wire [8:0] u_ca_in_253;
wire [8:0] u_ca_in_254;
wire [8:0] u_ca_in_255;
wire [8:0] u_ca_in_256;
wire [8:0] u_ca_in_257;
wire [8:0] u_ca_in_258;
wire [8:0] u_ca_in_259;
wire [8:0] u_ca_in_260;
wire [8:0] u_ca_in_261;
wire [8:0] u_ca_in_262;
wire [8:0] u_ca_in_263;
wire [8:0] u_ca_in_264;
wire [8:0] u_ca_in_265;
wire [8:0] u_ca_in_266;
wire [8:0] u_ca_in_267;
wire [8:0] u_ca_in_268;
wire [8:0] u_ca_in_269;
wire [8:0] u_ca_in_270;
wire [8:0] u_ca_in_271;
wire [8:0] u_ca_in_272;
wire [8:0] u_ca_in_273;
wire [8:0] u_ca_in_274;
wire [8:0] u_ca_in_275;
wire [8:0] u_ca_in_276;
wire [8:0] u_ca_in_277;
wire [8:0] u_ca_in_278;
wire [8:0] u_ca_in_279;
wire [8:0] u_ca_in_280;
wire [8:0] u_ca_in_281;
wire [8:0] u_ca_in_282;
wire [8:0] u_ca_in_283;
wire [8:0] u_ca_in_284;
wire [8:0] u_ca_in_285;
wire [8:0] u_ca_in_286;
wire [8:0] u_ca_in_287;
wire [8:0] u_ca_in_288;
wire [8:0] u_ca_in_289;
wire [8:0] u_ca_in_290;
wire [8:0] u_ca_in_291;
wire [8:0] u_ca_in_292;
wire [8:0] u_ca_in_293;
wire [8:0] u_ca_in_294;
wire [8:0] u_ca_in_295;
wire [8:0] u_ca_in_296;
wire [8:0] u_ca_in_297;
wire [8:0] u_ca_in_298;
wire [8:0] u_ca_in_299;
wire [8:0] u_ca_in_300;
wire [8:0] u_ca_in_301;
wire [8:0] u_ca_in_302;
wire [8:0] u_ca_in_303;
wire [8:0] u_ca_in_304;
wire [8:0] u_ca_in_305;
wire [8:0] u_ca_in_306;
wire [8:0] u_ca_in_307;
wire [8:0] u_ca_in_308;
wire [8:0] u_ca_in_309;
wire [8:0] u_ca_in_310;
wire [8:0] u_ca_in_311;
wire [8:0] u_ca_in_312;
wire [8:0] u_ca_in_313;
wire [8:0] u_ca_in_314;
wire [8:0] u_ca_in_315;
wire [8:0] u_ca_in_316;
wire [8:0] u_ca_in_317;
wire [8:0] u_ca_in_318;
wire [8:0] u_ca_in_319;
wire [8:0] u_ca_in_320;
wire [8:0] u_ca_in_321;
wire [8:0] u_ca_in_322;
wire [8:0] u_ca_in_323;
wire [8:0] u_ca_in_324;
wire [8:0] u_ca_in_325;
wire [8:0] u_ca_in_326;
wire [8:0] u_ca_in_327;
wire [8:0] u_ca_in_328;
wire [8:0] u_ca_in_329;
wire [8:0] u_ca_in_330;
wire [8:0] u_ca_in_331;
wire [8:0] u_ca_in_332;
wire [8:0] u_ca_in_333;
wire [8:0] u_ca_in_334;
wire [8:0] u_ca_in_335;
wire [8:0] u_ca_in_336;
wire [8:0] u_ca_in_337;
wire [8:0] u_ca_in_338;
wire [8:0] u_ca_in_339;
wire [8:0] u_ca_in_340;
wire [8:0] u_ca_in_341;
wire [8:0] u_ca_in_342;
wire [8:0] u_ca_in_343;
wire [8:0] u_ca_in_344;
wire [8:0] u_ca_in_345;
wire [8:0] u_ca_in_346;
wire [8:0] u_ca_in_347;
wire [8:0] u_ca_in_348;
wire [8:0] u_ca_in_349;
wire [8:0] u_ca_in_350;
wire [8:0] u_ca_in_351;
wire [8:0] u_ca_in_352;
wire [8:0] u_ca_in_353;
wire [8:0] u_ca_in_354;
wire [8:0] u_ca_in_355;
wire [8:0] u_ca_in_356;
wire [8:0] u_ca_in_357;
wire [8:0] u_ca_in_358;
wire [8:0] u_ca_in_359;
wire [8:0] u_ca_in_360;
wire [8:0] u_ca_in_361;
wire [8:0] u_ca_in_362;
wire [8:0] u_ca_in_363;
wire [8:0] u_ca_in_364;
wire [8:0] u_ca_in_365;
wire [8:0] u_ca_in_366;
wire [8:0] u_ca_in_367;
wire [8:0] u_ca_in_368;
wire [8:0] u_ca_in_369;
wire [8:0] u_ca_in_370;
wire [8:0] u_ca_in_371;
wire [8:0] u_ca_in_372;
wire [8:0] u_ca_in_373;
wire [8:0] u_ca_in_374;
wire [8:0] u_ca_in_375;
wire [8:0] u_ca_in_376;
wire [8:0] u_ca_in_377;
wire [8:0] u_ca_in_378;
wire [8:0] u_ca_in_379;
wire [8:0] u_ca_in_380;
wire [8:0] u_ca_in_381;
wire [8:0] u_ca_in_382;
wire [8:0] u_ca_in_383;
wire [8:0] u_ca_in_384;
wire [8:0] u_ca_in_385;
wire [8:0] u_ca_in_386;
wire [8:0] u_ca_in_387;
wire [8:0] u_ca_in_388;
wire [8:0] u_ca_in_389;
wire [8:0] u_ca_in_390;
wire [8:0] u_ca_in_391;
wire [8:0] u_ca_in_392;
wire [8:0] u_ca_in_393;
wire [8:0] u_ca_in_394;
wire [8:0] u_ca_in_395;
wire [8:0] u_ca_in_396;
wire [8:0] u_ca_in_397;
wire [8:0] u_ca_in_398;
wire [8:0] u_ca_in_399;
wire [8:0] u_ca_in_400;
wire [8:0] u_ca_in_401;
wire [8:0] u_ca_in_402;
wire [8:0] u_ca_in_403;
wire [8:0] u_ca_in_404;
wire [8:0] u_ca_in_405;
wire [8:0] u_ca_in_406;
wire [8:0] u_ca_in_407;
wire [8:0] u_ca_in_408;
wire [8:0] u_ca_in_409;
wire [8:0] u_ca_in_410;
wire [8:0] u_ca_in_411;
wire [8:0] u_ca_in_412;
wire [8:0] u_ca_in_413;
wire [8:0] u_ca_in_414;
wire [8:0] u_ca_in_415;
wire [8:0] u_ca_in_416;
wire [8:0] u_ca_in_417;
wire [8:0] u_ca_in_418;
wire [8:0] u_ca_in_419;
wire [8:0] u_ca_in_420;
wire [8:0] u_ca_in_421;
wire [8:0] u_ca_in_422;
wire [8:0] u_ca_in_423;
wire [8:0] u_ca_in_424;
wire [8:0] u_ca_in_425;
wire [8:0] u_ca_in_426;
wire [8:0] u_ca_in_427;
wire [8:0] u_ca_in_428;
wire [8:0] u_ca_in_429;
wire [8:0] u_ca_in_430;
wire [8:0] u_ca_in_431;
wire [8:0] u_ca_in_432;
wire [8:0] u_ca_in_433;
wire [8:0] u_ca_in_434;
wire [8:0] u_ca_in_435;
wire [8:0] u_ca_in_436;
wire [8:0] u_ca_in_437;
wire [8:0] u_ca_in_438;
wire [8:0] u_ca_in_439;
wire [8:0] u_ca_in_440;
wire [8:0] u_ca_in_441;
wire [8:0] u_ca_in_442;
wire [8:0] u_ca_in_443;
wire [8:0] u_ca_in_444;
wire [8:0] u_ca_in_445;
wire [8:0] u_ca_in_446;
wire [8:0] u_ca_in_447;
wire [8:0] u_ca_in_448;
wire [8:0] u_ca_in_449;
wire [8:0] u_ca_in_450;
wire [8:0] u_ca_in_451;
wire [8:0] u_ca_in_452;
wire [8:0] u_ca_in_453;
wire [8:0] u_ca_in_454;
wire [8:0] u_ca_in_455;
wire [8:0] u_ca_in_456;
wire [8:0] u_ca_in_457;
wire [8:0] u_ca_in_458;
wire [8:0] u_ca_in_459;
wire [8:0] u_ca_in_460;
wire [8:0] u_ca_in_461;
wire [8:0] u_ca_in_462;
wire [8:0] u_ca_in_463;
wire [8:0] u_ca_in_464;
wire [8:0] u_ca_in_465;
wire [8:0] u_ca_in_466;
wire [8:0] u_ca_in_467;
wire [8:0] u_ca_in_468;
wire [8:0] u_ca_in_469;
wire [8:0] u_ca_in_470;
wire [8:0] u_ca_in_471;
wire [8:0] u_ca_in_472;
wire [8:0] u_ca_in_473;
wire [8:0] u_ca_in_474;
wire [8:0] u_ca_in_475;
wire [8:0] u_ca_in_476;
wire [8:0] u_ca_in_477;
wire [8:0] u_ca_in_478;
wire [8:0] u_ca_in_479;
wire [8:0] u_ca_in_480;
wire [8:0] u_ca_in_481;
wire [8:0] u_ca_in_482;
wire [8:0] u_ca_in_483;
wire [8:0] u_ca_in_484;
wire [8:0] u_ca_in_485;
wire [8:0] u_ca_in_486;
wire [8:0] u_ca_in_487;
wire [8:0] u_ca_in_488;
wire [8:0] u_ca_in_489;
wire [8:0] u_ca_in_490;
wire [8:0] u_ca_in_491;
wire [8:0] u_ca_in_492;
wire [8:0] u_ca_in_493;
wire [8:0] u_ca_in_494;
wire [8:0] u_ca_in_495;
wire [8:0] u_ca_in_496;
wire [8:0] u_ca_in_497;
wire [8:0] u_ca_in_498;
wire [8:0] u_ca_in_499;
wire [8:0] u_ca_in_500;
wire [8:0] u_ca_in_501;
wire [8:0] u_ca_in_502;
wire [8:0] u_ca_in_503;
wire [8:0] u_ca_in_504;
wire [8:0] u_ca_in_505;
wire [8:0] u_ca_in_506;
wire [8:0] u_ca_in_507;
wire [8:0] u_ca_in_508;
wire [8:0] u_ca_in_509;
wire [8:0] u_ca_in_510;
wire [8:0] u_ca_in_511;
wire [8:0] u_ca_in_512;
wire [8:0] u_ca_in_513;
wire [8:0] u_ca_in_514;
wire [8:0] u_ca_in_515;
wire [8:0] u_ca_in_516;
wire [8:0] u_ca_in_517;
wire [8:0] u_ca_in_518;
wire [8:0] u_ca_in_519;
wire [8:0] u_ca_in_520;
wire [8:0] u_ca_in_521;
wire [8:0] u_ca_in_522;
wire [8:0] u_ca_in_523;
wire [8:0] u_ca_in_524;
wire [8:0] u_ca_in_525;
wire [8:0] u_ca_in_526;
wire [8:0] u_ca_in_527;
wire [8:0] u_ca_in_528;
wire [8:0] u_ca_in_529;
wire [8:0] u_ca_in_530;
wire [8:0] u_ca_in_531;
wire [8:0] u_ca_in_532;
wire [8:0] u_ca_in_533;
wire [8:0] u_ca_in_534;
wire [8:0] u_ca_in_535;
wire [8:0] u_ca_in_536;
wire [8:0] u_ca_in_537;
wire [8:0] u_ca_in_538;
wire [8:0] u_ca_in_539;
wire [8:0] u_ca_in_540;
wire [8:0] u_ca_in_541;
wire [8:0] u_ca_in_542;
wire [8:0] u_ca_in_543;
wire [8:0] u_ca_in_544;
wire [8:0] u_ca_in_545;
wire [8:0] u_ca_in_546;
wire [8:0] u_ca_in_547;
wire [8:0] u_ca_in_548;
wire [8:0] u_ca_in_549;
wire [8:0] u_ca_in_550;
wire [8:0] u_ca_in_551;
wire [8:0] u_ca_in_552;
wire [8:0] u_ca_in_553;
wire [8:0] u_ca_in_554;
wire [8:0] u_ca_in_555;
wire [8:0] u_ca_in_556;
wire [8:0] u_ca_in_557;
wire [8:0] u_ca_in_558;
wire [8:0] u_ca_in_559;
wire [8:0] u_ca_in_560;
wire [8:0] u_ca_in_561;
wire [8:0] u_ca_in_562;
wire [8:0] u_ca_in_563;
wire [8:0] u_ca_in_564;
wire [8:0] u_ca_in_565;
wire [8:0] u_ca_in_566;
wire [8:0] u_ca_in_567;
wire [8:0] u_ca_in_568;
wire [8:0] u_ca_in_569;
wire [8:0] u_ca_in_570;
wire [8:0] u_ca_in_571;
wire [8:0] u_ca_in_572;
wire [8:0] u_ca_in_573;
wire [8:0] u_ca_in_574;
wire [8:0] u_ca_in_575;
wire [8:0] u_ca_in_576;
wire [8:0] u_ca_in_577;
wire [8:0] u_ca_in_578;
wire [8:0] u_ca_in_579;
wire [8:0] u_ca_in_580;
wire [8:0] u_ca_in_581;
wire [8:0] u_ca_in_582;
wire [8:0] u_ca_in_583;
wire [8:0] u_ca_in_584;
wire [8:0] u_ca_in_585;
wire [8:0] u_ca_in_586;
wire [8:0] u_ca_in_587;
wire [8:0] u_ca_in_588;
wire [8:0] u_ca_in_589;
wire [8:0] u_ca_in_590;
wire [8:0] u_ca_in_591;
wire [8:0] u_ca_in_592;
wire [8:0] u_ca_in_593;
wire [8:0] u_ca_in_594;
wire [8:0] u_ca_in_595;
wire [8:0] u_ca_in_596;
wire [8:0] u_ca_in_597;
wire [8:0] u_ca_in_598;
wire [8:0] u_ca_in_599;
wire [8:0] u_ca_in_600;
wire [8:0] u_ca_in_601;
wire [8:0] u_ca_in_602;
wire [8:0] u_ca_in_603;
wire [8:0] u_ca_in_604;
wire [8:0] u_ca_in_605;
wire [8:0] u_ca_in_606;
wire [8:0] u_ca_in_607;
wire [8:0] u_ca_in_608;
wire [8:0] u_ca_in_609;
wire [8:0] u_ca_in_610;
wire [8:0] u_ca_in_611;
wire [8:0] u_ca_in_612;
wire [8:0] u_ca_in_613;
wire [8:0] u_ca_in_614;
wire [8:0] u_ca_in_615;
wire [8:0] u_ca_in_616;
wire [8:0] u_ca_in_617;
wire [8:0] u_ca_in_618;
wire [8:0] u_ca_in_619;
wire [8:0] u_ca_in_620;
wire [8:0] u_ca_in_621;
wire [8:0] u_ca_in_622;
wire [8:0] u_ca_in_623;
wire [8:0] u_ca_in_624;
wire [8:0] u_ca_in_625;
wire [8:0] u_ca_in_626;
wire [8:0] u_ca_in_627;
wire [8:0] u_ca_in_628;
wire [8:0] u_ca_in_629;
wire [8:0] u_ca_in_630;
wire [8:0] u_ca_in_631;
wire [8:0] u_ca_in_632;
wire [8:0] u_ca_in_633;
wire [8:0] u_ca_in_634;
wire [8:0] u_ca_in_635;
wire [8:0] u_ca_in_636;
wire [8:0] u_ca_in_637;
wire [8:0] u_ca_in_638;
wire [8:0] u_ca_in_639;
wire [8:0] u_ca_in_640;
wire [8:0] u_ca_in_641;
wire [8:0] u_ca_in_642;
wire [8:0] u_ca_in_643;
wire [8:0] u_ca_in_644;
wire [8:0] u_ca_in_645;
wire [8:0] u_ca_in_646;
wire [8:0] u_ca_in_647;
wire [8:0] u_ca_in_648;
wire [8:0] u_ca_in_649;
wire [8:0] u_ca_in_650;
wire [8:0] u_ca_in_651;
wire [8:0] u_ca_in_652;
wire [8:0] u_ca_in_653;
wire [8:0] u_ca_in_654;
wire [8:0] u_ca_in_655;
wire [8:0] u_ca_in_656;
wire [8:0] u_ca_in_657;
wire [8:0] u_ca_in_658;
wire [8:0] u_ca_in_659;
wire [8:0] u_ca_in_660;
wire [8:0] u_ca_in_661;
wire [8:0] u_ca_in_662;
wire [8:0] u_ca_in_663;
wire [8:0] u_ca_in_664;
wire [8:0] u_ca_in_665;
wire [8:0] u_ca_in_666;
wire [8:0] u_ca_in_667;
wire [8:0] u_ca_in_668;
wire [8:0] u_ca_in_669;
wire [8:0] u_ca_in_670;
wire [8:0] u_ca_in_671;
wire [8:0] u_ca_in_672;
wire [8:0] u_ca_in_673;
wire [8:0] u_ca_in_674;
wire [8:0] u_ca_in_675;
wire [8:0] u_ca_in_676;
wire [8:0] u_ca_in_677;
wire [8:0] u_ca_in_678;
wire [8:0] u_ca_in_679;
wire [8:0] u_ca_in_680;
wire [8:0] u_ca_in_681;
wire [8:0] u_ca_in_682;
wire [8:0] u_ca_in_683;
wire [8:0] u_ca_in_684;
wire [8:0] u_ca_in_685;
wire [8:0] u_ca_in_686;
wire [8:0] u_ca_in_687;
wire [8:0] u_ca_in_688;
wire [8:0] u_ca_in_689;
wire [8:0] u_ca_in_690;
wire [8:0] u_ca_in_691;
wire [8:0] u_ca_in_692;
wire [8:0] u_ca_in_693;
wire [8:0] u_ca_in_694;
wire [8:0] u_ca_in_695;
wire [8:0] u_ca_in_696;
wire [8:0] u_ca_in_697;
wire [8:0] u_ca_in_698;
wire [8:0] u_ca_in_699;
wire [8:0] u_ca_in_700;
wire [8:0] u_ca_in_701;
wire [8:0] u_ca_in_702;
wire [8:0] u_ca_in_703;
wire [8:0] u_ca_in_704;
wire [8:0] u_ca_in_705;
wire [8:0] u_ca_in_706;
wire [8:0] u_ca_in_707;
wire [8:0] u_ca_in_708;
wire [8:0] u_ca_in_709;
wire [8:0] u_ca_in_710;
wire [8:0] u_ca_in_711;
wire [8:0] u_ca_in_712;
wire [8:0] u_ca_in_713;
wire [8:0] u_ca_in_714;
wire [8:0] u_ca_in_715;
wire [8:0] u_ca_in_716;
wire [8:0] u_ca_in_717;
wire [8:0] u_ca_in_718;
wire [8:0] u_ca_in_719;
wire [8:0] u_ca_in_720;
wire [8:0] u_ca_in_721;
wire [8:0] u_ca_in_722;
wire [8:0] u_ca_in_723;
wire [8:0] u_ca_in_724;
wire [8:0] u_ca_in_725;
wire [8:0] u_ca_in_726;
wire [8:0] u_ca_in_727;
wire [8:0] u_ca_in_728;
wire [8:0] u_ca_in_729;
wire [8:0] u_ca_in_730;
wire [8:0] u_ca_in_731;
wire [8:0] u_ca_in_732;
wire [8:0] u_ca_in_733;
wire [8:0] u_ca_in_734;
wire [8:0] u_ca_in_735;
wire [8:0] u_ca_in_736;
wire [8:0] u_ca_in_737;
wire [8:0] u_ca_in_738;
wire [8:0] u_ca_in_739;
wire [8:0] u_ca_in_740;
wire [8:0] u_ca_in_741;
wire [8:0] u_ca_in_742;
wire [8:0] u_ca_in_743;
wire [8:0] u_ca_in_744;
wire [8:0] u_ca_in_745;
wire [8:0] u_ca_in_746;
wire [8:0] u_ca_in_747;
wire [8:0] u_ca_in_748;
wire [8:0] u_ca_in_749;
wire [8:0] u_ca_in_750;
wire [8:0] u_ca_in_751;
wire [8:0] u_ca_in_752;
wire [8:0] u_ca_in_753;
wire [8:0] u_ca_in_754;
wire [8:0] u_ca_in_755;
wire [8:0] u_ca_in_756;
wire [8:0] u_ca_in_757;
wire [8:0] u_ca_in_758;
wire [8:0] u_ca_in_759;
wire [8:0] u_ca_in_760;
wire [8:0] u_ca_in_761;
wire [8:0] u_ca_in_762;
wire [8:0] u_ca_in_763;
wire [8:0] u_ca_in_764;
wire [8:0] u_ca_in_765;
wire [8:0] u_ca_in_766;
wire [8:0] u_ca_in_767;
wire [8:0] u_ca_in_768;
wire [8:0] u_ca_in_769;
wire [8:0] u_ca_in_770;
wire [8:0] u_ca_in_771;
wire [8:0] u_ca_in_772;
wire [8:0] u_ca_in_773;
wire [8:0] u_ca_in_774;
wire [8:0] u_ca_in_775;
wire [8:0] u_ca_in_776;
wire [8:0] u_ca_in_777;
wire [8:0] u_ca_in_778;
wire [8:0] u_ca_in_779;
wire [8:0] u_ca_in_780;
wire [8:0] u_ca_in_781;
wire [8:0] u_ca_in_782;
wire [8:0] u_ca_in_783;
wire [8:0] u_ca_in_784;
wire [8:0] u_ca_in_785;
wire [8:0] u_ca_in_786;
wire [8:0] u_ca_in_787;
wire [8:0] u_ca_in_788;
wire [8:0] u_ca_in_789;
wire [8:0] u_ca_in_790;
wire [8:0] u_ca_in_791;
wire [8:0] u_ca_in_792;
wire [8:0] u_ca_in_793;
wire [8:0] u_ca_in_794;
wire [8:0] u_ca_in_795;
wire [8:0] u_ca_in_796;
wire [8:0] u_ca_in_797;
wire [8:0] u_ca_in_798;
wire [8:0] u_ca_in_799;
wire [8:0] u_ca_in_800;
wire [8:0] u_ca_in_801;
wire [8:0] u_ca_in_802;
wire [8:0] u_ca_in_803;
wire [8:0] u_ca_in_804;
wire [8:0] u_ca_in_805;
wire [8:0] u_ca_in_806;
wire [8:0] u_ca_in_807;
wire [8:0] u_ca_in_808;
wire [8:0] u_ca_in_809;
wire [8:0] u_ca_in_810;
wire [8:0] u_ca_in_811;
wire [8:0] u_ca_in_812;
wire [8:0] u_ca_in_813;
wire [8:0] u_ca_in_814;
wire [8:0] u_ca_in_815;
wire [8:0] u_ca_in_816;
wire [8:0] u_ca_in_817;
wire [8:0] u_ca_in_818;
wire [8:0] u_ca_in_819;
wire [8:0] u_ca_in_820;
wire [8:0] u_ca_in_821;
wire [8:0] u_ca_in_822;
wire [8:0] u_ca_in_823;
wire [8:0] u_ca_in_824;
wire [8:0] u_ca_in_825;
wire [8:0] u_ca_in_826;
wire [8:0] u_ca_in_827;
wire [8:0] u_ca_in_828;
wire [8:0] u_ca_in_829;
wire [8:0] u_ca_in_830;
wire [8:0] u_ca_in_831;
wire [8:0] u_ca_in_832;
wire [8:0] u_ca_in_833;
wire [8:0] u_ca_in_834;
wire [8:0] u_ca_in_835;
wire [8:0] u_ca_in_836;
wire [8:0] u_ca_in_837;
wire [8:0] u_ca_in_838;
wire [8:0] u_ca_in_839;
wire [8:0] u_ca_in_840;
wire [8:0] u_ca_in_841;
wire [8:0] u_ca_in_842;
wire [8:0] u_ca_in_843;
wire [8:0] u_ca_in_844;
wire [8:0] u_ca_in_845;
wire [8:0] u_ca_in_846;
wire [8:0] u_ca_in_847;
wire [8:0] u_ca_in_848;
wire [8:0] u_ca_in_849;
wire [8:0] u_ca_in_850;
wire [8:0] u_ca_in_851;
wire [8:0] u_ca_in_852;
wire [8:0] u_ca_in_853;
wire [8:0] u_ca_in_854;
wire [8:0] u_ca_in_855;
wire [8:0] u_ca_in_856;
wire [8:0] u_ca_in_857;
wire [8:0] u_ca_in_858;
wire [8:0] u_ca_in_859;
wire [8:0] u_ca_in_860;
wire [8:0] u_ca_in_861;
wire [8:0] u_ca_in_862;
wire [8:0] u_ca_in_863;
wire [8:0] u_ca_in_864;
wire [8:0] u_ca_in_865;
wire [8:0] u_ca_in_866;
wire [8:0] u_ca_in_867;
wire [8:0] u_ca_in_868;
wire [8:0] u_ca_in_869;
wire [8:0] u_ca_in_870;
wire [8:0] u_ca_in_871;
wire [8:0] u_ca_in_872;
wire [8:0] u_ca_in_873;
wire [8:0] u_ca_in_874;
wire [8:0] u_ca_in_875;
wire [8:0] u_ca_in_876;
wire [8:0] u_ca_in_877;
wire [8:0] u_ca_in_878;
wire [8:0] u_ca_in_879;
wire [8:0] u_ca_in_880;
wire [8:0] u_ca_in_881;
wire [8:0] u_ca_in_882;
wire [8:0] u_ca_in_883;
wire [8:0] u_ca_in_884;
wire [8:0] u_ca_in_885;
wire [8:0] u_ca_in_886;
wire [8:0] u_ca_in_887;
wire [8:0] u_ca_in_888;
wire [8:0] u_ca_in_889;
wire [8:0] u_ca_in_890;
wire [8:0] u_ca_in_891;
wire [8:0] u_ca_in_892;
wire [8:0] u_ca_in_893;
wire [8:0] u_ca_in_894;
wire [8:0] u_ca_in_895;
wire [8:0] u_ca_in_896;
wire [8:0] u_ca_in_897;
wire [8:0] u_ca_in_898;
wire [8:0] u_ca_in_899;
wire [8:0] u_ca_in_900;
wire [8:0] u_ca_in_901;
wire [8:0] u_ca_in_902;
wire [8:0] u_ca_in_903;
wire [8:0] u_ca_in_904;
wire [8:0] u_ca_in_905;
wire [8:0] u_ca_in_906;
wire [8:0] u_ca_in_907;
wire [8:0] u_ca_in_908;
wire [8:0] u_ca_in_909;
wire [8:0] u_ca_in_910;
wire [8:0] u_ca_in_911;
wire [8:0] u_ca_in_912;
wire [8:0] u_ca_in_913;
wire [8:0] u_ca_in_914;
wire [8:0] u_ca_in_915;
wire [8:0] u_ca_in_916;
wire [8:0] u_ca_in_917;
wire [8:0] u_ca_in_918;
wire [8:0] u_ca_in_919;
wire [8:0] u_ca_in_920;
wire [8:0] u_ca_in_921;
wire [8:0] u_ca_in_922;
wire [8:0] u_ca_in_923;
wire [8:0] u_ca_in_924;
wire [8:0] u_ca_in_925;
wire [8:0] u_ca_in_926;
wire [8:0] u_ca_in_927;
wire [8:0] u_ca_in_928;
wire [8:0] u_ca_in_929;
wire [8:0] u_ca_in_930;
wire [8:0] u_ca_in_931;
wire [8:0] u_ca_in_932;
wire [8:0] u_ca_in_933;
wire [8:0] u_ca_in_934;
wire [8:0] u_ca_in_935;
wire [8:0] u_ca_in_936;
wire [8:0] u_ca_in_937;
wire [8:0] u_ca_in_938;
wire [8:0] u_ca_in_939;
wire [8:0] u_ca_in_940;
wire [8:0] u_ca_in_941;
wire [8:0] u_ca_in_942;
wire [8:0] u_ca_in_943;
wire [8:0] u_ca_in_944;
wire [8:0] u_ca_in_945;
wire [8:0] u_ca_in_946;
wire [8:0] u_ca_in_947;
wire [8:0] u_ca_in_948;
wire [8:0] u_ca_in_949;
wire [8:0] u_ca_in_950;
wire [8:0] u_ca_in_951;
wire [8:0] u_ca_in_952;
wire [8:0] u_ca_in_953;
wire [8:0] u_ca_in_954;
wire [8:0] u_ca_in_955;
wire [8:0] u_ca_in_956;
wire [8:0] u_ca_in_957;
wire [8:0] u_ca_in_958;
wire [8:0] u_ca_in_959;
wire [8:0] u_ca_in_960;
wire [8:0] u_ca_in_961;
wire [8:0] u_ca_in_962;
wire [8:0] u_ca_in_963;
wire [8:0] u_ca_in_964;
wire [8:0] u_ca_in_965;
wire [8:0] u_ca_in_966;
wire [8:0] u_ca_in_967;
wire [8:0] u_ca_in_968;
wire [8:0] u_ca_in_969;
wire [8:0] u_ca_in_970;
wire [8:0] u_ca_in_971;
wire [8:0] u_ca_in_972;
wire [8:0] u_ca_in_973;
wire [8:0] u_ca_in_974;
wire [8:0] u_ca_in_975;
wire [8:0] u_ca_in_976;
wire [8:0] u_ca_in_977;
wire [8:0] u_ca_in_978;
wire [8:0] u_ca_in_979;
wire [8:0] u_ca_in_980;
wire [8:0] u_ca_in_981;
wire [8:0] u_ca_in_982;
wire [8:0] u_ca_in_983;
wire [8:0] u_ca_in_984;
wire [8:0] u_ca_in_985;
wire [8:0] u_ca_in_986;
wire [8:0] u_ca_in_987;
wire [8:0] u_ca_in_988;
wire [8:0] u_ca_in_989;
wire [8:0] u_ca_in_990;
wire [8:0] u_ca_in_991;
wire [8:0] u_ca_in_992;
wire [8:0] u_ca_in_993;
wire [8:0] u_ca_in_994;
wire [8:0] u_ca_in_995;
wire [8:0] u_ca_in_996;
wire [8:0] u_ca_in_997;
wire [8:0] u_ca_in_998;
wire [8:0] u_ca_in_999;
wire [8:0] u_ca_in_1000;
wire [8:0] u_ca_in_1001;
wire [8:0] u_ca_in_1002;
wire [8:0] u_ca_in_1003;
wire [8:0] u_ca_in_1004;
wire [8:0] u_ca_in_1005;
wire [8:0] u_ca_in_1006;
wire [8:0] u_ca_in_1007;
wire [8:0] u_ca_in_1008;
wire [8:0] u_ca_in_1009;
wire [8:0] u_ca_in_1010;
wire [8:0] u_ca_in_1011;
wire [8:0] u_ca_in_1012;
wire [8:0] u_ca_in_1013;
wire [8:0] u_ca_in_1014;
wire [8:0] u_ca_in_1015;
wire [8:0] u_ca_in_1016;
wire [8:0] u_ca_in_1017;
wire [8:0] u_ca_in_1018;
wire [8:0] u_ca_in_1019;
wire [8:0] u_ca_in_1020;
wire [8:0] u_ca_in_1021;
wire [8:0] u_ca_in_1022;
wire [8:0] u_ca_in_1023;
wire [8:0] u_ca_in_1024;
wire [8:0] u_ca_in_1025;
wire [8:0] u_ca_in_1026;
wire [8:0] u_ca_in_1027;
wire [8:0] u_ca_in_1028;
wire [8:0] u_ca_in_1029;
wire [8:0] u_ca_in_1030;
wire [8:0] u_ca_in_1031;
wire [8:0] u_ca_in_1032;
wire [8:0] u_ca_in_1033;
wire [8:0] u_ca_in_1034;
wire [8:0] u_ca_in_1035;
wire [8:0] u_ca_in_1036;
wire [8:0] u_ca_in_1037;
wire [8:0] u_ca_in_1038;
wire [8:0] u_ca_in_1039;
wire [8:0] u_ca_in_1040;
wire [8:0] u_ca_in_1041;
wire [8:0] u_ca_in_1042;
wire [8:0] u_ca_in_1043;
wire [8:0] u_ca_in_1044;
wire [8:0] u_ca_in_1045;
wire [8:0] u_ca_in_1046;
wire [8:0] u_ca_in_1047;
wire [8:0] u_ca_in_1048;
wire [8:0] u_ca_in_1049;
wire [8:0] u_ca_in_1050;
wire [8:0] u_ca_in_1051;
wire [8:0] u_ca_in_1052;
wire [8:0] u_ca_in_1053;
wire [8:0] u_ca_in_1054;
wire [8:0] u_ca_in_1055;
wire [8:0] u_ca_in_1056;
wire [8:0] u_ca_in_1057;
wire [8:0] u_ca_in_1058;
wire [8:0] u_ca_in_1059;
wire [8:0] u_ca_in_1060;
wire [8:0] u_ca_in_1061;
wire [8:0] u_ca_in_1062;
wire [8:0] u_ca_in_1063;
wire [8:0] u_ca_in_1064;
wire [8:0] u_ca_in_1065;
wire [8:0] u_ca_in_1066;
wire [8:0] u_ca_in_1067;
wire [8:0] u_ca_in_1068;
wire [8:0] u_ca_in_1069;
wire [8:0] u_ca_in_1070;
wire [8:0] u_ca_in_1071;
wire [8:0] u_ca_in_1072;
wire [8:0] u_ca_in_1073;
wire [8:0] u_ca_in_1074;
wire [8:0] u_ca_in_1075;
wire [8:0] u_ca_in_1076;
wire [8:0] u_ca_in_1077;
wire [8:0] u_ca_in_1078;
wire [8:0] u_ca_in_1079;
wire [8:0] u_ca_in_1080;
wire [8:0] u_ca_in_1081;
wire [8:0] u_ca_in_1082;
wire [8:0] u_ca_in_1083;
wire [8:0] u_ca_in_1084;
wire [8:0] u_ca_in_1085;
wire [8:0] u_ca_in_1086;
wire [8:0] u_ca_in_1087;
wire [8:0] u_ca_in_1088;
wire [8:0] u_ca_in_1089;
wire [8:0] u_ca_in_1090;
wire [8:0] u_ca_in_1091;
wire [8:0] u_ca_in_1092;
wire [8:0] u_ca_in_1093;
wire [8:0] u_ca_in_1094;
wire [8:0] u_ca_in_1095;
wire [8:0] u_ca_in_1096;
wire [8:0] u_ca_in_1097;
wire [8:0] u_ca_in_1098;
wire [8:0] u_ca_in_1099;
wire [8:0] u_ca_in_1100;
wire [8:0] u_ca_in_1101;
wire [8:0] u_ca_in_1102;
wire [8:0] u_ca_in_1103;
wire [8:0] u_ca_in_1104;
wire [8:0] u_ca_in_1105;
wire [8:0] u_ca_in_1106;
wire [8:0] u_ca_in_1107;
wire [8:0] u_ca_in_1108;
wire [8:0] u_ca_in_1109;
wire [8:0] u_ca_in_1110;
wire [8:0] u_ca_in_1111;
wire [8:0] u_ca_in_1112;
wire [8:0] u_ca_in_1113;
wire [8:0] u_ca_in_1114;
wire [8:0] u_ca_in_1115;
wire [8:0] u_ca_in_1116;
wire [8:0] u_ca_in_1117;
wire [8:0] u_ca_in_1118;
wire [8:0] u_ca_in_1119;
wire [8:0] u_ca_in_1120;
wire [8:0] u_ca_in_1121;
wire [8:0] u_ca_in_1122;
wire [8:0] u_ca_in_1123;
wire [8:0] u_ca_in_1124;
wire [8:0] u_ca_in_1125;
wire [8:0] u_ca_in_1126;
wire [8:0] u_ca_in_1127;
wire [8:0] u_ca_in_1128;
wire [8:0] u_ca_in_1129;
wire [8:0] u_ca_in_1130;
wire [8:0] u_ca_in_1131;
wire [8:0] u_ca_in_1132;
wire [8:0] u_ca_in_1133;
wire [8:0] u_ca_in_1134;
wire [8:0] u_ca_in_1135;
wire [8:0] u_ca_in_1136;
wire [8:0] u_ca_in_1137;
wire [8:0] u_ca_in_1138;
wire [8:0] u_ca_in_1139;
wire [8:0] u_ca_in_1140;
wire [8:0] u_ca_in_1141;
wire [8:0] u_ca_in_1142;
wire [8:0] u_ca_in_1143;
wire [8:0] u_ca_in_1144;
wire [8:0] u_ca_in_1145;
wire [8:0] u_ca_in_1146;
wire [8:0] u_ca_in_1147;
wire [8:0] u_ca_in_1148;
wire [8:0] u_ca_in_1149;
wire [8:0] u_ca_in_1150;
wire [8:0] u_ca_in_1151;
wire [8:0] u_ca_in_1152;
wire [8:0] u_ca_in_1153;
wire [8:0] u_ca_in_1154;
wire [8:0] u_ca_in_1155;
wire [8:0] u_ca_in_1156;
wire [8:0] u_ca_in_1157;
wire [8:0] u_ca_in_1158;
wire [8:0] u_ca_in_1159;
wire [8:0] u_ca_in_1160;
wire [8:0] u_ca_in_1161;
wire [8:0] u_ca_in_1162;
wire [8:0] u_ca_in_1163;
wire [8:0] u_ca_in_1164;
wire [8:0] u_ca_in_1165;
wire [8:0] u_ca_in_1166;
wire [8:0] u_ca_in_1167;
wire [8:0] u_ca_in_1168;
wire [8:0] u_ca_in_1169;
wire [8:0] u_ca_in_1170;
wire [8:0] u_ca_in_1171;
wire [8:0] u_ca_in_1172;
wire [8:0] u_ca_in_1173;
wire [8:0] u_ca_in_1174;
wire [8:0] u_ca_in_1175;
wire [8:0] u_ca_in_1176;
wire [8:0] u_ca_in_1177;
wire [8:0] u_ca_in_1178;
wire [8:0] u_ca_in_1179;
wire [8:0] u_ca_in_1180;
wire [8:0] u_ca_in_1181;
wire [8:0] u_ca_in_1182;
wire [8:0] u_ca_in_1183;
wire [8:0] u_ca_in_1184;
wire [8:0] u_ca_in_1185;
wire [8:0] u_ca_in_1186;
wire [8:0] u_ca_in_1187;
wire [8:0] u_ca_in_1188;
wire [8:0] u_ca_in_1189;
wire [8:0] u_ca_in_1190;
wire [8:0] u_ca_in_1191;
wire [8:0] u_ca_in_1192;
wire [8:0] u_ca_in_1193;
wire [8:0] u_ca_in_1194;
wire [8:0] u_ca_in_1195;
wire [8:0] u_ca_in_1196;
wire [8:0] u_ca_in_1197;
wire [8:0] u_ca_in_1198;
wire [8:0] u_ca_in_1199;
wire [8:0] u_ca_in_1200;
wire [8:0] u_ca_in_1201;
wire [8:0] u_ca_in_1202;
wire [8:0] u_ca_in_1203;
wire [8:0] u_ca_in_1204;
wire [8:0] u_ca_in_1205;
wire [8:0] u_ca_in_1206;
wire [8:0] u_ca_in_1207;
wire [8:0] u_ca_in_1208;
wire [8:0] u_ca_in_1209;
wire [8:0] u_ca_in_1210;
wire [8:0] u_ca_in_1211;
wire [8:0] u_ca_in_1212;
wire [8:0] u_ca_in_1213;
wire [8:0] u_ca_in_1214;
wire [8:0] u_ca_in_1215;
wire [8:0] u_ca_in_1216;
wire [8:0] u_ca_in_1217;
wire [8:0] u_ca_in_1218;
wire [8:0] u_ca_in_1219;
wire [8:0] u_ca_in_1220;
wire [8:0] u_ca_in_1221;
wire [8:0] u_ca_in_1222;
wire [8:0] u_ca_in_1223;
wire [8:0] u_ca_in_1224;
wire [8:0] u_ca_in_1225;
wire [8:0] u_ca_in_1226;
wire [8:0] u_ca_in_1227;
wire [8:0] u_ca_in_1228;
wire [8:0] u_ca_in_1229;
wire [8:0] u_ca_in_1230;
wire [8:0] u_ca_in_1231;
wire [8:0] u_ca_in_1232;
wire [8:0] u_ca_in_1233;
wire [8:0] u_ca_in_1234;
wire [8:0] u_ca_in_1235;
wire [8:0] u_ca_in_1236;
wire [8:0] u_ca_in_1237;
wire [8:0] u_ca_in_1238;
wire [8:0] u_ca_in_1239;
wire [8:0] u_ca_in_1240;
wire [8:0] u_ca_in_1241;
wire [8:0] u_ca_in_1242;
wire [8:0] u_ca_in_1243;
wire [8:0] u_ca_in_1244;
wire [8:0] u_ca_in_1245;
wire [8:0] u_ca_in_1246;
wire [8:0] u_ca_in_1247;
wire [8:0] u_ca_in_1248;
wire [8:0] u_ca_in_1249;
wire [8:0] u_ca_in_1250;
wire [8:0] u_ca_in_1251;
wire [8:0] u_ca_in_1252;
wire [8:0] u_ca_in_1253;
wire [8:0] u_ca_in_1254;
wire [8:0] u_ca_in_1255;
wire [8:0] u_ca_in_1256;
wire [8:0] u_ca_in_1257;
wire [8:0] u_ca_in_1258;
wire [8:0] u_ca_in_1259;
wire [8:0] u_ca_in_1260;
wire [8:0] u_ca_in_1261;
wire [8:0] u_ca_in_1262;
wire [8:0] u_ca_in_1263;
wire [8:0] u_ca_in_1264;
wire [8:0] u_ca_in_1265;
wire [8:0] u_ca_in_1266;
wire [8:0] u_ca_in_1267;
wire [8:0] u_ca_in_1268;
wire [8:0] u_ca_in_1269;
wire [8:0] u_ca_in_1270;
wire [8:0] u_ca_in_1271;
wire [8:0] u_ca_in_1272;
wire [8:0] u_ca_in_1273;
wire [8:0] u_ca_in_1274;
wire [8:0] u_ca_in_1275;
wire [8:0] u_ca_in_1276;
wire [8:0] u_ca_in_1277;
wire [8:0] u_ca_in_1278;
wire [8:0] u_ca_in_1279;
wire [8:0] u_ca_in_1280;
wire [8:0] u_ca_in_1281;
wire [8:0] u_ca_in_1282;
wire [8:0] u_ca_in_1283;
wire [8:0] u_ca_in_1284;
wire [8:0] u_ca_in_1285;
wire [8:0] u_ca_in_1286;
wire [8:0] u_ca_in_1287;


wire [5:0] u_ca_out_0;
wire [5:0] u_ca_out_1;
wire [5:0] u_ca_out_2;
wire [5:0] u_ca_out_3;
wire [5:0] u_ca_out_4;
wire [5:0] u_ca_out_5;
wire [5:0] u_ca_out_6;
wire [5:0] u_ca_out_7;
wire [5:0] u_ca_out_8;
wire [5:0] u_ca_out_9;
wire [5:0] u_ca_out_10;
wire [5:0] u_ca_out_11;
wire [5:0] u_ca_out_12;
wire [5:0] u_ca_out_13;
wire [5:0] u_ca_out_14;
wire [5:0] u_ca_out_15;
wire [5:0] u_ca_out_16;
wire [5:0] u_ca_out_17;
wire [5:0] u_ca_out_18;
wire [5:0] u_ca_out_19;
wire [5:0] u_ca_out_20;
wire [5:0] u_ca_out_21;
wire [5:0] u_ca_out_22;
wire [5:0] u_ca_out_23;
wire [5:0] u_ca_out_24;
wire [5:0] u_ca_out_25;
wire [5:0] u_ca_out_26;
wire [5:0] u_ca_out_27;
wire [5:0] u_ca_out_28;
wire [5:0] u_ca_out_29;
wire [5:0] u_ca_out_30;
wire [5:0] u_ca_out_31;
wire [5:0] u_ca_out_32;
wire [5:0] u_ca_out_33;
wire [5:0] u_ca_out_34;
wire [5:0] u_ca_out_35;
wire [5:0] u_ca_out_36;
wire [5:0] u_ca_out_37;
wire [5:0] u_ca_out_38;
wire [5:0] u_ca_out_39;
wire [5:0] u_ca_out_40;
wire [5:0] u_ca_out_41;
wire [5:0] u_ca_out_42;
wire [5:0] u_ca_out_43;
wire [5:0] u_ca_out_44;
wire [5:0] u_ca_out_45;
wire [5:0] u_ca_out_46;
wire [5:0] u_ca_out_47;
wire [5:0] u_ca_out_48;
wire [5:0] u_ca_out_49;
wire [5:0] u_ca_out_50;
wire [5:0] u_ca_out_51;
wire [5:0] u_ca_out_52;
wire [5:0] u_ca_out_53;
wire [5:0] u_ca_out_54;
wire [5:0] u_ca_out_55;
wire [5:0] u_ca_out_56;
wire [5:0] u_ca_out_57;
wire [5:0] u_ca_out_58;
wire [5:0] u_ca_out_59;
wire [5:0] u_ca_out_60;
wire [5:0] u_ca_out_61;
wire [5:0] u_ca_out_62;
wire [5:0] u_ca_out_63;
wire [5:0] u_ca_out_64;
wire [5:0] u_ca_out_65;
wire [5:0] u_ca_out_66;
wire [5:0] u_ca_out_67;
wire [5:0] u_ca_out_68;
wire [5:0] u_ca_out_69;
wire [5:0] u_ca_out_70;
wire [5:0] u_ca_out_71;
wire [5:0] u_ca_out_72;
wire [5:0] u_ca_out_73;
wire [5:0] u_ca_out_74;
wire [5:0] u_ca_out_75;
wire [5:0] u_ca_out_76;
wire [5:0] u_ca_out_77;
wire [5:0] u_ca_out_78;
wire [5:0] u_ca_out_79;
wire [5:0] u_ca_out_80;
wire [5:0] u_ca_out_81;
wire [5:0] u_ca_out_82;
wire [5:0] u_ca_out_83;
wire [5:0] u_ca_out_84;
wire [5:0] u_ca_out_85;
wire [5:0] u_ca_out_86;
wire [5:0] u_ca_out_87;
wire [5:0] u_ca_out_88;
wire [5:0] u_ca_out_89;
wire [5:0] u_ca_out_90;
wire [5:0] u_ca_out_91;
wire [5:0] u_ca_out_92;
wire [5:0] u_ca_out_93;
wire [5:0] u_ca_out_94;
wire [5:0] u_ca_out_95;
wire [5:0] u_ca_out_96;
wire [5:0] u_ca_out_97;
wire [5:0] u_ca_out_98;
wire [5:0] u_ca_out_99;
wire [5:0] u_ca_out_100;
wire [5:0] u_ca_out_101;
wire [5:0] u_ca_out_102;
wire [5:0] u_ca_out_103;
wire [5:0] u_ca_out_104;
wire [5:0] u_ca_out_105;
wire [5:0] u_ca_out_106;
wire [5:0] u_ca_out_107;
wire [5:0] u_ca_out_108;
wire [5:0] u_ca_out_109;
wire [5:0] u_ca_out_110;
wire [5:0] u_ca_out_111;
wire [5:0] u_ca_out_112;
wire [5:0] u_ca_out_113;
wire [5:0] u_ca_out_114;
wire [5:0] u_ca_out_115;
wire [5:0] u_ca_out_116;
wire [5:0] u_ca_out_117;
wire [5:0] u_ca_out_118;
wire [5:0] u_ca_out_119;
wire [5:0] u_ca_out_120;
wire [5:0] u_ca_out_121;
wire [5:0] u_ca_out_122;
wire [5:0] u_ca_out_123;
wire [5:0] u_ca_out_124;
wire [5:0] u_ca_out_125;
wire [5:0] u_ca_out_126;
wire [5:0] u_ca_out_127;
wire [5:0] u_ca_out_128;
wire [5:0] u_ca_out_129;
wire [5:0] u_ca_out_130;
wire [5:0] u_ca_out_131;
wire [5:0] u_ca_out_132;
wire [5:0] u_ca_out_133;
wire [5:0] u_ca_out_134;
wire [5:0] u_ca_out_135;
wire [5:0] u_ca_out_136;
wire [5:0] u_ca_out_137;
wire [5:0] u_ca_out_138;
wire [5:0] u_ca_out_139;
wire [5:0] u_ca_out_140;
wire [5:0] u_ca_out_141;
wire [5:0] u_ca_out_142;
wire [5:0] u_ca_out_143;
wire [5:0] u_ca_out_144;
wire [5:0] u_ca_out_145;
wire [5:0] u_ca_out_146;
wire [5:0] u_ca_out_147;
wire [5:0] u_ca_out_148;
wire [5:0] u_ca_out_149;
wire [5:0] u_ca_out_150;
wire [5:0] u_ca_out_151;
wire [5:0] u_ca_out_152;
wire [5:0] u_ca_out_153;
wire [5:0] u_ca_out_154;
wire [5:0] u_ca_out_155;
wire [5:0] u_ca_out_156;
wire [5:0] u_ca_out_157;
wire [5:0] u_ca_out_158;
wire [5:0] u_ca_out_159;
wire [5:0] u_ca_out_160;
wire [5:0] u_ca_out_161;
wire [5:0] u_ca_out_162;
wire [5:0] u_ca_out_163;
wire [5:0] u_ca_out_164;
wire [5:0] u_ca_out_165;
wire [5:0] u_ca_out_166;
wire [5:0] u_ca_out_167;
wire [5:0] u_ca_out_168;
wire [5:0] u_ca_out_169;
wire [5:0] u_ca_out_170;
wire [5:0] u_ca_out_171;
wire [5:0] u_ca_out_172;
wire [5:0] u_ca_out_173;
wire [5:0] u_ca_out_174;
wire [5:0] u_ca_out_175;
wire [5:0] u_ca_out_176;
wire [5:0] u_ca_out_177;
wire [5:0] u_ca_out_178;
wire [5:0] u_ca_out_179;
wire [5:0] u_ca_out_180;
wire [5:0] u_ca_out_181;
wire [5:0] u_ca_out_182;
wire [5:0] u_ca_out_183;
wire [5:0] u_ca_out_184;
wire [5:0] u_ca_out_185;
wire [5:0] u_ca_out_186;
wire [5:0] u_ca_out_187;
wire [5:0] u_ca_out_188;
wire [5:0] u_ca_out_189;
wire [5:0] u_ca_out_190;
wire [5:0] u_ca_out_191;
wire [5:0] u_ca_out_192;
wire [5:0] u_ca_out_193;
wire [5:0] u_ca_out_194;
wire [5:0] u_ca_out_195;
wire [5:0] u_ca_out_196;
wire [5:0] u_ca_out_197;
wire [5:0] u_ca_out_198;
wire [5:0] u_ca_out_199;
wire [5:0] u_ca_out_200;
wire [5:0] u_ca_out_201;
wire [5:0] u_ca_out_202;
wire [5:0] u_ca_out_203;
wire [5:0] u_ca_out_204;
wire [5:0] u_ca_out_205;
wire [5:0] u_ca_out_206;
wire [5:0] u_ca_out_207;
wire [5:0] u_ca_out_208;
wire [5:0] u_ca_out_209;
wire [5:0] u_ca_out_210;
wire [5:0] u_ca_out_211;
wire [5:0] u_ca_out_212;
wire [5:0] u_ca_out_213;
wire [5:0] u_ca_out_214;
wire [5:0] u_ca_out_215;
wire [5:0] u_ca_out_216;
wire [5:0] u_ca_out_217;
wire [5:0] u_ca_out_218;
wire [5:0] u_ca_out_219;
wire [5:0] u_ca_out_220;
wire [5:0] u_ca_out_221;
wire [5:0] u_ca_out_222;
wire [5:0] u_ca_out_223;
wire [5:0] u_ca_out_224;
wire [5:0] u_ca_out_225;
wire [5:0] u_ca_out_226;
wire [5:0] u_ca_out_227;
wire [5:0] u_ca_out_228;
wire [5:0] u_ca_out_229;
wire [5:0] u_ca_out_230;
wire [5:0] u_ca_out_231;
wire [5:0] u_ca_out_232;
wire [5:0] u_ca_out_233;
wire [5:0] u_ca_out_234;
wire [5:0] u_ca_out_235;
wire [5:0] u_ca_out_236;
wire [5:0] u_ca_out_237;
wire [5:0] u_ca_out_238;
wire [5:0] u_ca_out_239;
wire [5:0] u_ca_out_240;
wire [5:0] u_ca_out_241;
wire [5:0] u_ca_out_242;
wire [5:0] u_ca_out_243;
wire [5:0] u_ca_out_244;
wire [5:0] u_ca_out_245;
wire [5:0] u_ca_out_246;
wire [5:0] u_ca_out_247;
wire [5:0] u_ca_out_248;
wire [5:0] u_ca_out_249;
wire [5:0] u_ca_out_250;
wire [5:0] u_ca_out_251;
wire [5:0] u_ca_out_252;
wire [5:0] u_ca_out_253;
wire [5:0] u_ca_out_254;
wire [5:0] u_ca_out_255;
wire [5:0] u_ca_out_256;
wire [5:0] u_ca_out_257;
wire [5:0] u_ca_out_258;
wire [5:0] u_ca_out_259;
wire [5:0] u_ca_out_260;
wire [5:0] u_ca_out_261;
wire [5:0] u_ca_out_262;
wire [5:0] u_ca_out_263;
wire [5:0] u_ca_out_264;
wire [5:0] u_ca_out_265;
wire [5:0] u_ca_out_266;
wire [5:0] u_ca_out_267;
wire [5:0] u_ca_out_268;
wire [5:0] u_ca_out_269;
wire [5:0] u_ca_out_270;
wire [5:0] u_ca_out_271;
wire [5:0] u_ca_out_272;
wire [5:0] u_ca_out_273;
wire [5:0] u_ca_out_274;
wire [5:0] u_ca_out_275;
wire [5:0] u_ca_out_276;
wire [5:0] u_ca_out_277;
wire [5:0] u_ca_out_278;
wire [5:0] u_ca_out_279;
wire [5:0] u_ca_out_280;
wire [5:0] u_ca_out_281;
wire [5:0] u_ca_out_282;
wire [5:0] u_ca_out_283;
wire [5:0] u_ca_out_284;
wire [5:0] u_ca_out_285;
wire [5:0] u_ca_out_286;
wire [5:0] u_ca_out_287;
wire [5:0] u_ca_out_288;
wire [5:0] u_ca_out_289;
wire [5:0] u_ca_out_290;
wire [5:0] u_ca_out_291;
wire [5:0] u_ca_out_292;
wire [5:0] u_ca_out_293;
wire [5:0] u_ca_out_294;
wire [5:0] u_ca_out_295;
wire [5:0] u_ca_out_296;
wire [5:0] u_ca_out_297;
wire [5:0] u_ca_out_298;
wire [5:0] u_ca_out_299;
wire [5:0] u_ca_out_300;
wire [5:0] u_ca_out_301;
wire [5:0] u_ca_out_302;
wire [5:0] u_ca_out_303;
wire [5:0] u_ca_out_304;
wire [5:0] u_ca_out_305;
wire [5:0] u_ca_out_306;
wire [5:0] u_ca_out_307;
wire [5:0] u_ca_out_308;
wire [5:0] u_ca_out_309;
wire [5:0] u_ca_out_310;
wire [5:0] u_ca_out_311;
wire [5:0] u_ca_out_312;
wire [5:0] u_ca_out_313;
wire [5:0] u_ca_out_314;
wire [5:0] u_ca_out_315;
wire [5:0] u_ca_out_316;
wire [5:0] u_ca_out_317;
wire [5:0] u_ca_out_318;
wire [5:0] u_ca_out_319;
wire [5:0] u_ca_out_320;
wire [5:0] u_ca_out_321;
wire [5:0] u_ca_out_322;
wire [5:0] u_ca_out_323;
wire [5:0] u_ca_out_324;
wire [5:0] u_ca_out_325;
wire [5:0] u_ca_out_326;
wire [5:0] u_ca_out_327;
wire [5:0] u_ca_out_328;
wire [5:0] u_ca_out_329;
wire [5:0] u_ca_out_330;
wire [5:0] u_ca_out_331;
wire [5:0] u_ca_out_332;
wire [5:0] u_ca_out_333;
wire [5:0] u_ca_out_334;
wire [5:0] u_ca_out_335;
wire [5:0] u_ca_out_336;
wire [5:0] u_ca_out_337;
wire [5:0] u_ca_out_338;
wire [5:0] u_ca_out_339;
wire [5:0] u_ca_out_340;
wire [5:0] u_ca_out_341;
wire [5:0] u_ca_out_342;
wire [5:0] u_ca_out_343;
wire [5:0] u_ca_out_344;
wire [5:0] u_ca_out_345;
wire [5:0] u_ca_out_346;
wire [5:0] u_ca_out_347;
wire [5:0] u_ca_out_348;
wire [5:0] u_ca_out_349;
wire [5:0] u_ca_out_350;
wire [5:0] u_ca_out_351;
wire [5:0] u_ca_out_352;
wire [5:0] u_ca_out_353;
wire [5:0] u_ca_out_354;
wire [5:0] u_ca_out_355;
wire [5:0] u_ca_out_356;
wire [5:0] u_ca_out_357;
wire [5:0] u_ca_out_358;
wire [5:0] u_ca_out_359;
wire [5:0] u_ca_out_360;
wire [5:0] u_ca_out_361;
wire [5:0] u_ca_out_362;
wire [5:0] u_ca_out_363;
wire [5:0] u_ca_out_364;
wire [5:0] u_ca_out_365;
wire [5:0] u_ca_out_366;
wire [5:0] u_ca_out_367;
wire [5:0] u_ca_out_368;
wire [5:0] u_ca_out_369;
wire [5:0] u_ca_out_370;
wire [5:0] u_ca_out_371;
wire [5:0] u_ca_out_372;
wire [5:0] u_ca_out_373;
wire [5:0] u_ca_out_374;
wire [5:0] u_ca_out_375;
wire [5:0] u_ca_out_376;
wire [5:0] u_ca_out_377;
wire [5:0] u_ca_out_378;
wire [5:0] u_ca_out_379;
wire [5:0] u_ca_out_380;
wire [5:0] u_ca_out_381;
wire [5:0] u_ca_out_382;
wire [5:0] u_ca_out_383;
wire [5:0] u_ca_out_384;
wire [5:0] u_ca_out_385;
wire [5:0] u_ca_out_386;
wire [5:0] u_ca_out_387;
wire [5:0] u_ca_out_388;
wire [5:0] u_ca_out_389;
wire [5:0] u_ca_out_390;
wire [5:0] u_ca_out_391;
wire [5:0] u_ca_out_392;
wire [5:0] u_ca_out_393;
wire [5:0] u_ca_out_394;
wire [5:0] u_ca_out_395;
wire [5:0] u_ca_out_396;
wire [5:0] u_ca_out_397;
wire [5:0] u_ca_out_398;
wire [5:0] u_ca_out_399;
wire [5:0] u_ca_out_400;
wire [5:0] u_ca_out_401;
wire [5:0] u_ca_out_402;
wire [5:0] u_ca_out_403;
wire [5:0] u_ca_out_404;
wire [5:0] u_ca_out_405;
wire [5:0] u_ca_out_406;
wire [5:0] u_ca_out_407;
wire [5:0] u_ca_out_408;
wire [5:0] u_ca_out_409;
wire [5:0] u_ca_out_410;
wire [5:0] u_ca_out_411;
wire [5:0] u_ca_out_412;
wire [5:0] u_ca_out_413;
wire [5:0] u_ca_out_414;
wire [5:0] u_ca_out_415;
wire [5:0] u_ca_out_416;
wire [5:0] u_ca_out_417;
wire [5:0] u_ca_out_418;
wire [5:0] u_ca_out_419;
wire [5:0] u_ca_out_420;
wire [5:0] u_ca_out_421;
wire [5:0] u_ca_out_422;
wire [5:0] u_ca_out_423;
wire [5:0] u_ca_out_424;
wire [5:0] u_ca_out_425;
wire [5:0] u_ca_out_426;
wire [5:0] u_ca_out_427;
wire [5:0] u_ca_out_428;
wire [5:0] u_ca_out_429;
wire [5:0] u_ca_out_430;
wire [5:0] u_ca_out_431;
wire [5:0] u_ca_out_432;
wire [5:0] u_ca_out_433;
wire [5:0] u_ca_out_434;
wire [5:0] u_ca_out_435;
wire [5:0] u_ca_out_436;
wire [5:0] u_ca_out_437;
wire [5:0] u_ca_out_438;
wire [5:0] u_ca_out_439;
wire [5:0] u_ca_out_440;
wire [5:0] u_ca_out_441;
wire [5:0] u_ca_out_442;
wire [5:0] u_ca_out_443;
wire [5:0] u_ca_out_444;
wire [5:0] u_ca_out_445;
wire [5:0] u_ca_out_446;
wire [5:0] u_ca_out_447;
wire [5:0] u_ca_out_448;
wire [5:0] u_ca_out_449;
wire [5:0] u_ca_out_450;
wire [5:0] u_ca_out_451;
wire [5:0] u_ca_out_452;
wire [5:0] u_ca_out_453;
wire [5:0] u_ca_out_454;
wire [5:0] u_ca_out_455;
wire [5:0] u_ca_out_456;
wire [5:0] u_ca_out_457;
wire [5:0] u_ca_out_458;
wire [5:0] u_ca_out_459;
wire [5:0] u_ca_out_460;
wire [5:0] u_ca_out_461;
wire [5:0] u_ca_out_462;
wire [5:0] u_ca_out_463;
wire [5:0] u_ca_out_464;
wire [5:0] u_ca_out_465;
wire [5:0] u_ca_out_466;
wire [5:0] u_ca_out_467;
wire [5:0] u_ca_out_468;
wire [5:0] u_ca_out_469;
wire [5:0] u_ca_out_470;
wire [5:0] u_ca_out_471;
wire [5:0] u_ca_out_472;
wire [5:0] u_ca_out_473;
wire [5:0] u_ca_out_474;
wire [5:0] u_ca_out_475;
wire [5:0] u_ca_out_476;
wire [5:0] u_ca_out_477;
wire [5:0] u_ca_out_478;
wire [5:0] u_ca_out_479;
wire [5:0] u_ca_out_480;
wire [5:0] u_ca_out_481;
wire [5:0] u_ca_out_482;
wire [5:0] u_ca_out_483;
wire [5:0] u_ca_out_484;
wire [5:0] u_ca_out_485;
wire [5:0] u_ca_out_486;
wire [5:0] u_ca_out_487;
wire [5:0] u_ca_out_488;
wire [5:0] u_ca_out_489;
wire [5:0] u_ca_out_490;
wire [5:0] u_ca_out_491;
wire [5:0] u_ca_out_492;
wire [5:0] u_ca_out_493;
wire [5:0] u_ca_out_494;
wire [5:0] u_ca_out_495;
wire [5:0] u_ca_out_496;
wire [5:0] u_ca_out_497;
wire [5:0] u_ca_out_498;
wire [5:0] u_ca_out_499;
wire [5:0] u_ca_out_500;
wire [5:0] u_ca_out_501;
wire [5:0] u_ca_out_502;
wire [5:0] u_ca_out_503;
wire [5:0] u_ca_out_504;
wire [5:0] u_ca_out_505;
wire [5:0] u_ca_out_506;
wire [5:0] u_ca_out_507;
wire [5:0] u_ca_out_508;
wire [5:0] u_ca_out_509;
wire [5:0] u_ca_out_510;
wire [5:0] u_ca_out_511;
wire [5:0] u_ca_out_512;
wire [5:0] u_ca_out_513;
wire [5:0] u_ca_out_514;
wire [5:0] u_ca_out_515;
wire [5:0] u_ca_out_516;
wire [5:0] u_ca_out_517;
wire [5:0] u_ca_out_518;
wire [5:0] u_ca_out_519;
wire [5:0] u_ca_out_520;
wire [5:0] u_ca_out_521;
wire [5:0] u_ca_out_522;
wire [5:0] u_ca_out_523;
wire [5:0] u_ca_out_524;
wire [5:0] u_ca_out_525;
wire [5:0] u_ca_out_526;
wire [5:0] u_ca_out_527;
wire [5:0] u_ca_out_528;
wire [5:0] u_ca_out_529;
wire [5:0] u_ca_out_530;
wire [5:0] u_ca_out_531;
wire [5:0] u_ca_out_532;
wire [5:0] u_ca_out_533;
wire [5:0] u_ca_out_534;
wire [5:0] u_ca_out_535;
wire [5:0] u_ca_out_536;
wire [5:0] u_ca_out_537;
wire [5:0] u_ca_out_538;
wire [5:0] u_ca_out_539;
wire [5:0] u_ca_out_540;
wire [5:0] u_ca_out_541;
wire [5:0] u_ca_out_542;
wire [5:0] u_ca_out_543;
wire [5:0] u_ca_out_544;
wire [5:0] u_ca_out_545;
wire [5:0] u_ca_out_546;
wire [5:0] u_ca_out_547;
wire [5:0] u_ca_out_548;
wire [5:0] u_ca_out_549;
wire [5:0] u_ca_out_550;
wire [5:0] u_ca_out_551;
wire [5:0] u_ca_out_552;
wire [5:0] u_ca_out_553;
wire [5:0] u_ca_out_554;
wire [5:0] u_ca_out_555;
wire [5:0] u_ca_out_556;
wire [5:0] u_ca_out_557;
wire [5:0] u_ca_out_558;
wire [5:0] u_ca_out_559;
wire [5:0] u_ca_out_560;
wire [5:0] u_ca_out_561;
wire [5:0] u_ca_out_562;
wire [5:0] u_ca_out_563;
wire [5:0] u_ca_out_564;
wire [5:0] u_ca_out_565;
wire [5:0] u_ca_out_566;
wire [5:0] u_ca_out_567;
wire [5:0] u_ca_out_568;
wire [5:0] u_ca_out_569;
wire [5:0] u_ca_out_570;
wire [5:0] u_ca_out_571;
wire [5:0] u_ca_out_572;
wire [5:0] u_ca_out_573;
wire [5:0] u_ca_out_574;
wire [5:0] u_ca_out_575;
wire [5:0] u_ca_out_576;
wire [5:0] u_ca_out_577;
wire [5:0] u_ca_out_578;
wire [5:0] u_ca_out_579;
wire [5:0] u_ca_out_580;
wire [5:0] u_ca_out_581;
wire [5:0] u_ca_out_582;
wire [5:0] u_ca_out_583;
wire [5:0] u_ca_out_584;
wire [5:0] u_ca_out_585;
wire [5:0] u_ca_out_586;
wire [5:0] u_ca_out_587;
wire [5:0] u_ca_out_588;
wire [5:0] u_ca_out_589;
wire [5:0] u_ca_out_590;
wire [5:0] u_ca_out_591;
wire [5:0] u_ca_out_592;
wire [5:0] u_ca_out_593;
wire [5:0] u_ca_out_594;
wire [5:0] u_ca_out_595;
wire [5:0] u_ca_out_596;
wire [5:0] u_ca_out_597;
wire [5:0] u_ca_out_598;
wire [5:0] u_ca_out_599;
wire [5:0] u_ca_out_600;
wire [5:0] u_ca_out_601;
wire [5:0] u_ca_out_602;
wire [5:0] u_ca_out_603;
wire [5:0] u_ca_out_604;
wire [5:0] u_ca_out_605;
wire [5:0] u_ca_out_606;
wire [5:0] u_ca_out_607;
wire [5:0] u_ca_out_608;
wire [5:0] u_ca_out_609;
wire [5:0] u_ca_out_610;
wire [5:0] u_ca_out_611;
wire [5:0] u_ca_out_612;
wire [5:0] u_ca_out_613;
wire [5:0] u_ca_out_614;
wire [5:0] u_ca_out_615;
wire [5:0] u_ca_out_616;
wire [5:0] u_ca_out_617;
wire [5:0] u_ca_out_618;
wire [5:0] u_ca_out_619;
wire [5:0] u_ca_out_620;
wire [5:0] u_ca_out_621;
wire [5:0] u_ca_out_622;
wire [5:0] u_ca_out_623;
wire [5:0] u_ca_out_624;
wire [5:0] u_ca_out_625;
wire [5:0] u_ca_out_626;
wire [5:0] u_ca_out_627;
wire [5:0] u_ca_out_628;
wire [5:0] u_ca_out_629;
wire [5:0] u_ca_out_630;
wire [5:0] u_ca_out_631;
wire [5:0] u_ca_out_632;
wire [5:0] u_ca_out_633;
wire [5:0] u_ca_out_634;
wire [5:0] u_ca_out_635;
wire [5:0] u_ca_out_636;
wire [5:0] u_ca_out_637;
wire [5:0] u_ca_out_638;
wire [5:0] u_ca_out_639;
wire [5:0] u_ca_out_640;
wire [5:0] u_ca_out_641;
wire [5:0] u_ca_out_642;
wire [5:0] u_ca_out_643;
wire [5:0] u_ca_out_644;
wire [5:0] u_ca_out_645;
wire [5:0] u_ca_out_646;
wire [5:0] u_ca_out_647;
wire [5:0] u_ca_out_648;
wire [5:0] u_ca_out_649;
wire [5:0] u_ca_out_650;
wire [5:0] u_ca_out_651;
wire [5:0] u_ca_out_652;
wire [5:0] u_ca_out_653;
wire [5:0] u_ca_out_654;
wire [5:0] u_ca_out_655;
wire [5:0] u_ca_out_656;
wire [5:0] u_ca_out_657;
wire [5:0] u_ca_out_658;
wire [5:0] u_ca_out_659;
wire [5:0] u_ca_out_660;
wire [5:0] u_ca_out_661;
wire [5:0] u_ca_out_662;
wire [5:0] u_ca_out_663;
wire [5:0] u_ca_out_664;
wire [5:0] u_ca_out_665;
wire [5:0] u_ca_out_666;
wire [5:0] u_ca_out_667;
wire [5:0] u_ca_out_668;
wire [5:0] u_ca_out_669;
wire [5:0] u_ca_out_670;
wire [5:0] u_ca_out_671;
wire [5:0] u_ca_out_672;
wire [5:0] u_ca_out_673;
wire [5:0] u_ca_out_674;
wire [5:0] u_ca_out_675;
wire [5:0] u_ca_out_676;
wire [5:0] u_ca_out_677;
wire [5:0] u_ca_out_678;
wire [5:0] u_ca_out_679;
wire [5:0] u_ca_out_680;
wire [5:0] u_ca_out_681;
wire [5:0] u_ca_out_682;
wire [5:0] u_ca_out_683;
wire [5:0] u_ca_out_684;
wire [5:0] u_ca_out_685;
wire [5:0] u_ca_out_686;
wire [5:0] u_ca_out_687;
wire [5:0] u_ca_out_688;
wire [5:0] u_ca_out_689;
wire [5:0] u_ca_out_690;
wire [5:0] u_ca_out_691;
wire [5:0] u_ca_out_692;
wire [5:0] u_ca_out_693;
wire [5:0] u_ca_out_694;
wire [5:0] u_ca_out_695;
wire [5:0] u_ca_out_696;
wire [5:0] u_ca_out_697;
wire [5:0] u_ca_out_698;
wire [5:0] u_ca_out_699;
wire [5:0] u_ca_out_700;
wire [5:0] u_ca_out_701;
wire [5:0] u_ca_out_702;
wire [5:0] u_ca_out_703;
wire [5:0] u_ca_out_704;
wire [5:0] u_ca_out_705;
wire [5:0] u_ca_out_706;
wire [5:0] u_ca_out_707;
wire [5:0] u_ca_out_708;
wire [5:0] u_ca_out_709;
wire [5:0] u_ca_out_710;
wire [5:0] u_ca_out_711;
wire [5:0] u_ca_out_712;
wire [5:0] u_ca_out_713;
wire [5:0] u_ca_out_714;
wire [5:0] u_ca_out_715;
wire [5:0] u_ca_out_716;
wire [5:0] u_ca_out_717;
wire [5:0] u_ca_out_718;
wire [5:0] u_ca_out_719;
wire [5:0] u_ca_out_720;
wire [5:0] u_ca_out_721;
wire [5:0] u_ca_out_722;
wire [5:0] u_ca_out_723;
wire [5:0] u_ca_out_724;
wire [5:0] u_ca_out_725;
wire [5:0] u_ca_out_726;
wire [5:0] u_ca_out_727;
wire [5:0] u_ca_out_728;
wire [5:0] u_ca_out_729;
wire [5:0] u_ca_out_730;
wire [5:0] u_ca_out_731;
wire [5:0] u_ca_out_732;
wire [5:0] u_ca_out_733;
wire [5:0] u_ca_out_734;
wire [5:0] u_ca_out_735;
wire [5:0] u_ca_out_736;
wire [5:0] u_ca_out_737;
wire [5:0] u_ca_out_738;
wire [5:0] u_ca_out_739;
wire [5:0] u_ca_out_740;
wire [5:0] u_ca_out_741;
wire [5:0] u_ca_out_742;
wire [5:0] u_ca_out_743;
wire [5:0] u_ca_out_744;
wire [5:0] u_ca_out_745;
wire [5:0] u_ca_out_746;
wire [5:0] u_ca_out_747;
wire [5:0] u_ca_out_748;
wire [5:0] u_ca_out_749;
wire [5:0] u_ca_out_750;
wire [5:0] u_ca_out_751;
wire [5:0] u_ca_out_752;
wire [5:0] u_ca_out_753;
wire [5:0] u_ca_out_754;
wire [5:0] u_ca_out_755;
wire [5:0] u_ca_out_756;
wire [5:0] u_ca_out_757;
wire [5:0] u_ca_out_758;
wire [5:0] u_ca_out_759;
wire [5:0] u_ca_out_760;
wire [5:0] u_ca_out_761;
wire [5:0] u_ca_out_762;
wire [5:0] u_ca_out_763;
wire [5:0] u_ca_out_764;
wire [5:0] u_ca_out_765;
wire [5:0] u_ca_out_766;
wire [5:0] u_ca_out_767;
wire [5:0] u_ca_out_768;
wire [5:0] u_ca_out_769;
wire [5:0] u_ca_out_770;
wire [5:0] u_ca_out_771;
wire [5:0] u_ca_out_772;
wire [5:0] u_ca_out_773;
wire [5:0] u_ca_out_774;
wire [5:0] u_ca_out_775;
wire [5:0] u_ca_out_776;
wire [5:0] u_ca_out_777;
wire [5:0] u_ca_out_778;
wire [5:0] u_ca_out_779;
wire [5:0] u_ca_out_780;
wire [5:0] u_ca_out_781;
wire [5:0] u_ca_out_782;
wire [5:0] u_ca_out_783;
wire [5:0] u_ca_out_784;
wire [5:0] u_ca_out_785;
wire [5:0] u_ca_out_786;
wire [5:0] u_ca_out_787;
wire [5:0] u_ca_out_788;
wire [5:0] u_ca_out_789;
wire [5:0] u_ca_out_790;
wire [5:0] u_ca_out_791;
wire [5:0] u_ca_out_792;
wire [5:0] u_ca_out_793;
wire [5:0] u_ca_out_794;
wire [5:0] u_ca_out_795;
wire [5:0] u_ca_out_796;
wire [5:0] u_ca_out_797;
wire [5:0] u_ca_out_798;
wire [5:0] u_ca_out_799;
wire [5:0] u_ca_out_800;
wire [5:0] u_ca_out_801;
wire [5:0] u_ca_out_802;
wire [5:0] u_ca_out_803;
wire [5:0] u_ca_out_804;
wire [5:0] u_ca_out_805;
wire [5:0] u_ca_out_806;
wire [5:0] u_ca_out_807;
wire [5:0] u_ca_out_808;
wire [5:0] u_ca_out_809;
wire [5:0] u_ca_out_810;
wire [5:0] u_ca_out_811;
wire [5:0] u_ca_out_812;
wire [5:0] u_ca_out_813;
wire [5:0] u_ca_out_814;
wire [5:0] u_ca_out_815;
wire [5:0] u_ca_out_816;
wire [5:0] u_ca_out_817;
wire [5:0] u_ca_out_818;
wire [5:0] u_ca_out_819;
wire [5:0] u_ca_out_820;
wire [5:0] u_ca_out_821;
wire [5:0] u_ca_out_822;
wire [5:0] u_ca_out_823;
wire [5:0] u_ca_out_824;
wire [5:0] u_ca_out_825;
wire [5:0] u_ca_out_826;
wire [5:0] u_ca_out_827;
wire [5:0] u_ca_out_828;
wire [5:0] u_ca_out_829;
wire [5:0] u_ca_out_830;
wire [5:0] u_ca_out_831;
wire [5:0] u_ca_out_832;
wire [5:0] u_ca_out_833;
wire [5:0] u_ca_out_834;
wire [5:0] u_ca_out_835;
wire [5:0] u_ca_out_836;
wire [5:0] u_ca_out_837;
wire [5:0] u_ca_out_838;
wire [5:0] u_ca_out_839;
wire [5:0] u_ca_out_840;
wire [5:0] u_ca_out_841;
wire [5:0] u_ca_out_842;
wire [5:0] u_ca_out_843;
wire [5:0] u_ca_out_844;
wire [5:0] u_ca_out_845;
wire [5:0] u_ca_out_846;
wire [5:0] u_ca_out_847;
wire [5:0] u_ca_out_848;
wire [5:0] u_ca_out_849;
wire [5:0] u_ca_out_850;
wire [5:0] u_ca_out_851;
wire [5:0] u_ca_out_852;
wire [5:0] u_ca_out_853;
wire [5:0] u_ca_out_854;
wire [5:0] u_ca_out_855;
wire [5:0] u_ca_out_856;
wire [5:0] u_ca_out_857;
wire [5:0] u_ca_out_858;
wire [5:0] u_ca_out_859;
wire [5:0] u_ca_out_860;
wire [5:0] u_ca_out_861;
wire [5:0] u_ca_out_862;
wire [5:0] u_ca_out_863;
wire [5:0] u_ca_out_864;
wire [5:0] u_ca_out_865;
wire [5:0] u_ca_out_866;
wire [5:0] u_ca_out_867;
wire [5:0] u_ca_out_868;
wire [5:0] u_ca_out_869;
wire [5:0] u_ca_out_870;
wire [5:0] u_ca_out_871;
wire [5:0] u_ca_out_872;
wire [5:0] u_ca_out_873;
wire [5:0] u_ca_out_874;
wire [5:0] u_ca_out_875;
wire [5:0] u_ca_out_876;
wire [5:0] u_ca_out_877;
wire [5:0] u_ca_out_878;
wire [5:0] u_ca_out_879;
wire [5:0] u_ca_out_880;
wire [5:0] u_ca_out_881;
wire [5:0] u_ca_out_882;
wire [5:0] u_ca_out_883;
wire [5:0] u_ca_out_884;
wire [5:0] u_ca_out_885;
wire [5:0] u_ca_out_886;
wire [5:0] u_ca_out_887;
wire [5:0] u_ca_out_888;
wire [5:0] u_ca_out_889;
wire [5:0] u_ca_out_890;
wire [5:0] u_ca_out_891;
wire [5:0] u_ca_out_892;
wire [5:0] u_ca_out_893;
wire [5:0] u_ca_out_894;
wire [5:0] u_ca_out_895;
wire [5:0] u_ca_out_896;
wire [5:0] u_ca_out_897;
wire [5:0] u_ca_out_898;
wire [5:0] u_ca_out_899;
wire [5:0] u_ca_out_900;
wire [5:0] u_ca_out_901;
wire [5:0] u_ca_out_902;
wire [5:0] u_ca_out_903;
wire [5:0] u_ca_out_904;
wire [5:0] u_ca_out_905;
wire [5:0] u_ca_out_906;
wire [5:0] u_ca_out_907;
wire [5:0] u_ca_out_908;
wire [5:0] u_ca_out_909;
wire [5:0] u_ca_out_910;
wire [5:0] u_ca_out_911;
wire [5:0] u_ca_out_912;
wire [5:0] u_ca_out_913;
wire [5:0] u_ca_out_914;
wire [5:0] u_ca_out_915;
wire [5:0] u_ca_out_916;
wire [5:0] u_ca_out_917;
wire [5:0] u_ca_out_918;
wire [5:0] u_ca_out_919;
wire [5:0] u_ca_out_920;
wire [5:0] u_ca_out_921;
wire [5:0] u_ca_out_922;
wire [5:0] u_ca_out_923;
wire [5:0] u_ca_out_924;
wire [5:0] u_ca_out_925;
wire [5:0] u_ca_out_926;
wire [5:0] u_ca_out_927;
wire [5:0] u_ca_out_928;
wire [5:0] u_ca_out_929;
wire [5:0] u_ca_out_930;
wire [5:0] u_ca_out_931;
wire [5:0] u_ca_out_932;
wire [5:0] u_ca_out_933;
wire [5:0] u_ca_out_934;
wire [5:0] u_ca_out_935;
wire [5:0] u_ca_out_936;
wire [5:0] u_ca_out_937;
wire [5:0] u_ca_out_938;
wire [5:0] u_ca_out_939;
wire [5:0] u_ca_out_940;
wire [5:0] u_ca_out_941;
wire [5:0] u_ca_out_942;
wire [5:0] u_ca_out_943;
wire [5:0] u_ca_out_944;
wire [5:0] u_ca_out_945;
wire [5:0] u_ca_out_946;
wire [5:0] u_ca_out_947;
wire [5:0] u_ca_out_948;
wire [5:0] u_ca_out_949;
wire [5:0] u_ca_out_950;
wire [5:0] u_ca_out_951;
wire [5:0] u_ca_out_952;
wire [5:0] u_ca_out_953;
wire [5:0] u_ca_out_954;
wire [5:0] u_ca_out_955;
wire [5:0] u_ca_out_956;
wire [5:0] u_ca_out_957;
wire [5:0] u_ca_out_958;
wire [5:0] u_ca_out_959;
wire [5:0] u_ca_out_960;
wire [5:0] u_ca_out_961;
wire [5:0] u_ca_out_962;
wire [5:0] u_ca_out_963;
wire [5:0] u_ca_out_964;
wire [5:0] u_ca_out_965;
wire [5:0] u_ca_out_966;
wire [5:0] u_ca_out_967;
wire [5:0] u_ca_out_968;
wire [5:0] u_ca_out_969;
wire [5:0] u_ca_out_970;
wire [5:0] u_ca_out_971;
wire [5:0] u_ca_out_972;
wire [5:0] u_ca_out_973;
wire [5:0] u_ca_out_974;
wire [5:0] u_ca_out_975;
wire [5:0] u_ca_out_976;
wire [5:0] u_ca_out_977;
wire [5:0] u_ca_out_978;
wire [5:0] u_ca_out_979;
wire [5:0] u_ca_out_980;
wire [5:0] u_ca_out_981;
wire [5:0] u_ca_out_982;
wire [5:0] u_ca_out_983;
wire [5:0] u_ca_out_984;
wire [5:0] u_ca_out_985;
wire [5:0] u_ca_out_986;
wire [5:0] u_ca_out_987;
wire [5:0] u_ca_out_988;
wire [5:0] u_ca_out_989;
wire [5:0] u_ca_out_990;
wire [5:0] u_ca_out_991;
wire [5:0] u_ca_out_992;
wire [5:0] u_ca_out_993;
wire [5:0] u_ca_out_994;
wire [5:0] u_ca_out_995;
wire [5:0] u_ca_out_996;
wire [5:0] u_ca_out_997;
wire [5:0] u_ca_out_998;
wire [5:0] u_ca_out_999;
wire [5:0] u_ca_out_1000;
wire [5:0] u_ca_out_1001;
wire [5:0] u_ca_out_1002;
wire [5:0] u_ca_out_1003;
wire [5:0] u_ca_out_1004;
wire [5:0] u_ca_out_1005;
wire [5:0] u_ca_out_1006;
wire [5:0] u_ca_out_1007;
wire [5:0] u_ca_out_1008;
wire [5:0] u_ca_out_1009;
wire [5:0] u_ca_out_1010;
wire [5:0] u_ca_out_1011;
wire [5:0] u_ca_out_1012;
wire [5:0] u_ca_out_1013;
wire [5:0] u_ca_out_1014;
wire [5:0] u_ca_out_1015;
wire [5:0] u_ca_out_1016;
wire [5:0] u_ca_out_1017;
wire [5:0] u_ca_out_1018;
wire [5:0] u_ca_out_1019;
wire [5:0] u_ca_out_1020;
wire [5:0] u_ca_out_1021;
wire [5:0] u_ca_out_1022;
wire [5:0] u_ca_out_1023;
wire [5:0] u_ca_out_1024;
wire [5:0] u_ca_out_1025;
wire [5:0] u_ca_out_1026;
wire [5:0] u_ca_out_1027;
wire [5:0] u_ca_out_1028;
wire [5:0] u_ca_out_1029;
wire [5:0] u_ca_out_1030;
wire [5:0] u_ca_out_1031;
wire [5:0] u_ca_out_1032;
wire [5:0] u_ca_out_1033;
wire [5:0] u_ca_out_1034;
wire [5:0] u_ca_out_1035;
wire [5:0] u_ca_out_1036;
wire [5:0] u_ca_out_1037;
wire [5:0] u_ca_out_1038;
wire [5:0] u_ca_out_1039;
wire [5:0] u_ca_out_1040;
wire [5:0] u_ca_out_1041;
wire [5:0] u_ca_out_1042;
wire [5:0] u_ca_out_1043;
wire [5:0] u_ca_out_1044;
wire [5:0] u_ca_out_1045;
wire [5:0] u_ca_out_1046;
wire [5:0] u_ca_out_1047;
wire [5:0] u_ca_out_1048;
wire [5:0] u_ca_out_1049;
wire [5:0] u_ca_out_1050;
wire [5:0] u_ca_out_1051;
wire [5:0] u_ca_out_1052;
wire [5:0] u_ca_out_1053;
wire [5:0] u_ca_out_1054;
wire [5:0] u_ca_out_1055;
wire [5:0] u_ca_out_1056;
wire [5:0] u_ca_out_1057;
wire [5:0] u_ca_out_1058;
wire [5:0] u_ca_out_1059;
wire [5:0] u_ca_out_1060;
wire [5:0] u_ca_out_1061;
wire [5:0] u_ca_out_1062;
wire [5:0] u_ca_out_1063;
wire [5:0] u_ca_out_1064;
wire [5:0] u_ca_out_1065;
wire [5:0] u_ca_out_1066;
wire [5:0] u_ca_out_1067;
wire [5:0] u_ca_out_1068;
wire [5:0] u_ca_out_1069;
wire [5:0] u_ca_out_1070;
wire [5:0] u_ca_out_1071;
wire [5:0] u_ca_out_1072;
wire [5:0] u_ca_out_1073;
wire [5:0] u_ca_out_1074;
wire [5:0] u_ca_out_1075;
wire [5:0] u_ca_out_1076;
wire [5:0] u_ca_out_1077;
wire [5:0] u_ca_out_1078;
wire [5:0] u_ca_out_1079;
wire [5:0] u_ca_out_1080;
wire [5:0] u_ca_out_1081;
wire [5:0] u_ca_out_1082;
wire [5:0] u_ca_out_1083;
wire [5:0] u_ca_out_1084;
wire [5:0] u_ca_out_1085;
wire [5:0] u_ca_out_1086;
wire [5:0] u_ca_out_1087;
wire [5:0] u_ca_out_1088;
wire [5:0] u_ca_out_1089;
wire [5:0] u_ca_out_1090;
wire [5:0] u_ca_out_1091;
wire [5:0] u_ca_out_1092;
wire [5:0] u_ca_out_1093;
wire [5:0] u_ca_out_1094;
wire [5:0] u_ca_out_1095;
wire [5:0] u_ca_out_1096;
wire [5:0] u_ca_out_1097;
wire [5:0] u_ca_out_1098;
wire [5:0] u_ca_out_1099;
wire [5:0] u_ca_out_1100;
wire [5:0] u_ca_out_1101;
wire [5:0] u_ca_out_1102;
wire [5:0] u_ca_out_1103;
wire [5:0] u_ca_out_1104;
wire [5:0] u_ca_out_1105;
wire [5:0] u_ca_out_1106;
wire [5:0] u_ca_out_1107;
wire [5:0] u_ca_out_1108;
wire [5:0] u_ca_out_1109;
wire [5:0] u_ca_out_1110;
wire [5:0] u_ca_out_1111;
wire [5:0] u_ca_out_1112;
wire [5:0] u_ca_out_1113;
wire [5:0] u_ca_out_1114;
wire [5:0] u_ca_out_1115;
wire [5:0] u_ca_out_1116;
wire [5:0] u_ca_out_1117;
wire [5:0] u_ca_out_1118;
wire [5:0] u_ca_out_1119;
wire [5:0] u_ca_out_1120;
wire [5:0] u_ca_out_1121;
wire [5:0] u_ca_out_1122;
wire [5:0] u_ca_out_1123;
wire [5:0] u_ca_out_1124;
wire [5:0] u_ca_out_1125;
wire [5:0] u_ca_out_1126;
wire [5:0] u_ca_out_1127;
wire [5:0] u_ca_out_1128;
wire [5:0] u_ca_out_1129;
wire [5:0] u_ca_out_1130;
wire [5:0] u_ca_out_1131;
wire [5:0] u_ca_out_1132;
wire [5:0] u_ca_out_1133;
wire [5:0] u_ca_out_1134;
wire [5:0] u_ca_out_1135;
wire [5:0] u_ca_out_1136;
wire [5:0] u_ca_out_1137;
wire [5:0] u_ca_out_1138;
wire [5:0] u_ca_out_1139;
wire [5:0] u_ca_out_1140;
wire [5:0] u_ca_out_1141;
wire [5:0] u_ca_out_1142;
wire [5:0] u_ca_out_1143;
wire [5:0] u_ca_out_1144;
wire [5:0] u_ca_out_1145;
wire [5:0] u_ca_out_1146;
wire [5:0] u_ca_out_1147;
wire [5:0] u_ca_out_1148;
wire [5:0] u_ca_out_1149;
wire [5:0] u_ca_out_1150;
wire [5:0] u_ca_out_1151;
wire [5:0] u_ca_out_1152;
wire [5:0] u_ca_out_1153;
wire [5:0] u_ca_out_1154;
wire [5:0] u_ca_out_1155;
wire [5:0] u_ca_out_1156;
wire [5:0] u_ca_out_1157;
wire [5:0] u_ca_out_1158;
wire [5:0] u_ca_out_1159;
wire [5:0] u_ca_out_1160;
wire [5:0] u_ca_out_1161;
wire [5:0] u_ca_out_1162;
wire [5:0] u_ca_out_1163;
wire [5:0] u_ca_out_1164;
wire [5:0] u_ca_out_1165;
wire [5:0] u_ca_out_1166;
wire [5:0] u_ca_out_1167;
wire [5:0] u_ca_out_1168;
wire [5:0] u_ca_out_1169;
wire [5:0] u_ca_out_1170;
wire [5:0] u_ca_out_1171;
wire [5:0] u_ca_out_1172;
wire [5:0] u_ca_out_1173;
wire [5:0] u_ca_out_1174;
wire [5:0] u_ca_out_1175;
wire [5:0] u_ca_out_1176;
wire [5:0] u_ca_out_1177;
wire [5:0] u_ca_out_1178;
wire [5:0] u_ca_out_1179;
wire [5:0] u_ca_out_1180;
wire [5:0] u_ca_out_1181;
wire [5:0] u_ca_out_1182;
wire [5:0] u_ca_out_1183;
wire [5:0] u_ca_out_1184;
wire [5:0] u_ca_out_1185;
wire [5:0] u_ca_out_1186;
wire [5:0] u_ca_out_1187;
wire [5:0] u_ca_out_1188;
wire [5:0] u_ca_out_1189;
wire [5:0] u_ca_out_1190;
wire [5:0] u_ca_out_1191;
wire [5:0] u_ca_out_1192;
wire [5:0] u_ca_out_1193;
wire [5:0] u_ca_out_1194;
wire [5:0] u_ca_out_1195;
wire [5:0] u_ca_out_1196;
wire [5:0] u_ca_out_1197;
wire [5:0] u_ca_out_1198;
wire [5:0] u_ca_out_1199;
wire [5:0] u_ca_out_1200;
wire [5:0] u_ca_out_1201;
wire [5:0] u_ca_out_1202;
wire [5:0] u_ca_out_1203;
wire [5:0] u_ca_out_1204;
wire [5:0] u_ca_out_1205;
wire [5:0] u_ca_out_1206;
wire [5:0] u_ca_out_1207;
wire [5:0] u_ca_out_1208;
wire [5:0] u_ca_out_1209;
wire [5:0] u_ca_out_1210;
wire [5:0] u_ca_out_1211;
wire [5:0] u_ca_out_1212;
wire [5:0] u_ca_out_1213;
wire [5:0] u_ca_out_1214;
wire [5:0] u_ca_out_1215;
wire [5:0] u_ca_out_1216;
wire [5:0] u_ca_out_1217;
wire [5:0] u_ca_out_1218;
wire [5:0] u_ca_out_1219;
wire [5:0] u_ca_out_1220;
wire [5:0] u_ca_out_1221;
wire [5:0] u_ca_out_1222;
wire [5:0] u_ca_out_1223;
wire [5:0] u_ca_out_1224;
wire [5:0] u_ca_out_1225;
wire [5:0] u_ca_out_1226;
wire [5:0] u_ca_out_1227;
wire [5:0] u_ca_out_1228;
wire [5:0] u_ca_out_1229;
wire [5:0] u_ca_out_1230;
wire [5:0] u_ca_out_1231;
wire [5:0] u_ca_out_1232;
wire [5:0] u_ca_out_1233;
wire [5:0] u_ca_out_1234;
wire [5:0] u_ca_out_1235;
wire [5:0] u_ca_out_1236;
wire [5:0] u_ca_out_1237;
wire [5:0] u_ca_out_1238;
wire [5:0] u_ca_out_1239;
wire [5:0] u_ca_out_1240;
wire [5:0] u_ca_out_1241;
wire [5:0] u_ca_out_1242;
wire [5:0] u_ca_out_1243;
wire [5:0] u_ca_out_1244;
wire [5:0] u_ca_out_1245;
wire [5:0] u_ca_out_1246;
wire [5:0] u_ca_out_1247;
wire [5:0] u_ca_out_1248;
wire [5:0] u_ca_out_1249;
wire [5:0] u_ca_out_1250;
wire [5:0] u_ca_out_1251;
wire [5:0] u_ca_out_1252;
wire [5:0] u_ca_out_1253;
wire [5:0] u_ca_out_1254;
wire [5:0] u_ca_out_1255;
wire [5:0] u_ca_out_1256;
wire [5:0] u_ca_out_1257;
wire [5:0] u_ca_out_1258;
wire [5:0] u_ca_out_1259;
wire [5:0] u_ca_out_1260;
wire [5:0] u_ca_out_1261;
wire [5:0] u_ca_out_1262;
wire [5:0] u_ca_out_1263;
wire [5:0] u_ca_out_1264;
wire [5:0] u_ca_out_1265;
wire [5:0] u_ca_out_1266;
wire [5:0] u_ca_out_1267;
wire [5:0] u_ca_out_1268;
wire [5:0] u_ca_out_1269;
wire [5:0] u_ca_out_1270;
wire [5:0] u_ca_out_1271;
wire [5:0] u_ca_out_1272;
wire [5:0] u_ca_out_1273;
wire [5:0] u_ca_out_1274;
wire [5:0] u_ca_out_1275;
wire [5:0] u_ca_out_1276;
wire [5:0] u_ca_out_1277;
wire [5:0] u_ca_out_1278;
wire [5:0] u_ca_out_1279;
wire [5:0] u_ca_out_1280;
wire [5:0] u_ca_out_1281;
wire [5:0] u_ca_out_1282;
wire [5:0] u_ca_out_1283;
wire [5:0] u_ca_out_1284;
wire [5:0] u_ca_out_1285;
wire [5:0] u_ca_out_1286;
wire [5:0] u_ca_out_1287;

assign u_ca_in_0 = {{1{1'b0}}, col_in_0};
assign u_ca_in_1 = {{1{1'b0}}, col_in_1};
assign u_ca_in_2 = {{1{1'b0}}, col_in_2};
assign u_ca_in_3 = {{1{1'b0}}, col_in_3};
assign u_ca_in_4 = {{1{1'b0}}, col_in_4};
assign u_ca_in_5 = {{1{1'b0}}, col_in_5};
assign u_ca_in_6 = {{1{1'b0}}, col_in_6};
assign u_ca_in_7 = {{1{1'b0}}, col_in_7};
assign u_ca_in_8 = {{1{1'b0}}, col_in_8};
assign u_ca_in_9 = {{1{1'b0}}, col_in_9};
assign u_ca_in_10 = {{1{1'b0}}, col_in_10};
assign u_ca_in_11 = {{1{1'b0}}, col_in_11};
assign u_ca_in_12 = {{1{1'b0}}, col_in_12};
assign u_ca_in_13 = {{1{1'b0}}, col_in_13};
assign u_ca_in_14 = {{1{1'b0}}, col_in_14};
assign u_ca_in_15 = {{1{1'b0}}, col_in_15};
assign u_ca_in_16 = {{1{1'b0}}, col_in_16};
assign u_ca_in_17 = {{1{1'b0}}, col_in_17};
assign u_ca_in_18 = {{1{1'b0}}, col_in_18};
assign u_ca_in_19 = {{1{1'b0}}, col_in_19};
assign u_ca_in_20 = {{1{1'b0}}, col_in_20};
assign u_ca_in_21 = {{1{1'b0}}, col_in_21};
assign u_ca_in_22 = {{1{1'b0}}, col_in_22};
assign u_ca_in_23 = {{1{1'b0}}, col_in_23};
assign u_ca_in_24 = {{1{1'b0}}, col_in_24};
assign u_ca_in_25 = {{1{1'b0}}, col_in_25};
assign u_ca_in_26 = {{1{1'b0}}, col_in_26};
assign u_ca_in_27 = {{1{1'b0}}, col_in_27};
assign u_ca_in_28 = {{1{1'b0}}, col_in_28};
assign u_ca_in_29 = {{1{1'b0}}, col_in_29};
assign u_ca_in_30 = {{1{1'b0}}, col_in_30};
assign u_ca_in_31 = {{1{1'b0}}, col_in_31};
assign u_ca_in_32 = {{1{1'b0}}, col_in_32};
assign u_ca_in_33 = {{1{1'b0}}, col_in_33};
assign u_ca_in_34 = {{1{1'b0}}, col_in_34};
assign u_ca_in_35 = {{1{1'b0}}, col_in_35};
assign u_ca_in_36 = {{1{1'b0}}, col_in_36};
assign u_ca_in_37 = {{1{1'b0}}, col_in_37};
assign u_ca_in_38 = {{1{1'b0}}, col_in_38};
assign u_ca_in_39 = {{1{1'b0}}, col_in_39};
assign u_ca_in_40 = {{1{1'b0}}, col_in_40};
assign u_ca_in_41 = {{1{1'b0}}, col_in_41};
assign u_ca_in_42 = {{1{1'b0}}, col_in_42};
assign u_ca_in_43 = {{1{1'b0}}, col_in_43};
assign u_ca_in_44 = {{1{1'b0}}, col_in_44};
assign u_ca_in_45 = {{1{1'b0}}, col_in_45};
assign u_ca_in_46 = {{1{1'b0}}, col_in_46};
assign u_ca_in_47 = {{1{1'b0}}, col_in_47};
assign u_ca_in_48 = {{1{1'b0}}, col_in_48};
assign u_ca_in_49 = {{1{1'b0}}, col_in_49};
assign u_ca_in_50 = {{1{1'b0}}, col_in_50};
assign u_ca_in_51 = {{1{1'b0}}, col_in_51};
assign u_ca_in_52 = {{1{1'b0}}, col_in_52};
assign u_ca_in_53 = {{1{1'b0}}, col_in_53};
assign u_ca_in_54 = {{1{1'b0}}, col_in_54};
assign u_ca_in_55 = {{1{1'b0}}, col_in_55};
assign u_ca_in_56 = {{1{1'b0}}, col_in_56};
assign u_ca_in_57 = {{1{1'b0}}, col_in_57};
assign u_ca_in_58 = {{1{1'b0}}, col_in_58};
assign u_ca_in_59 = {{1{1'b0}}, col_in_59};
assign u_ca_in_60 = {{1{1'b0}}, col_in_60};
assign u_ca_in_61 = {{1{1'b0}}, col_in_61};
assign u_ca_in_62 = {{1{1'b0}}, col_in_62};
assign u_ca_in_63 = {{1{1'b0}}, col_in_63};
assign u_ca_in_64 = {{1{1'b0}}, col_in_64};
assign u_ca_in_65 = {{1{1'b0}}, col_in_65};
assign u_ca_in_66 = {{1{1'b0}}, col_in_66};
assign u_ca_in_67 = {{1{1'b0}}, col_in_67};
assign u_ca_in_68 = {{1{1'b0}}, col_in_68};
assign u_ca_in_69 = {{1{1'b0}}, col_in_69};
assign u_ca_in_70 = {{1{1'b0}}, col_in_70};
assign u_ca_in_71 = {{1{1'b0}}, col_in_71};
assign u_ca_in_72 = {{1{1'b0}}, col_in_72};
assign u_ca_in_73 = {{1{1'b0}}, col_in_73};
assign u_ca_in_74 = {{1{1'b0}}, col_in_74};
assign u_ca_in_75 = {{1{1'b0}}, col_in_75};
assign u_ca_in_76 = {{1{1'b0}}, col_in_76};
assign u_ca_in_77 = {{1{1'b0}}, col_in_77};
assign u_ca_in_78 = {{1{1'b0}}, col_in_78};
assign u_ca_in_79 = {{1{1'b0}}, col_in_79};
assign u_ca_in_80 = {{1{1'b0}}, col_in_80};
assign u_ca_in_81 = {{1{1'b0}}, col_in_81};
assign u_ca_in_82 = {{1{1'b0}}, col_in_82};
assign u_ca_in_83 = {{1{1'b0}}, col_in_83};
assign u_ca_in_84 = {{1{1'b0}}, col_in_84};
assign u_ca_in_85 = {{1{1'b0}}, col_in_85};
assign u_ca_in_86 = {{1{1'b0}}, col_in_86};
assign u_ca_in_87 = {{1{1'b0}}, col_in_87};
assign u_ca_in_88 = {{1{1'b0}}, col_in_88};
assign u_ca_in_89 = {{1{1'b0}}, col_in_89};
assign u_ca_in_90 = {{1{1'b0}}, col_in_90};
assign u_ca_in_91 = {{1{1'b0}}, col_in_91};
assign u_ca_in_92 = {{1{1'b0}}, col_in_92};
assign u_ca_in_93 = {{1{1'b0}}, col_in_93};
assign u_ca_in_94 = {{1{1'b0}}, col_in_94};
assign u_ca_in_95 = {{1{1'b0}}, col_in_95};
assign u_ca_in_96 = {{1{1'b0}}, col_in_96};
assign u_ca_in_97 = {{1{1'b0}}, col_in_97};
assign u_ca_in_98 = {{1{1'b0}}, col_in_98};
assign u_ca_in_99 = {{1{1'b0}}, col_in_99};
assign u_ca_in_100 = {{1{1'b0}}, col_in_100};
assign u_ca_in_101 = {{1{1'b0}}, col_in_101};
assign u_ca_in_102 = {{1{1'b0}}, col_in_102};
assign u_ca_in_103 = {{1{1'b0}}, col_in_103};
assign u_ca_in_104 = {{1{1'b0}}, col_in_104};
assign u_ca_in_105 = {{1{1'b0}}, col_in_105};
assign u_ca_in_106 = {{1{1'b0}}, col_in_106};
assign u_ca_in_107 = {{1{1'b0}}, col_in_107};
assign u_ca_in_108 = {{1{1'b0}}, col_in_108};
assign u_ca_in_109 = {{1{1'b0}}, col_in_109};
assign u_ca_in_110 = {{1{1'b0}}, col_in_110};
assign u_ca_in_111 = {{1{1'b0}}, col_in_111};
assign u_ca_in_112 = {{1{1'b0}}, col_in_112};
assign u_ca_in_113 = {{1{1'b0}}, col_in_113};
assign u_ca_in_114 = {{1{1'b0}}, col_in_114};
assign u_ca_in_115 = {{1{1'b0}}, col_in_115};
assign u_ca_in_116 = {{1{1'b0}}, col_in_116};
assign u_ca_in_117 = {{1{1'b0}}, col_in_117};
assign u_ca_in_118 = {{1{1'b0}}, col_in_118};
assign u_ca_in_119 = {{1{1'b0}}, col_in_119};
assign u_ca_in_120 = {{1{1'b0}}, col_in_120};
assign u_ca_in_121 = {{1{1'b0}}, col_in_121};
assign u_ca_in_122 = {{1{1'b0}}, col_in_122};
assign u_ca_in_123 = {{1{1'b0}}, col_in_123};
assign u_ca_in_124 = {{1{1'b0}}, col_in_124};
assign u_ca_in_125 = {{1{1'b0}}, col_in_125};
assign u_ca_in_126 = {{1{1'b0}}, col_in_126};
assign u_ca_in_127 = {{1{1'b0}}, col_in_127};
assign u_ca_in_128 = {{1{1'b0}}, col_in_128};
assign u_ca_in_129 = {{1{1'b0}}, col_in_129};
assign u_ca_in_130 = {{1{1'b0}}, col_in_130};
assign u_ca_in_131 = {{1{1'b0}}, col_in_131};
assign u_ca_in_132 = {{1{1'b0}}, col_in_132};
assign u_ca_in_133 = {{1{1'b0}}, col_in_133};
assign u_ca_in_134 = {{1{1'b0}}, col_in_134};
assign u_ca_in_135 = {{1{1'b0}}, col_in_135};
assign u_ca_in_136 = {{1{1'b0}}, col_in_136};
assign u_ca_in_137 = {{1{1'b0}}, col_in_137};
assign u_ca_in_138 = {{1{1'b0}}, col_in_138};
assign u_ca_in_139 = {{1{1'b0}}, col_in_139};
assign u_ca_in_140 = {{1{1'b0}}, col_in_140};
assign u_ca_in_141 = {{1{1'b0}}, col_in_141};
assign u_ca_in_142 = {{1{1'b0}}, col_in_142};
assign u_ca_in_143 = {{1{1'b0}}, col_in_143};
assign u_ca_in_144 = {{1{1'b0}}, col_in_144};
assign u_ca_in_145 = {{1{1'b0}}, col_in_145};
assign u_ca_in_146 = {{1{1'b0}}, col_in_146};
assign u_ca_in_147 = {{1{1'b0}}, col_in_147};
assign u_ca_in_148 = {{1{1'b0}}, col_in_148};
assign u_ca_in_149 = {{1{1'b0}}, col_in_149};
assign u_ca_in_150 = {{1{1'b0}}, col_in_150};
assign u_ca_in_151 = {{1{1'b0}}, col_in_151};
assign u_ca_in_152 = {{1{1'b0}}, col_in_152};
assign u_ca_in_153 = {{1{1'b0}}, col_in_153};
assign u_ca_in_154 = {{1{1'b0}}, col_in_154};
assign u_ca_in_155 = {{1{1'b0}}, col_in_155};
assign u_ca_in_156 = {{1{1'b0}}, col_in_156};
assign u_ca_in_157 = {{1{1'b0}}, col_in_157};
assign u_ca_in_158 = {{1{1'b0}}, col_in_158};
assign u_ca_in_159 = {{1{1'b0}}, col_in_159};
assign u_ca_in_160 = {{1{1'b0}}, col_in_160};
assign u_ca_in_161 = {{1{1'b0}}, col_in_161};
assign u_ca_in_162 = {{1{1'b0}}, col_in_162};
assign u_ca_in_163 = {{1{1'b0}}, col_in_163};
assign u_ca_in_164 = {{1{1'b0}}, col_in_164};
assign u_ca_in_165 = {{1{1'b0}}, col_in_165};
assign u_ca_in_166 = {{1{1'b0}}, col_in_166};
assign u_ca_in_167 = {{1{1'b0}}, col_in_167};
assign u_ca_in_168 = {{1{1'b0}}, col_in_168};
assign u_ca_in_169 = {{1{1'b0}}, col_in_169};
assign u_ca_in_170 = {{1{1'b0}}, col_in_170};
assign u_ca_in_171 = {{1{1'b0}}, col_in_171};
assign u_ca_in_172 = {{1{1'b0}}, col_in_172};
assign u_ca_in_173 = {{1{1'b0}}, col_in_173};
assign u_ca_in_174 = {{1{1'b0}}, col_in_174};
assign u_ca_in_175 = {{1{1'b0}}, col_in_175};
assign u_ca_in_176 = {{1{1'b0}}, col_in_176};
assign u_ca_in_177 = {{1{1'b0}}, col_in_177};
assign u_ca_in_178 = {{1{1'b0}}, col_in_178};
assign u_ca_in_179 = {{1{1'b0}}, col_in_179};
assign u_ca_in_180 = {{1{1'b0}}, col_in_180};
assign u_ca_in_181 = {{1{1'b0}}, col_in_181};
assign u_ca_in_182 = {{1{1'b0}}, col_in_182};
assign u_ca_in_183 = {{1{1'b0}}, col_in_183};
assign u_ca_in_184 = {{1{1'b0}}, col_in_184};
assign u_ca_in_185 = {{1{1'b0}}, col_in_185};
assign u_ca_in_186 = {{1{1'b0}}, col_in_186};
assign u_ca_in_187 = {{1{1'b0}}, col_in_187};
assign u_ca_in_188 = {{1{1'b0}}, col_in_188};
assign u_ca_in_189 = {{1{1'b0}}, col_in_189};
assign u_ca_in_190 = {{1{1'b0}}, col_in_190};
assign u_ca_in_191 = {{1{1'b0}}, col_in_191};
assign u_ca_in_192 = {{1{1'b0}}, col_in_192};
assign u_ca_in_193 = {{1{1'b0}}, col_in_193};
assign u_ca_in_194 = {{1{1'b0}}, col_in_194};
assign u_ca_in_195 = {{1{1'b0}}, col_in_195};
assign u_ca_in_196 = {{1{1'b0}}, col_in_196};
assign u_ca_in_197 = {{1{1'b0}}, col_in_197};
assign u_ca_in_198 = {{1{1'b0}}, col_in_198};
assign u_ca_in_199 = {{1{1'b0}}, col_in_199};
assign u_ca_in_200 = {{1{1'b0}}, col_in_200};
assign u_ca_in_201 = {{1{1'b0}}, col_in_201};
assign u_ca_in_202 = {{1{1'b0}}, col_in_202};
assign u_ca_in_203 = {{1{1'b0}}, col_in_203};
assign u_ca_in_204 = {{1{1'b0}}, col_in_204};
assign u_ca_in_205 = {{1{1'b0}}, col_in_205};
assign u_ca_in_206 = {{1{1'b0}}, col_in_206};
assign u_ca_in_207 = {{1{1'b0}}, col_in_207};
assign u_ca_in_208 = {{1{1'b0}}, col_in_208};
assign u_ca_in_209 = {{1{1'b0}}, col_in_209};
assign u_ca_in_210 = {{1{1'b0}}, col_in_210};
assign u_ca_in_211 = {{1{1'b0}}, col_in_211};
assign u_ca_in_212 = {{1{1'b0}}, col_in_212};
assign u_ca_in_213 = {{1{1'b0}}, col_in_213};
assign u_ca_in_214 = {{1{1'b0}}, col_in_214};
assign u_ca_in_215 = {{1{1'b0}}, col_in_215};
assign u_ca_in_216 = {{1{1'b0}}, col_in_216};
assign u_ca_in_217 = {{1{1'b0}}, col_in_217};
assign u_ca_in_218 = {{1{1'b0}}, col_in_218};
assign u_ca_in_219 = {{1{1'b0}}, col_in_219};
assign u_ca_in_220 = {{1{1'b0}}, col_in_220};
assign u_ca_in_221 = {{1{1'b0}}, col_in_221};
assign u_ca_in_222 = {{1{1'b0}}, col_in_222};
assign u_ca_in_223 = {{1{1'b0}}, col_in_223};
assign u_ca_in_224 = {{1{1'b0}}, col_in_224};
assign u_ca_in_225 = {{1{1'b0}}, col_in_225};
assign u_ca_in_226 = {{1{1'b0}}, col_in_226};
assign u_ca_in_227 = {{1{1'b0}}, col_in_227};
assign u_ca_in_228 = {{1{1'b0}}, col_in_228};
assign u_ca_in_229 = {{1{1'b0}}, col_in_229};
assign u_ca_in_230 = {{1{1'b0}}, col_in_230};
assign u_ca_in_231 = {{1{1'b0}}, col_in_231};
assign u_ca_in_232 = {{1{1'b0}}, col_in_232};
assign u_ca_in_233 = {{1{1'b0}}, col_in_233};
assign u_ca_in_234 = {{1{1'b0}}, col_in_234};
assign u_ca_in_235 = {{1{1'b0}}, col_in_235};
assign u_ca_in_236 = {{1{1'b0}}, col_in_236};
assign u_ca_in_237 = {{1{1'b0}}, col_in_237};
assign u_ca_in_238 = {{1{1'b0}}, col_in_238};
assign u_ca_in_239 = {{1{1'b0}}, col_in_239};
assign u_ca_in_240 = {{1{1'b0}}, col_in_240};
assign u_ca_in_241 = {{1{1'b0}}, col_in_241};
assign u_ca_in_242 = {{1{1'b0}}, col_in_242};
assign u_ca_in_243 = {{1{1'b0}}, col_in_243};
assign u_ca_in_244 = {{1{1'b0}}, col_in_244};
assign u_ca_in_245 = {{1{1'b0}}, col_in_245};
assign u_ca_in_246 = {{1{1'b0}}, col_in_246};
assign u_ca_in_247 = {{1{1'b0}}, col_in_247};
assign u_ca_in_248 = {{1{1'b0}}, col_in_248};
assign u_ca_in_249 = {{1{1'b0}}, col_in_249};
assign u_ca_in_250 = {{1{1'b0}}, col_in_250};
assign u_ca_in_251 = {{1{1'b0}}, col_in_251};
assign u_ca_in_252 = {{1{1'b0}}, col_in_252};
assign u_ca_in_253 = {{1{1'b0}}, col_in_253};
assign u_ca_in_254 = {{1{1'b0}}, col_in_254};
assign u_ca_in_255 = {{1{1'b0}}, col_in_255};
assign u_ca_in_256 = {{1{1'b0}}, col_in_256};
assign u_ca_in_257 = {{1{1'b0}}, col_in_257};
assign u_ca_in_258 = {{1{1'b0}}, col_in_258};
assign u_ca_in_259 = {{1{1'b0}}, col_in_259};
assign u_ca_in_260 = {{1{1'b0}}, col_in_260};
assign u_ca_in_261 = {{1{1'b0}}, col_in_261};
assign u_ca_in_262 = {{1{1'b0}}, col_in_262};
assign u_ca_in_263 = {{1{1'b0}}, col_in_263};
assign u_ca_in_264 = {{1{1'b0}}, col_in_264};
assign u_ca_in_265 = {{1{1'b0}}, col_in_265};
assign u_ca_in_266 = {{1{1'b0}}, col_in_266};
assign u_ca_in_267 = {{1{1'b0}}, col_in_267};
assign u_ca_in_268 = {{1{1'b0}}, col_in_268};
assign u_ca_in_269 = {{1{1'b0}}, col_in_269};
assign u_ca_in_270 = {{1{1'b0}}, col_in_270};
assign u_ca_in_271 = {{1{1'b0}}, col_in_271};
assign u_ca_in_272 = {{1{1'b0}}, col_in_272};
assign u_ca_in_273 = {{1{1'b0}}, col_in_273};
assign u_ca_in_274 = {{1{1'b0}}, col_in_274};
assign u_ca_in_275 = {{1{1'b0}}, col_in_275};
assign u_ca_in_276 = {{1{1'b0}}, col_in_276};
assign u_ca_in_277 = {{1{1'b0}}, col_in_277};
assign u_ca_in_278 = {{1{1'b0}}, col_in_278};
assign u_ca_in_279 = {{1{1'b0}}, col_in_279};
assign u_ca_in_280 = {{1{1'b0}}, col_in_280};
assign u_ca_in_281 = {{1{1'b0}}, col_in_281};
assign u_ca_in_282 = {{1{1'b0}}, col_in_282};
assign u_ca_in_283 = {{1{1'b0}}, col_in_283};
assign u_ca_in_284 = {{1{1'b0}}, col_in_284};
assign u_ca_in_285 = {{1{1'b0}}, col_in_285};
assign u_ca_in_286 = {{1{1'b0}}, col_in_286};
assign u_ca_in_287 = {{1{1'b0}}, col_in_287};
assign u_ca_in_288 = {{1{1'b0}}, col_in_288};
assign u_ca_in_289 = {{1{1'b0}}, col_in_289};
assign u_ca_in_290 = {{1{1'b0}}, col_in_290};
assign u_ca_in_291 = {{1{1'b0}}, col_in_291};
assign u_ca_in_292 = {{1{1'b0}}, col_in_292};
assign u_ca_in_293 = {{1{1'b0}}, col_in_293};
assign u_ca_in_294 = {{1{1'b0}}, col_in_294};
assign u_ca_in_295 = {{1{1'b0}}, col_in_295};
assign u_ca_in_296 = {{1{1'b0}}, col_in_296};
assign u_ca_in_297 = {{1{1'b0}}, col_in_297};
assign u_ca_in_298 = {{1{1'b0}}, col_in_298};
assign u_ca_in_299 = {{1{1'b0}}, col_in_299};
assign u_ca_in_300 = {{1{1'b0}}, col_in_300};
assign u_ca_in_301 = {{1{1'b0}}, col_in_301};
assign u_ca_in_302 = {{1{1'b0}}, col_in_302};
assign u_ca_in_303 = {{1{1'b0}}, col_in_303};
assign u_ca_in_304 = {{1{1'b0}}, col_in_304};
assign u_ca_in_305 = {{1{1'b0}}, col_in_305};
assign u_ca_in_306 = {{1{1'b0}}, col_in_306};
assign u_ca_in_307 = {{1{1'b0}}, col_in_307};
assign u_ca_in_308 = {{1{1'b0}}, col_in_308};
assign u_ca_in_309 = {{1{1'b0}}, col_in_309};
assign u_ca_in_310 = {{1{1'b0}}, col_in_310};
assign u_ca_in_311 = {{1{1'b0}}, col_in_311};
assign u_ca_in_312 = {{1{1'b0}}, col_in_312};
assign u_ca_in_313 = {{1{1'b0}}, col_in_313};
assign u_ca_in_314 = {{1{1'b0}}, col_in_314};
assign u_ca_in_315 = {{1{1'b0}}, col_in_315};
assign u_ca_in_316 = {{1{1'b0}}, col_in_316};
assign u_ca_in_317 = {{1{1'b0}}, col_in_317};
assign u_ca_in_318 = {{1{1'b0}}, col_in_318};
assign u_ca_in_319 = {{1{1'b0}}, col_in_319};
assign u_ca_in_320 = {{1{1'b0}}, col_in_320};
assign u_ca_in_321 = {{1{1'b0}}, col_in_321};
assign u_ca_in_322 = {{1{1'b0}}, col_in_322};
assign u_ca_in_323 = {{1{1'b0}}, col_in_323};
assign u_ca_in_324 = {{1{1'b0}}, col_in_324};
assign u_ca_in_325 = {{1{1'b0}}, col_in_325};
assign u_ca_in_326 = {{1{1'b0}}, col_in_326};
assign u_ca_in_327 = {{1{1'b0}}, col_in_327};
assign u_ca_in_328 = {{1{1'b0}}, col_in_328};
assign u_ca_in_329 = {{1{1'b0}}, col_in_329};
assign u_ca_in_330 = {{1{1'b0}}, col_in_330};
assign u_ca_in_331 = {{1{1'b0}}, col_in_331};
assign u_ca_in_332 = {{1{1'b0}}, col_in_332};
assign u_ca_in_333 = {{1{1'b0}}, col_in_333};
assign u_ca_in_334 = {{1{1'b0}}, col_in_334};
assign u_ca_in_335 = {{1{1'b0}}, col_in_335};
assign u_ca_in_336 = {{1{1'b0}}, col_in_336};
assign u_ca_in_337 = {{1{1'b0}}, col_in_337};
assign u_ca_in_338 = {{1{1'b0}}, col_in_338};
assign u_ca_in_339 = {{1{1'b0}}, col_in_339};
assign u_ca_in_340 = {{1{1'b0}}, col_in_340};
assign u_ca_in_341 = {{1{1'b0}}, col_in_341};
assign u_ca_in_342 = {{1{1'b0}}, col_in_342};
assign u_ca_in_343 = {{1{1'b0}}, col_in_343};
assign u_ca_in_344 = {{1{1'b0}}, col_in_344};
assign u_ca_in_345 = {{1{1'b0}}, col_in_345};
assign u_ca_in_346 = {{1{1'b0}}, col_in_346};
assign u_ca_in_347 = {{1{1'b0}}, col_in_347};
assign u_ca_in_348 = {{1{1'b0}}, col_in_348};
assign u_ca_in_349 = {{1{1'b0}}, col_in_349};
assign u_ca_in_350 = {{1{1'b0}}, col_in_350};
assign u_ca_in_351 = {{1{1'b0}}, col_in_351};
assign u_ca_in_352 = {{1{1'b0}}, col_in_352};
assign u_ca_in_353 = {{1{1'b0}}, col_in_353};
assign u_ca_in_354 = {{1{1'b0}}, col_in_354};
assign u_ca_in_355 = {{1{1'b0}}, col_in_355};
assign u_ca_in_356 = {{1{1'b0}}, col_in_356};
assign u_ca_in_357 = {{1{1'b0}}, col_in_357};
assign u_ca_in_358 = {{1{1'b0}}, col_in_358};
assign u_ca_in_359 = {{1{1'b0}}, col_in_359};
assign u_ca_in_360 = {{1{1'b0}}, col_in_360};
assign u_ca_in_361 = {{1{1'b0}}, col_in_361};
assign u_ca_in_362 = {{1{1'b0}}, col_in_362};
assign u_ca_in_363 = {{1{1'b0}}, col_in_363};
assign u_ca_in_364 = {{1{1'b0}}, col_in_364};
assign u_ca_in_365 = {{1{1'b0}}, col_in_365};
assign u_ca_in_366 = {{1{1'b0}}, col_in_366};
assign u_ca_in_367 = {{1{1'b0}}, col_in_367};
assign u_ca_in_368 = {{1{1'b0}}, col_in_368};
assign u_ca_in_369 = {{1{1'b0}}, col_in_369};
assign u_ca_in_370 = {{1{1'b0}}, col_in_370};
assign u_ca_in_371 = {{1{1'b0}}, col_in_371};
assign u_ca_in_372 = {{1{1'b0}}, col_in_372};
assign u_ca_in_373 = {{1{1'b0}}, col_in_373};
assign u_ca_in_374 = {{1{1'b0}}, col_in_374};
assign u_ca_in_375 = {{1{1'b0}}, col_in_375};
assign u_ca_in_376 = {{1{1'b0}}, col_in_376};
assign u_ca_in_377 = {{1{1'b0}}, col_in_377};
assign u_ca_in_378 = {{1{1'b0}}, col_in_378};
assign u_ca_in_379 = {{1{1'b0}}, col_in_379};
assign u_ca_in_380 = {{1{1'b0}}, col_in_380};
assign u_ca_in_381 = {{1{1'b0}}, col_in_381};
assign u_ca_in_382 = {{1{1'b0}}, col_in_382};
assign u_ca_in_383 = {{1{1'b0}}, col_in_383};
assign u_ca_in_384 = {{1{1'b0}}, col_in_384};
assign u_ca_in_385 = {{1{1'b0}}, col_in_385};
assign u_ca_in_386 = {{1{1'b0}}, col_in_386};
assign u_ca_in_387 = {{1{1'b0}}, col_in_387};
assign u_ca_in_388 = {{1{1'b0}}, col_in_388};
assign u_ca_in_389 = {{1{1'b0}}, col_in_389};
assign u_ca_in_390 = {{1{1'b0}}, col_in_390};
assign u_ca_in_391 = {{1{1'b0}}, col_in_391};
assign u_ca_in_392 = {{1{1'b0}}, col_in_392};
assign u_ca_in_393 = {{1{1'b0}}, col_in_393};
assign u_ca_in_394 = {{1{1'b0}}, col_in_394};
assign u_ca_in_395 = {{1{1'b0}}, col_in_395};
assign u_ca_in_396 = {{1{1'b0}}, col_in_396};
assign u_ca_in_397 = {{1{1'b0}}, col_in_397};
assign u_ca_in_398 = {{1{1'b0}}, col_in_398};
assign u_ca_in_399 = {{1{1'b0}}, col_in_399};
assign u_ca_in_400 = {{1{1'b0}}, col_in_400};
assign u_ca_in_401 = {{1{1'b0}}, col_in_401};
assign u_ca_in_402 = {{1{1'b0}}, col_in_402};
assign u_ca_in_403 = {{1{1'b0}}, col_in_403};
assign u_ca_in_404 = {{1{1'b0}}, col_in_404};
assign u_ca_in_405 = {{1{1'b0}}, col_in_405};
assign u_ca_in_406 = {{1{1'b0}}, col_in_406};
assign u_ca_in_407 = {{1{1'b0}}, col_in_407};
assign u_ca_in_408 = {{1{1'b0}}, col_in_408};
assign u_ca_in_409 = {{1{1'b0}}, col_in_409};
assign u_ca_in_410 = {{1{1'b0}}, col_in_410};
assign u_ca_in_411 = {{1{1'b0}}, col_in_411};
assign u_ca_in_412 = {{1{1'b0}}, col_in_412};
assign u_ca_in_413 = {{1{1'b0}}, col_in_413};
assign u_ca_in_414 = {{1{1'b0}}, col_in_414};
assign u_ca_in_415 = {{1{1'b0}}, col_in_415};
assign u_ca_in_416 = {{1{1'b0}}, col_in_416};
assign u_ca_in_417 = {{1{1'b0}}, col_in_417};
assign u_ca_in_418 = {{1{1'b0}}, col_in_418};
assign u_ca_in_419 = {{1{1'b0}}, col_in_419};
assign u_ca_in_420 = {{1{1'b0}}, col_in_420};
assign u_ca_in_421 = {{1{1'b0}}, col_in_421};
assign u_ca_in_422 = {{1{1'b0}}, col_in_422};
assign u_ca_in_423 = {{1{1'b0}}, col_in_423};
assign u_ca_in_424 = {{1{1'b0}}, col_in_424};
assign u_ca_in_425 = {{1{1'b0}}, col_in_425};
assign u_ca_in_426 = {{1{1'b0}}, col_in_426};
assign u_ca_in_427 = {{1{1'b0}}, col_in_427};
assign u_ca_in_428 = {{1{1'b0}}, col_in_428};
assign u_ca_in_429 = {{1{1'b0}}, col_in_429};
assign u_ca_in_430 = {{1{1'b0}}, col_in_430};
assign u_ca_in_431 = {{1{1'b0}}, col_in_431};
assign u_ca_in_432 = {{1{1'b0}}, col_in_432};
assign u_ca_in_433 = {{1{1'b0}}, col_in_433};
assign u_ca_in_434 = {{1{1'b0}}, col_in_434};
assign u_ca_in_435 = {{1{1'b0}}, col_in_435};
assign u_ca_in_436 = {{1{1'b0}}, col_in_436};
assign u_ca_in_437 = {{1{1'b0}}, col_in_437};
assign u_ca_in_438 = {{1{1'b0}}, col_in_438};
assign u_ca_in_439 = {{1{1'b0}}, col_in_439};
assign u_ca_in_440 = {{1{1'b0}}, col_in_440};
assign u_ca_in_441 = {{1{1'b0}}, col_in_441};
assign u_ca_in_442 = {{1{1'b0}}, col_in_442};
assign u_ca_in_443 = {{1{1'b0}}, col_in_443};
assign u_ca_in_444 = {{1{1'b0}}, col_in_444};
assign u_ca_in_445 = {{1{1'b0}}, col_in_445};
assign u_ca_in_446 = {{1{1'b0}}, col_in_446};
assign u_ca_in_447 = {{1{1'b0}}, col_in_447};
assign u_ca_in_448 = {{1{1'b0}}, col_in_448};
assign u_ca_in_449 = {{1{1'b0}}, col_in_449};
assign u_ca_in_450 = {{1{1'b0}}, col_in_450};
assign u_ca_in_451 = {{1{1'b0}}, col_in_451};
assign u_ca_in_452 = {{1{1'b0}}, col_in_452};
assign u_ca_in_453 = {{1{1'b0}}, col_in_453};
assign u_ca_in_454 = {{1{1'b0}}, col_in_454};
assign u_ca_in_455 = {{1{1'b0}}, col_in_455};
assign u_ca_in_456 = {{1{1'b0}}, col_in_456};
assign u_ca_in_457 = {{1{1'b0}}, col_in_457};
assign u_ca_in_458 = {{1{1'b0}}, col_in_458};
assign u_ca_in_459 = {{1{1'b0}}, col_in_459};
assign u_ca_in_460 = {{1{1'b0}}, col_in_460};
assign u_ca_in_461 = {{1{1'b0}}, col_in_461};
assign u_ca_in_462 = {{1{1'b0}}, col_in_462};
assign u_ca_in_463 = {{1{1'b0}}, col_in_463};
assign u_ca_in_464 = {{1{1'b0}}, col_in_464};
assign u_ca_in_465 = {{1{1'b0}}, col_in_465};
assign u_ca_in_466 = {{1{1'b0}}, col_in_466};
assign u_ca_in_467 = {{1{1'b0}}, col_in_467};
assign u_ca_in_468 = {{1{1'b0}}, col_in_468};
assign u_ca_in_469 = {{1{1'b0}}, col_in_469};
assign u_ca_in_470 = {{1{1'b0}}, col_in_470};
assign u_ca_in_471 = {{1{1'b0}}, col_in_471};
assign u_ca_in_472 = {{1{1'b0}}, col_in_472};
assign u_ca_in_473 = {{1{1'b0}}, col_in_473};
assign u_ca_in_474 = {{1{1'b0}}, col_in_474};
assign u_ca_in_475 = {{1{1'b0}}, col_in_475};
assign u_ca_in_476 = {{1{1'b0}}, col_in_476};
assign u_ca_in_477 = {{1{1'b0}}, col_in_477};
assign u_ca_in_478 = {{1{1'b0}}, col_in_478};
assign u_ca_in_479 = {{1{1'b0}}, col_in_479};
assign u_ca_in_480 = {{1{1'b0}}, col_in_480};
assign u_ca_in_481 = {{1{1'b0}}, col_in_481};
assign u_ca_in_482 = {{1{1'b0}}, col_in_482};
assign u_ca_in_483 = {{1{1'b0}}, col_in_483};
assign u_ca_in_484 = {{1{1'b0}}, col_in_484};
assign u_ca_in_485 = {{1{1'b0}}, col_in_485};
assign u_ca_in_486 = {{1{1'b0}}, col_in_486};
assign u_ca_in_487 = {{1{1'b0}}, col_in_487};
assign u_ca_in_488 = {{1{1'b0}}, col_in_488};
assign u_ca_in_489 = {{1{1'b0}}, col_in_489};
assign u_ca_in_490 = {{1{1'b0}}, col_in_490};
assign u_ca_in_491 = {{1{1'b0}}, col_in_491};
assign u_ca_in_492 = {{1{1'b0}}, col_in_492};
assign u_ca_in_493 = {{1{1'b0}}, col_in_493};
assign u_ca_in_494 = {{1{1'b0}}, col_in_494};
assign u_ca_in_495 = {{1{1'b0}}, col_in_495};
assign u_ca_in_496 = {{1{1'b0}}, col_in_496};
assign u_ca_in_497 = {{1{1'b0}}, col_in_497};
assign u_ca_in_498 = {{1{1'b0}}, col_in_498};
assign u_ca_in_499 = {{1{1'b0}}, col_in_499};
assign u_ca_in_500 = {{1{1'b0}}, col_in_500};
assign u_ca_in_501 = {{1{1'b0}}, col_in_501};
assign u_ca_in_502 = {{1{1'b0}}, col_in_502};
assign u_ca_in_503 = {{1{1'b0}}, col_in_503};
assign u_ca_in_504 = {{1{1'b0}}, col_in_504};
assign u_ca_in_505 = {{1{1'b0}}, col_in_505};
assign u_ca_in_506 = {{1{1'b0}}, col_in_506};
assign u_ca_in_507 = {{1{1'b0}}, col_in_507};
assign u_ca_in_508 = {{1{1'b0}}, col_in_508};
assign u_ca_in_509 = {{1{1'b0}}, col_in_509};
assign u_ca_in_510 = {{1{1'b0}}, col_in_510};
assign u_ca_in_511 = {{1{1'b0}}, col_in_511};
assign u_ca_in_512 = {{1{1'b0}}, col_in_512};
assign u_ca_in_513 = {{1{1'b0}}, col_in_513};
assign u_ca_in_514 = {{1{1'b0}}, col_in_514};
assign u_ca_in_515 = {{1{1'b0}}, col_in_515};
assign u_ca_in_516 = {{1{1'b0}}, col_in_516};
assign u_ca_in_517 = {{1{1'b0}}, col_in_517};
assign u_ca_in_518 = {{1{1'b0}}, col_in_518};
assign u_ca_in_519 = {{1{1'b0}}, col_in_519};
assign u_ca_in_520 = {{1{1'b0}}, col_in_520};
assign u_ca_in_521 = {{1{1'b0}}, col_in_521};
assign u_ca_in_522 = {{1{1'b0}}, col_in_522};
assign u_ca_in_523 = {{1{1'b0}}, col_in_523};
assign u_ca_in_524 = {{1{1'b0}}, col_in_524};
assign u_ca_in_525 = {{1{1'b0}}, col_in_525};
assign u_ca_in_526 = {{1{1'b0}}, col_in_526};
assign u_ca_in_527 = {{1{1'b0}}, col_in_527};
assign u_ca_in_528 = {{1{1'b0}}, col_in_528};
assign u_ca_in_529 = {{1{1'b0}}, col_in_529};
assign u_ca_in_530 = {{1{1'b0}}, col_in_530};
assign u_ca_in_531 = {{1{1'b0}}, col_in_531};
assign u_ca_in_532 = {{1{1'b0}}, col_in_532};
assign u_ca_in_533 = {{1{1'b0}}, col_in_533};
assign u_ca_in_534 = {{1{1'b0}}, col_in_534};
assign u_ca_in_535 = {{1{1'b0}}, col_in_535};
assign u_ca_in_536 = {{1{1'b0}}, col_in_536};
assign u_ca_in_537 = {{1{1'b0}}, col_in_537};
assign u_ca_in_538 = {{1{1'b0}}, col_in_538};
assign u_ca_in_539 = {{1{1'b0}}, col_in_539};
assign u_ca_in_540 = {{1{1'b0}}, col_in_540};
assign u_ca_in_541 = {{1{1'b0}}, col_in_541};
assign u_ca_in_542 = {{1{1'b0}}, col_in_542};
assign u_ca_in_543 = {{1{1'b0}}, col_in_543};
assign u_ca_in_544 = {{1{1'b0}}, col_in_544};
assign u_ca_in_545 = {{1{1'b0}}, col_in_545};
assign u_ca_in_546 = {{1{1'b0}}, col_in_546};
assign u_ca_in_547 = {{1{1'b0}}, col_in_547};
assign u_ca_in_548 = {{1{1'b0}}, col_in_548};
assign u_ca_in_549 = {{1{1'b0}}, col_in_549};
assign u_ca_in_550 = {{1{1'b0}}, col_in_550};
assign u_ca_in_551 = {{1{1'b0}}, col_in_551};
assign u_ca_in_552 = {{1{1'b0}}, col_in_552};
assign u_ca_in_553 = {{1{1'b0}}, col_in_553};
assign u_ca_in_554 = {{1{1'b0}}, col_in_554};
assign u_ca_in_555 = {{1{1'b0}}, col_in_555};
assign u_ca_in_556 = {{1{1'b0}}, col_in_556};
assign u_ca_in_557 = {{1{1'b0}}, col_in_557};
assign u_ca_in_558 = {{1{1'b0}}, col_in_558};
assign u_ca_in_559 = {{1{1'b0}}, col_in_559};
assign u_ca_in_560 = {{1{1'b0}}, col_in_560};
assign u_ca_in_561 = {{1{1'b0}}, col_in_561};
assign u_ca_in_562 = {{1{1'b0}}, col_in_562};
assign u_ca_in_563 = {{1{1'b0}}, col_in_563};
assign u_ca_in_564 = {{1{1'b0}}, col_in_564};
assign u_ca_in_565 = {{1{1'b0}}, col_in_565};
assign u_ca_in_566 = {{1{1'b0}}, col_in_566};
assign u_ca_in_567 = {{1{1'b0}}, col_in_567};
assign u_ca_in_568 = {{1{1'b0}}, col_in_568};
assign u_ca_in_569 = {{1{1'b0}}, col_in_569};
assign u_ca_in_570 = {{1{1'b0}}, col_in_570};
assign u_ca_in_571 = {{1{1'b0}}, col_in_571};
assign u_ca_in_572 = {{1{1'b0}}, col_in_572};
assign u_ca_in_573 = {{1{1'b0}}, col_in_573};
assign u_ca_in_574 = {{1{1'b0}}, col_in_574};
assign u_ca_in_575 = {{1{1'b0}}, col_in_575};
assign u_ca_in_576 = {{1{1'b0}}, col_in_576};
assign u_ca_in_577 = {{1{1'b0}}, col_in_577};
assign u_ca_in_578 = {{1{1'b0}}, col_in_578};
assign u_ca_in_579 = {{1{1'b0}}, col_in_579};
assign u_ca_in_580 = {{1{1'b0}}, col_in_580};
assign u_ca_in_581 = {{1{1'b0}}, col_in_581};
assign u_ca_in_582 = {{1{1'b0}}, col_in_582};
assign u_ca_in_583 = {{1{1'b0}}, col_in_583};
assign u_ca_in_584 = {{1{1'b0}}, col_in_584};
assign u_ca_in_585 = {{1{1'b0}}, col_in_585};
assign u_ca_in_586 = {{1{1'b0}}, col_in_586};
assign u_ca_in_587 = {{1{1'b0}}, col_in_587};
assign u_ca_in_588 = {{1{1'b0}}, col_in_588};
assign u_ca_in_589 = {{1{1'b0}}, col_in_589};
assign u_ca_in_590 = {{1{1'b0}}, col_in_590};
assign u_ca_in_591 = {{1{1'b0}}, col_in_591};
assign u_ca_in_592 = {{1{1'b0}}, col_in_592};
assign u_ca_in_593 = {{1{1'b0}}, col_in_593};
assign u_ca_in_594 = {{1{1'b0}}, col_in_594};
assign u_ca_in_595 = {{1{1'b0}}, col_in_595};
assign u_ca_in_596 = {{1{1'b0}}, col_in_596};
assign u_ca_in_597 = {{1{1'b0}}, col_in_597};
assign u_ca_in_598 = {{1{1'b0}}, col_in_598};
assign u_ca_in_599 = {{1{1'b0}}, col_in_599};
assign u_ca_in_600 = {{1{1'b0}}, col_in_600};
assign u_ca_in_601 = {{1{1'b0}}, col_in_601};
assign u_ca_in_602 = {{1{1'b0}}, col_in_602};
assign u_ca_in_603 = {{1{1'b0}}, col_in_603};
assign u_ca_in_604 = {{1{1'b0}}, col_in_604};
assign u_ca_in_605 = {{1{1'b0}}, col_in_605};
assign u_ca_in_606 = {{1{1'b0}}, col_in_606};
assign u_ca_in_607 = {{1{1'b0}}, col_in_607};
assign u_ca_in_608 = {{1{1'b0}}, col_in_608};
assign u_ca_in_609 = {{1{1'b0}}, col_in_609};
assign u_ca_in_610 = {{1{1'b0}}, col_in_610};
assign u_ca_in_611 = {{1{1'b0}}, col_in_611};
assign u_ca_in_612 = {{1{1'b0}}, col_in_612};
assign u_ca_in_613 = {{1{1'b0}}, col_in_613};
assign u_ca_in_614 = {{1{1'b0}}, col_in_614};
assign u_ca_in_615 = {{1{1'b0}}, col_in_615};
assign u_ca_in_616 = {{1{1'b0}}, col_in_616};
assign u_ca_in_617 = {{1{1'b0}}, col_in_617};
assign u_ca_in_618 = {{1{1'b0}}, col_in_618};
assign u_ca_in_619 = {{1{1'b0}}, col_in_619};
assign u_ca_in_620 = {{1{1'b0}}, col_in_620};
assign u_ca_in_621 = {{1{1'b0}}, col_in_621};
assign u_ca_in_622 = {{1{1'b0}}, col_in_622};
assign u_ca_in_623 = {{1{1'b0}}, col_in_623};
assign u_ca_in_624 = {{1{1'b0}}, col_in_624};
assign u_ca_in_625 = {{1{1'b0}}, col_in_625};
assign u_ca_in_626 = {{1{1'b0}}, col_in_626};
assign u_ca_in_627 = {{1{1'b0}}, col_in_627};
assign u_ca_in_628 = {{1{1'b0}}, col_in_628};
assign u_ca_in_629 = {{1{1'b0}}, col_in_629};
assign u_ca_in_630 = {{1{1'b0}}, col_in_630};
assign u_ca_in_631 = {{1{1'b0}}, col_in_631};
assign u_ca_in_632 = {{1{1'b0}}, col_in_632};
assign u_ca_in_633 = {{1{1'b0}}, col_in_633};
assign u_ca_in_634 = {{1{1'b0}}, col_in_634};
assign u_ca_in_635 = {{1{1'b0}}, col_in_635};
assign u_ca_in_636 = {{1{1'b0}}, col_in_636};
assign u_ca_in_637 = {{1{1'b0}}, col_in_637};
assign u_ca_in_638 = {{1{1'b0}}, col_in_638};
assign u_ca_in_639 = {{1{1'b0}}, col_in_639};
assign u_ca_in_640 = {{1{1'b0}}, col_in_640};
assign u_ca_in_641 = {{1{1'b0}}, col_in_641};
assign u_ca_in_642 = {{1{1'b0}}, col_in_642};
assign u_ca_in_643 = {{1{1'b0}}, col_in_643};
assign u_ca_in_644 = {{1{1'b0}}, col_in_644};
assign u_ca_in_645 = {{1{1'b0}}, col_in_645};
assign u_ca_in_646 = {{1{1'b0}}, col_in_646};
assign u_ca_in_647 = {{1{1'b0}}, col_in_647};
assign u_ca_in_648 = {{1{1'b0}}, col_in_648};
assign u_ca_in_649 = {{1{1'b0}}, col_in_649};
assign u_ca_in_650 = {{1{1'b0}}, col_in_650};
assign u_ca_in_651 = {{1{1'b0}}, col_in_651};
assign u_ca_in_652 = {{1{1'b0}}, col_in_652};
assign u_ca_in_653 = {{1{1'b0}}, col_in_653};
assign u_ca_in_654 = {{1{1'b0}}, col_in_654};
assign u_ca_in_655 = {{1{1'b0}}, col_in_655};
assign u_ca_in_656 = {{1{1'b0}}, col_in_656};
assign u_ca_in_657 = {{1{1'b0}}, col_in_657};
assign u_ca_in_658 = {{1{1'b0}}, col_in_658};
assign u_ca_in_659 = {{1{1'b0}}, col_in_659};
assign u_ca_in_660 = {{1{1'b0}}, col_in_660};
assign u_ca_in_661 = {{1{1'b0}}, col_in_661};
assign u_ca_in_662 = {{1{1'b0}}, col_in_662};
assign u_ca_in_663 = {{1{1'b0}}, col_in_663};
assign u_ca_in_664 = {{1{1'b0}}, col_in_664};
assign u_ca_in_665 = {{1{1'b0}}, col_in_665};
assign u_ca_in_666 = {{1{1'b0}}, col_in_666};
assign u_ca_in_667 = {{1{1'b0}}, col_in_667};
assign u_ca_in_668 = {{1{1'b0}}, col_in_668};
assign u_ca_in_669 = {{1{1'b0}}, col_in_669};
assign u_ca_in_670 = {{1{1'b0}}, col_in_670};
assign u_ca_in_671 = {{1{1'b0}}, col_in_671};
assign u_ca_in_672 = {{1{1'b0}}, col_in_672};
assign u_ca_in_673 = {{1{1'b0}}, col_in_673};
assign u_ca_in_674 = {{1{1'b0}}, col_in_674};
assign u_ca_in_675 = {{1{1'b0}}, col_in_675};
assign u_ca_in_676 = {{1{1'b0}}, col_in_676};
assign u_ca_in_677 = {{1{1'b0}}, col_in_677};
assign u_ca_in_678 = {{1{1'b0}}, col_in_678};
assign u_ca_in_679 = {{1{1'b0}}, col_in_679};
assign u_ca_in_680 = {{1{1'b0}}, col_in_680};
assign u_ca_in_681 = {{1{1'b0}}, col_in_681};
assign u_ca_in_682 = {{1{1'b0}}, col_in_682};
assign u_ca_in_683 = {{1{1'b0}}, col_in_683};
assign u_ca_in_684 = {{1{1'b0}}, col_in_684};
assign u_ca_in_685 = {{1{1'b0}}, col_in_685};
assign u_ca_in_686 = {{1{1'b0}}, col_in_686};
assign u_ca_in_687 = {{1{1'b0}}, col_in_687};
assign u_ca_in_688 = {{1{1'b0}}, col_in_688};
assign u_ca_in_689 = {{1{1'b0}}, col_in_689};
assign u_ca_in_690 = {{1{1'b0}}, col_in_690};
assign u_ca_in_691 = {{1{1'b0}}, col_in_691};
assign u_ca_in_692 = {{1{1'b0}}, col_in_692};
assign u_ca_in_693 = {{1{1'b0}}, col_in_693};
assign u_ca_in_694 = {{1{1'b0}}, col_in_694};
assign u_ca_in_695 = {{1{1'b0}}, col_in_695};
assign u_ca_in_696 = {{1{1'b0}}, col_in_696};
assign u_ca_in_697 = {{1{1'b0}}, col_in_697};
assign u_ca_in_698 = {{1{1'b0}}, col_in_698};
assign u_ca_in_699 = {{1{1'b0}}, col_in_699};
assign u_ca_in_700 = {{1{1'b0}}, col_in_700};
assign u_ca_in_701 = {{1{1'b0}}, col_in_701};
assign u_ca_in_702 = {{1{1'b0}}, col_in_702};
assign u_ca_in_703 = {{1{1'b0}}, col_in_703};
assign u_ca_in_704 = {{1{1'b0}}, col_in_704};
assign u_ca_in_705 = {{1{1'b0}}, col_in_705};
assign u_ca_in_706 = {{1{1'b0}}, col_in_706};
assign u_ca_in_707 = {{1{1'b0}}, col_in_707};
assign u_ca_in_708 = {{1{1'b0}}, col_in_708};
assign u_ca_in_709 = {{1{1'b0}}, col_in_709};
assign u_ca_in_710 = {{1{1'b0}}, col_in_710};
assign u_ca_in_711 = {{1{1'b0}}, col_in_711};
assign u_ca_in_712 = {{1{1'b0}}, col_in_712};
assign u_ca_in_713 = {{1{1'b0}}, col_in_713};
assign u_ca_in_714 = {{1{1'b0}}, col_in_714};
assign u_ca_in_715 = {{1{1'b0}}, col_in_715};
assign u_ca_in_716 = {{1{1'b0}}, col_in_716};
assign u_ca_in_717 = {{1{1'b0}}, col_in_717};
assign u_ca_in_718 = {{1{1'b0}}, col_in_718};
assign u_ca_in_719 = {{1{1'b0}}, col_in_719};
assign u_ca_in_720 = {{1{1'b0}}, col_in_720};
assign u_ca_in_721 = {{1{1'b0}}, col_in_721};
assign u_ca_in_722 = {{1{1'b0}}, col_in_722};
assign u_ca_in_723 = {{1{1'b0}}, col_in_723};
assign u_ca_in_724 = {{1{1'b0}}, col_in_724};
assign u_ca_in_725 = {{1{1'b0}}, col_in_725};
assign u_ca_in_726 = {{1{1'b0}}, col_in_726};
assign u_ca_in_727 = {{1{1'b0}}, col_in_727};
assign u_ca_in_728 = {{1{1'b0}}, col_in_728};
assign u_ca_in_729 = {{1{1'b0}}, col_in_729};
assign u_ca_in_730 = {{1{1'b0}}, col_in_730};
assign u_ca_in_731 = {{1{1'b0}}, col_in_731};
assign u_ca_in_732 = {{1{1'b0}}, col_in_732};
assign u_ca_in_733 = {{1{1'b0}}, col_in_733};
assign u_ca_in_734 = {{1{1'b0}}, col_in_734};
assign u_ca_in_735 = {{1{1'b0}}, col_in_735};
assign u_ca_in_736 = {{1{1'b0}}, col_in_736};
assign u_ca_in_737 = {{1{1'b0}}, col_in_737};
assign u_ca_in_738 = {{1{1'b0}}, col_in_738};
assign u_ca_in_739 = {{1{1'b0}}, col_in_739};
assign u_ca_in_740 = {{1{1'b0}}, col_in_740};
assign u_ca_in_741 = {{1{1'b0}}, col_in_741};
assign u_ca_in_742 = {{1{1'b0}}, col_in_742};
assign u_ca_in_743 = {{1{1'b0}}, col_in_743};
assign u_ca_in_744 = {{1{1'b0}}, col_in_744};
assign u_ca_in_745 = {{1{1'b0}}, col_in_745};
assign u_ca_in_746 = {{1{1'b0}}, col_in_746};
assign u_ca_in_747 = {{1{1'b0}}, col_in_747};
assign u_ca_in_748 = {{1{1'b0}}, col_in_748};
assign u_ca_in_749 = {{1{1'b0}}, col_in_749};
assign u_ca_in_750 = {{1{1'b0}}, col_in_750};
assign u_ca_in_751 = {{1{1'b0}}, col_in_751};
assign u_ca_in_752 = {{1{1'b0}}, col_in_752};
assign u_ca_in_753 = {{1{1'b0}}, col_in_753};
assign u_ca_in_754 = {{1{1'b0}}, col_in_754};
assign u_ca_in_755 = {{1{1'b0}}, col_in_755};
assign u_ca_in_756 = {{1{1'b0}}, col_in_756};
assign u_ca_in_757 = {{1{1'b0}}, col_in_757};
assign u_ca_in_758 = {{1{1'b0}}, col_in_758};
assign u_ca_in_759 = {{1{1'b0}}, col_in_759};
assign u_ca_in_760 = {{1{1'b0}}, col_in_760};
assign u_ca_in_761 = {{1{1'b0}}, col_in_761};
assign u_ca_in_762 = {{1{1'b0}}, col_in_762};
assign u_ca_in_763 = {{1{1'b0}}, col_in_763};
assign u_ca_in_764 = {{1{1'b0}}, col_in_764};
assign u_ca_in_765 = {{1{1'b0}}, col_in_765};
assign u_ca_in_766 = {{1{1'b0}}, col_in_766};
assign u_ca_in_767 = {{1{1'b0}}, col_in_767};
assign u_ca_in_768 = {{1{1'b0}}, col_in_768};
assign u_ca_in_769 = {{1{1'b0}}, col_in_769};
assign u_ca_in_770 = {{1{1'b0}}, col_in_770};
assign u_ca_in_771 = {{1{1'b0}}, col_in_771};
assign u_ca_in_772 = {{1{1'b0}}, col_in_772};
assign u_ca_in_773 = {{1{1'b0}}, col_in_773};
assign u_ca_in_774 = {{1{1'b0}}, col_in_774};
assign u_ca_in_775 = {{1{1'b0}}, col_in_775};
assign u_ca_in_776 = {{1{1'b0}}, col_in_776};
assign u_ca_in_777 = {{1{1'b0}}, col_in_777};
assign u_ca_in_778 = {{1{1'b0}}, col_in_778};
assign u_ca_in_779 = {{1{1'b0}}, col_in_779};
assign u_ca_in_780 = {{1{1'b0}}, col_in_780};
assign u_ca_in_781 = {{1{1'b0}}, col_in_781};
assign u_ca_in_782 = {{1{1'b0}}, col_in_782};
assign u_ca_in_783 = {{1{1'b0}}, col_in_783};
assign u_ca_in_784 = {{1{1'b0}}, col_in_784};
assign u_ca_in_785 = {{1{1'b0}}, col_in_785};
assign u_ca_in_786 = {{1{1'b0}}, col_in_786};
assign u_ca_in_787 = {{1{1'b0}}, col_in_787};
assign u_ca_in_788 = {{1{1'b0}}, col_in_788};
assign u_ca_in_789 = {{1{1'b0}}, col_in_789};
assign u_ca_in_790 = {{1{1'b0}}, col_in_790};
assign u_ca_in_791 = {{1{1'b0}}, col_in_791};
assign u_ca_in_792 = {{1{1'b0}}, col_in_792};
assign u_ca_in_793 = {{1{1'b0}}, col_in_793};
assign u_ca_in_794 = {{1{1'b0}}, col_in_794};
assign u_ca_in_795 = {{1{1'b0}}, col_in_795};
assign u_ca_in_796 = {{1{1'b0}}, col_in_796};
assign u_ca_in_797 = {{1{1'b0}}, col_in_797};
assign u_ca_in_798 = {{1{1'b0}}, col_in_798};
assign u_ca_in_799 = {{1{1'b0}}, col_in_799};
assign u_ca_in_800 = {{1{1'b0}}, col_in_800};
assign u_ca_in_801 = {{1{1'b0}}, col_in_801};
assign u_ca_in_802 = {{1{1'b0}}, col_in_802};
assign u_ca_in_803 = {{1{1'b0}}, col_in_803};
assign u_ca_in_804 = {{1{1'b0}}, col_in_804};
assign u_ca_in_805 = {{1{1'b0}}, col_in_805};
assign u_ca_in_806 = {{1{1'b0}}, col_in_806};
assign u_ca_in_807 = {{1{1'b0}}, col_in_807};
assign u_ca_in_808 = {{1{1'b0}}, col_in_808};
assign u_ca_in_809 = {{1{1'b0}}, col_in_809};
assign u_ca_in_810 = {{1{1'b0}}, col_in_810};
assign u_ca_in_811 = {{1{1'b0}}, col_in_811};
assign u_ca_in_812 = {{1{1'b0}}, col_in_812};
assign u_ca_in_813 = {{1{1'b0}}, col_in_813};
assign u_ca_in_814 = {{1{1'b0}}, col_in_814};
assign u_ca_in_815 = {{1{1'b0}}, col_in_815};
assign u_ca_in_816 = {{1{1'b0}}, col_in_816};
assign u_ca_in_817 = {{1{1'b0}}, col_in_817};
assign u_ca_in_818 = {{1{1'b0}}, col_in_818};
assign u_ca_in_819 = {{1{1'b0}}, col_in_819};
assign u_ca_in_820 = {{1{1'b0}}, col_in_820};
assign u_ca_in_821 = {{1{1'b0}}, col_in_821};
assign u_ca_in_822 = {{1{1'b0}}, col_in_822};
assign u_ca_in_823 = {{1{1'b0}}, col_in_823};
assign u_ca_in_824 = {{1{1'b0}}, col_in_824};
assign u_ca_in_825 = {{1{1'b0}}, col_in_825};
assign u_ca_in_826 = {{1{1'b0}}, col_in_826};
assign u_ca_in_827 = {{1{1'b0}}, col_in_827};
assign u_ca_in_828 = {{1{1'b0}}, col_in_828};
assign u_ca_in_829 = {{1{1'b0}}, col_in_829};
assign u_ca_in_830 = {{1{1'b0}}, col_in_830};
assign u_ca_in_831 = {{1{1'b0}}, col_in_831};
assign u_ca_in_832 = {{1{1'b0}}, col_in_832};
assign u_ca_in_833 = {{1{1'b0}}, col_in_833};
assign u_ca_in_834 = {{1{1'b0}}, col_in_834};
assign u_ca_in_835 = {{1{1'b0}}, col_in_835};
assign u_ca_in_836 = {{1{1'b0}}, col_in_836};
assign u_ca_in_837 = {{1{1'b0}}, col_in_837};
assign u_ca_in_838 = {{1{1'b0}}, col_in_838};
assign u_ca_in_839 = {{1{1'b0}}, col_in_839};
assign u_ca_in_840 = {{1{1'b0}}, col_in_840};
assign u_ca_in_841 = {{1{1'b0}}, col_in_841};
assign u_ca_in_842 = {{1{1'b0}}, col_in_842};
assign u_ca_in_843 = {{1{1'b0}}, col_in_843};
assign u_ca_in_844 = {{1{1'b0}}, col_in_844};
assign u_ca_in_845 = {{1{1'b0}}, col_in_845};
assign u_ca_in_846 = {{1{1'b0}}, col_in_846};
assign u_ca_in_847 = {{1{1'b0}}, col_in_847};
assign u_ca_in_848 = {{1{1'b0}}, col_in_848};
assign u_ca_in_849 = {{1{1'b0}}, col_in_849};
assign u_ca_in_850 = {{1{1'b0}}, col_in_850};
assign u_ca_in_851 = {{1{1'b0}}, col_in_851};
assign u_ca_in_852 = {{1{1'b0}}, col_in_852};
assign u_ca_in_853 = {{1{1'b0}}, col_in_853};
assign u_ca_in_854 = {{1{1'b0}}, col_in_854};
assign u_ca_in_855 = {{1{1'b0}}, col_in_855};
assign u_ca_in_856 = {{1{1'b0}}, col_in_856};
assign u_ca_in_857 = {{1{1'b0}}, col_in_857};
assign u_ca_in_858 = {{1{1'b0}}, col_in_858};
assign u_ca_in_859 = {{1{1'b0}}, col_in_859};
assign u_ca_in_860 = {{1{1'b0}}, col_in_860};
assign u_ca_in_861 = {{1{1'b0}}, col_in_861};
assign u_ca_in_862 = {{1{1'b0}}, col_in_862};
assign u_ca_in_863 = {{1{1'b0}}, col_in_863};
assign u_ca_in_864 = {{1{1'b0}}, col_in_864};
assign u_ca_in_865 = {{1{1'b0}}, col_in_865};
assign u_ca_in_866 = {{1{1'b0}}, col_in_866};
assign u_ca_in_867 = {{1{1'b0}}, col_in_867};
assign u_ca_in_868 = {{1{1'b0}}, col_in_868};
assign u_ca_in_869 = {{1{1'b0}}, col_in_869};
assign u_ca_in_870 = {{1{1'b0}}, col_in_870};
assign u_ca_in_871 = {{1{1'b0}}, col_in_871};
assign u_ca_in_872 = {{1{1'b0}}, col_in_872};
assign u_ca_in_873 = {{1{1'b0}}, col_in_873};
assign u_ca_in_874 = {{1{1'b0}}, col_in_874};
assign u_ca_in_875 = {{1{1'b0}}, col_in_875};
assign u_ca_in_876 = {{1{1'b0}}, col_in_876};
assign u_ca_in_877 = {{1{1'b0}}, col_in_877};
assign u_ca_in_878 = {{1{1'b0}}, col_in_878};
assign u_ca_in_879 = {{1{1'b0}}, col_in_879};
assign u_ca_in_880 = {{1{1'b0}}, col_in_880};
assign u_ca_in_881 = {{1{1'b0}}, col_in_881};
assign u_ca_in_882 = {{1{1'b0}}, col_in_882};
assign u_ca_in_883 = {{1{1'b0}}, col_in_883};
assign u_ca_in_884 = {{1{1'b0}}, col_in_884};
assign u_ca_in_885 = {{1{1'b0}}, col_in_885};
assign u_ca_in_886 = {{1{1'b0}}, col_in_886};
assign u_ca_in_887 = {{1{1'b0}}, col_in_887};
assign u_ca_in_888 = {{1{1'b0}}, col_in_888};
assign u_ca_in_889 = {{1{1'b0}}, col_in_889};
assign u_ca_in_890 = {{1{1'b0}}, col_in_890};
assign u_ca_in_891 = {{1{1'b0}}, col_in_891};
assign u_ca_in_892 = {{1{1'b0}}, col_in_892};
assign u_ca_in_893 = {{1{1'b0}}, col_in_893};
assign u_ca_in_894 = {{1{1'b0}}, col_in_894};
assign u_ca_in_895 = {{1{1'b0}}, col_in_895};
assign u_ca_in_896 = {{1{1'b0}}, col_in_896};
assign u_ca_in_897 = {{1{1'b0}}, col_in_897};
assign u_ca_in_898 = {{1{1'b0}}, col_in_898};
assign u_ca_in_899 = {{1{1'b0}}, col_in_899};
assign u_ca_in_900 = {{1{1'b0}}, col_in_900};
assign u_ca_in_901 = {{1{1'b0}}, col_in_901};
assign u_ca_in_902 = {{1{1'b0}}, col_in_902};
assign u_ca_in_903 = {{1{1'b0}}, col_in_903};
assign u_ca_in_904 = {{1{1'b0}}, col_in_904};
assign u_ca_in_905 = {{1{1'b0}}, col_in_905};
assign u_ca_in_906 = {{1{1'b0}}, col_in_906};
assign u_ca_in_907 = {{1{1'b0}}, col_in_907};
assign u_ca_in_908 = {{1{1'b0}}, col_in_908};
assign u_ca_in_909 = {{1{1'b0}}, col_in_909};
assign u_ca_in_910 = {{1{1'b0}}, col_in_910};
assign u_ca_in_911 = {{1{1'b0}}, col_in_911};
assign u_ca_in_912 = {{1{1'b0}}, col_in_912};
assign u_ca_in_913 = {{1{1'b0}}, col_in_913};
assign u_ca_in_914 = {{1{1'b0}}, col_in_914};
assign u_ca_in_915 = {{1{1'b0}}, col_in_915};
assign u_ca_in_916 = {{1{1'b0}}, col_in_916};
assign u_ca_in_917 = {{1{1'b0}}, col_in_917};
assign u_ca_in_918 = {{1{1'b0}}, col_in_918};
assign u_ca_in_919 = {{1{1'b0}}, col_in_919};
assign u_ca_in_920 = {{1{1'b0}}, col_in_920};
assign u_ca_in_921 = {{1{1'b0}}, col_in_921};
assign u_ca_in_922 = {{1{1'b0}}, col_in_922};
assign u_ca_in_923 = {{1{1'b0}}, col_in_923};
assign u_ca_in_924 = {{1{1'b0}}, col_in_924};
assign u_ca_in_925 = {{1{1'b0}}, col_in_925};
assign u_ca_in_926 = {{1{1'b0}}, col_in_926};
assign u_ca_in_927 = {{1{1'b0}}, col_in_927};
assign u_ca_in_928 = {{1{1'b0}}, col_in_928};
assign u_ca_in_929 = {{1{1'b0}}, col_in_929};
assign u_ca_in_930 = {{1{1'b0}}, col_in_930};
assign u_ca_in_931 = {{1{1'b0}}, col_in_931};
assign u_ca_in_932 = {{1{1'b0}}, col_in_932};
assign u_ca_in_933 = {{1{1'b0}}, col_in_933};
assign u_ca_in_934 = {{1{1'b0}}, col_in_934};
assign u_ca_in_935 = {{1{1'b0}}, col_in_935};
assign u_ca_in_936 = {{1{1'b0}}, col_in_936};
assign u_ca_in_937 = {{1{1'b0}}, col_in_937};
assign u_ca_in_938 = {{1{1'b0}}, col_in_938};
assign u_ca_in_939 = {{1{1'b0}}, col_in_939};
assign u_ca_in_940 = {{1{1'b0}}, col_in_940};
assign u_ca_in_941 = {{1{1'b0}}, col_in_941};
assign u_ca_in_942 = {{1{1'b0}}, col_in_942};
assign u_ca_in_943 = {{1{1'b0}}, col_in_943};
assign u_ca_in_944 = {{1{1'b0}}, col_in_944};
assign u_ca_in_945 = {{1{1'b0}}, col_in_945};
assign u_ca_in_946 = {{1{1'b0}}, col_in_946};
assign u_ca_in_947 = {{1{1'b0}}, col_in_947};
assign u_ca_in_948 = {{1{1'b0}}, col_in_948};
assign u_ca_in_949 = {{1{1'b0}}, col_in_949};
assign u_ca_in_950 = {{1{1'b0}}, col_in_950};
assign u_ca_in_951 = {{1{1'b0}}, col_in_951};
assign u_ca_in_952 = {{1{1'b0}}, col_in_952};
assign u_ca_in_953 = {{1{1'b0}}, col_in_953};
assign u_ca_in_954 = {{1{1'b0}}, col_in_954};
assign u_ca_in_955 = {{1{1'b0}}, col_in_955};
assign u_ca_in_956 = {{1{1'b0}}, col_in_956};
assign u_ca_in_957 = {{1{1'b0}}, col_in_957};
assign u_ca_in_958 = {{1{1'b0}}, col_in_958};
assign u_ca_in_959 = {{1{1'b0}}, col_in_959};
assign u_ca_in_960 = {{1{1'b0}}, col_in_960};
assign u_ca_in_961 = {{1{1'b0}}, col_in_961};
assign u_ca_in_962 = {{1{1'b0}}, col_in_962};
assign u_ca_in_963 = {{1{1'b0}}, col_in_963};
assign u_ca_in_964 = {{1{1'b0}}, col_in_964};
assign u_ca_in_965 = {{1{1'b0}}, col_in_965};
assign u_ca_in_966 = {{1{1'b0}}, col_in_966};
assign u_ca_in_967 = {{1{1'b0}}, col_in_967};
assign u_ca_in_968 = {{1{1'b0}}, col_in_968};
assign u_ca_in_969 = {{1{1'b0}}, col_in_969};
assign u_ca_in_970 = {{1{1'b0}}, col_in_970};
assign u_ca_in_971 = {{1{1'b0}}, col_in_971};
assign u_ca_in_972 = {{1{1'b0}}, col_in_972};
assign u_ca_in_973 = {{1{1'b0}}, col_in_973};
assign u_ca_in_974 = {{1{1'b0}}, col_in_974};
assign u_ca_in_975 = {{1{1'b0}}, col_in_975};
assign u_ca_in_976 = {{1{1'b0}}, col_in_976};
assign u_ca_in_977 = {{1{1'b0}}, col_in_977};
assign u_ca_in_978 = {{1{1'b0}}, col_in_978};
assign u_ca_in_979 = {{1{1'b0}}, col_in_979};
assign u_ca_in_980 = {{1{1'b0}}, col_in_980};
assign u_ca_in_981 = {{1{1'b0}}, col_in_981};
assign u_ca_in_982 = {{1{1'b0}}, col_in_982};
assign u_ca_in_983 = {{1{1'b0}}, col_in_983};
assign u_ca_in_984 = {{1{1'b0}}, col_in_984};
assign u_ca_in_985 = {{1{1'b0}}, col_in_985};
assign u_ca_in_986 = {{1{1'b0}}, col_in_986};
assign u_ca_in_987 = {{1{1'b0}}, col_in_987};
assign u_ca_in_988 = {{1{1'b0}}, col_in_988};
assign u_ca_in_989 = {{1{1'b0}}, col_in_989};
assign u_ca_in_990 = {{1{1'b0}}, col_in_990};
assign u_ca_in_991 = {{1{1'b0}}, col_in_991};
assign u_ca_in_992 = {{1{1'b0}}, col_in_992};
assign u_ca_in_993 = {{1{1'b0}}, col_in_993};
assign u_ca_in_994 = {{1{1'b0}}, col_in_994};
assign u_ca_in_995 = {{1{1'b0}}, col_in_995};
assign u_ca_in_996 = {{1{1'b0}}, col_in_996};
assign u_ca_in_997 = {{1{1'b0}}, col_in_997};
assign u_ca_in_998 = {{1{1'b0}}, col_in_998};
assign u_ca_in_999 = {{1{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{1{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{1{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{1{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{1{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{1{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{1{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{1{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{1{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{1{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{1{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{1{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{1{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{1{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{1{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{1{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{1{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{1{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{1{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{1{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{1{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{1{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{1{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{1{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{1{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{1{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{1{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{1{1'b0}}, col_in_1026};
assign u_ca_in_1027 = {{1{1'b0}}, col_in_1027};
assign u_ca_in_1028 = {{1{1'b0}}, col_in_1028};
assign u_ca_in_1029 = {{1{1'b0}}, col_in_1029};
assign u_ca_in_1030 = {{1{1'b0}}, col_in_1030};
assign u_ca_in_1031 = {{1{1'b0}}, col_in_1031};
assign u_ca_in_1032 = {{1{1'b0}}, col_in_1032};
assign u_ca_in_1033 = {{1{1'b0}}, col_in_1033};
assign u_ca_in_1034 = {{1{1'b0}}, col_in_1034};
assign u_ca_in_1035 = {{1{1'b0}}, col_in_1035};
assign u_ca_in_1036 = {{1{1'b0}}, col_in_1036};
assign u_ca_in_1037 = {{1{1'b0}}, col_in_1037};
assign u_ca_in_1038 = {{1{1'b0}}, col_in_1038};
assign u_ca_in_1039 = {{1{1'b0}}, col_in_1039};
assign u_ca_in_1040 = {{1{1'b0}}, col_in_1040};
assign u_ca_in_1041 = {{1{1'b0}}, col_in_1041};
assign u_ca_in_1042 = {{1{1'b0}}, col_in_1042};
assign u_ca_in_1043 = {{1{1'b0}}, col_in_1043};
assign u_ca_in_1044 = {{1{1'b0}}, col_in_1044};
assign u_ca_in_1045 = {{1{1'b0}}, col_in_1045};
assign u_ca_in_1046 = {{1{1'b0}}, col_in_1046};
assign u_ca_in_1047 = {{1{1'b0}}, col_in_1047};
assign u_ca_in_1048 = {{1{1'b0}}, col_in_1048};
assign u_ca_in_1049 = {{1{1'b0}}, col_in_1049};
assign u_ca_in_1050 = {{1{1'b0}}, col_in_1050};
assign u_ca_in_1051 = {{1{1'b0}}, col_in_1051};
assign u_ca_in_1052 = {{1{1'b0}}, col_in_1052};
assign u_ca_in_1053 = {{1{1'b0}}, col_in_1053};
assign u_ca_in_1054 = {{1{1'b0}}, col_in_1054};
assign u_ca_in_1055 = {{1{1'b0}}, col_in_1055};
assign u_ca_in_1056 = {{1{1'b0}}, col_in_1056};
assign u_ca_in_1057 = {{1{1'b0}}, col_in_1057};
assign u_ca_in_1058 = {{1{1'b0}}, col_in_1058};
assign u_ca_in_1059 = {{1{1'b0}}, col_in_1059};
assign u_ca_in_1060 = {{1{1'b0}}, col_in_1060};
assign u_ca_in_1061 = {{1{1'b0}}, col_in_1061};
assign u_ca_in_1062 = {{1{1'b0}}, col_in_1062};
assign u_ca_in_1063 = {{1{1'b0}}, col_in_1063};
assign u_ca_in_1064 = {{1{1'b0}}, col_in_1064};
assign u_ca_in_1065 = {{1{1'b0}}, col_in_1065};
assign u_ca_in_1066 = {{1{1'b0}}, col_in_1066};
assign u_ca_in_1067 = {{1{1'b0}}, col_in_1067};
assign u_ca_in_1068 = {{1{1'b0}}, col_in_1068};
assign u_ca_in_1069 = {{1{1'b0}}, col_in_1069};
assign u_ca_in_1070 = {{1{1'b0}}, col_in_1070};
assign u_ca_in_1071 = {{1{1'b0}}, col_in_1071};
assign u_ca_in_1072 = {{1{1'b0}}, col_in_1072};
assign u_ca_in_1073 = {{1{1'b0}}, col_in_1073};
assign u_ca_in_1074 = {{1{1'b0}}, col_in_1074};
assign u_ca_in_1075 = {{1{1'b0}}, col_in_1075};
assign u_ca_in_1076 = {{1{1'b0}}, col_in_1076};
assign u_ca_in_1077 = {{1{1'b0}}, col_in_1077};
assign u_ca_in_1078 = {{1{1'b0}}, col_in_1078};
assign u_ca_in_1079 = {{1{1'b0}}, col_in_1079};
assign u_ca_in_1080 = {{1{1'b0}}, col_in_1080};
assign u_ca_in_1081 = {{1{1'b0}}, col_in_1081};
assign u_ca_in_1082 = {{1{1'b0}}, col_in_1082};
assign u_ca_in_1083 = {{1{1'b0}}, col_in_1083};
assign u_ca_in_1084 = {{1{1'b0}}, col_in_1084};
assign u_ca_in_1085 = {{1{1'b0}}, col_in_1085};
assign u_ca_in_1086 = {{1{1'b0}}, col_in_1086};
assign u_ca_in_1087 = {{1{1'b0}}, col_in_1087};
assign u_ca_in_1088 = {{1{1'b0}}, col_in_1088};
assign u_ca_in_1089 = {{1{1'b0}}, col_in_1089};
assign u_ca_in_1090 = {{1{1'b0}}, col_in_1090};
assign u_ca_in_1091 = {{1{1'b0}}, col_in_1091};
assign u_ca_in_1092 = {{1{1'b0}}, col_in_1092};
assign u_ca_in_1093 = {{1{1'b0}}, col_in_1093};
assign u_ca_in_1094 = {{1{1'b0}}, col_in_1094};
assign u_ca_in_1095 = {{1{1'b0}}, col_in_1095};
assign u_ca_in_1096 = {{1{1'b0}}, col_in_1096};
assign u_ca_in_1097 = {{1{1'b0}}, col_in_1097};
assign u_ca_in_1098 = {{1{1'b0}}, col_in_1098};
assign u_ca_in_1099 = {{1{1'b0}}, col_in_1099};
assign u_ca_in_1100 = {{1{1'b0}}, col_in_1100};
assign u_ca_in_1101 = {{1{1'b0}}, col_in_1101};
assign u_ca_in_1102 = {{1{1'b0}}, col_in_1102};
assign u_ca_in_1103 = {{1{1'b0}}, col_in_1103};
assign u_ca_in_1104 = {{1{1'b0}}, col_in_1104};
assign u_ca_in_1105 = {{1{1'b0}}, col_in_1105};
assign u_ca_in_1106 = {{1{1'b0}}, col_in_1106};
assign u_ca_in_1107 = {{1{1'b0}}, col_in_1107};
assign u_ca_in_1108 = {{1{1'b0}}, col_in_1108};
assign u_ca_in_1109 = {{1{1'b0}}, col_in_1109};
assign u_ca_in_1110 = {{1{1'b0}}, col_in_1110};
assign u_ca_in_1111 = {{1{1'b0}}, col_in_1111};
assign u_ca_in_1112 = {{1{1'b0}}, col_in_1112};
assign u_ca_in_1113 = {{1{1'b0}}, col_in_1113};
assign u_ca_in_1114 = {{1{1'b0}}, col_in_1114};
assign u_ca_in_1115 = {{1{1'b0}}, col_in_1115};
assign u_ca_in_1116 = {{1{1'b0}}, col_in_1116};
assign u_ca_in_1117 = {{1{1'b0}}, col_in_1117};
assign u_ca_in_1118 = {{1{1'b0}}, col_in_1118};
assign u_ca_in_1119 = {{1{1'b0}}, col_in_1119};
assign u_ca_in_1120 = {{1{1'b0}}, col_in_1120};
assign u_ca_in_1121 = {{1{1'b0}}, col_in_1121};
assign u_ca_in_1122 = {{1{1'b0}}, col_in_1122};
assign u_ca_in_1123 = {{1{1'b0}}, col_in_1123};
assign u_ca_in_1124 = {{1{1'b0}}, col_in_1124};
assign u_ca_in_1125 = {{1{1'b0}}, col_in_1125};
assign u_ca_in_1126 = {{1{1'b0}}, col_in_1126};
assign u_ca_in_1127 = {{1{1'b0}}, col_in_1127};
assign u_ca_in_1128 = {{1{1'b0}}, col_in_1128};
assign u_ca_in_1129 = {{1{1'b0}}, col_in_1129};
assign u_ca_in_1130 = {{1{1'b0}}, col_in_1130};
assign u_ca_in_1131 = {{1{1'b0}}, col_in_1131};
assign u_ca_in_1132 = {{1{1'b0}}, col_in_1132};
assign u_ca_in_1133 = {{1{1'b0}}, col_in_1133};
assign u_ca_in_1134 = {{1{1'b0}}, col_in_1134};
assign u_ca_in_1135 = {{1{1'b0}}, col_in_1135};
assign u_ca_in_1136 = {{1{1'b0}}, col_in_1136};
assign u_ca_in_1137 = {{1{1'b0}}, col_in_1137};
assign u_ca_in_1138 = {{1{1'b0}}, col_in_1138};
assign u_ca_in_1139 = {{1{1'b0}}, col_in_1139};
assign u_ca_in_1140 = {{1{1'b0}}, col_in_1140};
assign u_ca_in_1141 = {{1{1'b0}}, col_in_1141};
assign u_ca_in_1142 = {{1{1'b0}}, col_in_1142};
assign u_ca_in_1143 = {{1{1'b0}}, col_in_1143};
assign u_ca_in_1144 = {{1{1'b0}}, col_in_1144};
assign u_ca_in_1145 = {{1{1'b0}}, col_in_1145};
assign u_ca_in_1146 = {{1{1'b0}}, col_in_1146};
assign u_ca_in_1147 = {{1{1'b0}}, col_in_1147};
assign u_ca_in_1148 = {{1{1'b0}}, col_in_1148};
assign u_ca_in_1149 = {{1{1'b0}}, col_in_1149};
assign u_ca_in_1150 = {{1{1'b0}}, col_in_1150};
assign u_ca_in_1151 = {{1{1'b0}}, col_in_1151};
assign u_ca_in_1152 = {{1{1'b0}}, col_in_1152};
assign u_ca_in_1153 = {{1{1'b0}}, col_in_1153};
assign u_ca_in_1154 = {{1{1'b0}}, col_in_1154};
assign u_ca_in_1155 = {{1{1'b0}}, col_in_1155};
assign u_ca_in_1156 = {{1{1'b0}}, col_in_1156};
assign u_ca_in_1157 = {{1{1'b0}}, col_in_1157};
assign u_ca_in_1158 = {{1{1'b0}}, col_in_1158};
assign u_ca_in_1159 = {{1{1'b0}}, col_in_1159};
assign u_ca_in_1160 = {{1{1'b0}}, col_in_1160};
assign u_ca_in_1161 = {{1{1'b0}}, col_in_1161};
assign u_ca_in_1162 = {{1{1'b0}}, col_in_1162};
assign u_ca_in_1163 = {{1{1'b0}}, col_in_1163};
assign u_ca_in_1164 = {{1{1'b0}}, col_in_1164};
assign u_ca_in_1165 = {{1{1'b0}}, col_in_1165};
assign u_ca_in_1166 = {{1{1'b0}}, col_in_1166};
assign u_ca_in_1167 = {{1{1'b0}}, col_in_1167};
assign u_ca_in_1168 = {{1{1'b0}}, col_in_1168};
assign u_ca_in_1169 = {{1{1'b0}}, col_in_1169};
assign u_ca_in_1170 = {{1{1'b0}}, col_in_1170};
assign u_ca_in_1171 = {{1{1'b0}}, col_in_1171};
assign u_ca_in_1172 = {{1{1'b0}}, col_in_1172};
assign u_ca_in_1173 = {{1{1'b0}}, col_in_1173};
assign u_ca_in_1174 = {{1{1'b0}}, col_in_1174};
assign u_ca_in_1175 = {{1{1'b0}}, col_in_1175};
assign u_ca_in_1176 = {{1{1'b0}}, col_in_1176};
assign u_ca_in_1177 = {{1{1'b0}}, col_in_1177};
assign u_ca_in_1178 = {{1{1'b0}}, col_in_1178};
assign u_ca_in_1179 = {{1{1'b0}}, col_in_1179};
assign u_ca_in_1180 = {{1{1'b0}}, col_in_1180};
assign u_ca_in_1181 = {{1{1'b0}}, col_in_1181};
assign u_ca_in_1182 = {{1{1'b0}}, col_in_1182};
assign u_ca_in_1183 = {{1{1'b0}}, col_in_1183};
assign u_ca_in_1184 = {{1{1'b0}}, col_in_1184};
assign u_ca_in_1185 = {{1{1'b0}}, col_in_1185};
assign u_ca_in_1186 = {{1{1'b0}}, col_in_1186};
assign u_ca_in_1187 = {{1{1'b0}}, col_in_1187};
assign u_ca_in_1188 = {{1{1'b0}}, col_in_1188};
assign u_ca_in_1189 = {{1{1'b0}}, col_in_1189};
assign u_ca_in_1190 = {{1{1'b0}}, col_in_1190};
assign u_ca_in_1191 = {{1{1'b0}}, col_in_1191};
assign u_ca_in_1192 = {{1{1'b0}}, col_in_1192};
assign u_ca_in_1193 = {{1{1'b0}}, col_in_1193};
assign u_ca_in_1194 = {{1{1'b0}}, col_in_1194};
assign u_ca_in_1195 = {{1{1'b0}}, col_in_1195};
assign u_ca_in_1196 = {{1{1'b0}}, col_in_1196};
assign u_ca_in_1197 = {{1{1'b0}}, col_in_1197};
assign u_ca_in_1198 = {{1{1'b0}}, col_in_1198};
assign u_ca_in_1199 = {{1{1'b0}}, col_in_1199};
assign u_ca_in_1200 = {{1{1'b0}}, col_in_1200};
assign u_ca_in_1201 = {{1{1'b0}}, col_in_1201};
assign u_ca_in_1202 = {{1{1'b0}}, col_in_1202};
assign u_ca_in_1203 = {{1{1'b0}}, col_in_1203};
assign u_ca_in_1204 = {{1{1'b0}}, col_in_1204};
assign u_ca_in_1205 = {{1{1'b0}}, col_in_1205};
assign u_ca_in_1206 = {{1{1'b0}}, col_in_1206};
assign u_ca_in_1207 = {{1{1'b0}}, col_in_1207};
assign u_ca_in_1208 = {{1{1'b0}}, col_in_1208};
assign u_ca_in_1209 = {{1{1'b0}}, col_in_1209};
assign u_ca_in_1210 = {{1{1'b0}}, col_in_1210};
assign u_ca_in_1211 = {{1{1'b0}}, col_in_1211};
assign u_ca_in_1212 = {{1{1'b0}}, col_in_1212};
assign u_ca_in_1213 = {{1{1'b0}}, col_in_1213};
assign u_ca_in_1214 = {{1{1'b0}}, col_in_1214};
assign u_ca_in_1215 = {{1{1'b0}}, col_in_1215};
assign u_ca_in_1216 = {{1{1'b0}}, col_in_1216};
assign u_ca_in_1217 = {{1{1'b0}}, col_in_1217};
assign u_ca_in_1218 = {{1{1'b0}}, col_in_1218};
assign u_ca_in_1219 = {{1{1'b0}}, col_in_1219};
assign u_ca_in_1220 = {{1{1'b0}}, col_in_1220};
assign u_ca_in_1221 = {{1{1'b0}}, col_in_1221};
assign u_ca_in_1222 = {{1{1'b0}}, col_in_1222};
assign u_ca_in_1223 = {{1{1'b0}}, col_in_1223};
assign u_ca_in_1224 = {{1{1'b0}}, col_in_1224};
assign u_ca_in_1225 = {{1{1'b0}}, col_in_1225};
assign u_ca_in_1226 = {{1{1'b0}}, col_in_1226};
assign u_ca_in_1227 = {{1{1'b0}}, col_in_1227};
assign u_ca_in_1228 = {{1{1'b0}}, col_in_1228};
assign u_ca_in_1229 = {{1{1'b0}}, col_in_1229};
assign u_ca_in_1230 = {{1{1'b0}}, col_in_1230};
assign u_ca_in_1231 = {{1{1'b0}}, col_in_1231};
assign u_ca_in_1232 = {{1{1'b0}}, col_in_1232};
assign u_ca_in_1233 = {{1{1'b0}}, col_in_1233};
assign u_ca_in_1234 = {{1{1'b0}}, col_in_1234};
assign u_ca_in_1235 = {{1{1'b0}}, col_in_1235};
assign u_ca_in_1236 = {{1{1'b0}}, col_in_1236};
assign u_ca_in_1237 = {{1{1'b0}}, col_in_1237};
assign u_ca_in_1238 = {{1{1'b0}}, col_in_1238};
assign u_ca_in_1239 = {{1{1'b0}}, col_in_1239};
assign u_ca_in_1240 = {{1{1'b0}}, col_in_1240};
assign u_ca_in_1241 = {{1{1'b0}}, col_in_1241};
assign u_ca_in_1242 = {{1{1'b0}}, col_in_1242};
assign u_ca_in_1243 = {{1{1'b0}}, col_in_1243};
assign u_ca_in_1244 = {{1{1'b0}}, col_in_1244};
assign u_ca_in_1245 = {{1{1'b0}}, col_in_1245};
assign u_ca_in_1246 = {{1{1'b0}}, col_in_1246};
assign u_ca_in_1247 = {{1{1'b0}}, col_in_1247};
assign u_ca_in_1248 = {{1{1'b0}}, col_in_1248};
assign u_ca_in_1249 = {{1{1'b0}}, col_in_1249};
assign u_ca_in_1250 = {{1{1'b0}}, col_in_1250};
assign u_ca_in_1251 = {{1{1'b0}}, col_in_1251};
assign u_ca_in_1252 = {{1{1'b0}}, col_in_1252};
assign u_ca_in_1253 = {{1{1'b0}}, col_in_1253};
assign u_ca_in_1254 = {{1{1'b0}}, col_in_1254};
assign u_ca_in_1255 = {{1{1'b0}}, col_in_1255};
assign u_ca_in_1256 = {{1{1'b0}}, col_in_1256};
assign u_ca_in_1257 = {{1{1'b0}}, col_in_1257};
assign u_ca_in_1258 = {{1{1'b0}}, col_in_1258};
assign u_ca_in_1259 = {{1{1'b0}}, col_in_1259};
assign u_ca_in_1260 = {{1{1'b0}}, col_in_1260};
assign u_ca_in_1261 = {{1{1'b0}}, col_in_1261};
assign u_ca_in_1262 = {{1{1'b0}}, col_in_1262};
assign u_ca_in_1263 = {{1{1'b0}}, col_in_1263};
assign u_ca_in_1264 = {{1{1'b0}}, col_in_1264};
assign u_ca_in_1265 = {{1{1'b0}}, col_in_1265};
assign u_ca_in_1266 = {{1{1'b0}}, col_in_1266};
assign u_ca_in_1267 = {{1{1'b0}}, col_in_1267};
assign u_ca_in_1268 = {{1{1'b0}}, col_in_1268};
assign u_ca_in_1269 = {{1{1'b0}}, col_in_1269};
assign u_ca_in_1270 = {{1{1'b0}}, col_in_1270};
assign u_ca_in_1271 = {{1{1'b0}}, col_in_1271};
assign u_ca_in_1272 = {{1{1'b0}}, col_in_1272};
assign u_ca_in_1273 = {{1{1'b0}}, col_in_1273};
assign u_ca_in_1274 = {{1{1'b0}}, col_in_1274};
assign u_ca_in_1275 = {{1{1'b0}}, col_in_1275};
assign u_ca_in_1276 = {{1{1'b0}}, col_in_1276};
assign u_ca_in_1277 = {{1{1'b0}}, col_in_1277};
assign u_ca_in_1278 = {{1{1'b0}}, col_in_1278};
assign u_ca_in_1279 = {{1{1'b0}}, col_in_1279};
assign u_ca_in_1280 = {{1{1'b0}}, col_in_1280};
assign u_ca_in_1281 = {{1{1'b0}}, col_in_1281};
assign u_ca_in_1282 = {{1{1'b0}}, col_in_1282};
assign u_ca_in_1283 = {{1{1'b0}}, col_in_1283};
assign u_ca_in_1284 = {{1{1'b0}}, col_in_1284};
assign u_ca_in_1285 = {{1{1'b0}}, col_in_1285};
assign u_ca_in_1286 = {{1{1'b0}}, col_in_1286};
assign u_ca_in_1287 = {{1{1'b0}}, col_in_1287};

//---------------------------------------------------------


compressor_9_6 u_ca_9_6_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_9_6 u_ca_9_6_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_9_6 u_ca_9_6_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_9_6 u_ca_9_6_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_9_6 u_ca_9_6_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_9_6 u_ca_9_6_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_9_6 u_ca_9_6_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_9_6 u_ca_9_6_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_9_6 u_ca_9_6_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_9_6 u_ca_9_6_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_9_6 u_ca_9_6_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_9_6 u_ca_9_6_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_9_6 u_ca_9_6_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_9_6 u_ca_9_6_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_9_6 u_ca_9_6_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_9_6 u_ca_9_6_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_9_6 u_ca_9_6_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_9_6 u_ca_9_6_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_9_6 u_ca_9_6_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_9_6 u_ca_9_6_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_9_6 u_ca_9_6_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_9_6 u_ca_9_6_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_9_6 u_ca_9_6_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_9_6 u_ca_9_6_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_9_6 u_ca_9_6_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_9_6 u_ca_9_6_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_9_6 u_ca_9_6_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_9_6 u_ca_9_6_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_9_6 u_ca_9_6_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_9_6 u_ca_9_6_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_9_6 u_ca_9_6_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_9_6 u_ca_9_6_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_9_6 u_ca_9_6_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_9_6 u_ca_9_6_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_9_6 u_ca_9_6_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_9_6 u_ca_9_6_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_9_6 u_ca_9_6_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_9_6 u_ca_9_6_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_9_6 u_ca_9_6_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_9_6 u_ca_9_6_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_9_6 u_ca_9_6_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_9_6 u_ca_9_6_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_9_6 u_ca_9_6_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_9_6 u_ca_9_6_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_9_6 u_ca_9_6_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_9_6 u_ca_9_6_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_9_6 u_ca_9_6_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_9_6 u_ca_9_6_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_9_6 u_ca_9_6_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_9_6 u_ca_9_6_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_9_6 u_ca_9_6_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_9_6 u_ca_9_6_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_9_6 u_ca_9_6_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_9_6 u_ca_9_6_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_9_6 u_ca_9_6_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_9_6 u_ca_9_6_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_9_6 u_ca_9_6_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_9_6 u_ca_9_6_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_9_6 u_ca_9_6_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_9_6 u_ca_9_6_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_9_6 u_ca_9_6_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_9_6 u_ca_9_6_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_9_6 u_ca_9_6_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_9_6 u_ca_9_6_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_9_6 u_ca_9_6_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_9_6 u_ca_9_6_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_9_6 u_ca_9_6_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_9_6 u_ca_9_6_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_9_6 u_ca_9_6_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_9_6 u_ca_9_6_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_9_6 u_ca_9_6_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_9_6 u_ca_9_6_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_9_6 u_ca_9_6_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_9_6 u_ca_9_6_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_9_6 u_ca_9_6_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_9_6 u_ca_9_6_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_9_6 u_ca_9_6_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_9_6 u_ca_9_6_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_9_6 u_ca_9_6_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_9_6 u_ca_9_6_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_9_6 u_ca_9_6_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_9_6 u_ca_9_6_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_9_6 u_ca_9_6_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_9_6 u_ca_9_6_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_9_6 u_ca_9_6_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_9_6 u_ca_9_6_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_9_6 u_ca_9_6_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_9_6 u_ca_9_6_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_9_6 u_ca_9_6_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_9_6 u_ca_9_6_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_9_6 u_ca_9_6_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_9_6 u_ca_9_6_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_9_6 u_ca_9_6_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_9_6 u_ca_9_6_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_9_6 u_ca_9_6_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_9_6 u_ca_9_6_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_9_6 u_ca_9_6_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_9_6 u_ca_9_6_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_9_6 u_ca_9_6_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_9_6 u_ca_9_6_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_9_6 u_ca_9_6_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_9_6 u_ca_9_6_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_9_6 u_ca_9_6_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_9_6 u_ca_9_6_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_9_6 u_ca_9_6_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_9_6 u_ca_9_6_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_9_6 u_ca_9_6_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_9_6 u_ca_9_6_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_9_6 u_ca_9_6_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_9_6 u_ca_9_6_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_9_6 u_ca_9_6_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_9_6 u_ca_9_6_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_9_6 u_ca_9_6_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_9_6 u_ca_9_6_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_9_6 u_ca_9_6_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_9_6 u_ca_9_6_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_9_6 u_ca_9_6_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_9_6 u_ca_9_6_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_9_6 u_ca_9_6_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_9_6 u_ca_9_6_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_9_6 u_ca_9_6_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_9_6 u_ca_9_6_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_9_6 u_ca_9_6_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_9_6 u_ca_9_6_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_9_6 u_ca_9_6_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_9_6 u_ca_9_6_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_9_6 u_ca_9_6_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_9_6 u_ca_9_6_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_9_6 u_ca_9_6_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_9_6 u_ca_9_6_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_9_6 u_ca_9_6_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_9_6 u_ca_9_6_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_9_6 u_ca_9_6_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_9_6 u_ca_9_6_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_9_6 u_ca_9_6_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_9_6 u_ca_9_6_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_9_6 u_ca_9_6_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_9_6 u_ca_9_6_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_9_6 u_ca_9_6_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_9_6 u_ca_9_6_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_9_6 u_ca_9_6_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_9_6 u_ca_9_6_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_9_6 u_ca_9_6_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_9_6 u_ca_9_6_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_9_6 u_ca_9_6_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_9_6 u_ca_9_6_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_9_6 u_ca_9_6_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_9_6 u_ca_9_6_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_9_6 u_ca_9_6_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_9_6 u_ca_9_6_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_9_6 u_ca_9_6_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_9_6 u_ca_9_6_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_9_6 u_ca_9_6_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_9_6 u_ca_9_6_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_9_6 u_ca_9_6_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_9_6 u_ca_9_6_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_9_6 u_ca_9_6_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_9_6 u_ca_9_6_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_9_6 u_ca_9_6_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_9_6 u_ca_9_6_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_9_6 u_ca_9_6_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_9_6 u_ca_9_6_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_9_6 u_ca_9_6_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_9_6 u_ca_9_6_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_9_6 u_ca_9_6_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_9_6 u_ca_9_6_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_9_6 u_ca_9_6_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_9_6 u_ca_9_6_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_9_6 u_ca_9_6_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_9_6 u_ca_9_6_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_9_6 u_ca_9_6_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_9_6 u_ca_9_6_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_9_6 u_ca_9_6_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_9_6 u_ca_9_6_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_9_6 u_ca_9_6_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_9_6 u_ca_9_6_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_9_6 u_ca_9_6_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_9_6 u_ca_9_6_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_9_6 u_ca_9_6_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_9_6 u_ca_9_6_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_9_6 u_ca_9_6_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_9_6 u_ca_9_6_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_9_6 u_ca_9_6_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_9_6 u_ca_9_6_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_9_6 u_ca_9_6_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_9_6 u_ca_9_6_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_9_6 u_ca_9_6_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_9_6 u_ca_9_6_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_9_6 u_ca_9_6_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_9_6 u_ca_9_6_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_9_6 u_ca_9_6_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_9_6 u_ca_9_6_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_9_6 u_ca_9_6_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_9_6 u_ca_9_6_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_9_6 u_ca_9_6_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_9_6 u_ca_9_6_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_9_6 u_ca_9_6_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_9_6 u_ca_9_6_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_9_6 u_ca_9_6_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_9_6 u_ca_9_6_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_9_6 u_ca_9_6_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_9_6 u_ca_9_6_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_9_6 u_ca_9_6_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_9_6 u_ca_9_6_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_9_6 u_ca_9_6_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_9_6 u_ca_9_6_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_9_6 u_ca_9_6_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_9_6 u_ca_9_6_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_9_6 u_ca_9_6_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_9_6 u_ca_9_6_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_9_6 u_ca_9_6_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_9_6 u_ca_9_6_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_9_6 u_ca_9_6_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_9_6 u_ca_9_6_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_9_6 u_ca_9_6_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_9_6 u_ca_9_6_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_9_6 u_ca_9_6_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_9_6 u_ca_9_6_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_9_6 u_ca_9_6_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_9_6 u_ca_9_6_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_9_6 u_ca_9_6_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_9_6 u_ca_9_6_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_9_6 u_ca_9_6_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_9_6 u_ca_9_6_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_9_6 u_ca_9_6_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_9_6 u_ca_9_6_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_9_6 u_ca_9_6_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_9_6 u_ca_9_6_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_9_6 u_ca_9_6_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_9_6 u_ca_9_6_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_9_6 u_ca_9_6_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_9_6 u_ca_9_6_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_9_6 u_ca_9_6_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_9_6 u_ca_9_6_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_9_6 u_ca_9_6_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_9_6 u_ca_9_6_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_9_6 u_ca_9_6_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_9_6 u_ca_9_6_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_9_6 u_ca_9_6_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_9_6 u_ca_9_6_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_9_6 u_ca_9_6_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_9_6 u_ca_9_6_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_9_6 u_ca_9_6_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_9_6 u_ca_9_6_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_9_6 u_ca_9_6_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_9_6 u_ca_9_6_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_9_6 u_ca_9_6_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_9_6 u_ca_9_6_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_9_6 u_ca_9_6_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_9_6 u_ca_9_6_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_9_6 u_ca_9_6_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_9_6 u_ca_9_6_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_9_6 u_ca_9_6_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_9_6 u_ca_9_6_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_9_6 u_ca_9_6_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_9_6 u_ca_9_6_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_9_6 u_ca_9_6_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_9_6 u_ca_9_6_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_9_6 u_ca_9_6_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_9_6 u_ca_9_6_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_9_6 u_ca_9_6_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_9_6 u_ca_9_6_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_9_6 u_ca_9_6_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_9_6 u_ca_9_6_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_9_6 u_ca_9_6_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_9_6 u_ca_9_6_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_9_6 u_ca_9_6_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_9_6 u_ca_9_6_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_9_6 u_ca_9_6_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_9_6 u_ca_9_6_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_9_6 u_ca_9_6_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_9_6 u_ca_9_6_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_9_6 u_ca_9_6_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_9_6 u_ca_9_6_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_9_6 u_ca_9_6_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_9_6 u_ca_9_6_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_9_6 u_ca_9_6_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_9_6 u_ca_9_6_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_9_6 u_ca_9_6_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_9_6 u_ca_9_6_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_9_6 u_ca_9_6_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_9_6 u_ca_9_6_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_9_6 u_ca_9_6_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_9_6 u_ca_9_6_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_9_6 u_ca_9_6_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_9_6 u_ca_9_6_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_9_6 u_ca_9_6_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_9_6 u_ca_9_6_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_9_6 u_ca_9_6_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_9_6 u_ca_9_6_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_9_6 u_ca_9_6_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_9_6 u_ca_9_6_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_9_6 u_ca_9_6_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_9_6 u_ca_9_6_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_9_6 u_ca_9_6_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_9_6 u_ca_9_6_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_9_6 u_ca_9_6_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_9_6 u_ca_9_6_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_9_6 u_ca_9_6_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_9_6 u_ca_9_6_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_9_6 u_ca_9_6_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_9_6 u_ca_9_6_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_9_6 u_ca_9_6_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_9_6 u_ca_9_6_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_9_6 u_ca_9_6_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_9_6 u_ca_9_6_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_9_6 u_ca_9_6_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_9_6 u_ca_9_6_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_9_6 u_ca_9_6_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_9_6 u_ca_9_6_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_9_6 u_ca_9_6_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_9_6 u_ca_9_6_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_9_6 u_ca_9_6_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_9_6 u_ca_9_6_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_9_6 u_ca_9_6_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_9_6 u_ca_9_6_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_9_6 u_ca_9_6_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_9_6 u_ca_9_6_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_9_6 u_ca_9_6_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_9_6 u_ca_9_6_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_9_6 u_ca_9_6_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_9_6 u_ca_9_6_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_9_6 u_ca_9_6_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_9_6 u_ca_9_6_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_9_6 u_ca_9_6_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_9_6 u_ca_9_6_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_9_6 u_ca_9_6_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_9_6 u_ca_9_6_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_9_6 u_ca_9_6_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_9_6 u_ca_9_6_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_9_6 u_ca_9_6_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_9_6 u_ca_9_6_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_9_6 u_ca_9_6_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_9_6 u_ca_9_6_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_9_6 u_ca_9_6_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_9_6 u_ca_9_6_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_9_6 u_ca_9_6_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_9_6 u_ca_9_6_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_9_6 u_ca_9_6_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_9_6 u_ca_9_6_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_9_6 u_ca_9_6_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_9_6 u_ca_9_6_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_9_6 u_ca_9_6_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_9_6 u_ca_9_6_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_9_6 u_ca_9_6_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_9_6 u_ca_9_6_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_9_6 u_ca_9_6_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_9_6 u_ca_9_6_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_9_6 u_ca_9_6_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_9_6 u_ca_9_6_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_9_6 u_ca_9_6_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_9_6 u_ca_9_6_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_9_6 u_ca_9_6_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_9_6 u_ca_9_6_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_9_6 u_ca_9_6_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_9_6 u_ca_9_6_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_9_6 u_ca_9_6_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_9_6 u_ca_9_6_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_9_6 u_ca_9_6_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_9_6 u_ca_9_6_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_9_6 u_ca_9_6_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_9_6 u_ca_9_6_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_9_6 u_ca_9_6_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_9_6 u_ca_9_6_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_9_6 u_ca_9_6_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_9_6 u_ca_9_6_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_9_6 u_ca_9_6_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_9_6 u_ca_9_6_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_9_6 u_ca_9_6_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_9_6 u_ca_9_6_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_9_6 u_ca_9_6_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_9_6 u_ca_9_6_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_9_6 u_ca_9_6_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_9_6 u_ca_9_6_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_9_6 u_ca_9_6_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_9_6 u_ca_9_6_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_9_6 u_ca_9_6_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_9_6 u_ca_9_6_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_9_6 u_ca_9_6_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_9_6 u_ca_9_6_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_9_6 u_ca_9_6_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_9_6 u_ca_9_6_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_9_6 u_ca_9_6_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_9_6 u_ca_9_6_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_9_6 u_ca_9_6_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_9_6 u_ca_9_6_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_9_6 u_ca_9_6_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_9_6 u_ca_9_6_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_9_6 u_ca_9_6_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_9_6 u_ca_9_6_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_9_6 u_ca_9_6_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_9_6 u_ca_9_6_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_9_6 u_ca_9_6_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_9_6 u_ca_9_6_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_9_6 u_ca_9_6_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_9_6 u_ca_9_6_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_9_6 u_ca_9_6_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_9_6 u_ca_9_6_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_9_6 u_ca_9_6_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_9_6 u_ca_9_6_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_9_6 u_ca_9_6_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_9_6 u_ca_9_6_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_9_6 u_ca_9_6_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_9_6 u_ca_9_6_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_9_6 u_ca_9_6_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_9_6 u_ca_9_6_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_9_6 u_ca_9_6_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_9_6 u_ca_9_6_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_9_6 u_ca_9_6_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_9_6 u_ca_9_6_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_9_6 u_ca_9_6_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_9_6 u_ca_9_6_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_9_6 u_ca_9_6_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_9_6 u_ca_9_6_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_9_6 u_ca_9_6_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_9_6 u_ca_9_6_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_9_6 u_ca_9_6_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_9_6 u_ca_9_6_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_9_6 u_ca_9_6_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_9_6 u_ca_9_6_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_9_6 u_ca_9_6_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_9_6 u_ca_9_6_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_9_6 u_ca_9_6_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_9_6 u_ca_9_6_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_9_6 u_ca_9_6_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_9_6 u_ca_9_6_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_9_6 u_ca_9_6_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_9_6 u_ca_9_6_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_9_6 u_ca_9_6_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_9_6 u_ca_9_6_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_9_6 u_ca_9_6_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_9_6 u_ca_9_6_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_9_6 u_ca_9_6_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_9_6 u_ca_9_6_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_9_6 u_ca_9_6_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_9_6 u_ca_9_6_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_9_6 u_ca_9_6_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_9_6 u_ca_9_6_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_9_6 u_ca_9_6_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_9_6 u_ca_9_6_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_9_6 u_ca_9_6_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_9_6 u_ca_9_6_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_9_6 u_ca_9_6_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_9_6 u_ca_9_6_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_9_6 u_ca_9_6_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_9_6 u_ca_9_6_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_9_6 u_ca_9_6_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_9_6 u_ca_9_6_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_9_6 u_ca_9_6_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_9_6 u_ca_9_6_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_9_6 u_ca_9_6_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_9_6 u_ca_9_6_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_9_6 u_ca_9_6_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_9_6 u_ca_9_6_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_9_6 u_ca_9_6_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_9_6 u_ca_9_6_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_9_6 u_ca_9_6_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_9_6 u_ca_9_6_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_9_6 u_ca_9_6_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_9_6 u_ca_9_6_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_9_6 u_ca_9_6_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_9_6 u_ca_9_6_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_9_6 u_ca_9_6_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_9_6 u_ca_9_6_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_9_6 u_ca_9_6_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_9_6 u_ca_9_6_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_9_6 u_ca_9_6_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_9_6 u_ca_9_6_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_9_6 u_ca_9_6_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_9_6 u_ca_9_6_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_9_6 u_ca_9_6_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_9_6 u_ca_9_6_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_9_6 u_ca_9_6_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_9_6 u_ca_9_6_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_9_6 u_ca_9_6_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_9_6 u_ca_9_6_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_9_6 u_ca_9_6_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_9_6 u_ca_9_6_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_9_6 u_ca_9_6_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_9_6 u_ca_9_6_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_9_6 u_ca_9_6_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_9_6 u_ca_9_6_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_9_6 u_ca_9_6_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_9_6 u_ca_9_6_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_9_6 u_ca_9_6_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_9_6 u_ca_9_6_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_9_6 u_ca_9_6_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_9_6 u_ca_9_6_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_9_6 u_ca_9_6_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_9_6 u_ca_9_6_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_9_6 u_ca_9_6_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_9_6 u_ca_9_6_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_9_6 u_ca_9_6_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_9_6 u_ca_9_6_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_9_6 u_ca_9_6_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_9_6 u_ca_9_6_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_9_6 u_ca_9_6_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_9_6 u_ca_9_6_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_9_6 u_ca_9_6_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_9_6 u_ca_9_6_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_9_6 u_ca_9_6_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_9_6 u_ca_9_6_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_9_6 u_ca_9_6_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_9_6 u_ca_9_6_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_9_6 u_ca_9_6_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_9_6 u_ca_9_6_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_9_6 u_ca_9_6_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_9_6 u_ca_9_6_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_9_6 u_ca_9_6_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_9_6 u_ca_9_6_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_9_6 u_ca_9_6_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_9_6 u_ca_9_6_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_9_6 u_ca_9_6_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_9_6 u_ca_9_6_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_9_6 u_ca_9_6_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_9_6 u_ca_9_6_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_9_6 u_ca_9_6_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_9_6 u_ca_9_6_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_9_6 u_ca_9_6_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_9_6 u_ca_9_6_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_9_6 u_ca_9_6_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_9_6 u_ca_9_6_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_9_6 u_ca_9_6_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_9_6 u_ca_9_6_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_9_6 u_ca_9_6_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_9_6 u_ca_9_6_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_9_6 u_ca_9_6_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_9_6 u_ca_9_6_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_9_6 u_ca_9_6_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_9_6 u_ca_9_6_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_9_6 u_ca_9_6_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_9_6 u_ca_9_6_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_9_6 u_ca_9_6_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_9_6 u_ca_9_6_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_9_6 u_ca_9_6_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_9_6 u_ca_9_6_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_9_6 u_ca_9_6_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_9_6 u_ca_9_6_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_9_6 u_ca_9_6_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_9_6 u_ca_9_6_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_9_6 u_ca_9_6_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_9_6 u_ca_9_6_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_9_6 u_ca_9_6_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_9_6 u_ca_9_6_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_9_6 u_ca_9_6_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_9_6 u_ca_9_6_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_9_6 u_ca_9_6_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_9_6 u_ca_9_6_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_9_6 u_ca_9_6_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_9_6 u_ca_9_6_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_9_6 u_ca_9_6_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_9_6 u_ca_9_6_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_9_6 u_ca_9_6_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_9_6 u_ca_9_6_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_9_6 u_ca_9_6_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_9_6 u_ca_9_6_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_9_6 u_ca_9_6_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_9_6 u_ca_9_6_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_9_6 u_ca_9_6_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_9_6 u_ca_9_6_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_9_6 u_ca_9_6_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_9_6 u_ca_9_6_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_9_6 u_ca_9_6_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_9_6 u_ca_9_6_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_9_6 u_ca_9_6_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_9_6 u_ca_9_6_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_9_6 u_ca_9_6_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_9_6 u_ca_9_6_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_9_6 u_ca_9_6_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_9_6 u_ca_9_6_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_9_6 u_ca_9_6_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_9_6 u_ca_9_6_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_9_6 u_ca_9_6_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_9_6 u_ca_9_6_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_9_6 u_ca_9_6_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_9_6 u_ca_9_6_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_9_6 u_ca_9_6_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_9_6 u_ca_9_6_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_9_6 u_ca_9_6_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_9_6 u_ca_9_6_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_9_6 u_ca_9_6_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_9_6 u_ca_9_6_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_9_6 u_ca_9_6_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_9_6 u_ca_9_6_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_9_6 u_ca_9_6_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_9_6 u_ca_9_6_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_9_6 u_ca_9_6_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_9_6 u_ca_9_6_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_9_6 u_ca_9_6_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_9_6 u_ca_9_6_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_9_6 u_ca_9_6_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_9_6 u_ca_9_6_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_9_6 u_ca_9_6_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_9_6 u_ca_9_6_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_9_6 u_ca_9_6_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_9_6 u_ca_9_6_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_9_6 u_ca_9_6_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_9_6 u_ca_9_6_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_9_6 u_ca_9_6_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_9_6 u_ca_9_6_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_9_6 u_ca_9_6_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_9_6 u_ca_9_6_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_9_6 u_ca_9_6_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_9_6 u_ca_9_6_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_9_6 u_ca_9_6_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_9_6 u_ca_9_6_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_9_6 u_ca_9_6_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_9_6 u_ca_9_6_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_9_6 u_ca_9_6_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_9_6 u_ca_9_6_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_9_6 u_ca_9_6_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_9_6 u_ca_9_6_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_9_6 u_ca_9_6_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_9_6 u_ca_9_6_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_9_6 u_ca_9_6_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_9_6 u_ca_9_6_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_9_6 u_ca_9_6_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_9_6 u_ca_9_6_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_9_6 u_ca_9_6_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_9_6 u_ca_9_6_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_9_6 u_ca_9_6_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_9_6 u_ca_9_6_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_9_6 u_ca_9_6_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_9_6 u_ca_9_6_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_9_6 u_ca_9_6_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_9_6 u_ca_9_6_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_9_6 u_ca_9_6_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_9_6 u_ca_9_6_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_9_6 u_ca_9_6_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_9_6 u_ca_9_6_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_9_6 u_ca_9_6_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_9_6 u_ca_9_6_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_9_6 u_ca_9_6_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_9_6 u_ca_9_6_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_9_6 u_ca_9_6_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_9_6 u_ca_9_6_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_9_6 u_ca_9_6_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_9_6 u_ca_9_6_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_9_6 u_ca_9_6_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_9_6 u_ca_9_6_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_9_6 u_ca_9_6_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_9_6 u_ca_9_6_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_9_6 u_ca_9_6_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_9_6 u_ca_9_6_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_9_6 u_ca_9_6_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_9_6 u_ca_9_6_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_9_6 u_ca_9_6_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_9_6 u_ca_9_6_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_9_6 u_ca_9_6_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_9_6 u_ca_9_6_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_9_6 u_ca_9_6_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_9_6 u_ca_9_6_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_9_6 u_ca_9_6_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_9_6 u_ca_9_6_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_9_6 u_ca_9_6_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_9_6 u_ca_9_6_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_9_6 u_ca_9_6_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_9_6 u_ca_9_6_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_9_6 u_ca_9_6_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_9_6 u_ca_9_6_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_9_6 u_ca_9_6_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_9_6 u_ca_9_6_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_9_6 u_ca_9_6_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_9_6 u_ca_9_6_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_9_6 u_ca_9_6_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_9_6 u_ca_9_6_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_9_6 u_ca_9_6_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_9_6 u_ca_9_6_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_9_6 u_ca_9_6_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_9_6 u_ca_9_6_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_9_6 u_ca_9_6_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_9_6 u_ca_9_6_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_9_6 u_ca_9_6_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_9_6 u_ca_9_6_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_9_6 u_ca_9_6_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_9_6 u_ca_9_6_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_9_6 u_ca_9_6_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_9_6 u_ca_9_6_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_9_6 u_ca_9_6_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_9_6 u_ca_9_6_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_9_6 u_ca_9_6_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_9_6 u_ca_9_6_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_9_6 u_ca_9_6_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_9_6 u_ca_9_6_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_9_6 u_ca_9_6_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_9_6 u_ca_9_6_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_9_6 u_ca_9_6_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_9_6 u_ca_9_6_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_9_6 u_ca_9_6_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_9_6 u_ca_9_6_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_9_6 u_ca_9_6_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_9_6 u_ca_9_6_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_9_6 u_ca_9_6_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_9_6 u_ca_9_6_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_9_6 u_ca_9_6_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_9_6 u_ca_9_6_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_9_6 u_ca_9_6_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_9_6 u_ca_9_6_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_9_6 u_ca_9_6_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_9_6 u_ca_9_6_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_9_6 u_ca_9_6_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_9_6 u_ca_9_6_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_9_6 u_ca_9_6_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_9_6 u_ca_9_6_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_9_6 u_ca_9_6_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_9_6 u_ca_9_6_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_9_6 u_ca_9_6_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_9_6 u_ca_9_6_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_9_6 u_ca_9_6_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_9_6 u_ca_9_6_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_9_6 u_ca_9_6_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_9_6 u_ca_9_6_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_9_6 u_ca_9_6_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_9_6 u_ca_9_6_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_9_6 u_ca_9_6_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_9_6 u_ca_9_6_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_9_6 u_ca_9_6_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_9_6 u_ca_9_6_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_9_6 u_ca_9_6_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_9_6 u_ca_9_6_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_9_6 u_ca_9_6_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_9_6 u_ca_9_6_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_9_6 u_ca_9_6_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_9_6 u_ca_9_6_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_9_6 u_ca_9_6_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_9_6 u_ca_9_6_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_9_6 u_ca_9_6_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_9_6 u_ca_9_6_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_9_6 u_ca_9_6_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_9_6 u_ca_9_6_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_9_6 u_ca_9_6_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_9_6 u_ca_9_6_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_9_6 u_ca_9_6_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_9_6 u_ca_9_6_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_9_6 u_ca_9_6_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_9_6 u_ca_9_6_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_9_6 u_ca_9_6_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_9_6 u_ca_9_6_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_9_6 u_ca_9_6_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_9_6 u_ca_9_6_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_9_6 u_ca_9_6_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_9_6 u_ca_9_6_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_9_6 u_ca_9_6_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_9_6 u_ca_9_6_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_9_6 u_ca_9_6_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_9_6 u_ca_9_6_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_9_6 u_ca_9_6_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_9_6 u_ca_9_6_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_9_6 u_ca_9_6_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_9_6 u_ca_9_6_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_9_6 u_ca_9_6_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_9_6 u_ca_9_6_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_9_6 u_ca_9_6_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_9_6 u_ca_9_6_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_9_6 u_ca_9_6_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_9_6 u_ca_9_6_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_9_6 u_ca_9_6_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_9_6 u_ca_9_6_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_9_6 u_ca_9_6_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_9_6 u_ca_9_6_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_9_6 u_ca_9_6_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_9_6 u_ca_9_6_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_9_6 u_ca_9_6_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_9_6 u_ca_9_6_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_9_6 u_ca_9_6_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_9_6 u_ca_9_6_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_9_6 u_ca_9_6_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_9_6 u_ca_9_6_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_9_6 u_ca_9_6_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_9_6 u_ca_9_6_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_9_6 u_ca_9_6_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_9_6 u_ca_9_6_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_9_6 u_ca_9_6_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_9_6 u_ca_9_6_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_9_6 u_ca_9_6_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_9_6 u_ca_9_6_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_9_6 u_ca_9_6_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_9_6 u_ca_9_6_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_9_6 u_ca_9_6_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_9_6 u_ca_9_6_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_9_6 u_ca_9_6_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_9_6 u_ca_9_6_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_9_6 u_ca_9_6_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_9_6 u_ca_9_6_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_9_6 u_ca_9_6_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_9_6 u_ca_9_6_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_9_6 u_ca_9_6_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_9_6 u_ca_9_6_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_9_6 u_ca_9_6_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_9_6 u_ca_9_6_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_9_6 u_ca_9_6_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_9_6 u_ca_9_6_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_9_6 u_ca_9_6_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_9_6 u_ca_9_6_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_9_6 u_ca_9_6_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_9_6 u_ca_9_6_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_9_6 u_ca_9_6_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_9_6 u_ca_9_6_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_9_6 u_ca_9_6_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_9_6 u_ca_9_6_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_9_6 u_ca_9_6_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_9_6 u_ca_9_6_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_9_6 u_ca_9_6_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_9_6 u_ca_9_6_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_9_6 u_ca_9_6_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_9_6 u_ca_9_6_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_9_6 u_ca_9_6_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_9_6 u_ca_9_6_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_9_6 u_ca_9_6_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_9_6 u_ca_9_6_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_9_6 u_ca_9_6_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_9_6 u_ca_9_6_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_9_6 u_ca_9_6_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_9_6 u_ca_9_6_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_9_6 u_ca_9_6_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_9_6 u_ca_9_6_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_9_6 u_ca_9_6_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_9_6 u_ca_9_6_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_9_6 u_ca_9_6_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_9_6 u_ca_9_6_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_9_6 u_ca_9_6_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_9_6 u_ca_9_6_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_9_6 u_ca_9_6_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_9_6 u_ca_9_6_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_9_6 u_ca_9_6_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_9_6 u_ca_9_6_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_9_6 u_ca_9_6_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_9_6 u_ca_9_6_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_9_6 u_ca_9_6_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_9_6 u_ca_9_6_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_9_6 u_ca_9_6_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_9_6 u_ca_9_6_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_9_6 u_ca_9_6_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_9_6 u_ca_9_6_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_9_6 u_ca_9_6_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_9_6 u_ca_9_6_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_9_6 u_ca_9_6_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_9_6 u_ca_9_6_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_9_6 u_ca_9_6_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_9_6 u_ca_9_6_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_9_6 u_ca_9_6_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_9_6 u_ca_9_6_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_9_6 u_ca_9_6_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_9_6 u_ca_9_6_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_9_6 u_ca_9_6_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_9_6 u_ca_9_6_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_9_6 u_ca_9_6_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_9_6 u_ca_9_6_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_9_6 u_ca_9_6_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_9_6 u_ca_9_6_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_9_6 u_ca_9_6_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_9_6 u_ca_9_6_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_9_6 u_ca_9_6_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_9_6 u_ca_9_6_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_9_6 u_ca_9_6_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_9_6 u_ca_9_6_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_9_6 u_ca_9_6_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_9_6 u_ca_9_6_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_9_6 u_ca_9_6_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_9_6 u_ca_9_6_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_9_6 u_ca_9_6_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_9_6 u_ca_9_6_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_9_6 u_ca_9_6_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_9_6 u_ca_9_6_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_9_6 u_ca_9_6_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_9_6 u_ca_9_6_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_9_6 u_ca_9_6_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_9_6 u_ca_9_6_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_9_6 u_ca_9_6_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_9_6 u_ca_9_6_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_9_6 u_ca_9_6_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_9_6 u_ca_9_6_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_9_6 u_ca_9_6_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_9_6 u_ca_9_6_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_9_6 u_ca_9_6_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_9_6 u_ca_9_6_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_9_6 u_ca_9_6_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_9_6 u_ca_9_6_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_9_6 u_ca_9_6_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_9_6 u_ca_9_6_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_9_6 u_ca_9_6_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_9_6 u_ca_9_6_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_9_6 u_ca_9_6_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_9_6 u_ca_9_6_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_9_6 u_ca_9_6_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_9_6 u_ca_9_6_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_9_6 u_ca_9_6_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_9_6 u_ca_9_6_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_9_6 u_ca_9_6_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_9_6 u_ca_9_6_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_9_6 u_ca_9_6_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_9_6 u_ca_9_6_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_9_6 u_ca_9_6_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_9_6 u_ca_9_6_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_9_6 u_ca_9_6_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_9_6 u_ca_9_6_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_9_6 u_ca_9_6_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_9_6 u_ca_9_6_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_9_6 u_ca_9_6_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_9_6 u_ca_9_6_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_9_6 u_ca_9_6_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_9_6 u_ca_9_6_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_9_6 u_ca_9_6_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_9_6 u_ca_9_6_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_9_6 u_ca_9_6_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_9_6 u_ca_9_6_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_9_6 u_ca_9_6_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_9_6 u_ca_9_6_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_9_6 u_ca_9_6_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_9_6 u_ca_9_6_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_9_6 u_ca_9_6_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_9_6 u_ca_9_6_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_9_6 u_ca_9_6_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_9_6 u_ca_9_6_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_9_6 u_ca_9_6_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_9_6 u_ca_9_6_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_9_6 u_ca_9_6_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_9_6 u_ca_9_6_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_9_6 u_ca_9_6_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_9_6 u_ca_9_6_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_9_6 u_ca_9_6_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_9_6 u_ca_9_6_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_9_6 u_ca_9_6_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_9_6 u_ca_9_6_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_9_6 u_ca_9_6_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_9_6 u_ca_9_6_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_9_6 u_ca_9_6_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_9_6 u_ca_9_6_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_9_6 u_ca_9_6_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_9_6 u_ca_9_6_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_9_6 u_ca_9_6_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_9_6 u_ca_9_6_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_9_6 u_ca_9_6_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_9_6 u_ca_9_6_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_9_6 u_ca_9_6_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_9_6 u_ca_9_6_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_9_6 u_ca_9_6_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_9_6 u_ca_9_6_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_9_6 u_ca_9_6_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_9_6 u_ca_9_6_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_9_6 u_ca_9_6_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_9_6 u_ca_9_6_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_9_6 u_ca_9_6_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_9_6 u_ca_9_6_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_9_6 u_ca_9_6_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_9_6 u_ca_9_6_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_9_6 u_ca_9_6_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_9_6 u_ca_9_6_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_9_6 u_ca_9_6_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_9_6 u_ca_9_6_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_9_6 u_ca_9_6_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_9_6 u_ca_9_6_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_9_6 u_ca_9_6_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_9_6 u_ca_9_6_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_9_6 u_ca_9_6_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_9_6 u_ca_9_6_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_9_6 u_ca_9_6_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_9_6 u_ca_9_6_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_9_6 u_ca_9_6_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_9_6 u_ca_9_6_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_9_6 u_ca_9_6_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_9_6 u_ca_9_6_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_9_6 u_ca_9_6_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_9_6 u_ca_9_6_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_9_6 u_ca_9_6_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_9_6 u_ca_9_6_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_9_6 u_ca_9_6_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_9_6 u_ca_9_6_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_9_6 u_ca_9_6_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_9_6 u_ca_9_6_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_9_6 u_ca_9_6_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_9_6 u_ca_9_6_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_9_6 u_ca_9_6_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_9_6 u_ca_9_6_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_9_6 u_ca_9_6_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_9_6 u_ca_9_6_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_9_6 u_ca_9_6_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_9_6 u_ca_9_6_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_9_6 u_ca_9_6_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_9_6 u_ca_9_6_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_9_6 u_ca_9_6_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_9_6 u_ca_9_6_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_9_6 u_ca_9_6_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_9_6 u_ca_9_6_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_9_6 u_ca_9_6_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_9_6 u_ca_9_6_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_9_6 u_ca_9_6_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_9_6 u_ca_9_6_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_9_6 u_ca_9_6_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_9_6 u_ca_9_6_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_9_6 u_ca_9_6_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_9_6 u_ca_9_6_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_9_6 u_ca_9_6_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_9_6 u_ca_9_6_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_9_6 u_ca_9_6_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_9_6 u_ca_9_6_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_9_6 u_ca_9_6_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_9_6 u_ca_9_6_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_9_6 u_ca_9_6_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_9_6 u_ca_9_6_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_9_6 u_ca_9_6_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_9_6 u_ca_9_6_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_9_6 u_ca_9_6_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_9_6 u_ca_9_6_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_9_6 u_ca_9_6_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_9_6 u_ca_9_6_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_9_6 u_ca_9_6_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_9_6 u_ca_9_6_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_9_6 u_ca_9_6_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_9_6 u_ca_9_6_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_9_6 u_ca_9_6_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_9_6 u_ca_9_6_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_9_6 u_ca_9_6_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_9_6 u_ca_9_6_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_9_6 u_ca_9_6_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_9_6 u_ca_9_6_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_9_6 u_ca_9_6_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_9_6 u_ca_9_6_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_9_6 u_ca_9_6_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_9_6 u_ca_9_6_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_9_6 u_ca_9_6_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_9_6 u_ca_9_6_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_9_6 u_ca_9_6_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_9_6 u_ca_9_6_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_9_6 u_ca_9_6_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_9_6 u_ca_9_6_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_9_6 u_ca_9_6_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_9_6 u_ca_9_6_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_9_6 u_ca_9_6_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_9_6 u_ca_9_6_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));
compressor_9_6 u_ca_9_6_1030(.d_in(u_ca_in_1030), .d_out(u_ca_out_1030));
compressor_9_6 u_ca_9_6_1031(.d_in(u_ca_in_1031), .d_out(u_ca_out_1031));
compressor_9_6 u_ca_9_6_1032(.d_in(u_ca_in_1032), .d_out(u_ca_out_1032));
compressor_9_6 u_ca_9_6_1033(.d_in(u_ca_in_1033), .d_out(u_ca_out_1033));
compressor_9_6 u_ca_9_6_1034(.d_in(u_ca_in_1034), .d_out(u_ca_out_1034));
compressor_9_6 u_ca_9_6_1035(.d_in(u_ca_in_1035), .d_out(u_ca_out_1035));
compressor_9_6 u_ca_9_6_1036(.d_in(u_ca_in_1036), .d_out(u_ca_out_1036));
compressor_9_6 u_ca_9_6_1037(.d_in(u_ca_in_1037), .d_out(u_ca_out_1037));
compressor_9_6 u_ca_9_6_1038(.d_in(u_ca_in_1038), .d_out(u_ca_out_1038));
compressor_9_6 u_ca_9_6_1039(.d_in(u_ca_in_1039), .d_out(u_ca_out_1039));
compressor_9_6 u_ca_9_6_1040(.d_in(u_ca_in_1040), .d_out(u_ca_out_1040));
compressor_9_6 u_ca_9_6_1041(.d_in(u_ca_in_1041), .d_out(u_ca_out_1041));
compressor_9_6 u_ca_9_6_1042(.d_in(u_ca_in_1042), .d_out(u_ca_out_1042));
compressor_9_6 u_ca_9_6_1043(.d_in(u_ca_in_1043), .d_out(u_ca_out_1043));
compressor_9_6 u_ca_9_6_1044(.d_in(u_ca_in_1044), .d_out(u_ca_out_1044));
compressor_9_6 u_ca_9_6_1045(.d_in(u_ca_in_1045), .d_out(u_ca_out_1045));
compressor_9_6 u_ca_9_6_1046(.d_in(u_ca_in_1046), .d_out(u_ca_out_1046));
compressor_9_6 u_ca_9_6_1047(.d_in(u_ca_in_1047), .d_out(u_ca_out_1047));
compressor_9_6 u_ca_9_6_1048(.d_in(u_ca_in_1048), .d_out(u_ca_out_1048));
compressor_9_6 u_ca_9_6_1049(.d_in(u_ca_in_1049), .d_out(u_ca_out_1049));
compressor_9_6 u_ca_9_6_1050(.d_in(u_ca_in_1050), .d_out(u_ca_out_1050));
compressor_9_6 u_ca_9_6_1051(.d_in(u_ca_in_1051), .d_out(u_ca_out_1051));
compressor_9_6 u_ca_9_6_1052(.d_in(u_ca_in_1052), .d_out(u_ca_out_1052));
compressor_9_6 u_ca_9_6_1053(.d_in(u_ca_in_1053), .d_out(u_ca_out_1053));
compressor_9_6 u_ca_9_6_1054(.d_in(u_ca_in_1054), .d_out(u_ca_out_1054));
compressor_9_6 u_ca_9_6_1055(.d_in(u_ca_in_1055), .d_out(u_ca_out_1055));
compressor_9_6 u_ca_9_6_1056(.d_in(u_ca_in_1056), .d_out(u_ca_out_1056));
compressor_9_6 u_ca_9_6_1057(.d_in(u_ca_in_1057), .d_out(u_ca_out_1057));
compressor_9_6 u_ca_9_6_1058(.d_in(u_ca_in_1058), .d_out(u_ca_out_1058));
compressor_9_6 u_ca_9_6_1059(.d_in(u_ca_in_1059), .d_out(u_ca_out_1059));
compressor_9_6 u_ca_9_6_1060(.d_in(u_ca_in_1060), .d_out(u_ca_out_1060));
compressor_9_6 u_ca_9_6_1061(.d_in(u_ca_in_1061), .d_out(u_ca_out_1061));
compressor_9_6 u_ca_9_6_1062(.d_in(u_ca_in_1062), .d_out(u_ca_out_1062));
compressor_9_6 u_ca_9_6_1063(.d_in(u_ca_in_1063), .d_out(u_ca_out_1063));
compressor_9_6 u_ca_9_6_1064(.d_in(u_ca_in_1064), .d_out(u_ca_out_1064));
compressor_9_6 u_ca_9_6_1065(.d_in(u_ca_in_1065), .d_out(u_ca_out_1065));
compressor_9_6 u_ca_9_6_1066(.d_in(u_ca_in_1066), .d_out(u_ca_out_1066));
compressor_9_6 u_ca_9_6_1067(.d_in(u_ca_in_1067), .d_out(u_ca_out_1067));
compressor_9_6 u_ca_9_6_1068(.d_in(u_ca_in_1068), .d_out(u_ca_out_1068));
compressor_9_6 u_ca_9_6_1069(.d_in(u_ca_in_1069), .d_out(u_ca_out_1069));
compressor_9_6 u_ca_9_6_1070(.d_in(u_ca_in_1070), .d_out(u_ca_out_1070));
compressor_9_6 u_ca_9_6_1071(.d_in(u_ca_in_1071), .d_out(u_ca_out_1071));
compressor_9_6 u_ca_9_6_1072(.d_in(u_ca_in_1072), .d_out(u_ca_out_1072));
compressor_9_6 u_ca_9_6_1073(.d_in(u_ca_in_1073), .d_out(u_ca_out_1073));
compressor_9_6 u_ca_9_6_1074(.d_in(u_ca_in_1074), .d_out(u_ca_out_1074));
compressor_9_6 u_ca_9_6_1075(.d_in(u_ca_in_1075), .d_out(u_ca_out_1075));
compressor_9_6 u_ca_9_6_1076(.d_in(u_ca_in_1076), .d_out(u_ca_out_1076));
compressor_9_6 u_ca_9_6_1077(.d_in(u_ca_in_1077), .d_out(u_ca_out_1077));
compressor_9_6 u_ca_9_6_1078(.d_in(u_ca_in_1078), .d_out(u_ca_out_1078));
compressor_9_6 u_ca_9_6_1079(.d_in(u_ca_in_1079), .d_out(u_ca_out_1079));
compressor_9_6 u_ca_9_6_1080(.d_in(u_ca_in_1080), .d_out(u_ca_out_1080));
compressor_9_6 u_ca_9_6_1081(.d_in(u_ca_in_1081), .d_out(u_ca_out_1081));
compressor_9_6 u_ca_9_6_1082(.d_in(u_ca_in_1082), .d_out(u_ca_out_1082));
compressor_9_6 u_ca_9_6_1083(.d_in(u_ca_in_1083), .d_out(u_ca_out_1083));
compressor_9_6 u_ca_9_6_1084(.d_in(u_ca_in_1084), .d_out(u_ca_out_1084));
compressor_9_6 u_ca_9_6_1085(.d_in(u_ca_in_1085), .d_out(u_ca_out_1085));
compressor_9_6 u_ca_9_6_1086(.d_in(u_ca_in_1086), .d_out(u_ca_out_1086));
compressor_9_6 u_ca_9_6_1087(.d_in(u_ca_in_1087), .d_out(u_ca_out_1087));
compressor_9_6 u_ca_9_6_1088(.d_in(u_ca_in_1088), .d_out(u_ca_out_1088));
compressor_9_6 u_ca_9_6_1089(.d_in(u_ca_in_1089), .d_out(u_ca_out_1089));
compressor_9_6 u_ca_9_6_1090(.d_in(u_ca_in_1090), .d_out(u_ca_out_1090));
compressor_9_6 u_ca_9_6_1091(.d_in(u_ca_in_1091), .d_out(u_ca_out_1091));
compressor_9_6 u_ca_9_6_1092(.d_in(u_ca_in_1092), .d_out(u_ca_out_1092));
compressor_9_6 u_ca_9_6_1093(.d_in(u_ca_in_1093), .d_out(u_ca_out_1093));
compressor_9_6 u_ca_9_6_1094(.d_in(u_ca_in_1094), .d_out(u_ca_out_1094));
compressor_9_6 u_ca_9_6_1095(.d_in(u_ca_in_1095), .d_out(u_ca_out_1095));
compressor_9_6 u_ca_9_6_1096(.d_in(u_ca_in_1096), .d_out(u_ca_out_1096));
compressor_9_6 u_ca_9_6_1097(.d_in(u_ca_in_1097), .d_out(u_ca_out_1097));
compressor_9_6 u_ca_9_6_1098(.d_in(u_ca_in_1098), .d_out(u_ca_out_1098));
compressor_9_6 u_ca_9_6_1099(.d_in(u_ca_in_1099), .d_out(u_ca_out_1099));
compressor_9_6 u_ca_9_6_1100(.d_in(u_ca_in_1100), .d_out(u_ca_out_1100));
compressor_9_6 u_ca_9_6_1101(.d_in(u_ca_in_1101), .d_out(u_ca_out_1101));
compressor_9_6 u_ca_9_6_1102(.d_in(u_ca_in_1102), .d_out(u_ca_out_1102));
compressor_9_6 u_ca_9_6_1103(.d_in(u_ca_in_1103), .d_out(u_ca_out_1103));
compressor_9_6 u_ca_9_6_1104(.d_in(u_ca_in_1104), .d_out(u_ca_out_1104));
compressor_9_6 u_ca_9_6_1105(.d_in(u_ca_in_1105), .d_out(u_ca_out_1105));
compressor_9_6 u_ca_9_6_1106(.d_in(u_ca_in_1106), .d_out(u_ca_out_1106));
compressor_9_6 u_ca_9_6_1107(.d_in(u_ca_in_1107), .d_out(u_ca_out_1107));
compressor_9_6 u_ca_9_6_1108(.d_in(u_ca_in_1108), .d_out(u_ca_out_1108));
compressor_9_6 u_ca_9_6_1109(.d_in(u_ca_in_1109), .d_out(u_ca_out_1109));
compressor_9_6 u_ca_9_6_1110(.d_in(u_ca_in_1110), .d_out(u_ca_out_1110));
compressor_9_6 u_ca_9_6_1111(.d_in(u_ca_in_1111), .d_out(u_ca_out_1111));
compressor_9_6 u_ca_9_6_1112(.d_in(u_ca_in_1112), .d_out(u_ca_out_1112));
compressor_9_6 u_ca_9_6_1113(.d_in(u_ca_in_1113), .d_out(u_ca_out_1113));
compressor_9_6 u_ca_9_6_1114(.d_in(u_ca_in_1114), .d_out(u_ca_out_1114));
compressor_9_6 u_ca_9_6_1115(.d_in(u_ca_in_1115), .d_out(u_ca_out_1115));
compressor_9_6 u_ca_9_6_1116(.d_in(u_ca_in_1116), .d_out(u_ca_out_1116));
compressor_9_6 u_ca_9_6_1117(.d_in(u_ca_in_1117), .d_out(u_ca_out_1117));
compressor_9_6 u_ca_9_6_1118(.d_in(u_ca_in_1118), .d_out(u_ca_out_1118));
compressor_9_6 u_ca_9_6_1119(.d_in(u_ca_in_1119), .d_out(u_ca_out_1119));
compressor_9_6 u_ca_9_6_1120(.d_in(u_ca_in_1120), .d_out(u_ca_out_1120));
compressor_9_6 u_ca_9_6_1121(.d_in(u_ca_in_1121), .d_out(u_ca_out_1121));
compressor_9_6 u_ca_9_6_1122(.d_in(u_ca_in_1122), .d_out(u_ca_out_1122));
compressor_9_6 u_ca_9_6_1123(.d_in(u_ca_in_1123), .d_out(u_ca_out_1123));
compressor_9_6 u_ca_9_6_1124(.d_in(u_ca_in_1124), .d_out(u_ca_out_1124));
compressor_9_6 u_ca_9_6_1125(.d_in(u_ca_in_1125), .d_out(u_ca_out_1125));
compressor_9_6 u_ca_9_6_1126(.d_in(u_ca_in_1126), .d_out(u_ca_out_1126));
compressor_9_6 u_ca_9_6_1127(.d_in(u_ca_in_1127), .d_out(u_ca_out_1127));
compressor_9_6 u_ca_9_6_1128(.d_in(u_ca_in_1128), .d_out(u_ca_out_1128));
compressor_9_6 u_ca_9_6_1129(.d_in(u_ca_in_1129), .d_out(u_ca_out_1129));
compressor_9_6 u_ca_9_6_1130(.d_in(u_ca_in_1130), .d_out(u_ca_out_1130));
compressor_9_6 u_ca_9_6_1131(.d_in(u_ca_in_1131), .d_out(u_ca_out_1131));
compressor_9_6 u_ca_9_6_1132(.d_in(u_ca_in_1132), .d_out(u_ca_out_1132));
compressor_9_6 u_ca_9_6_1133(.d_in(u_ca_in_1133), .d_out(u_ca_out_1133));
compressor_9_6 u_ca_9_6_1134(.d_in(u_ca_in_1134), .d_out(u_ca_out_1134));
compressor_9_6 u_ca_9_6_1135(.d_in(u_ca_in_1135), .d_out(u_ca_out_1135));
compressor_9_6 u_ca_9_6_1136(.d_in(u_ca_in_1136), .d_out(u_ca_out_1136));
compressor_9_6 u_ca_9_6_1137(.d_in(u_ca_in_1137), .d_out(u_ca_out_1137));
compressor_9_6 u_ca_9_6_1138(.d_in(u_ca_in_1138), .d_out(u_ca_out_1138));
compressor_9_6 u_ca_9_6_1139(.d_in(u_ca_in_1139), .d_out(u_ca_out_1139));
compressor_9_6 u_ca_9_6_1140(.d_in(u_ca_in_1140), .d_out(u_ca_out_1140));
compressor_9_6 u_ca_9_6_1141(.d_in(u_ca_in_1141), .d_out(u_ca_out_1141));
compressor_9_6 u_ca_9_6_1142(.d_in(u_ca_in_1142), .d_out(u_ca_out_1142));
compressor_9_6 u_ca_9_6_1143(.d_in(u_ca_in_1143), .d_out(u_ca_out_1143));
compressor_9_6 u_ca_9_6_1144(.d_in(u_ca_in_1144), .d_out(u_ca_out_1144));
compressor_9_6 u_ca_9_6_1145(.d_in(u_ca_in_1145), .d_out(u_ca_out_1145));
compressor_9_6 u_ca_9_6_1146(.d_in(u_ca_in_1146), .d_out(u_ca_out_1146));
compressor_9_6 u_ca_9_6_1147(.d_in(u_ca_in_1147), .d_out(u_ca_out_1147));
compressor_9_6 u_ca_9_6_1148(.d_in(u_ca_in_1148), .d_out(u_ca_out_1148));
compressor_9_6 u_ca_9_6_1149(.d_in(u_ca_in_1149), .d_out(u_ca_out_1149));
compressor_9_6 u_ca_9_6_1150(.d_in(u_ca_in_1150), .d_out(u_ca_out_1150));
compressor_9_6 u_ca_9_6_1151(.d_in(u_ca_in_1151), .d_out(u_ca_out_1151));
compressor_9_6 u_ca_9_6_1152(.d_in(u_ca_in_1152), .d_out(u_ca_out_1152));
compressor_9_6 u_ca_9_6_1153(.d_in(u_ca_in_1153), .d_out(u_ca_out_1153));
compressor_9_6 u_ca_9_6_1154(.d_in(u_ca_in_1154), .d_out(u_ca_out_1154));
compressor_9_6 u_ca_9_6_1155(.d_in(u_ca_in_1155), .d_out(u_ca_out_1155));
compressor_9_6 u_ca_9_6_1156(.d_in(u_ca_in_1156), .d_out(u_ca_out_1156));
compressor_9_6 u_ca_9_6_1157(.d_in(u_ca_in_1157), .d_out(u_ca_out_1157));
compressor_9_6 u_ca_9_6_1158(.d_in(u_ca_in_1158), .d_out(u_ca_out_1158));
compressor_9_6 u_ca_9_6_1159(.d_in(u_ca_in_1159), .d_out(u_ca_out_1159));
compressor_9_6 u_ca_9_6_1160(.d_in(u_ca_in_1160), .d_out(u_ca_out_1160));
compressor_9_6 u_ca_9_6_1161(.d_in(u_ca_in_1161), .d_out(u_ca_out_1161));
compressor_9_6 u_ca_9_6_1162(.d_in(u_ca_in_1162), .d_out(u_ca_out_1162));
compressor_9_6 u_ca_9_6_1163(.d_in(u_ca_in_1163), .d_out(u_ca_out_1163));
compressor_9_6 u_ca_9_6_1164(.d_in(u_ca_in_1164), .d_out(u_ca_out_1164));
compressor_9_6 u_ca_9_6_1165(.d_in(u_ca_in_1165), .d_out(u_ca_out_1165));
compressor_9_6 u_ca_9_6_1166(.d_in(u_ca_in_1166), .d_out(u_ca_out_1166));
compressor_9_6 u_ca_9_6_1167(.d_in(u_ca_in_1167), .d_out(u_ca_out_1167));
compressor_9_6 u_ca_9_6_1168(.d_in(u_ca_in_1168), .d_out(u_ca_out_1168));
compressor_9_6 u_ca_9_6_1169(.d_in(u_ca_in_1169), .d_out(u_ca_out_1169));
compressor_9_6 u_ca_9_6_1170(.d_in(u_ca_in_1170), .d_out(u_ca_out_1170));
compressor_9_6 u_ca_9_6_1171(.d_in(u_ca_in_1171), .d_out(u_ca_out_1171));
compressor_9_6 u_ca_9_6_1172(.d_in(u_ca_in_1172), .d_out(u_ca_out_1172));
compressor_9_6 u_ca_9_6_1173(.d_in(u_ca_in_1173), .d_out(u_ca_out_1173));
compressor_9_6 u_ca_9_6_1174(.d_in(u_ca_in_1174), .d_out(u_ca_out_1174));
compressor_9_6 u_ca_9_6_1175(.d_in(u_ca_in_1175), .d_out(u_ca_out_1175));
compressor_9_6 u_ca_9_6_1176(.d_in(u_ca_in_1176), .d_out(u_ca_out_1176));
compressor_9_6 u_ca_9_6_1177(.d_in(u_ca_in_1177), .d_out(u_ca_out_1177));
compressor_9_6 u_ca_9_6_1178(.d_in(u_ca_in_1178), .d_out(u_ca_out_1178));
compressor_9_6 u_ca_9_6_1179(.d_in(u_ca_in_1179), .d_out(u_ca_out_1179));
compressor_9_6 u_ca_9_6_1180(.d_in(u_ca_in_1180), .d_out(u_ca_out_1180));
compressor_9_6 u_ca_9_6_1181(.d_in(u_ca_in_1181), .d_out(u_ca_out_1181));
compressor_9_6 u_ca_9_6_1182(.d_in(u_ca_in_1182), .d_out(u_ca_out_1182));
compressor_9_6 u_ca_9_6_1183(.d_in(u_ca_in_1183), .d_out(u_ca_out_1183));
compressor_9_6 u_ca_9_6_1184(.d_in(u_ca_in_1184), .d_out(u_ca_out_1184));
compressor_9_6 u_ca_9_6_1185(.d_in(u_ca_in_1185), .d_out(u_ca_out_1185));
compressor_9_6 u_ca_9_6_1186(.d_in(u_ca_in_1186), .d_out(u_ca_out_1186));
compressor_9_6 u_ca_9_6_1187(.d_in(u_ca_in_1187), .d_out(u_ca_out_1187));
compressor_9_6 u_ca_9_6_1188(.d_in(u_ca_in_1188), .d_out(u_ca_out_1188));
compressor_9_6 u_ca_9_6_1189(.d_in(u_ca_in_1189), .d_out(u_ca_out_1189));
compressor_9_6 u_ca_9_6_1190(.d_in(u_ca_in_1190), .d_out(u_ca_out_1190));
compressor_9_6 u_ca_9_6_1191(.d_in(u_ca_in_1191), .d_out(u_ca_out_1191));
compressor_9_6 u_ca_9_6_1192(.d_in(u_ca_in_1192), .d_out(u_ca_out_1192));
compressor_9_6 u_ca_9_6_1193(.d_in(u_ca_in_1193), .d_out(u_ca_out_1193));
compressor_9_6 u_ca_9_6_1194(.d_in(u_ca_in_1194), .d_out(u_ca_out_1194));
compressor_9_6 u_ca_9_6_1195(.d_in(u_ca_in_1195), .d_out(u_ca_out_1195));
compressor_9_6 u_ca_9_6_1196(.d_in(u_ca_in_1196), .d_out(u_ca_out_1196));
compressor_9_6 u_ca_9_6_1197(.d_in(u_ca_in_1197), .d_out(u_ca_out_1197));
compressor_9_6 u_ca_9_6_1198(.d_in(u_ca_in_1198), .d_out(u_ca_out_1198));
compressor_9_6 u_ca_9_6_1199(.d_in(u_ca_in_1199), .d_out(u_ca_out_1199));
compressor_9_6 u_ca_9_6_1200(.d_in(u_ca_in_1200), .d_out(u_ca_out_1200));
compressor_9_6 u_ca_9_6_1201(.d_in(u_ca_in_1201), .d_out(u_ca_out_1201));
compressor_9_6 u_ca_9_6_1202(.d_in(u_ca_in_1202), .d_out(u_ca_out_1202));
compressor_9_6 u_ca_9_6_1203(.d_in(u_ca_in_1203), .d_out(u_ca_out_1203));
compressor_9_6 u_ca_9_6_1204(.d_in(u_ca_in_1204), .d_out(u_ca_out_1204));
compressor_9_6 u_ca_9_6_1205(.d_in(u_ca_in_1205), .d_out(u_ca_out_1205));
compressor_9_6 u_ca_9_6_1206(.d_in(u_ca_in_1206), .d_out(u_ca_out_1206));
compressor_9_6 u_ca_9_6_1207(.d_in(u_ca_in_1207), .d_out(u_ca_out_1207));
compressor_9_6 u_ca_9_6_1208(.d_in(u_ca_in_1208), .d_out(u_ca_out_1208));
compressor_9_6 u_ca_9_6_1209(.d_in(u_ca_in_1209), .d_out(u_ca_out_1209));
compressor_9_6 u_ca_9_6_1210(.d_in(u_ca_in_1210), .d_out(u_ca_out_1210));
compressor_9_6 u_ca_9_6_1211(.d_in(u_ca_in_1211), .d_out(u_ca_out_1211));
compressor_9_6 u_ca_9_6_1212(.d_in(u_ca_in_1212), .d_out(u_ca_out_1212));
compressor_9_6 u_ca_9_6_1213(.d_in(u_ca_in_1213), .d_out(u_ca_out_1213));
compressor_9_6 u_ca_9_6_1214(.d_in(u_ca_in_1214), .d_out(u_ca_out_1214));
compressor_9_6 u_ca_9_6_1215(.d_in(u_ca_in_1215), .d_out(u_ca_out_1215));
compressor_9_6 u_ca_9_6_1216(.d_in(u_ca_in_1216), .d_out(u_ca_out_1216));
compressor_9_6 u_ca_9_6_1217(.d_in(u_ca_in_1217), .d_out(u_ca_out_1217));
compressor_9_6 u_ca_9_6_1218(.d_in(u_ca_in_1218), .d_out(u_ca_out_1218));
compressor_9_6 u_ca_9_6_1219(.d_in(u_ca_in_1219), .d_out(u_ca_out_1219));
compressor_9_6 u_ca_9_6_1220(.d_in(u_ca_in_1220), .d_out(u_ca_out_1220));
compressor_9_6 u_ca_9_6_1221(.d_in(u_ca_in_1221), .d_out(u_ca_out_1221));
compressor_9_6 u_ca_9_6_1222(.d_in(u_ca_in_1222), .d_out(u_ca_out_1222));
compressor_9_6 u_ca_9_6_1223(.d_in(u_ca_in_1223), .d_out(u_ca_out_1223));
compressor_9_6 u_ca_9_6_1224(.d_in(u_ca_in_1224), .d_out(u_ca_out_1224));
compressor_9_6 u_ca_9_6_1225(.d_in(u_ca_in_1225), .d_out(u_ca_out_1225));
compressor_9_6 u_ca_9_6_1226(.d_in(u_ca_in_1226), .d_out(u_ca_out_1226));
compressor_9_6 u_ca_9_6_1227(.d_in(u_ca_in_1227), .d_out(u_ca_out_1227));
compressor_9_6 u_ca_9_6_1228(.d_in(u_ca_in_1228), .d_out(u_ca_out_1228));
compressor_9_6 u_ca_9_6_1229(.d_in(u_ca_in_1229), .d_out(u_ca_out_1229));
compressor_9_6 u_ca_9_6_1230(.d_in(u_ca_in_1230), .d_out(u_ca_out_1230));
compressor_9_6 u_ca_9_6_1231(.d_in(u_ca_in_1231), .d_out(u_ca_out_1231));
compressor_9_6 u_ca_9_6_1232(.d_in(u_ca_in_1232), .d_out(u_ca_out_1232));
compressor_9_6 u_ca_9_6_1233(.d_in(u_ca_in_1233), .d_out(u_ca_out_1233));
compressor_9_6 u_ca_9_6_1234(.d_in(u_ca_in_1234), .d_out(u_ca_out_1234));
compressor_9_6 u_ca_9_6_1235(.d_in(u_ca_in_1235), .d_out(u_ca_out_1235));
compressor_9_6 u_ca_9_6_1236(.d_in(u_ca_in_1236), .d_out(u_ca_out_1236));
compressor_9_6 u_ca_9_6_1237(.d_in(u_ca_in_1237), .d_out(u_ca_out_1237));
compressor_9_6 u_ca_9_6_1238(.d_in(u_ca_in_1238), .d_out(u_ca_out_1238));
compressor_9_6 u_ca_9_6_1239(.d_in(u_ca_in_1239), .d_out(u_ca_out_1239));
compressor_9_6 u_ca_9_6_1240(.d_in(u_ca_in_1240), .d_out(u_ca_out_1240));
compressor_9_6 u_ca_9_6_1241(.d_in(u_ca_in_1241), .d_out(u_ca_out_1241));
compressor_9_6 u_ca_9_6_1242(.d_in(u_ca_in_1242), .d_out(u_ca_out_1242));
compressor_9_6 u_ca_9_6_1243(.d_in(u_ca_in_1243), .d_out(u_ca_out_1243));
compressor_9_6 u_ca_9_6_1244(.d_in(u_ca_in_1244), .d_out(u_ca_out_1244));
compressor_9_6 u_ca_9_6_1245(.d_in(u_ca_in_1245), .d_out(u_ca_out_1245));
compressor_9_6 u_ca_9_6_1246(.d_in(u_ca_in_1246), .d_out(u_ca_out_1246));
compressor_9_6 u_ca_9_6_1247(.d_in(u_ca_in_1247), .d_out(u_ca_out_1247));
compressor_9_6 u_ca_9_6_1248(.d_in(u_ca_in_1248), .d_out(u_ca_out_1248));
compressor_9_6 u_ca_9_6_1249(.d_in(u_ca_in_1249), .d_out(u_ca_out_1249));
compressor_9_6 u_ca_9_6_1250(.d_in(u_ca_in_1250), .d_out(u_ca_out_1250));
compressor_9_6 u_ca_9_6_1251(.d_in(u_ca_in_1251), .d_out(u_ca_out_1251));
compressor_9_6 u_ca_9_6_1252(.d_in(u_ca_in_1252), .d_out(u_ca_out_1252));
compressor_9_6 u_ca_9_6_1253(.d_in(u_ca_in_1253), .d_out(u_ca_out_1253));
compressor_9_6 u_ca_9_6_1254(.d_in(u_ca_in_1254), .d_out(u_ca_out_1254));
compressor_9_6 u_ca_9_6_1255(.d_in(u_ca_in_1255), .d_out(u_ca_out_1255));
compressor_9_6 u_ca_9_6_1256(.d_in(u_ca_in_1256), .d_out(u_ca_out_1256));
compressor_9_6 u_ca_9_6_1257(.d_in(u_ca_in_1257), .d_out(u_ca_out_1257));
compressor_9_6 u_ca_9_6_1258(.d_in(u_ca_in_1258), .d_out(u_ca_out_1258));
compressor_9_6 u_ca_9_6_1259(.d_in(u_ca_in_1259), .d_out(u_ca_out_1259));
compressor_9_6 u_ca_9_6_1260(.d_in(u_ca_in_1260), .d_out(u_ca_out_1260));
compressor_9_6 u_ca_9_6_1261(.d_in(u_ca_in_1261), .d_out(u_ca_out_1261));
compressor_9_6 u_ca_9_6_1262(.d_in(u_ca_in_1262), .d_out(u_ca_out_1262));
compressor_9_6 u_ca_9_6_1263(.d_in(u_ca_in_1263), .d_out(u_ca_out_1263));
compressor_9_6 u_ca_9_6_1264(.d_in(u_ca_in_1264), .d_out(u_ca_out_1264));
compressor_9_6 u_ca_9_6_1265(.d_in(u_ca_in_1265), .d_out(u_ca_out_1265));
compressor_9_6 u_ca_9_6_1266(.d_in(u_ca_in_1266), .d_out(u_ca_out_1266));
compressor_9_6 u_ca_9_6_1267(.d_in(u_ca_in_1267), .d_out(u_ca_out_1267));
compressor_9_6 u_ca_9_6_1268(.d_in(u_ca_in_1268), .d_out(u_ca_out_1268));
compressor_9_6 u_ca_9_6_1269(.d_in(u_ca_in_1269), .d_out(u_ca_out_1269));
compressor_9_6 u_ca_9_6_1270(.d_in(u_ca_in_1270), .d_out(u_ca_out_1270));
compressor_9_6 u_ca_9_6_1271(.d_in(u_ca_in_1271), .d_out(u_ca_out_1271));
compressor_9_6 u_ca_9_6_1272(.d_in(u_ca_in_1272), .d_out(u_ca_out_1272));
compressor_9_6 u_ca_9_6_1273(.d_in(u_ca_in_1273), .d_out(u_ca_out_1273));
compressor_9_6 u_ca_9_6_1274(.d_in(u_ca_in_1274), .d_out(u_ca_out_1274));
compressor_9_6 u_ca_9_6_1275(.d_in(u_ca_in_1275), .d_out(u_ca_out_1275));
compressor_9_6 u_ca_9_6_1276(.d_in(u_ca_in_1276), .d_out(u_ca_out_1276));
compressor_9_6 u_ca_9_6_1277(.d_in(u_ca_in_1277), .d_out(u_ca_out_1277));
compressor_9_6 u_ca_9_6_1278(.d_in(u_ca_in_1278), .d_out(u_ca_out_1278));
compressor_9_6 u_ca_9_6_1279(.d_in(u_ca_in_1279), .d_out(u_ca_out_1279));
compressor_9_6 u_ca_9_6_1280(.d_in(u_ca_in_1280), .d_out(u_ca_out_1280));
compressor_9_6 u_ca_9_6_1281(.d_in(u_ca_in_1281), .d_out(u_ca_out_1281));
compressor_9_6 u_ca_9_6_1282(.d_in(u_ca_in_1282), .d_out(u_ca_out_1282));
compressor_9_6 u_ca_9_6_1283(.d_in(u_ca_in_1283), .d_out(u_ca_out_1283));
compressor_9_6 u_ca_9_6_1284(.d_in(u_ca_in_1284), .d_out(u_ca_out_1284));
compressor_9_6 u_ca_9_6_1285(.d_in(u_ca_in_1285), .d_out(u_ca_out_1285));
compressor_9_6 u_ca_9_6_1286(.d_in(u_ca_in_1286), .d_out(u_ca_out_1286));
compressor_9_6 u_ca_9_6_1287(.d_in(u_ca_in_1287), .d_out(u_ca_out_1287));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{3{1'b0}}, u_ca_out_0[2:0]};
assign col_out_1 = {u_ca_out_1[2:0], u_ca_out_0[5:3]};
assign col_out_2 = {u_ca_out_2[2:0], u_ca_out_1[5:3]};
assign col_out_3 = {u_ca_out_3[2:0], u_ca_out_2[5:3]};
assign col_out_4 = {u_ca_out_4[2:0], u_ca_out_3[5:3]};
assign col_out_5 = {u_ca_out_5[2:0], u_ca_out_4[5:3]};
assign col_out_6 = {u_ca_out_6[2:0], u_ca_out_5[5:3]};
assign col_out_7 = {u_ca_out_7[2:0], u_ca_out_6[5:3]};
assign col_out_8 = {u_ca_out_8[2:0], u_ca_out_7[5:3]};
assign col_out_9 = {u_ca_out_9[2:0], u_ca_out_8[5:3]};
assign col_out_10 = {u_ca_out_10[2:0], u_ca_out_9[5:3]};
assign col_out_11 = {u_ca_out_11[2:0], u_ca_out_10[5:3]};
assign col_out_12 = {u_ca_out_12[2:0], u_ca_out_11[5:3]};
assign col_out_13 = {u_ca_out_13[2:0], u_ca_out_12[5:3]};
assign col_out_14 = {u_ca_out_14[2:0], u_ca_out_13[5:3]};
assign col_out_15 = {u_ca_out_15[2:0], u_ca_out_14[5:3]};
assign col_out_16 = {u_ca_out_16[2:0], u_ca_out_15[5:3]};
assign col_out_17 = {u_ca_out_17[2:0], u_ca_out_16[5:3]};
assign col_out_18 = {u_ca_out_18[2:0], u_ca_out_17[5:3]};
assign col_out_19 = {u_ca_out_19[2:0], u_ca_out_18[5:3]};
assign col_out_20 = {u_ca_out_20[2:0], u_ca_out_19[5:3]};
assign col_out_21 = {u_ca_out_21[2:0], u_ca_out_20[5:3]};
assign col_out_22 = {u_ca_out_22[2:0], u_ca_out_21[5:3]};
assign col_out_23 = {u_ca_out_23[2:0], u_ca_out_22[5:3]};
assign col_out_24 = {u_ca_out_24[2:0], u_ca_out_23[5:3]};
assign col_out_25 = {u_ca_out_25[2:0], u_ca_out_24[5:3]};
assign col_out_26 = {u_ca_out_26[2:0], u_ca_out_25[5:3]};
assign col_out_27 = {u_ca_out_27[2:0], u_ca_out_26[5:3]};
assign col_out_28 = {u_ca_out_28[2:0], u_ca_out_27[5:3]};
assign col_out_29 = {u_ca_out_29[2:0], u_ca_out_28[5:3]};
assign col_out_30 = {u_ca_out_30[2:0], u_ca_out_29[5:3]};
assign col_out_31 = {u_ca_out_31[2:0], u_ca_out_30[5:3]};
assign col_out_32 = {u_ca_out_32[2:0], u_ca_out_31[5:3]};
assign col_out_33 = {u_ca_out_33[2:0], u_ca_out_32[5:3]};
assign col_out_34 = {u_ca_out_34[2:0], u_ca_out_33[5:3]};
assign col_out_35 = {u_ca_out_35[2:0], u_ca_out_34[5:3]};
assign col_out_36 = {u_ca_out_36[2:0], u_ca_out_35[5:3]};
assign col_out_37 = {u_ca_out_37[2:0], u_ca_out_36[5:3]};
assign col_out_38 = {u_ca_out_38[2:0], u_ca_out_37[5:3]};
assign col_out_39 = {u_ca_out_39[2:0], u_ca_out_38[5:3]};
assign col_out_40 = {u_ca_out_40[2:0], u_ca_out_39[5:3]};
assign col_out_41 = {u_ca_out_41[2:0], u_ca_out_40[5:3]};
assign col_out_42 = {u_ca_out_42[2:0], u_ca_out_41[5:3]};
assign col_out_43 = {u_ca_out_43[2:0], u_ca_out_42[5:3]};
assign col_out_44 = {u_ca_out_44[2:0], u_ca_out_43[5:3]};
assign col_out_45 = {u_ca_out_45[2:0], u_ca_out_44[5:3]};
assign col_out_46 = {u_ca_out_46[2:0], u_ca_out_45[5:3]};
assign col_out_47 = {u_ca_out_47[2:0], u_ca_out_46[5:3]};
assign col_out_48 = {u_ca_out_48[2:0], u_ca_out_47[5:3]};
assign col_out_49 = {u_ca_out_49[2:0], u_ca_out_48[5:3]};
assign col_out_50 = {u_ca_out_50[2:0], u_ca_out_49[5:3]};
assign col_out_51 = {u_ca_out_51[2:0], u_ca_out_50[5:3]};
assign col_out_52 = {u_ca_out_52[2:0], u_ca_out_51[5:3]};
assign col_out_53 = {u_ca_out_53[2:0], u_ca_out_52[5:3]};
assign col_out_54 = {u_ca_out_54[2:0], u_ca_out_53[5:3]};
assign col_out_55 = {u_ca_out_55[2:0], u_ca_out_54[5:3]};
assign col_out_56 = {u_ca_out_56[2:0], u_ca_out_55[5:3]};
assign col_out_57 = {u_ca_out_57[2:0], u_ca_out_56[5:3]};
assign col_out_58 = {u_ca_out_58[2:0], u_ca_out_57[5:3]};
assign col_out_59 = {u_ca_out_59[2:0], u_ca_out_58[5:3]};
assign col_out_60 = {u_ca_out_60[2:0], u_ca_out_59[5:3]};
assign col_out_61 = {u_ca_out_61[2:0], u_ca_out_60[5:3]};
assign col_out_62 = {u_ca_out_62[2:0], u_ca_out_61[5:3]};
assign col_out_63 = {u_ca_out_63[2:0], u_ca_out_62[5:3]};
assign col_out_64 = {u_ca_out_64[2:0], u_ca_out_63[5:3]};
assign col_out_65 = {u_ca_out_65[2:0], u_ca_out_64[5:3]};
assign col_out_66 = {u_ca_out_66[2:0], u_ca_out_65[5:3]};
assign col_out_67 = {u_ca_out_67[2:0], u_ca_out_66[5:3]};
assign col_out_68 = {u_ca_out_68[2:0], u_ca_out_67[5:3]};
assign col_out_69 = {u_ca_out_69[2:0], u_ca_out_68[5:3]};
assign col_out_70 = {u_ca_out_70[2:0], u_ca_out_69[5:3]};
assign col_out_71 = {u_ca_out_71[2:0], u_ca_out_70[5:3]};
assign col_out_72 = {u_ca_out_72[2:0], u_ca_out_71[5:3]};
assign col_out_73 = {u_ca_out_73[2:0], u_ca_out_72[5:3]};
assign col_out_74 = {u_ca_out_74[2:0], u_ca_out_73[5:3]};
assign col_out_75 = {u_ca_out_75[2:0], u_ca_out_74[5:3]};
assign col_out_76 = {u_ca_out_76[2:0], u_ca_out_75[5:3]};
assign col_out_77 = {u_ca_out_77[2:0], u_ca_out_76[5:3]};
assign col_out_78 = {u_ca_out_78[2:0], u_ca_out_77[5:3]};
assign col_out_79 = {u_ca_out_79[2:0], u_ca_out_78[5:3]};
assign col_out_80 = {u_ca_out_80[2:0], u_ca_out_79[5:3]};
assign col_out_81 = {u_ca_out_81[2:0], u_ca_out_80[5:3]};
assign col_out_82 = {u_ca_out_82[2:0], u_ca_out_81[5:3]};
assign col_out_83 = {u_ca_out_83[2:0], u_ca_out_82[5:3]};
assign col_out_84 = {u_ca_out_84[2:0], u_ca_out_83[5:3]};
assign col_out_85 = {u_ca_out_85[2:0], u_ca_out_84[5:3]};
assign col_out_86 = {u_ca_out_86[2:0], u_ca_out_85[5:3]};
assign col_out_87 = {u_ca_out_87[2:0], u_ca_out_86[5:3]};
assign col_out_88 = {u_ca_out_88[2:0], u_ca_out_87[5:3]};
assign col_out_89 = {u_ca_out_89[2:0], u_ca_out_88[5:3]};
assign col_out_90 = {u_ca_out_90[2:0], u_ca_out_89[5:3]};
assign col_out_91 = {u_ca_out_91[2:0], u_ca_out_90[5:3]};
assign col_out_92 = {u_ca_out_92[2:0], u_ca_out_91[5:3]};
assign col_out_93 = {u_ca_out_93[2:0], u_ca_out_92[5:3]};
assign col_out_94 = {u_ca_out_94[2:0], u_ca_out_93[5:3]};
assign col_out_95 = {u_ca_out_95[2:0], u_ca_out_94[5:3]};
assign col_out_96 = {u_ca_out_96[2:0], u_ca_out_95[5:3]};
assign col_out_97 = {u_ca_out_97[2:0], u_ca_out_96[5:3]};
assign col_out_98 = {u_ca_out_98[2:0], u_ca_out_97[5:3]};
assign col_out_99 = {u_ca_out_99[2:0], u_ca_out_98[5:3]};
assign col_out_100 = {u_ca_out_100[2:0], u_ca_out_99[5:3]};
assign col_out_101 = {u_ca_out_101[2:0], u_ca_out_100[5:3]};
assign col_out_102 = {u_ca_out_102[2:0], u_ca_out_101[5:3]};
assign col_out_103 = {u_ca_out_103[2:0], u_ca_out_102[5:3]};
assign col_out_104 = {u_ca_out_104[2:0], u_ca_out_103[5:3]};
assign col_out_105 = {u_ca_out_105[2:0], u_ca_out_104[5:3]};
assign col_out_106 = {u_ca_out_106[2:0], u_ca_out_105[5:3]};
assign col_out_107 = {u_ca_out_107[2:0], u_ca_out_106[5:3]};
assign col_out_108 = {u_ca_out_108[2:0], u_ca_out_107[5:3]};
assign col_out_109 = {u_ca_out_109[2:0], u_ca_out_108[5:3]};
assign col_out_110 = {u_ca_out_110[2:0], u_ca_out_109[5:3]};
assign col_out_111 = {u_ca_out_111[2:0], u_ca_out_110[5:3]};
assign col_out_112 = {u_ca_out_112[2:0], u_ca_out_111[5:3]};
assign col_out_113 = {u_ca_out_113[2:0], u_ca_out_112[5:3]};
assign col_out_114 = {u_ca_out_114[2:0], u_ca_out_113[5:3]};
assign col_out_115 = {u_ca_out_115[2:0], u_ca_out_114[5:3]};
assign col_out_116 = {u_ca_out_116[2:0], u_ca_out_115[5:3]};
assign col_out_117 = {u_ca_out_117[2:0], u_ca_out_116[5:3]};
assign col_out_118 = {u_ca_out_118[2:0], u_ca_out_117[5:3]};
assign col_out_119 = {u_ca_out_119[2:0], u_ca_out_118[5:3]};
assign col_out_120 = {u_ca_out_120[2:0], u_ca_out_119[5:3]};
assign col_out_121 = {u_ca_out_121[2:0], u_ca_out_120[5:3]};
assign col_out_122 = {u_ca_out_122[2:0], u_ca_out_121[5:3]};
assign col_out_123 = {u_ca_out_123[2:0], u_ca_out_122[5:3]};
assign col_out_124 = {u_ca_out_124[2:0], u_ca_out_123[5:3]};
assign col_out_125 = {u_ca_out_125[2:0], u_ca_out_124[5:3]};
assign col_out_126 = {u_ca_out_126[2:0], u_ca_out_125[5:3]};
assign col_out_127 = {u_ca_out_127[2:0], u_ca_out_126[5:3]};
assign col_out_128 = {u_ca_out_128[2:0], u_ca_out_127[5:3]};
assign col_out_129 = {u_ca_out_129[2:0], u_ca_out_128[5:3]};
assign col_out_130 = {u_ca_out_130[2:0], u_ca_out_129[5:3]};
assign col_out_131 = {u_ca_out_131[2:0], u_ca_out_130[5:3]};
assign col_out_132 = {u_ca_out_132[2:0], u_ca_out_131[5:3]};
assign col_out_133 = {u_ca_out_133[2:0], u_ca_out_132[5:3]};
assign col_out_134 = {u_ca_out_134[2:0], u_ca_out_133[5:3]};
assign col_out_135 = {u_ca_out_135[2:0], u_ca_out_134[5:3]};
assign col_out_136 = {u_ca_out_136[2:0], u_ca_out_135[5:3]};
assign col_out_137 = {u_ca_out_137[2:0], u_ca_out_136[5:3]};
assign col_out_138 = {u_ca_out_138[2:0], u_ca_out_137[5:3]};
assign col_out_139 = {u_ca_out_139[2:0], u_ca_out_138[5:3]};
assign col_out_140 = {u_ca_out_140[2:0], u_ca_out_139[5:3]};
assign col_out_141 = {u_ca_out_141[2:0], u_ca_out_140[5:3]};
assign col_out_142 = {u_ca_out_142[2:0], u_ca_out_141[5:3]};
assign col_out_143 = {u_ca_out_143[2:0], u_ca_out_142[5:3]};
assign col_out_144 = {u_ca_out_144[2:0], u_ca_out_143[5:3]};
assign col_out_145 = {u_ca_out_145[2:0], u_ca_out_144[5:3]};
assign col_out_146 = {u_ca_out_146[2:0], u_ca_out_145[5:3]};
assign col_out_147 = {u_ca_out_147[2:0], u_ca_out_146[5:3]};
assign col_out_148 = {u_ca_out_148[2:0], u_ca_out_147[5:3]};
assign col_out_149 = {u_ca_out_149[2:0], u_ca_out_148[5:3]};
assign col_out_150 = {u_ca_out_150[2:0], u_ca_out_149[5:3]};
assign col_out_151 = {u_ca_out_151[2:0], u_ca_out_150[5:3]};
assign col_out_152 = {u_ca_out_152[2:0], u_ca_out_151[5:3]};
assign col_out_153 = {u_ca_out_153[2:0], u_ca_out_152[5:3]};
assign col_out_154 = {u_ca_out_154[2:0], u_ca_out_153[5:3]};
assign col_out_155 = {u_ca_out_155[2:0], u_ca_out_154[5:3]};
assign col_out_156 = {u_ca_out_156[2:0], u_ca_out_155[5:3]};
assign col_out_157 = {u_ca_out_157[2:0], u_ca_out_156[5:3]};
assign col_out_158 = {u_ca_out_158[2:0], u_ca_out_157[5:3]};
assign col_out_159 = {u_ca_out_159[2:0], u_ca_out_158[5:3]};
assign col_out_160 = {u_ca_out_160[2:0], u_ca_out_159[5:3]};
assign col_out_161 = {u_ca_out_161[2:0], u_ca_out_160[5:3]};
assign col_out_162 = {u_ca_out_162[2:0], u_ca_out_161[5:3]};
assign col_out_163 = {u_ca_out_163[2:0], u_ca_out_162[5:3]};
assign col_out_164 = {u_ca_out_164[2:0], u_ca_out_163[5:3]};
assign col_out_165 = {u_ca_out_165[2:0], u_ca_out_164[5:3]};
assign col_out_166 = {u_ca_out_166[2:0], u_ca_out_165[5:3]};
assign col_out_167 = {u_ca_out_167[2:0], u_ca_out_166[5:3]};
assign col_out_168 = {u_ca_out_168[2:0], u_ca_out_167[5:3]};
assign col_out_169 = {u_ca_out_169[2:0], u_ca_out_168[5:3]};
assign col_out_170 = {u_ca_out_170[2:0], u_ca_out_169[5:3]};
assign col_out_171 = {u_ca_out_171[2:0], u_ca_out_170[5:3]};
assign col_out_172 = {u_ca_out_172[2:0], u_ca_out_171[5:3]};
assign col_out_173 = {u_ca_out_173[2:0], u_ca_out_172[5:3]};
assign col_out_174 = {u_ca_out_174[2:0], u_ca_out_173[5:3]};
assign col_out_175 = {u_ca_out_175[2:0], u_ca_out_174[5:3]};
assign col_out_176 = {u_ca_out_176[2:0], u_ca_out_175[5:3]};
assign col_out_177 = {u_ca_out_177[2:0], u_ca_out_176[5:3]};
assign col_out_178 = {u_ca_out_178[2:0], u_ca_out_177[5:3]};
assign col_out_179 = {u_ca_out_179[2:0], u_ca_out_178[5:3]};
assign col_out_180 = {u_ca_out_180[2:0], u_ca_out_179[5:3]};
assign col_out_181 = {u_ca_out_181[2:0], u_ca_out_180[5:3]};
assign col_out_182 = {u_ca_out_182[2:0], u_ca_out_181[5:3]};
assign col_out_183 = {u_ca_out_183[2:0], u_ca_out_182[5:3]};
assign col_out_184 = {u_ca_out_184[2:0], u_ca_out_183[5:3]};
assign col_out_185 = {u_ca_out_185[2:0], u_ca_out_184[5:3]};
assign col_out_186 = {u_ca_out_186[2:0], u_ca_out_185[5:3]};
assign col_out_187 = {u_ca_out_187[2:0], u_ca_out_186[5:3]};
assign col_out_188 = {u_ca_out_188[2:0], u_ca_out_187[5:3]};
assign col_out_189 = {u_ca_out_189[2:0], u_ca_out_188[5:3]};
assign col_out_190 = {u_ca_out_190[2:0], u_ca_out_189[5:3]};
assign col_out_191 = {u_ca_out_191[2:0], u_ca_out_190[5:3]};
assign col_out_192 = {u_ca_out_192[2:0], u_ca_out_191[5:3]};
assign col_out_193 = {u_ca_out_193[2:0], u_ca_out_192[5:3]};
assign col_out_194 = {u_ca_out_194[2:0], u_ca_out_193[5:3]};
assign col_out_195 = {u_ca_out_195[2:0], u_ca_out_194[5:3]};
assign col_out_196 = {u_ca_out_196[2:0], u_ca_out_195[5:3]};
assign col_out_197 = {u_ca_out_197[2:0], u_ca_out_196[5:3]};
assign col_out_198 = {u_ca_out_198[2:0], u_ca_out_197[5:3]};
assign col_out_199 = {u_ca_out_199[2:0], u_ca_out_198[5:3]};
assign col_out_200 = {u_ca_out_200[2:0], u_ca_out_199[5:3]};
assign col_out_201 = {u_ca_out_201[2:0], u_ca_out_200[5:3]};
assign col_out_202 = {u_ca_out_202[2:0], u_ca_out_201[5:3]};
assign col_out_203 = {u_ca_out_203[2:0], u_ca_out_202[5:3]};
assign col_out_204 = {u_ca_out_204[2:0], u_ca_out_203[5:3]};
assign col_out_205 = {u_ca_out_205[2:0], u_ca_out_204[5:3]};
assign col_out_206 = {u_ca_out_206[2:0], u_ca_out_205[5:3]};
assign col_out_207 = {u_ca_out_207[2:0], u_ca_out_206[5:3]};
assign col_out_208 = {u_ca_out_208[2:0], u_ca_out_207[5:3]};
assign col_out_209 = {u_ca_out_209[2:0], u_ca_out_208[5:3]};
assign col_out_210 = {u_ca_out_210[2:0], u_ca_out_209[5:3]};
assign col_out_211 = {u_ca_out_211[2:0], u_ca_out_210[5:3]};
assign col_out_212 = {u_ca_out_212[2:0], u_ca_out_211[5:3]};
assign col_out_213 = {u_ca_out_213[2:0], u_ca_out_212[5:3]};
assign col_out_214 = {u_ca_out_214[2:0], u_ca_out_213[5:3]};
assign col_out_215 = {u_ca_out_215[2:0], u_ca_out_214[5:3]};
assign col_out_216 = {u_ca_out_216[2:0], u_ca_out_215[5:3]};
assign col_out_217 = {u_ca_out_217[2:0], u_ca_out_216[5:3]};
assign col_out_218 = {u_ca_out_218[2:0], u_ca_out_217[5:3]};
assign col_out_219 = {u_ca_out_219[2:0], u_ca_out_218[5:3]};
assign col_out_220 = {u_ca_out_220[2:0], u_ca_out_219[5:3]};
assign col_out_221 = {u_ca_out_221[2:0], u_ca_out_220[5:3]};
assign col_out_222 = {u_ca_out_222[2:0], u_ca_out_221[5:3]};
assign col_out_223 = {u_ca_out_223[2:0], u_ca_out_222[5:3]};
assign col_out_224 = {u_ca_out_224[2:0], u_ca_out_223[5:3]};
assign col_out_225 = {u_ca_out_225[2:0], u_ca_out_224[5:3]};
assign col_out_226 = {u_ca_out_226[2:0], u_ca_out_225[5:3]};
assign col_out_227 = {u_ca_out_227[2:0], u_ca_out_226[5:3]};
assign col_out_228 = {u_ca_out_228[2:0], u_ca_out_227[5:3]};
assign col_out_229 = {u_ca_out_229[2:0], u_ca_out_228[5:3]};
assign col_out_230 = {u_ca_out_230[2:0], u_ca_out_229[5:3]};
assign col_out_231 = {u_ca_out_231[2:0], u_ca_out_230[5:3]};
assign col_out_232 = {u_ca_out_232[2:0], u_ca_out_231[5:3]};
assign col_out_233 = {u_ca_out_233[2:0], u_ca_out_232[5:3]};
assign col_out_234 = {u_ca_out_234[2:0], u_ca_out_233[5:3]};
assign col_out_235 = {u_ca_out_235[2:0], u_ca_out_234[5:3]};
assign col_out_236 = {u_ca_out_236[2:0], u_ca_out_235[5:3]};
assign col_out_237 = {u_ca_out_237[2:0], u_ca_out_236[5:3]};
assign col_out_238 = {u_ca_out_238[2:0], u_ca_out_237[5:3]};
assign col_out_239 = {u_ca_out_239[2:0], u_ca_out_238[5:3]};
assign col_out_240 = {u_ca_out_240[2:0], u_ca_out_239[5:3]};
assign col_out_241 = {u_ca_out_241[2:0], u_ca_out_240[5:3]};
assign col_out_242 = {u_ca_out_242[2:0], u_ca_out_241[5:3]};
assign col_out_243 = {u_ca_out_243[2:0], u_ca_out_242[5:3]};
assign col_out_244 = {u_ca_out_244[2:0], u_ca_out_243[5:3]};
assign col_out_245 = {u_ca_out_245[2:0], u_ca_out_244[5:3]};
assign col_out_246 = {u_ca_out_246[2:0], u_ca_out_245[5:3]};
assign col_out_247 = {u_ca_out_247[2:0], u_ca_out_246[5:3]};
assign col_out_248 = {u_ca_out_248[2:0], u_ca_out_247[5:3]};
assign col_out_249 = {u_ca_out_249[2:0], u_ca_out_248[5:3]};
assign col_out_250 = {u_ca_out_250[2:0], u_ca_out_249[5:3]};
assign col_out_251 = {u_ca_out_251[2:0], u_ca_out_250[5:3]};
assign col_out_252 = {u_ca_out_252[2:0], u_ca_out_251[5:3]};
assign col_out_253 = {u_ca_out_253[2:0], u_ca_out_252[5:3]};
assign col_out_254 = {u_ca_out_254[2:0], u_ca_out_253[5:3]};
assign col_out_255 = {u_ca_out_255[2:0], u_ca_out_254[5:3]};
assign col_out_256 = {u_ca_out_256[2:0], u_ca_out_255[5:3]};
assign col_out_257 = {u_ca_out_257[2:0], u_ca_out_256[5:3]};
assign col_out_258 = {u_ca_out_258[2:0], u_ca_out_257[5:3]};
assign col_out_259 = {u_ca_out_259[2:0], u_ca_out_258[5:3]};
assign col_out_260 = {u_ca_out_260[2:0], u_ca_out_259[5:3]};
assign col_out_261 = {u_ca_out_261[2:0], u_ca_out_260[5:3]};
assign col_out_262 = {u_ca_out_262[2:0], u_ca_out_261[5:3]};
assign col_out_263 = {u_ca_out_263[2:0], u_ca_out_262[5:3]};
assign col_out_264 = {u_ca_out_264[2:0], u_ca_out_263[5:3]};
assign col_out_265 = {u_ca_out_265[2:0], u_ca_out_264[5:3]};
assign col_out_266 = {u_ca_out_266[2:0], u_ca_out_265[5:3]};
assign col_out_267 = {u_ca_out_267[2:0], u_ca_out_266[5:3]};
assign col_out_268 = {u_ca_out_268[2:0], u_ca_out_267[5:3]};
assign col_out_269 = {u_ca_out_269[2:0], u_ca_out_268[5:3]};
assign col_out_270 = {u_ca_out_270[2:0], u_ca_out_269[5:3]};
assign col_out_271 = {u_ca_out_271[2:0], u_ca_out_270[5:3]};
assign col_out_272 = {u_ca_out_272[2:0], u_ca_out_271[5:3]};
assign col_out_273 = {u_ca_out_273[2:0], u_ca_out_272[5:3]};
assign col_out_274 = {u_ca_out_274[2:0], u_ca_out_273[5:3]};
assign col_out_275 = {u_ca_out_275[2:0], u_ca_out_274[5:3]};
assign col_out_276 = {u_ca_out_276[2:0], u_ca_out_275[5:3]};
assign col_out_277 = {u_ca_out_277[2:0], u_ca_out_276[5:3]};
assign col_out_278 = {u_ca_out_278[2:0], u_ca_out_277[5:3]};
assign col_out_279 = {u_ca_out_279[2:0], u_ca_out_278[5:3]};
assign col_out_280 = {u_ca_out_280[2:0], u_ca_out_279[5:3]};
assign col_out_281 = {u_ca_out_281[2:0], u_ca_out_280[5:3]};
assign col_out_282 = {u_ca_out_282[2:0], u_ca_out_281[5:3]};
assign col_out_283 = {u_ca_out_283[2:0], u_ca_out_282[5:3]};
assign col_out_284 = {u_ca_out_284[2:0], u_ca_out_283[5:3]};
assign col_out_285 = {u_ca_out_285[2:0], u_ca_out_284[5:3]};
assign col_out_286 = {u_ca_out_286[2:0], u_ca_out_285[5:3]};
assign col_out_287 = {u_ca_out_287[2:0], u_ca_out_286[5:3]};
assign col_out_288 = {u_ca_out_288[2:0], u_ca_out_287[5:3]};
assign col_out_289 = {u_ca_out_289[2:0], u_ca_out_288[5:3]};
assign col_out_290 = {u_ca_out_290[2:0], u_ca_out_289[5:3]};
assign col_out_291 = {u_ca_out_291[2:0], u_ca_out_290[5:3]};
assign col_out_292 = {u_ca_out_292[2:0], u_ca_out_291[5:3]};
assign col_out_293 = {u_ca_out_293[2:0], u_ca_out_292[5:3]};
assign col_out_294 = {u_ca_out_294[2:0], u_ca_out_293[5:3]};
assign col_out_295 = {u_ca_out_295[2:0], u_ca_out_294[5:3]};
assign col_out_296 = {u_ca_out_296[2:0], u_ca_out_295[5:3]};
assign col_out_297 = {u_ca_out_297[2:0], u_ca_out_296[5:3]};
assign col_out_298 = {u_ca_out_298[2:0], u_ca_out_297[5:3]};
assign col_out_299 = {u_ca_out_299[2:0], u_ca_out_298[5:3]};
assign col_out_300 = {u_ca_out_300[2:0], u_ca_out_299[5:3]};
assign col_out_301 = {u_ca_out_301[2:0], u_ca_out_300[5:3]};
assign col_out_302 = {u_ca_out_302[2:0], u_ca_out_301[5:3]};
assign col_out_303 = {u_ca_out_303[2:0], u_ca_out_302[5:3]};
assign col_out_304 = {u_ca_out_304[2:0], u_ca_out_303[5:3]};
assign col_out_305 = {u_ca_out_305[2:0], u_ca_out_304[5:3]};
assign col_out_306 = {u_ca_out_306[2:0], u_ca_out_305[5:3]};
assign col_out_307 = {u_ca_out_307[2:0], u_ca_out_306[5:3]};
assign col_out_308 = {u_ca_out_308[2:0], u_ca_out_307[5:3]};
assign col_out_309 = {u_ca_out_309[2:0], u_ca_out_308[5:3]};
assign col_out_310 = {u_ca_out_310[2:0], u_ca_out_309[5:3]};
assign col_out_311 = {u_ca_out_311[2:0], u_ca_out_310[5:3]};
assign col_out_312 = {u_ca_out_312[2:0], u_ca_out_311[5:3]};
assign col_out_313 = {u_ca_out_313[2:0], u_ca_out_312[5:3]};
assign col_out_314 = {u_ca_out_314[2:0], u_ca_out_313[5:3]};
assign col_out_315 = {u_ca_out_315[2:0], u_ca_out_314[5:3]};
assign col_out_316 = {u_ca_out_316[2:0], u_ca_out_315[5:3]};
assign col_out_317 = {u_ca_out_317[2:0], u_ca_out_316[5:3]};
assign col_out_318 = {u_ca_out_318[2:0], u_ca_out_317[5:3]};
assign col_out_319 = {u_ca_out_319[2:0], u_ca_out_318[5:3]};
assign col_out_320 = {u_ca_out_320[2:0], u_ca_out_319[5:3]};
assign col_out_321 = {u_ca_out_321[2:0], u_ca_out_320[5:3]};
assign col_out_322 = {u_ca_out_322[2:0], u_ca_out_321[5:3]};
assign col_out_323 = {u_ca_out_323[2:0], u_ca_out_322[5:3]};
assign col_out_324 = {u_ca_out_324[2:0], u_ca_out_323[5:3]};
assign col_out_325 = {u_ca_out_325[2:0], u_ca_out_324[5:3]};
assign col_out_326 = {u_ca_out_326[2:0], u_ca_out_325[5:3]};
assign col_out_327 = {u_ca_out_327[2:0], u_ca_out_326[5:3]};
assign col_out_328 = {u_ca_out_328[2:0], u_ca_out_327[5:3]};
assign col_out_329 = {u_ca_out_329[2:0], u_ca_out_328[5:3]};
assign col_out_330 = {u_ca_out_330[2:0], u_ca_out_329[5:3]};
assign col_out_331 = {u_ca_out_331[2:0], u_ca_out_330[5:3]};
assign col_out_332 = {u_ca_out_332[2:0], u_ca_out_331[5:3]};
assign col_out_333 = {u_ca_out_333[2:0], u_ca_out_332[5:3]};
assign col_out_334 = {u_ca_out_334[2:0], u_ca_out_333[5:3]};
assign col_out_335 = {u_ca_out_335[2:0], u_ca_out_334[5:3]};
assign col_out_336 = {u_ca_out_336[2:0], u_ca_out_335[5:3]};
assign col_out_337 = {u_ca_out_337[2:0], u_ca_out_336[5:3]};
assign col_out_338 = {u_ca_out_338[2:0], u_ca_out_337[5:3]};
assign col_out_339 = {u_ca_out_339[2:0], u_ca_out_338[5:3]};
assign col_out_340 = {u_ca_out_340[2:0], u_ca_out_339[5:3]};
assign col_out_341 = {u_ca_out_341[2:0], u_ca_out_340[5:3]};
assign col_out_342 = {u_ca_out_342[2:0], u_ca_out_341[5:3]};
assign col_out_343 = {u_ca_out_343[2:0], u_ca_out_342[5:3]};
assign col_out_344 = {u_ca_out_344[2:0], u_ca_out_343[5:3]};
assign col_out_345 = {u_ca_out_345[2:0], u_ca_out_344[5:3]};
assign col_out_346 = {u_ca_out_346[2:0], u_ca_out_345[5:3]};
assign col_out_347 = {u_ca_out_347[2:0], u_ca_out_346[5:3]};
assign col_out_348 = {u_ca_out_348[2:0], u_ca_out_347[5:3]};
assign col_out_349 = {u_ca_out_349[2:0], u_ca_out_348[5:3]};
assign col_out_350 = {u_ca_out_350[2:0], u_ca_out_349[5:3]};
assign col_out_351 = {u_ca_out_351[2:0], u_ca_out_350[5:3]};
assign col_out_352 = {u_ca_out_352[2:0], u_ca_out_351[5:3]};
assign col_out_353 = {u_ca_out_353[2:0], u_ca_out_352[5:3]};
assign col_out_354 = {u_ca_out_354[2:0], u_ca_out_353[5:3]};
assign col_out_355 = {u_ca_out_355[2:0], u_ca_out_354[5:3]};
assign col_out_356 = {u_ca_out_356[2:0], u_ca_out_355[5:3]};
assign col_out_357 = {u_ca_out_357[2:0], u_ca_out_356[5:3]};
assign col_out_358 = {u_ca_out_358[2:0], u_ca_out_357[5:3]};
assign col_out_359 = {u_ca_out_359[2:0], u_ca_out_358[5:3]};
assign col_out_360 = {u_ca_out_360[2:0], u_ca_out_359[5:3]};
assign col_out_361 = {u_ca_out_361[2:0], u_ca_out_360[5:3]};
assign col_out_362 = {u_ca_out_362[2:0], u_ca_out_361[5:3]};
assign col_out_363 = {u_ca_out_363[2:0], u_ca_out_362[5:3]};
assign col_out_364 = {u_ca_out_364[2:0], u_ca_out_363[5:3]};
assign col_out_365 = {u_ca_out_365[2:0], u_ca_out_364[5:3]};
assign col_out_366 = {u_ca_out_366[2:0], u_ca_out_365[5:3]};
assign col_out_367 = {u_ca_out_367[2:0], u_ca_out_366[5:3]};
assign col_out_368 = {u_ca_out_368[2:0], u_ca_out_367[5:3]};
assign col_out_369 = {u_ca_out_369[2:0], u_ca_out_368[5:3]};
assign col_out_370 = {u_ca_out_370[2:0], u_ca_out_369[5:3]};
assign col_out_371 = {u_ca_out_371[2:0], u_ca_out_370[5:3]};
assign col_out_372 = {u_ca_out_372[2:0], u_ca_out_371[5:3]};
assign col_out_373 = {u_ca_out_373[2:0], u_ca_out_372[5:3]};
assign col_out_374 = {u_ca_out_374[2:0], u_ca_out_373[5:3]};
assign col_out_375 = {u_ca_out_375[2:0], u_ca_out_374[5:3]};
assign col_out_376 = {u_ca_out_376[2:0], u_ca_out_375[5:3]};
assign col_out_377 = {u_ca_out_377[2:0], u_ca_out_376[5:3]};
assign col_out_378 = {u_ca_out_378[2:0], u_ca_out_377[5:3]};
assign col_out_379 = {u_ca_out_379[2:0], u_ca_out_378[5:3]};
assign col_out_380 = {u_ca_out_380[2:0], u_ca_out_379[5:3]};
assign col_out_381 = {u_ca_out_381[2:0], u_ca_out_380[5:3]};
assign col_out_382 = {u_ca_out_382[2:0], u_ca_out_381[5:3]};
assign col_out_383 = {u_ca_out_383[2:0], u_ca_out_382[5:3]};
assign col_out_384 = {u_ca_out_384[2:0], u_ca_out_383[5:3]};
assign col_out_385 = {u_ca_out_385[2:0], u_ca_out_384[5:3]};
assign col_out_386 = {u_ca_out_386[2:0], u_ca_out_385[5:3]};
assign col_out_387 = {u_ca_out_387[2:0], u_ca_out_386[5:3]};
assign col_out_388 = {u_ca_out_388[2:0], u_ca_out_387[5:3]};
assign col_out_389 = {u_ca_out_389[2:0], u_ca_out_388[5:3]};
assign col_out_390 = {u_ca_out_390[2:0], u_ca_out_389[5:3]};
assign col_out_391 = {u_ca_out_391[2:0], u_ca_out_390[5:3]};
assign col_out_392 = {u_ca_out_392[2:0], u_ca_out_391[5:3]};
assign col_out_393 = {u_ca_out_393[2:0], u_ca_out_392[5:3]};
assign col_out_394 = {u_ca_out_394[2:0], u_ca_out_393[5:3]};
assign col_out_395 = {u_ca_out_395[2:0], u_ca_out_394[5:3]};
assign col_out_396 = {u_ca_out_396[2:0], u_ca_out_395[5:3]};
assign col_out_397 = {u_ca_out_397[2:0], u_ca_out_396[5:3]};
assign col_out_398 = {u_ca_out_398[2:0], u_ca_out_397[5:3]};
assign col_out_399 = {u_ca_out_399[2:0], u_ca_out_398[5:3]};
assign col_out_400 = {u_ca_out_400[2:0], u_ca_out_399[5:3]};
assign col_out_401 = {u_ca_out_401[2:0], u_ca_out_400[5:3]};
assign col_out_402 = {u_ca_out_402[2:0], u_ca_out_401[5:3]};
assign col_out_403 = {u_ca_out_403[2:0], u_ca_out_402[5:3]};
assign col_out_404 = {u_ca_out_404[2:0], u_ca_out_403[5:3]};
assign col_out_405 = {u_ca_out_405[2:0], u_ca_out_404[5:3]};
assign col_out_406 = {u_ca_out_406[2:0], u_ca_out_405[5:3]};
assign col_out_407 = {u_ca_out_407[2:0], u_ca_out_406[5:3]};
assign col_out_408 = {u_ca_out_408[2:0], u_ca_out_407[5:3]};
assign col_out_409 = {u_ca_out_409[2:0], u_ca_out_408[5:3]};
assign col_out_410 = {u_ca_out_410[2:0], u_ca_out_409[5:3]};
assign col_out_411 = {u_ca_out_411[2:0], u_ca_out_410[5:3]};
assign col_out_412 = {u_ca_out_412[2:0], u_ca_out_411[5:3]};
assign col_out_413 = {u_ca_out_413[2:0], u_ca_out_412[5:3]};
assign col_out_414 = {u_ca_out_414[2:0], u_ca_out_413[5:3]};
assign col_out_415 = {u_ca_out_415[2:0], u_ca_out_414[5:3]};
assign col_out_416 = {u_ca_out_416[2:0], u_ca_out_415[5:3]};
assign col_out_417 = {u_ca_out_417[2:0], u_ca_out_416[5:3]};
assign col_out_418 = {u_ca_out_418[2:0], u_ca_out_417[5:3]};
assign col_out_419 = {u_ca_out_419[2:0], u_ca_out_418[5:3]};
assign col_out_420 = {u_ca_out_420[2:0], u_ca_out_419[5:3]};
assign col_out_421 = {u_ca_out_421[2:0], u_ca_out_420[5:3]};
assign col_out_422 = {u_ca_out_422[2:0], u_ca_out_421[5:3]};
assign col_out_423 = {u_ca_out_423[2:0], u_ca_out_422[5:3]};
assign col_out_424 = {u_ca_out_424[2:0], u_ca_out_423[5:3]};
assign col_out_425 = {u_ca_out_425[2:0], u_ca_out_424[5:3]};
assign col_out_426 = {u_ca_out_426[2:0], u_ca_out_425[5:3]};
assign col_out_427 = {u_ca_out_427[2:0], u_ca_out_426[5:3]};
assign col_out_428 = {u_ca_out_428[2:0], u_ca_out_427[5:3]};
assign col_out_429 = {u_ca_out_429[2:0], u_ca_out_428[5:3]};
assign col_out_430 = {u_ca_out_430[2:0], u_ca_out_429[5:3]};
assign col_out_431 = {u_ca_out_431[2:0], u_ca_out_430[5:3]};
assign col_out_432 = {u_ca_out_432[2:0], u_ca_out_431[5:3]};
assign col_out_433 = {u_ca_out_433[2:0], u_ca_out_432[5:3]};
assign col_out_434 = {u_ca_out_434[2:0], u_ca_out_433[5:3]};
assign col_out_435 = {u_ca_out_435[2:0], u_ca_out_434[5:3]};
assign col_out_436 = {u_ca_out_436[2:0], u_ca_out_435[5:3]};
assign col_out_437 = {u_ca_out_437[2:0], u_ca_out_436[5:3]};
assign col_out_438 = {u_ca_out_438[2:0], u_ca_out_437[5:3]};
assign col_out_439 = {u_ca_out_439[2:0], u_ca_out_438[5:3]};
assign col_out_440 = {u_ca_out_440[2:0], u_ca_out_439[5:3]};
assign col_out_441 = {u_ca_out_441[2:0], u_ca_out_440[5:3]};
assign col_out_442 = {u_ca_out_442[2:0], u_ca_out_441[5:3]};
assign col_out_443 = {u_ca_out_443[2:0], u_ca_out_442[5:3]};
assign col_out_444 = {u_ca_out_444[2:0], u_ca_out_443[5:3]};
assign col_out_445 = {u_ca_out_445[2:0], u_ca_out_444[5:3]};
assign col_out_446 = {u_ca_out_446[2:0], u_ca_out_445[5:3]};
assign col_out_447 = {u_ca_out_447[2:0], u_ca_out_446[5:3]};
assign col_out_448 = {u_ca_out_448[2:0], u_ca_out_447[5:3]};
assign col_out_449 = {u_ca_out_449[2:0], u_ca_out_448[5:3]};
assign col_out_450 = {u_ca_out_450[2:0], u_ca_out_449[5:3]};
assign col_out_451 = {u_ca_out_451[2:0], u_ca_out_450[5:3]};
assign col_out_452 = {u_ca_out_452[2:0], u_ca_out_451[5:3]};
assign col_out_453 = {u_ca_out_453[2:0], u_ca_out_452[5:3]};
assign col_out_454 = {u_ca_out_454[2:0], u_ca_out_453[5:3]};
assign col_out_455 = {u_ca_out_455[2:0], u_ca_out_454[5:3]};
assign col_out_456 = {u_ca_out_456[2:0], u_ca_out_455[5:3]};
assign col_out_457 = {u_ca_out_457[2:0], u_ca_out_456[5:3]};
assign col_out_458 = {u_ca_out_458[2:0], u_ca_out_457[5:3]};
assign col_out_459 = {u_ca_out_459[2:0], u_ca_out_458[5:3]};
assign col_out_460 = {u_ca_out_460[2:0], u_ca_out_459[5:3]};
assign col_out_461 = {u_ca_out_461[2:0], u_ca_out_460[5:3]};
assign col_out_462 = {u_ca_out_462[2:0], u_ca_out_461[5:3]};
assign col_out_463 = {u_ca_out_463[2:0], u_ca_out_462[5:3]};
assign col_out_464 = {u_ca_out_464[2:0], u_ca_out_463[5:3]};
assign col_out_465 = {u_ca_out_465[2:0], u_ca_out_464[5:3]};
assign col_out_466 = {u_ca_out_466[2:0], u_ca_out_465[5:3]};
assign col_out_467 = {u_ca_out_467[2:0], u_ca_out_466[5:3]};
assign col_out_468 = {u_ca_out_468[2:0], u_ca_out_467[5:3]};
assign col_out_469 = {u_ca_out_469[2:0], u_ca_out_468[5:3]};
assign col_out_470 = {u_ca_out_470[2:0], u_ca_out_469[5:3]};
assign col_out_471 = {u_ca_out_471[2:0], u_ca_out_470[5:3]};
assign col_out_472 = {u_ca_out_472[2:0], u_ca_out_471[5:3]};
assign col_out_473 = {u_ca_out_473[2:0], u_ca_out_472[5:3]};
assign col_out_474 = {u_ca_out_474[2:0], u_ca_out_473[5:3]};
assign col_out_475 = {u_ca_out_475[2:0], u_ca_out_474[5:3]};
assign col_out_476 = {u_ca_out_476[2:0], u_ca_out_475[5:3]};
assign col_out_477 = {u_ca_out_477[2:0], u_ca_out_476[5:3]};
assign col_out_478 = {u_ca_out_478[2:0], u_ca_out_477[5:3]};
assign col_out_479 = {u_ca_out_479[2:0], u_ca_out_478[5:3]};
assign col_out_480 = {u_ca_out_480[2:0], u_ca_out_479[5:3]};
assign col_out_481 = {u_ca_out_481[2:0], u_ca_out_480[5:3]};
assign col_out_482 = {u_ca_out_482[2:0], u_ca_out_481[5:3]};
assign col_out_483 = {u_ca_out_483[2:0], u_ca_out_482[5:3]};
assign col_out_484 = {u_ca_out_484[2:0], u_ca_out_483[5:3]};
assign col_out_485 = {u_ca_out_485[2:0], u_ca_out_484[5:3]};
assign col_out_486 = {u_ca_out_486[2:0], u_ca_out_485[5:3]};
assign col_out_487 = {u_ca_out_487[2:0], u_ca_out_486[5:3]};
assign col_out_488 = {u_ca_out_488[2:0], u_ca_out_487[5:3]};
assign col_out_489 = {u_ca_out_489[2:0], u_ca_out_488[5:3]};
assign col_out_490 = {u_ca_out_490[2:0], u_ca_out_489[5:3]};
assign col_out_491 = {u_ca_out_491[2:0], u_ca_out_490[5:3]};
assign col_out_492 = {u_ca_out_492[2:0], u_ca_out_491[5:3]};
assign col_out_493 = {u_ca_out_493[2:0], u_ca_out_492[5:3]};
assign col_out_494 = {u_ca_out_494[2:0], u_ca_out_493[5:3]};
assign col_out_495 = {u_ca_out_495[2:0], u_ca_out_494[5:3]};
assign col_out_496 = {u_ca_out_496[2:0], u_ca_out_495[5:3]};
assign col_out_497 = {u_ca_out_497[2:0], u_ca_out_496[5:3]};
assign col_out_498 = {u_ca_out_498[2:0], u_ca_out_497[5:3]};
assign col_out_499 = {u_ca_out_499[2:0], u_ca_out_498[5:3]};
assign col_out_500 = {u_ca_out_500[2:0], u_ca_out_499[5:3]};
assign col_out_501 = {u_ca_out_501[2:0], u_ca_out_500[5:3]};
assign col_out_502 = {u_ca_out_502[2:0], u_ca_out_501[5:3]};
assign col_out_503 = {u_ca_out_503[2:0], u_ca_out_502[5:3]};
assign col_out_504 = {u_ca_out_504[2:0], u_ca_out_503[5:3]};
assign col_out_505 = {u_ca_out_505[2:0], u_ca_out_504[5:3]};
assign col_out_506 = {u_ca_out_506[2:0], u_ca_out_505[5:3]};
assign col_out_507 = {u_ca_out_507[2:0], u_ca_out_506[5:3]};
assign col_out_508 = {u_ca_out_508[2:0], u_ca_out_507[5:3]};
assign col_out_509 = {u_ca_out_509[2:0], u_ca_out_508[5:3]};
assign col_out_510 = {u_ca_out_510[2:0], u_ca_out_509[5:3]};
assign col_out_511 = {u_ca_out_511[2:0], u_ca_out_510[5:3]};
assign col_out_512 = {u_ca_out_512[2:0], u_ca_out_511[5:3]};
assign col_out_513 = {u_ca_out_513[2:0], u_ca_out_512[5:3]};
assign col_out_514 = {u_ca_out_514[2:0], u_ca_out_513[5:3]};
assign col_out_515 = {u_ca_out_515[2:0], u_ca_out_514[5:3]};
assign col_out_516 = {u_ca_out_516[2:0], u_ca_out_515[5:3]};
assign col_out_517 = {u_ca_out_517[2:0], u_ca_out_516[5:3]};
assign col_out_518 = {u_ca_out_518[2:0], u_ca_out_517[5:3]};
assign col_out_519 = {u_ca_out_519[2:0], u_ca_out_518[5:3]};
assign col_out_520 = {u_ca_out_520[2:0], u_ca_out_519[5:3]};
assign col_out_521 = {u_ca_out_521[2:0], u_ca_out_520[5:3]};
assign col_out_522 = {u_ca_out_522[2:0], u_ca_out_521[5:3]};
assign col_out_523 = {u_ca_out_523[2:0], u_ca_out_522[5:3]};
assign col_out_524 = {u_ca_out_524[2:0], u_ca_out_523[5:3]};
assign col_out_525 = {u_ca_out_525[2:0], u_ca_out_524[5:3]};
assign col_out_526 = {u_ca_out_526[2:0], u_ca_out_525[5:3]};
assign col_out_527 = {u_ca_out_527[2:0], u_ca_out_526[5:3]};
assign col_out_528 = {u_ca_out_528[2:0], u_ca_out_527[5:3]};
assign col_out_529 = {u_ca_out_529[2:0], u_ca_out_528[5:3]};
assign col_out_530 = {u_ca_out_530[2:0], u_ca_out_529[5:3]};
assign col_out_531 = {u_ca_out_531[2:0], u_ca_out_530[5:3]};
assign col_out_532 = {u_ca_out_532[2:0], u_ca_out_531[5:3]};
assign col_out_533 = {u_ca_out_533[2:0], u_ca_out_532[5:3]};
assign col_out_534 = {u_ca_out_534[2:0], u_ca_out_533[5:3]};
assign col_out_535 = {u_ca_out_535[2:0], u_ca_out_534[5:3]};
assign col_out_536 = {u_ca_out_536[2:0], u_ca_out_535[5:3]};
assign col_out_537 = {u_ca_out_537[2:0], u_ca_out_536[5:3]};
assign col_out_538 = {u_ca_out_538[2:0], u_ca_out_537[5:3]};
assign col_out_539 = {u_ca_out_539[2:0], u_ca_out_538[5:3]};
assign col_out_540 = {u_ca_out_540[2:0], u_ca_out_539[5:3]};
assign col_out_541 = {u_ca_out_541[2:0], u_ca_out_540[5:3]};
assign col_out_542 = {u_ca_out_542[2:0], u_ca_out_541[5:3]};
assign col_out_543 = {u_ca_out_543[2:0], u_ca_out_542[5:3]};
assign col_out_544 = {u_ca_out_544[2:0], u_ca_out_543[5:3]};
assign col_out_545 = {u_ca_out_545[2:0], u_ca_out_544[5:3]};
assign col_out_546 = {u_ca_out_546[2:0], u_ca_out_545[5:3]};
assign col_out_547 = {u_ca_out_547[2:0], u_ca_out_546[5:3]};
assign col_out_548 = {u_ca_out_548[2:0], u_ca_out_547[5:3]};
assign col_out_549 = {u_ca_out_549[2:0], u_ca_out_548[5:3]};
assign col_out_550 = {u_ca_out_550[2:0], u_ca_out_549[5:3]};
assign col_out_551 = {u_ca_out_551[2:0], u_ca_out_550[5:3]};
assign col_out_552 = {u_ca_out_552[2:0], u_ca_out_551[5:3]};
assign col_out_553 = {u_ca_out_553[2:0], u_ca_out_552[5:3]};
assign col_out_554 = {u_ca_out_554[2:0], u_ca_out_553[5:3]};
assign col_out_555 = {u_ca_out_555[2:0], u_ca_out_554[5:3]};
assign col_out_556 = {u_ca_out_556[2:0], u_ca_out_555[5:3]};
assign col_out_557 = {u_ca_out_557[2:0], u_ca_out_556[5:3]};
assign col_out_558 = {u_ca_out_558[2:0], u_ca_out_557[5:3]};
assign col_out_559 = {u_ca_out_559[2:0], u_ca_out_558[5:3]};
assign col_out_560 = {u_ca_out_560[2:0], u_ca_out_559[5:3]};
assign col_out_561 = {u_ca_out_561[2:0], u_ca_out_560[5:3]};
assign col_out_562 = {u_ca_out_562[2:0], u_ca_out_561[5:3]};
assign col_out_563 = {u_ca_out_563[2:0], u_ca_out_562[5:3]};
assign col_out_564 = {u_ca_out_564[2:0], u_ca_out_563[5:3]};
assign col_out_565 = {u_ca_out_565[2:0], u_ca_out_564[5:3]};
assign col_out_566 = {u_ca_out_566[2:0], u_ca_out_565[5:3]};
assign col_out_567 = {u_ca_out_567[2:0], u_ca_out_566[5:3]};
assign col_out_568 = {u_ca_out_568[2:0], u_ca_out_567[5:3]};
assign col_out_569 = {u_ca_out_569[2:0], u_ca_out_568[5:3]};
assign col_out_570 = {u_ca_out_570[2:0], u_ca_out_569[5:3]};
assign col_out_571 = {u_ca_out_571[2:0], u_ca_out_570[5:3]};
assign col_out_572 = {u_ca_out_572[2:0], u_ca_out_571[5:3]};
assign col_out_573 = {u_ca_out_573[2:0], u_ca_out_572[5:3]};
assign col_out_574 = {u_ca_out_574[2:0], u_ca_out_573[5:3]};
assign col_out_575 = {u_ca_out_575[2:0], u_ca_out_574[5:3]};
assign col_out_576 = {u_ca_out_576[2:0], u_ca_out_575[5:3]};
assign col_out_577 = {u_ca_out_577[2:0], u_ca_out_576[5:3]};
assign col_out_578 = {u_ca_out_578[2:0], u_ca_out_577[5:3]};
assign col_out_579 = {u_ca_out_579[2:0], u_ca_out_578[5:3]};
assign col_out_580 = {u_ca_out_580[2:0], u_ca_out_579[5:3]};
assign col_out_581 = {u_ca_out_581[2:0], u_ca_out_580[5:3]};
assign col_out_582 = {u_ca_out_582[2:0], u_ca_out_581[5:3]};
assign col_out_583 = {u_ca_out_583[2:0], u_ca_out_582[5:3]};
assign col_out_584 = {u_ca_out_584[2:0], u_ca_out_583[5:3]};
assign col_out_585 = {u_ca_out_585[2:0], u_ca_out_584[5:3]};
assign col_out_586 = {u_ca_out_586[2:0], u_ca_out_585[5:3]};
assign col_out_587 = {u_ca_out_587[2:0], u_ca_out_586[5:3]};
assign col_out_588 = {u_ca_out_588[2:0], u_ca_out_587[5:3]};
assign col_out_589 = {u_ca_out_589[2:0], u_ca_out_588[5:3]};
assign col_out_590 = {u_ca_out_590[2:0], u_ca_out_589[5:3]};
assign col_out_591 = {u_ca_out_591[2:0], u_ca_out_590[5:3]};
assign col_out_592 = {u_ca_out_592[2:0], u_ca_out_591[5:3]};
assign col_out_593 = {u_ca_out_593[2:0], u_ca_out_592[5:3]};
assign col_out_594 = {u_ca_out_594[2:0], u_ca_out_593[5:3]};
assign col_out_595 = {u_ca_out_595[2:0], u_ca_out_594[5:3]};
assign col_out_596 = {u_ca_out_596[2:0], u_ca_out_595[5:3]};
assign col_out_597 = {u_ca_out_597[2:0], u_ca_out_596[5:3]};
assign col_out_598 = {u_ca_out_598[2:0], u_ca_out_597[5:3]};
assign col_out_599 = {u_ca_out_599[2:0], u_ca_out_598[5:3]};
assign col_out_600 = {u_ca_out_600[2:0], u_ca_out_599[5:3]};
assign col_out_601 = {u_ca_out_601[2:0], u_ca_out_600[5:3]};
assign col_out_602 = {u_ca_out_602[2:0], u_ca_out_601[5:3]};
assign col_out_603 = {u_ca_out_603[2:0], u_ca_out_602[5:3]};
assign col_out_604 = {u_ca_out_604[2:0], u_ca_out_603[5:3]};
assign col_out_605 = {u_ca_out_605[2:0], u_ca_out_604[5:3]};
assign col_out_606 = {u_ca_out_606[2:0], u_ca_out_605[5:3]};
assign col_out_607 = {u_ca_out_607[2:0], u_ca_out_606[5:3]};
assign col_out_608 = {u_ca_out_608[2:0], u_ca_out_607[5:3]};
assign col_out_609 = {u_ca_out_609[2:0], u_ca_out_608[5:3]};
assign col_out_610 = {u_ca_out_610[2:0], u_ca_out_609[5:3]};
assign col_out_611 = {u_ca_out_611[2:0], u_ca_out_610[5:3]};
assign col_out_612 = {u_ca_out_612[2:0], u_ca_out_611[5:3]};
assign col_out_613 = {u_ca_out_613[2:0], u_ca_out_612[5:3]};
assign col_out_614 = {u_ca_out_614[2:0], u_ca_out_613[5:3]};
assign col_out_615 = {u_ca_out_615[2:0], u_ca_out_614[5:3]};
assign col_out_616 = {u_ca_out_616[2:0], u_ca_out_615[5:3]};
assign col_out_617 = {u_ca_out_617[2:0], u_ca_out_616[5:3]};
assign col_out_618 = {u_ca_out_618[2:0], u_ca_out_617[5:3]};
assign col_out_619 = {u_ca_out_619[2:0], u_ca_out_618[5:3]};
assign col_out_620 = {u_ca_out_620[2:0], u_ca_out_619[5:3]};
assign col_out_621 = {u_ca_out_621[2:0], u_ca_out_620[5:3]};
assign col_out_622 = {u_ca_out_622[2:0], u_ca_out_621[5:3]};
assign col_out_623 = {u_ca_out_623[2:0], u_ca_out_622[5:3]};
assign col_out_624 = {u_ca_out_624[2:0], u_ca_out_623[5:3]};
assign col_out_625 = {u_ca_out_625[2:0], u_ca_out_624[5:3]};
assign col_out_626 = {u_ca_out_626[2:0], u_ca_out_625[5:3]};
assign col_out_627 = {u_ca_out_627[2:0], u_ca_out_626[5:3]};
assign col_out_628 = {u_ca_out_628[2:0], u_ca_out_627[5:3]};
assign col_out_629 = {u_ca_out_629[2:0], u_ca_out_628[5:3]};
assign col_out_630 = {u_ca_out_630[2:0], u_ca_out_629[5:3]};
assign col_out_631 = {u_ca_out_631[2:0], u_ca_out_630[5:3]};
assign col_out_632 = {u_ca_out_632[2:0], u_ca_out_631[5:3]};
assign col_out_633 = {u_ca_out_633[2:0], u_ca_out_632[5:3]};
assign col_out_634 = {u_ca_out_634[2:0], u_ca_out_633[5:3]};
assign col_out_635 = {u_ca_out_635[2:0], u_ca_out_634[5:3]};
assign col_out_636 = {u_ca_out_636[2:0], u_ca_out_635[5:3]};
assign col_out_637 = {u_ca_out_637[2:0], u_ca_out_636[5:3]};
assign col_out_638 = {u_ca_out_638[2:0], u_ca_out_637[5:3]};
assign col_out_639 = {u_ca_out_639[2:0], u_ca_out_638[5:3]};
assign col_out_640 = {u_ca_out_640[2:0], u_ca_out_639[5:3]};
assign col_out_641 = {u_ca_out_641[2:0], u_ca_out_640[5:3]};
assign col_out_642 = {u_ca_out_642[2:0], u_ca_out_641[5:3]};
assign col_out_643 = {u_ca_out_643[2:0], u_ca_out_642[5:3]};
assign col_out_644 = {u_ca_out_644[2:0], u_ca_out_643[5:3]};
assign col_out_645 = {u_ca_out_645[2:0], u_ca_out_644[5:3]};
assign col_out_646 = {u_ca_out_646[2:0], u_ca_out_645[5:3]};
assign col_out_647 = {u_ca_out_647[2:0], u_ca_out_646[5:3]};
assign col_out_648 = {u_ca_out_648[2:0], u_ca_out_647[5:3]};
assign col_out_649 = {u_ca_out_649[2:0], u_ca_out_648[5:3]};
assign col_out_650 = {u_ca_out_650[2:0], u_ca_out_649[5:3]};
assign col_out_651 = {u_ca_out_651[2:0], u_ca_out_650[5:3]};
assign col_out_652 = {u_ca_out_652[2:0], u_ca_out_651[5:3]};
assign col_out_653 = {u_ca_out_653[2:0], u_ca_out_652[5:3]};
assign col_out_654 = {u_ca_out_654[2:0], u_ca_out_653[5:3]};
assign col_out_655 = {u_ca_out_655[2:0], u_ca_out_654[5:3]};
assign col_out_656 = {u_ca_out_656[2:0], u_ca_out_655[5:3]};
assign col_out_657 = {u_ca_out_657[2:0], u_ca_out_656[5:3]};
assign col_out_658 = {u_ca_out_658[2:0], u_ca_out_657[5:3]};
assign col_out_659 = {u_ca_out_659[2:0], u_ca_out_658[5:3]};
assign col_out_660 = {u_ca_out_660[2:0], u_ca_out_659[5:3]};
assign col_out_661 = {u_ca_out_661[2:0], u_ca_out_660[5:3]};
assign col_out_662 = {u_ca_out_662[2:0], u_ca_out_661[5:3]};
assign col_out_663 = {u_ca_out_663[2:0], u_ca_out_662[5:3]};
assign col_out_664 = {u_ca_out_664[2:0], u_ca_out_663[5:3]};
assign col_out_665 = {u_ca_out_665[2:0], u_ca_out_664[5:3]};
assign col_out_666 = {u_ca_out_666[2:0], u_ca_out_665[5:3]};
assign col_out_667 = {u_ca_out_667[2:0], u_ca_out_666[5:3]};
assign col_out_668 = {u_ca_out_668[2:0], u_ca_out_667[5:3]};
assign col_out_669 = {u_ca_out_669[2:0], u_ca_out_668[5:3]};
assign col_out_670 = {u_ca_out_670[2:0], u_ca_out_669[5:3]};
assign col_out_671 = {u_ca_out_671[2:0], u_ca_out_670[5:3]};
assign col_out_672 = {u_ca_out_672[2:0], u_ca_out_671[5:3]};
assign col_out_673 = {u_ca_out_673[2:0], u_ca_out_672[5:3]};
assign col_out_674 = {u_ca_out_674[2:0], u_ca_out_673[5:3]};
assign col_out_675 = {u_ca_out_675[2:0], u_ca_out_674[5:3]};
assign col_out_676 = {u_ca_out_676[2:0], u_ca_out_675[5:3]};
assign col_out_677 = {u_ca_out_677[2:0], u_ca_out_676[5:3]};
assign col_out_678 = {u_ca_out_678[2:0], u_ca_out_677[5:3]};
assign col_out_679 = {u_ca_out_679[2:0], u_ca_out_678[5:3]};
assign col_out_680 = {u_ca_out_680[2:0], u_ca_out_679[5:3]};
assign col_out_681 = {u_ca_out_681[2:0], u_ca_out_680[5:3]};
assign col_out_682 = {u_ca_out_682[2:0], u_ca_out_681[5:3]};
assign col_out_683 = {u_ca_out_683[2:0], u_ca_out_682[5:3]};
assign col_out_684 = {u_ca_out_684[2:0], u_ca_out_683[5:3]};
assign col_out_685 = {u_ca_out_685[2:0], u_ca_out_684[5:3]};
assign col_out_686 = {u_ca_out_686[2:0], u_ca_out_685[5:3]};
assign col_out_687 = {u_ca_out_687[2:0], u_ca_out_686[5:3]};
assign col_out_688 = {u_ca_out_688[2:0], u_ca_out_687[5:3]};
assign col_out_689 = {u_ca_out_689[2:0], u_ca_out_688[5:3]};
assign col_out_690 = {u_ca_out_690[2:0], u_ca_out_689[5:3]};
assign col_out_691 = {u_ca_out_691[2:0], u_ca_out_690[5:3]};
assign col_out_692 = {u_ca_out_692[2:0], u_ca_out_691[5:3]};
assign col_out_693 = {u_ca_out_693[2:0], u_ca_out_692[5:3]};
assign col_out_694 = {u_ca_out_694[2:0], u_ca_out_693[5:3]};
assign col_out_695 = {u_ca_out_695[2:0], u_ca_out_694[5:3]};
assign col_out_696 = {u_ca_out_696[2:0], u_ca_out_695[5:3]};
assign col_out_697 = {u_ca_out_697[2:0], u_ca_out_696[5:3]};
assign col_out_698 = {u_ca_out_698[2:0], u_ca_out_697[5:3]};
assign col_out_699 = {u_ca_out_699[2:0], u_ca_out_698[5:3]};
assign col_out_700 = {u_ca_out_700[2:0], u_ca_out_699[5:3]};
assign col_out_701 = {u_ca_out_701[2:0], u_ca_out_700[5:3]};
assign col_out_702 = {u_ca_out_702[2:0], u_ca_out_701[5:3]};
assign col_out_703 = {u_ca_out_703[2:0], u_ca_out_702[5:3]};
assign col_out_704 = {u_ca_out_704[2:0], u_ca_out_703[5:3]};
assign col_out_705 = {u_ca_out_705[2:0], u_ca_out_704[5:3]};
assign col_out_706 = {u_ca_out_706[2:0], u_ca_out_705[5:3]};
assign col_out_707 = {u_ca_out_707[2:0], u_ca_out_706[5:3]};
assign col_out_708 = {u_ca_out_708[2:0], u_ca_out_707[5:3]};
assign col_out_709 = {u_ca_out_709[2:0], u_ca_out_708[5:3]};
assign col_out_710 = {u_ca_out_710[2:0], u_ca_out_709[5:3]};
assign col_out_711 = {u_ca_out_711[2:0], u_ca_out_710[5:3]};
assign col_out_712 = {u_ca_out_712[2:0], u_ca_out_711[5:3]};
assign col_out_713 = {u_ca_out_713[2:0], u_ca_out_712[5:3]};
assign col_out_714 = {u_ca_out_714[2:0], u_ca_out_713[5:3]};
assign col_out_715 = {u_ca_out_715[2:0], u_ca_out_714[5:3]};
assign col_out_716 = {u_ca_out_716[2:0], u_ca_out_715[5:3]};
assign col_out_717 = {u_ca_out_717[2:0], u_ca_out_716[5:3]};
assign col_out_718 = {u_ca_out_718[2:0], u_ca_out_717[5:3]};
assign col_out_719 = {u_ca_out_719[2:0], u_ca_out_718[5:3]};
assign col_out_720 = {u_ca_out_720[2:0], u_ca_out_719[5:3]};
assign col_out_721 = {u_ca_out_721[2:0], u_ca_out_720[5:3]};
assign col_out_722 = {u_ca_out_722[2:0], u_ca_out_721[5:3]};
assign col_out_723 = {u_ca_out_723[2:0], u_ca_out_722[5:3]};
assign col_out_724 = {u_ca_out_724[2:0], u_ca_out_723[5:3]};
assign col_out_725 = {u_ca_out_725[2:0], u_ca_out_724[5:3]};
assign col_out_726 = {u_ca_out_726[2:0], u_ca_out_725[5:3]};
assign col_out_727 = {u_ca_out_727[2:0], u_ca_out_726[5:3]};
assign col_out_728 = {u_ca_out_728[2:0], u_ca_out_727[5:3]};
assign col_out_729 = {u_ca_out_729[2:0], u_ca_out_728[5:3]};
assign col_out_730 = {u_ca_out_730[2:0], u_ca_out_729[5:3]};
assign col_out_731 = {u_ca_out_731[2:0], u_ca_out_730[5:3]};
assign col_out_732 = {u_ca_out_732[2:0], u_ca_out_731[5:3]};
assign col_out_733 = {u_ca_out_733[2:0], u_ca_out_732[5:3]};
assign col_out_734 = {u_ca_out_734[2:0], u_ca_out_733[5:3]};
assign col_out_735 = {u_ca_out_735[2:0], u_ca_out_734[5:3]};
assign col_out_736 = {u_ca_out_736[2:0], u_ca_out_735[5:3]};
assign col_out_737 = {u_ca_out_737[2:0], u_ca_out_736[5:3]};
assign col_out_738 = {u_ca_out_738[2:0], u_ca_out_737[5:3]};
assign col_out_739 = {u_ca_out_739[2:0], u_ca_out_738[5:3]};
assign col_out_740 = {u_ca_out_740[2:0], u_ca_out_739[5:3]};
assign col_out_741 = {u_ca_out_741[2:0], u_ca_out_740[5:3]};
assign col_out_742 = {u_ca_out_742[2:0], u_ca_out_741[5:3]};
assign col_out_743 = {u_ca_out_743[2:0], u_ca_out_742[5:3]};
assign col_out_744 = {u_ca_out_744[2:0], u_ca_out_743[5:3]};
assign col_out_745 = {u_ca_out_745[2:0], u_ca_out_744[5:3]};
assign col_out_746 = {u_ca_out_746[2:0], u_ca_out_745[5:3]};
assign col_out_747 = {u_ca_out_747[2:0], u_ca_out_746[5:3]};
assign col_out_748 = {u_ca_out_748[2:0], u_ca_out_747[5:3]};
assign col_out_749 = {u_ca_out_749[2:0], u_ca_out_748[5:3]};
assign col_out_750 = {u_ca_out_750[2:0], u_ca_out_749[5:3]};
assign col_out_751 = {u_ca_out_751[2:0], u_ca_out_750[5:3]};
assign col_out_752 = {u_ca_out_752[2:0], u_ca_out_751[5:3]};
assign col_out_753 = {u_ca_out_753[2:0], u_ca_out_752[5:3]};
assign col_out_754 = {u_ca_out_754[2:0], u_ca_out_753[5:3]};
assign col_out_755 = {u_ca_out_755[2:0], u_ca_out_754[5:3]};
assign col_out_756 = {u_ca_out_756[2:0], u_ca_out_755[5:3]};
assign col_out_757 = {u_ca_out_757[2:0], u_ca_out_756[5:3]};
assign col_out_758 = {u_ca_out_758[2:0], u_ca_out_757[5:3]};
assign col_out_759 = {u_ca_out_759[2:0], u_ca_out_758[5:3]};
assign col_out_760 = {u_ca_out_760[2:0], u_ca_out_759[5:3]};
assign col_out_761 = {u_ca_out_761[2:0], u_ca_out_760[5:3]};
assign col_out_762 = {u_ca_out_762[2:0], u_ca_out_761[5:3]};
assign col_out_763 = {u_ca_out_763[2:0], u_ca_out_762[5:3]};
assign col_out_764 = {u_ca_out_764[2:0], u_ca_out_763[5:3]};
assign col_out_765 = {u_ca_out_765[2:0], u_ca_out_764[5:3]};
assign col_out_766 = {u_ca_out_766[2:0], u_ca_out_765[5:3]};
assign col_out_767 = {u_ca_out_767[2:0], u_ca_out_766[5:3]};
assign col_out_768 = {u_ca_out_768[2:0], u_ca_out_767[5:3]};
assign col_out_769 = {u_ca_out_769[2:0], u_ca_out_768[5:3]};
assign col_out_770 = {u_ca_out_770[2:0], u_ca_out_769[5:3]};
assign col_out_771 = {u_ca_out_771[2:0], u_ca_out_770[5:3]};
assign col_out_772 = {u_ca_out_772[2:0], u_ca_out_771[5:3]};
assign col_out_773 = {u_ca_out_773[2:0], u_ca_out_772[5:3]};
assign col_out_774 = {u_ca_out_774[2:0], u_ca_out_773[5:3]};
assign col_out_775 = {u_ca_out_775[2:0], u_ca_out_774[5:3]};
assign col_out_776 = {u_ca_out_776[2:0], u_ca_out_775[5:3]};
assign col_out_777 = {u_ca_out_777[2:0], u_ca_out_776[5:3]};
assign col_out_778 = {u_ca_out_778[2:0], u_ca_out_777[5:3]};
assign col_out_779 = {u_ca_out_779[2:0], u_ca_out_778[5:3]};
assign col_out_780 = {u_ca_out_780[2:0], u_ca_out_779[5:3]};
assign col_out_781 = {u_ca_out_781[2:0], u_ca_out_780[5:3]};
assign col_out_782 = {u_ca_out_782[2:0], u_ca_out_781[5:3]};
assign col_out_783 = {u_ca_out_783[2:0], u_ca_out_782[5:3]};
assign col_out_784 = {u_ca_out_784[2:0], u_ca_out_783[5:3]};
assign col_out_785 = {u_ca_out_785[2:0], u_ca_out_784[5:3]};
assign col_out_786 = {u_ca_out_786[2:0], u_ca_out_785[5:3]};
assign col_out_787 = {u_ca_out_787[2:0], u_ca_out_786[5:3]};
assign col_out_788 = {u_ca_out_788[2:0], u_ca_out_787[5:3]};
assign col_out_789 = {u_ca_out_789[2:0], u_ca_out_788[5:3]};
assign col_out_790 = {u_ca_out_790[2:0], u_ca_out_789[5:3]};
assign col_out_791 = {u_ca_out_791[2:0], u_ca_out_790[5:3]};
assign col_out_792 = {u_ca_out_792[2:0], u_ca_out_791[5:3]};
assign col_out_793 = {u_ca_out_793[2:0], u_ca_out_792[5:3]};
assign col_out_794 = {u_ca_out_794[2:0], u_ca_out_793[5:3]};
assign col_out_795 = {u_ca_out_795[2:0], u_ca_out_794[5:3]};
assign col_out_796 = {u_ca_out_796[2:0], u_ca_out_795[5:3]};
assign col_out_797 = {u_ca_out_797[2:0], u_ca_out_796[5:3]};
assign col_out_798 = {u_ca_out_798[2:0], u_ca_out_797[5:3]};
assign col_out_799 = {u_ca_out_799[2:0], u_ca_out_798[5:3]};
assign col_out_800 = {u_ca_out_800[2:0], u_ca_out_799[5:3]};
assign col_out_801 = {u_ca_out_801[2:0], u_ca_out_800[5:3]};
assign col_out_802 = {u_ca_out_802[2:0], u_ca_out_801[5:3]};
assign col_out_803 = {u_ca_out_803[2:0], u_ca_out_802[5:3]};
assign col_out_804 = {u_ca_out_804[2:0], u_ca_out_803[5:3]};
assign col_out_805 = {u_ca_out_805[2:0], u_ca_out_804[5:3]};
assign col_out_806 = {u_ca_out_806[2:0], u_ca_out_805[5:3]};
assign col_out_807 = {u_ca_out_807[2:0], u_ca_out_806[5:3]};
assign col_out_808 = {u_ca_out_808[2:0], u_ca_out_807[5:3]};
assign col_out_809 = {u_ca_out_809[2:0], u_ca_out_808[5:3]};
assign col_out_810 = {u_ca_out_810[2:0], u_ca_out_809[5:3]};
assign col_out_811 = {u_ca_out_811[2:0], u_ca_out_810[5:3]};
assign col_out_812 = {u_ca_out_812[2:0], u_ca_out_811[5:3]};
assign col_out_813 = {u_ca_out_813[2:0], u_ca_out_812[5:3]};
assign col_out_814 = {u_ca_out_814[2:0], u_ca_out_813[5:3]};
assign col_out_815 = {u_ca_out_815[2:0], u_ca_out_814[5:3]};
assign col_out_816 = {u_ca_out_816[2:0], u_ca_out_815[5:3]};
assign col_out_817 = {u_ca_out_817[2:0], u_ca_out_816[5:3]};
assign col_out_818 = {u_ca_out_818[2:0], u_ca_out_817[5:3]};
assign col_out_819 = {u_ca_out_819[2:0], u_ca_out_818[5:3]};
assign col_out_820 = {u_ca_out_820[2:0], u_ca_out_819[5:3]};
assign col_out_821 = {u_ca_out_821[2:0], u_ca_out_820[5:3]};
assign col_out_822 = {u_ca_out_822[2:0], u_ca_out_821[5:3]};
assign col_out_823 = {u_ca_out_823[2:0], u_ca_out_822[5:3]};
assign col_out_824 = {u_ca_out_824[2:0], u_ca_out_823[5:3]};
assign col_out_825 = {u_ca_out_825[2:0], u_ca_out_824[5:3]};
assign col_out_826 = {u_ca_out_826[2:0], u_ca_out_825[5:3]};
assign col_out_827 = {u_ca_out_827[2:0], u_ca_out_826[5:3]};
assign col_out_828 = {u_ca_out_828[2:0], u_ca_out_827[5:3]};
assign col_out_829 = {u_ca_out_829[2:0], u_ca_out_828[5:3]};
assign col_out_830 = {u_ca_out_830[2:0], u_ca_out_829[5:3]};
assign col_out_831 = {u_ca_out_831[2:0], u_ca_out_830[5:3]};
assign col_out_832 = {u_ca_out_832[2:0], u_ca_out_831[5:3]};
assign col_out_833 = {u_ca_out_833[2:0], u_ca_out_832[5:3]};
assign col_out_834 = {u_ca_out_834[2:0], u_ca_out_833[5:3]};
assign col_out_835 = {u_ca_out_835[2:0], u_ca_out_834[5:3]};
assign col_out_836 = {u_ca_out_836[2:0], u_ca_out_835[5:3]};
assign col_out_837 = {u_ca_out_837[2:0], u_ca_out_836[5:3]};
assign col_out_838 = {u_ca_out_838[2:0], u_ca_out_837[5:3]};
assign col_out_839 = {u_ca_out_839[2:0], u_ca_out_838[5:3]};
assign col_out_840 = {u_ca_out_840[2:0], u_ca_out_839[5:3]};
assign col_out_841 = {u_ca_out_841[2:0], u_ca_out_840[5:3]};
assign col_out_842 = {u_ca_out_842[2:0], u_ca_out_841[5:3]};
assign col_out_843 = {u_ca_out_843[2:0], u_ca_out_842[5:3]};
assign col_out_844 = {u_ca_out_844[2:0], u_ca_out_843[5:3]};
assign col_out_845 = {u_ca_out_845[2:0], u_ca_out_844[5:3]};
assign col_out_846 = {u_ca_out_846[2:0], u_ca_out_845[5:3]};
assign col_out_847 = {u_ca_out_847[2:0], u_ca_out_846[5:3]};
assign col_out_848 = {u_ca_out_848[2:0], u_ca_out_847[5:3]};
assign col_out_849 = {u_ca_out_849[2:0], u_ca_out_848[5:3]};
assign col_out_850 = {u_ca_out_850[2:0], u_ca_out_849[5:3]};
assign col_out_851 = {u_ca_out_851[2:0], u_ca_out_850[5:3]};
assign col_out_852 = {u_ca_out_852[2:0], u_ca_out_851[5:3]};
assign col_out_853 = {u_ca_out_853[2:0], u_ca_out_852[5:3]};
assign col_out_854 = {u_ca_out_854[2:0], u_ca_out_853[5:3]};
assign col_out_855 = {u_ca_out_855[2:0], u_ca_out_854[5:3]};
assign col_out_856 = {u_ca_out_856[2:0], u_ca_out_855[5:3]};
assign col_out_857 = {u_ca_out_857[2:0], u_ca_out_856[5:3]};
assign col_out_858 = {u_ca_out_858[2:0], u_ca_out_857[5:3]};
assign col_out_859 = {u_ca_out_859[2:0], u_ca_out_858[5:3]};
assign col_out_860 = {u_ca_out_860[2:0], u_ca_out_859[5:3]};
assign col_out_861 = {u_ca_out_861[2:0], u_ca_out_860[5:3]};
assign col_out_862 = {u_ca_out_862[2:0], u_ca_out_861[5:3]};
assign col_out_863 = {u_ca_out_863[2:0], u_ca_out_862[5:3]};
assign col_out_864 = {u_ca_out_864[2:0], u_ca_out_863[5:3]};
assign col_out_865 = {u_ca_out_865[2:0], u_ca_out_864[5:3]};
assign col_out_866 = {u_ca_out_866[2:0], u_ca_out_865[5:3]};
assign col_out_867 = {u_ca_out_867[2:0], u_ca_out_866[5:3]};
assign col_out_868 = {u_ca_out_868[2:0], u_ca_out_867[5:3]};
assign col_out_869 = {u_ca_out_869[2:0], u_ca_out_868[5:3]};
assign col_out_870 = {u_ca_out_870[2:0], u_ca_out_869[5:3]};
assign col_out_871 = {u_ca_out_871[2:0], u_ca_out_870[5:3]};
assign col_out_872 = {u_ca_out_872[2:0], u_ca_out_871[5:3]};
assign col_out_873 = {u_ca_out_873[2:0], u_ca_out_872[5:3]};
assign col_out_874 = {u_ca_out_874[2:0], u_ca_out_873[5:3]};
assign col_out_875 = {u_ca_out_875[2:0], u_ca_out_874[5:3]};
assign col_out_876 = {u_ca_out_876[2:0], u_ca_out_875[5:3]};
assign col_out_877 = {u_ca_out_877[2:0], u_ca_out_876[5:3]};
assign col_out_878 = {u_ca_out_878[2:0], u_ca_out_877[5:3]};
assign col_out_879 = {u_ca_out_879[2:0], u_ca_out_878[5:3]};
assign col_out_880 = {u_ca_out_880[2:0], u_ca_out_879[5:3]};
assign col_out_881 = {u_ca_out_881[2:0], u_ca_out_880[5:3]};
assign col_out_882 = {u_ca_out_882[2:0], u_ca_out_881[5:3]};
assign col_out_883 = {u_ca_out_883[2:0], u_ca_out_882[5:3]};
assign col_out_884 = {u_ca_out_884[2:0], u_ca_out_883[5:3]};
assign col_out_885 = {u_ca_out_885[2:0], u_ca_out_884[5:3]};
assign col_out_886 = {u_ca_out_886[2:0], u_ca_out_885[5:3]};
assign col_out_887 = {u_ca_out_887[2:0], u_ca_out_886[5:3]};
assign col_out_888 = {u_ca_out_888[2:0], u_ca_out_887[5:3]};
assign col_out_889 = {u_ca_out_889[2:0], u_ca_out_888[5:3]};
assign col_out_890 = {u_ca_out_890[2:0], u_ca_out_889[5:3]};
assign col_out_891 = {u_ca_out_891[2:0], u_ca_out_890[5:3]};
assign col_out_892 = {u_ca_out_892[2:0], u_ca_out_891[5:3]};
assign col_out_893 = {u_ca_out_893[2:0], u_ca_out_892[5:3]};
assign col_out_894 = {u_ca_out_894[2:0], u_ca_out_893[5:3]};
assign col_out_895 = {u_ca_out_895[2:0], u_ca_out_894[5:3]};
assign col_out_896 = {u_ca_out_896[2:0], u_ca_out_895[5:3]};
assign col_out_897 = {u_ca_out_897[2:0], u_ca_out_896[5:3]};
assign col_out_898 = {u_ca_out_898[2:0], u_ca_out_897[5:3]};
assign col_out_899 = {u_ca_out_899[2:0], u_ca_out_898[5:3]};
assign col_out_900 = {u_ca_out_900[2:0], u_ca_out_899[5:3]};
assign col_out_901 = {u_ca_out_901[2:0], u_ca_out_900[5:3]};
assign col_out_902 = {u_ca_out_902[2:0], u_ca_out_901[5:3]};
assign col_out_903 = {u_ca_out_903[2:0], u_ca_out_902[5:3]};
assign col_out_904 = {u_ca_out_904[2:0], u_ca_out_903[5:3]};
assign col_out_905 = {u_ca_out_905[2:0], u_ca_out_904[5:3]};
assign col_out_906 = {u_ca_out_906[2:0], u_ca_out_905[5:3]};
assign col_out_907 = {u_ca_out_907[2:0], u_ca_out_906[5:3]};
assign col_out_908 = {u_ca_out_908[2:0], u_ca_out_907[5:3]};
assign col_out_909 = {u_ca_out_909[2:0], u_ca_out_908[5:3]};
assign col_out_910 = {u_ca_out_910[2:0], u_ca_out_909[5:3]};
assign col_out_911 = {u_ca_out_911[2:0], u_ca_out_910[5:3]};
assign col_out_912 = {u_ca_out_912[2:0], u_ca_out_911[5:3]};
assign col_out_913 = {u_ca_out_913[2:0], u_ca_out_912[5:3]};
assign col_out_914 = {u_ca_out_914[2:0], u_ca_out_913[5:3]};
assign col_out_915 = {u_ca_out_915[2:0], u_ca_out_914[5:3]};
assign col_out_916 = {u_ca_out_916[2:0], u_ca_out_915[5:3]};
assign col_out_917 = {u_ca_out_917[2:0], u_ca_out_916[5:3]};
assign col_out_918 = {u_ca_out_918[2:0], u_ca_out_917[5:3]};
assign col_out_919 = {u_ca_out_919[2:0], u_ca_out_918[5:3]};
assign col_out_920 = {u_ca_out_920[2:0], u_ca_out_919[5:3]};
assign col_out_921 = {u_ca_out_921[2:0], u_ca_out_920[5:3]};
assign col_out_922 = {u_ca_out_922[2:0], u_ca_out_921[5:3]};
assign col_out_923 = {u_ca_out_923[2:0], u_ca_out_922[5:3]};
assign col_out_924 = {u_ca_out_924[2:0], u_ca_out_923[5:3]};
assign col_out_925 = {u_ca_out_925[2:0], u_ca_out_924[5:3]};
assign col_out_926 = {u_ca_out_926[2:0], u_ca_out_925[5:3]};
assign col_out_927 = {u_ca_out_927[2:0], u_ca_out_926[5:3]};
assign col_out_928 = {u_ca_out_928[2:0], u_ca_out_927[5:3]};
assign col_out_929 = {u_ca_out_929[2:0], u_ca_out_928[5:3]};
assign col_out_930 = {u_ca_out_930[2:0], u_ca_out_929[5:3]};
assign col_out_931 = {u_ca_out_931[2:0], u_ca_out_930[5:3]};
assign col_out_932 = {u_ca_out_932[2:0], u_ca_out_931[5:3]};
assign col_out_933 = {u_ca_out_933[2:0], u_ca_out_932[5:3]};
assign col_out_934 = {u_ca_out_934[2:0], u_ca_out_933[5:3]};
assign col_out_935 = {u_ca_out_935[2:0], u_ca_out_934[5:3]};
assign col_out_936 = {u_ca_out_936[2:0], u_ca_out_935[5:3]};
assign col_out_937 = {u_ca_out_937[2:0], u_ca_out_936[5:3]};
assign col_out_938 = {u_ca_out_938[2:0], u_ca_out_937[5:3]};
assign col_out_939 = {u_ca_out_939[2:0], u_ca_out_938[5:3]};
assign col_out_940 = {u_ca_out_940[2:0], u_ca_out_939[5:3]};
assign col_out_941 = {u_ca_out_941[2:0], u_ca_out_940[5:3]};
assign col_out_942 = {u_ca_out_942[2:0], u_ca_out_941[5:3]};
assign col_out_943 = {u_ca_out_943[2:0], u_ca_out_942[5:3]};
assign col_out_944 = {u_ca_out_944[2:0], u_ca_out_943[5:3]};
assign col_out_945 = {u_ca_out_945[2:0], u_ca_out_944[5:3]};
assign col_out_946 = {u_ca_out_946[2:0], u_ca_out_945[5:3]};
assign col_out_947 = {u_ca_out_947[2:0], u_ca_out_946[5:3]};
assign col_out_948 = {u_ca_out_948[2:0], u_ca_out_947[5:3]};
assign col_out_949 = {u_ca_out_949[2:0], u_ca_out_948[5:3]};
assign col_out_950 = {u_ca_out_950[2:0], u_ca_out_949[5:3]};
assign col_out_951 = {u_ca_out_951[2:0], u_ca_out_950[5:3]};
assign col_out_952 = {u_ca_out_952[2:0], u_ca_out_951[5:3]};
assign col_out_953 = {u_ca_out_953[2:0], u_ca_out_952[5:3]};
assign col_out_954 = {u_ca_out_954[2:0], u_ca_out_953[5:3]};
assign col_out_955 = {u_ca_out_955[2:0], u_ca_out_954[5:3]};
assign col_out_956 = {u_ca_out_956[2:0], u_ca_out_955[5:3]};
assign col_out_957 = {u_ca_out_957[2:0], u_ca_out_956[5:3]};
assign col_out_958 = {u_ca_out_958[2:0], u_ca_out_957[5:3]};
assign col_out_959 = {u_ca_out_959[2:0], u_ca_out_958[5:3]};
assign col_out_960 = {u_ca_out_960[2:0], u_ca_out_959[5:3]};
assign col_out_961 = {u_ca_out_961[2:0], u_ca_out_960[5:3]};
assign col_out_962 = {u_ca_out_962[2:0], u_ca_out_961[5:3]};
assign col_out_963 = {u_ca_out_963[2:0], u_ca_out_962[5:3]};
assign col_out_964 = {u_ca_out_964[2:0], u_ca_out_963[5:3]};
assign col_out_965 = {u_ca_out_965[2:0], u_ca_out_964[5:3]};
assign col_out_966 = {u_ca_out_966[2:0], u_ca_out_965[5:3]};
assign col_out_967 = {u_ca_out_967[2:0], u_ca_out_966[5:3]};
assign col_out_968 = {u_ca_out_968[2:0], u_ca_out_967[5:3]};
assign col_out_969 = {u_ca_out_969[2:0], u_ca_out_968[5:3]};
assign col_out_970 = {u_ca_out_970[2:0], u_ca_out_969[5:3]};
assign col_out_971 = {u_ca_out_971[2:0], u_ca_out_970[5:3]};
assign col_out_972 = {u_ca_out_972[2:0], u_ca_out_971[5:3]};
assign col_out_973 = {u_ca_out_973[2:0], u_ca_out_972[5:3]};
assign col_out_974 = {u_ca_out_974[2:0], u_ca_out_973[5:3]};
assign col_out_975 = {u_ca_out_975[2:0], u_ca_out_974[5:3]};
assign col_out_976 = {u_ca_out_976[2:0], u_ca_out_975[5:3]};
assign col_out_977 = {u_ca_out_977[2:0], u_ca_out_976[5:3]};
assign col_out_978 = {u_ca_out_978[2:0], u_ca_out_977[5:3]};
assign col_out_979 = {u_ca_out_979[2:0], u_ca_out_978[5:3]};
assign col_out_980 = {u_ca_out_980[2:0], u_ca_out_979[5:3]};
assign col_out_981 = {u_ca_out_981[2:0], u_ca_out_980[5:3]};
assign col_out_982 = {u_ca_out_982[2:0], u_ca_out_981[5:3]};
assign col_out_983 = {u_ca_out_983[2:0], u_ca_out_982[5:3]};
assign col_out_984 = {u_ca_out_984[2:0], u_ca_out_983[5:3]};
assign col_out_985 = {u_ca_out_985[2:0], u_ca_out_984[5:3]};
assign col_out_986 = {u_ca_out_986[2:0], u_ca_out_985[5:3]};
assign col_out_987 = {u_ca_out_987[2:0], u_ca_out_986[5:3]};
assign col_out_988 = {u_ca_out_988[2:0], u_ca_out_987[5:3]};
assign col_out_989 = {u_ca_out_989[2:0], u_ca_out_988[5:3]};
assign col_out_990 = {u_ca_out_990[2:0], u_ca_out_989[5:3]};
assign col_out_991 = {u_ca_out_991[2:0], u_ca_out_990[5:3]};
assign col_out_992 = {u_ca_out_992[2:0], u_ca_out_991[5:3]};
assign col_out_993 = {u_ca_out_993[2:0], u_ca_out_992[5:3]};
assign col_out_994 = {u_ca_out_994[2:0], u_ca_out_993[5:3]};
assign col_out_995 = {u_ca_out_995[2:0], u_ca_out_994[5:3]};
assign col_out_996 = {u_ca_out_996[2:0], u_ca_out_995[5:3]};
assign col_out_997 = {u_ca_out_997[2:0], u_ca_out_996[5:3]};
assign col_out_998 = {u_ca_out_998[2:0], u_ca_out_997[5:3]};
assign col_out_999 = {u_ca_out_999[2:0], u_ca_out_998[5:3]};
assign col_out_1000 = {u_ca_out_1000[2:0], u_ca_out_999[5:3]};
assign col_out_1001 = {u_ca_out_1001[2:0], u_ca_out_1000[5:3]};
assign col_out_1002 = {u_ca_out_1002[2:0], u_ca_out_1001[5:3]};
assign col_out_1003 = {u_ca_out_1003[2:0], u_ca_out_1002[5:3]};
assign col_out_1004 = {u_ca_out_1004[2:0], u_ca_out_1003[5:3]};
assign col_out_1005 = {u_ca_out_1005[2:0], u_ca_out_1004[5:3]};
assign col_out_1006 = {u_ca_out_1006[2:0], u_ca_out_1005[5:3]};
assign col_out_1007 = {u_ca_out_1007[2:0], u_ca_out_1006[5:3]};
assign col_out_1008 = {u_ca_out_1008[2:0], u_ca_out_1007[5:3]};
assign col_out_1009 = {u_ca_out_1009[2:0], u_ca_out_1008[5:3]};
assign col_out_1010 = {u_ca_out_1010[2:0], u_ca_out_1009[5:3]};
assign col_out_1011 = {u_ca_out_1011[2:0], u_ca_out_1010[5:3]};
assign col_out_1012 = {u_ca_out_1012[2:0], u_ca_out_1011[5:3]};
assign col_out_1013 = {u_ca_out_1013[2:0], u_ca_out_1012[5:3]};
assign col_out_1014 = {u_ca_out_1014[2:0], u_ca_out_1013[5:3]};
assign col_out_1015 = {u_ca_out_1015[2:0], u_ca_out_1014[5:3]};
assign col_out_1016 = {u_ca_out_1016[2:0], u_ca_out_1015[5:3]};
assign col_out_1017 = {u_ca_out_1017[2:0], u_ca_out_1016[5:3]};
assign col_out_1018 = {u_ca_out_1018[2:0], u_ca_out_1017[5:3]};
assign col_out_1019 = {u_ca_out_1019[2:0], u_ca_out_1018[5:3]};
assign col_out_1020 = {u_ca_out_1020[2:0], u_ca_out_1019[5:3]};
assign col_out_1021 = {u_ca_out_1021[2:0], u_ca_out_1020[5:3]};
assign col_out_1022 = {u_ca_out_1022[2:0], u_ca_out_1021[5:3]};
assign col_out_1023 = {u_ca_out_1023[2:0], u_ca_out_1022[5:3]};
assign col_out_1024 = {u_ca_out_1024[2:0], u_ca_out_1023[5:3]};
assign col_out_1025 = {u_ca_out_1025[2:0], u_ca_out_1024[5:3]};
assign col_out_1026 = {u_ca_out_1026[2:0], u_ca_out_1025[5:3]};
assign col_out_1027 = {u_ca_out_1027[2:0], u_ca_out_1026[5:3]};
assign col_out_1028 = {u_ca_out_1028[2:0], u_ca_out_1027[5:3]};
assign col_out_1029 = {u_ca_out_1029[2:0], u_ca_out_1028[5:3]};
assign col_out_1030 = {u_ca_out_1030[2:0], u_ca_out_1029[5:3]};
assign col_out_1031 = {u_ca_out_1031[2:0], u_ca_out_1030[5:3]};
assign col_out_1032 = {u_ca_out_1032[2:0], u_ca_out_1031[5:3]};
assign col_out_1033 = {u_ca_out_1033[2:0], u_ca_out_1032[5:3]};
assign col_out_1034 = {u_ca_out_1034[2:0], u_ca_out_1033[5:3]};
assign col_out_1035 = {u_ca_out_1035[2:0], u_ca_out_1034[5:3]};
assign col_out_1036 = {u_ca_out_1036[2:0], u_ca_out_1035[5:3]};
assign col_out_1037 = {u_ca_out_1037[2:0], u_ca_out_1036[5:3]};
assign col_out_1038 = {u_ca_out_1038[2:0], u_ca_out_1037[5:3]};
assign col_out_1039 = {u_ca_out_1039[2:0], u_ca_out_1038[5:3]};
assign col_out_1040 = {u_ca_out_1040[2:0], u_ca_out_1039[5:3]};
assign col_out_1041 = {u_ca_out_1041[2:0], u_ca_out_1040[5:3]};
assign col_out_1042 = {u_ca_out_1042[2:0], u_ca_out_1041[5:3]};
assign col_out_1043 = {u_ca_out_1043[2:0], u_ca_out_1042[5:3]};
assign col_out_1044 = {u_ca_out_1044[2:0], u_ca_out_1043[5:3]};
assign col_out_1045 = {u_ca_out_1045[2:0], u_ca_out_1044[5:3]};
assign col_out_1046 = {u_ca_out_1046[2:0], u_ca_out_1045[5:3]};
assign col_out_1047 = {u_ca_out_1047[2:0], u_ca_out_1046[5:3]};
assign col_out_1048 = {u_ca_out_1048[2:0], u_ca_out_1047[5:3]};
assign col_out_1049 = {u_ca_out_1049[2:0], u_ca_out_1048[5:3]};
assign col_out_1050 = {u_ca_out_1050[2:0], u_ca_out_1049[5:3]};
assign col_out_1051 = {u_ca_out_1051[2:0], u_ca_out_1050[5:3]};
assign col_out_1052 = {u_ca_out_1052[2:0], u_ca_out_1051[5:3]};
assign col_out_1053 = {u_ca_out_1053[2:0], u_ca_out_1052[5:3]};
assign col_out_1054 = {u_ca_out_1054[2:0], u_ca_out_1053[5:3]};
assign col_out_1055 = {u_ca_out_1055[2:0], u_ca_out_1054[5:3]};
assign col_out_1056 = {u_ca_out_1056[2:0], u_ca_out_1055[5:3]};
assign col_out_1057 = {u_ca_out_1057[2:0], u_ca_out_1056[5:3]};
assign col_out_1058 = {u_ca_out_1058[2:0], u_ca_out_1057[5:3]};
assign col_out_1059 = {u_ca_out_1059[2:0], u_ca_out_1058[5:3]};
assign col_out_1060 = {u_ca_out_1060[2:0], u_ca_out_1059[5:3]};
assign col_out_1061 = {u_ca_out_1061[2:0], u_ca_out_1060[5:3]};
assign col_out_1062 = {u_ca_out_1062[2:0], u_ca_out_1061[5:3]};
assign col_out_1063 = {u_ca_out_1063[2:0], u_ca_out_1062[5:3]};
assign col_out_1064 = {u_ca_out_1064[2:0], u_ca_out_1063[5:3]};
assign col_out_1065 = {u_ca_out_1065[2:0], u_ca_out_1064[5:3]};
assign col_out_1066 = {u_ca_out_1066[2:0], u_ca_out_1065[5:3]};
assign col_out_1067 = {u_ca_out_1067[2:0], u_ca_out_1066[5:3]};
assign col_out_1068 = {u_ca_out_1068[2:0], u_ca_out_1067[5:3]};
assign col_out_1069 = {u_ca_out_1069[2:0], u_ca_out_1068[5:3]};
assign col_out_1070 = {u_ca_out_1070[2:0], u_ca_out_1069[5:3]};
assign col_out_1071 = {u_ca_out_1071[2:0], u_ca_out_1070[5:3]};
assign col_out_1072 = {u_ca_out_1072[2:0], u_ca_out_1071[5:3]};
assign col_out_1073 = {u_ca_out_1073[2:0], u_ca_out_1072[5:3]};
assign col_out_1074 = {u_ca_out_1074[2:0], u_ca_out_1073[5:3]};
assign col_out_1075 = {u_ca_out_1075[2:0], u_ca_out_1074[5:3]};
assign col_out_1076 = {u_ca_out_1076[2:0], u_ca_out_1075[5:3]};
assign col_out_1077 = {u_ca_out_1077[2:0], u_ca_out_1076[5:3]};
assign col_out_1078 = {u_ca_out_1078[2:0], u_ca_out_1077[5:3]};
assign col_out_1079 = {u_ca_out_1079[2:0], u_ca_out_1078[5:3]};
assign col_out_1080 = {u_ca_out_1080[2:0], u_ca_out_1079[5:3]};
assign col_out_1081 = {u_ca_out_1081[2:0], u_ca_out_1080[5:3]};
assign col_out_1082 = {u_ca_out_1082[2:0], u_ca_out_1081[5:3]};
assign col_out_1083 = {u_ca_out_1083[2:0], u_ca_out_1082[5:3]};
assign col_out_1084 = {u_ca_out_1084[2:0], u_ca_out_1083[5:3]};
assign col_out_1085 = {u_ca_out_1085[2:0], u_ca_out_1084[5:3]};
assign col_out_1086 = {u_ca_out_1086[2:0], u_ca_out_1085[5:3]};
assign col_out_1087 = {u_ca_out_1087[2:0], u_ca_out_1086[5:3]};
assign col_out_1088 = {u_ca_out_1088[2:0], u_ca_out_1087[5:3]};
assign col_out_1089 = {u_ca_out_1089[2:0], u_ca_out_1088[5:3]};
assign col_out_1090 = {u_ca_out_1090[2:0], u_ca_out_1089[5:3]};
assign col_out_1091 = {u_ca_out_1091[2:0], u_ca_out_1090[5:3]};
assign col_out_1092 = {u_ca_out_1092[2:0], u_ca_out_1091[5:3]};
assign col_out_1093 = {u_ca_out_1093[2:0], u_ca_out_1092[5:3]};
assign col_out_1094 = {u_ca_out_1094[2:0], u_ca_out_1093[5:3]};
assign col_out_1095 = {u_ca_out_1095[2:0], u_ca_out_1094[5:3]};
assign col_out_1096 = {u_ca_out_1096[2:0], u_ca_out_1095[5:3]};
assign col_out_1097 = {u_ca_out_1097[2:0], u_ca_out_1096[5:3]};
assign col_out_1098 = {u_ca_out_1098[2:0], u_ca_out_1097[5:3]};
assign col_out_1099 = {u_ca_out_1099[2:0], u_ca_out_1098[5:3]};
assign col_out_1100 = {u_ca_out_1100[2:0], u_ca_out_1099[5:3]};
assign col_out_1101 = {u_ca_out_1101[2:0], u_ca_out_1100[5:3]};
assign col_out_1102 = {u_ca_out_1102[2:0], u_ca_out_1101[5:3]};
assign col_out_1103 = {u_ca_out_1103[2:0], u_ca_out_1102[5:3]};
assign col_out_1104 = {u_ca_out_1104[2:0], u_ca_out_1103[5:3]};
assign col_out_1105 = {u_ca_out_1105[2:0], u_ca_out_1104[5:3]};
assign col_out_1106 = {u_ca_out_1106[2:0], u_ca_out_1105[5:3]};
assign col_out_1107 = {u_ca_out_1107[2:0], u_ca_out_1106[5:3]};
assign col_out_1108 = {u_ca_out_1108[2:0], u_ca_out_1107[5:3]};
assign col_out_1109 = {u_ca_out_1109[2:0], u_ca_out_1108[5:3]};
assign col_out_1110 = {u_ca_out_1110[2:0], u_ca_out_1109[5:3]};
assign col_out_1111 = {u_ca_out_1111[2:0], u_ca_out_1110[5:3]};
assign col_out_1112 = {u_ca_out_1112[2:0], u_ca_out_1111[5:3]};
assign col_out_1113 = {u_ca_out_1113[2:0], u_ca_out_1112[5:3]};
assign col_out_1114 = {u_ca_out_1114[2:0], u_ca_out_1113[5:3]};
assign col_out_1115 = {u_ca_out_1115[2:0], u_ca_out_1114[5:3]};
assign col_out_1116 = {u_ca_out_1116[2:0], u_ca_out_1115[5:3]};
assign col_out_1117 = {u_ca_out_1117[2:0], u_ca_out_1116[5:3]};
assign col_out_1118 = {u_ca_out_1118[2:0], u_ca_out_1117[5:3]};
assign col_out_1119 = {u_ca_out_1119[2:0], u_ca_out_1118[5:3]};
assign col_out_1120 = {u_ca_out_1120[2:0], u_ca_out_1119[5:3]};
assign col_out_1121 = {u_ca_out_1121[2:0], u_ca_out_1120[5:3]};
assign col_out_1122 = {u_ca_out_1122[2:0], u_ca_out_1121[5:3]};
assign col_out_1123 = {u_ca_out_1123[2:0], u_ca_out_1122[5:3]};
assign col_out_1124 = {u_ca_out_1124[2:0], u_ca_out_1123[5:3]};
assign col_out_1125 = {u_ca_out_1125[2:0], u_ca_out_1124[5:3]};
assign col_out_1126 = {u_ca_out_1126[2:0], u_ca_out_1125[5:3]};
assign col_out_1127 = {u_ca_out_1127[2:0], u_ca_out_1126[5:3]};
assign col_out_1128 = {u_ca_out_1128[2:0], u_ca_out_1127[5:3]};
assign col_out_1129 = {u_ca_out_1129[2:0], u_ca_out_1128[5:3]};
assign col_out_1130 = {u_ca_out_1130[2:0], u_ca_out_1129[5:3]};
assign col_out_1131 = {u_ca_out_1131[2:0], u_ca_out_1130[5:3]};
assign col_out_1132 = {u_ca_out_1132[2:0], u_ca_out_1131[5:3]};
assign col_out_1133 = {u_ca_out_1133[2:0], u_ca_out_1132[5:3]};
assign col_out_1134 = {u_ca_out_1134[2:0], u_ca_out_1133[5:3]};
assign col_out_1135 = {u_ca_out_1135[2:0], u_ca_out_1134[5:3]};
assign col_out_1136 = {u_ca_out_1136[2:0], u_ca_out_1135[5:3]};
assign col_out_1137 = {u_ca_out_1137[2:0], u_ca_out_1136[5:3]};
assign col_out_1138 = {u_ca_out_1138[2:0], u_ca_out_1137[5:3]};
assign col_out_1139 = {u_ca_out_1139[2:0], u_ca_out_1138[5:3]};
assign col_out_1140 = {u_ca_out_1140[2:0], u_ca_out_1139[5:3]};
assign col_out_1141 = {u_ca_out_1141[2:0], u_ca_out_1140[5:3]};
assign col_out_1142 = {u_ca_out_1142[2:0], u_ca_out_1141[5:3]};
assign col_out_1143 = {u_ca_out_1143[2:0], u_ca_out_1142[5:3]};
assign col_out_1144 = {u_ca_out_1144[2:0], u_ca_out_1143[5:3]};
assign col_out_1145 = {u_ca_out_1145[2:0], u_ca_out_1144[5:3]};
assign col_out_1146 = {u_ca_out_1146[2:0], u_ca_out_1145[5:3]};
assign col_out_1147 = {u_ca_out_1147[2:0], u_ca_out_1146[5:3]};
assign col_out_1148 = {u_ca_out_1148[2:0], u_ca_out_1147[5:3]};
assign col_out_1149 = {u_ca_out_1149[2:0], u_ca_out_1148[5:3]};
assign col_out_1150 = {u_ca_out_1150[2:0], u_ca_out_1149[5:3]};
assign col_out_1151 = {u_ca_out_1151[2:0], u_ca_out_1150[5:3]};
assign col_out_1152 = {u_ca_out_1152[2:0], u_ca_out_1151[5:3]};
assign col_out_1153 = {u_ca_out_1153[2:0], u_ca_out_1152[5:3]};
assign col_out_1154 = {u_ca_out_1154[2:0], u_ca_out_1153[5:3]};
assign col_out_1155 = {u_ca_out_1155[2:0], u_ca_out_1154[5:3]};
assign col_out_1156 = {u_ca_out_1156[2:0], u_ca_out_1155[5:3]};
assign col_out_1157 = {u_ca_out_1157[2:0], u_ca_out_1156[5:3]};
assign col_out_1158 = {u_ca_out_1158[2:0], u_ca_out_1157[5:3]};
assign col_out_1159 = {u_ca_out_1159[2:0], u_ca_out_1158[5:3]};
assign col_out_1160 = {u_ca_out_1160[2:0], u_ca_out_1159[5:3]};
assign col_out_1161 = {u_ca_out_1161[2:0], u_ca_out_1160[5:3]};
assign col_out_1162 = {u_ca_out_1162[2:0], u_ca_out_1161[5:3]};
assign col_out_1163 = {u_ca_out_1163[2:0], u_ca_out_1162[5:3]};
assign col_out_1164 = {u_ca_out_1164[2:0], u_ca_out_1163[5:3]};
assign col_out_1165 = {u_ca_out_1165[2:0], u_ca_out_1164[5:3]};
assign col_out_1166 = {u_ca_out_1166[2:0], u_ca_out_1165[5:3]};
assign col_out_1167 = {u_ca_out_1167[2:0], u_ca_out_1166[5:3]};
assign col_out_1168 = {u_ca_out_1168[2:0], u_ca_out_1167[5:3]};
assign col_out_1169 = {u_ca_out_1169[2:0], u_ca_out_1168[5:3]};
assign col_out_1170 = {u_ca_out_1170[2:0], u_ca_out_1169[5:3]};
assign col_out_1171 = {u_ca_out_1171[2:0], u_ca_out_1170[5:3]};
assign col_out_1172 = {u_ca_out_1172[2:0], u_ca_out_1171[5:3]};
assign col_out_1173 = {u_ca_out_1173[2:0], u_ca_out_1172[5:3]};
assign col_out_1174 = {u_ca_out_1174[2:0], u_ca_out_1173[5:3]};
assign col_out_1175 = {u_ca_out_1175[2:0], u_ca_out_1174[5:3]};
assign col_out_1176 = {u_ca_out_1176[2:0], u_ca_out_1175[5:3]};
assign col_out_1177 = {u_ca_out_1177[2:0], u_ca_out_1176[5:3]};
assign col_out_1178 = {u_ca_out_1178[2:0], u_ca_out_1177[5:3]};
assign col_out_1179 = {u_ca_out_1179[2:0], u_ca_out_1178[5:3]};
assign col_out_1180 = {u_ca_out_1180[2:0], u_ca_out_1179[5:3]};
assign col_out_1181 = {u_ca_out_1181[2:0], u_ca_out_1180[5:3]};
assign col_out_1182 = {u_ca_out_1182[2:0], u_ca_out_1181[5:3]};
assign col_out_1183 = {u_ca_out_1183[2:0], u_ca_out_1182[5:3]};
assign col_out_1184 = {u_ca_out_1184[2:0], u_ca_out_1183[5:3]};
assign col_out_1185 = {u_ca_out_1185[2:0], u_ca_out_1184[5:3]};
assign col_out_1186 = {u_ca_out_1186[2:0], u_ca_out_1185[5:3]};
assign col_out_1187 = {u_ca_out_1187[2:0], u_ca_out_1186[5:3]};
assign col_out_1188 = {u_ca_out_1188[2:0], u_ca_out_1187[5:3]};
assign col_out_1189 = {u_ca_out_1189[2:0], u_ca_out_1188[5:3]};
assign col_out_1190 = {u_ca_out_1190[2:0], u_ca_out_1189[5:3]};
assign col_out_1191 = {u_ca_out_1191[2:0], u_ca_out_1190[5:3]};
assign col_out_1192 = {u_ca_out_1192[2:0], u_ca_out_1191[5:3]};
assign col_out_1193 = {u_ca_out_1193[2:0], u_ca_out_1192[5:3]};
assign col_out_1194 = {u_ca_out_1194[2:0], u_ca_out_1193[5:3]};
assign col_out_1195 = {u_ca_out_1195[2:0], u_ca_out_1194[5:3]};
assign col_out_1196 = {u_ca_out_1196[2:0], u_ca_out_1195[5:3]};
assign col_out_1197 = {u_ca_out_1197[2:0], u_ca_out_1196[5:3]};
assign col_out_1198 = {u_ca_out_1198[2:0], u_ca_out_1197[5:3]};
assign col_out_1199 = {u_ca_out_1199[2:0], u_ca_out_1198[5:3]};
assign col_out_1200 = {u_ca_out_1200[2:0], u_ca_out_1199[5:3]};
assign col_out_1201 = {u_ca_out_1201[2:0], u_ca_out_1200[5:3]};
assign col_out_1202 = {u_ca_out_1202[2:0], u_ca_out_1201[5:3]};
assign col_out_1203 = {u_ca_out_1203[2:0], u_ca_out_1202[5:3]};
assign col_out_1204 = {u_ca_out_1204[2:0], u_ca_out_1203[5:3]};
assign col_out_1205 = {u_ca_out_1205[2:0], u_ca_out_1204[5:3]};
assign col_out_1206 = {u_ca_out_1206[2:0], u_ca_out_1205[5:3]};
assign col_out_1207 = {u_ca_out_1207[2:0], u_ca_out_1206[5:3]};
assign col_out_1208 = {u_ca_out_1208[2:0], u_ca_out_1207[5:3]};
assign col_out_1209 = {u_ca_out_1209[2:0], u_ca_out_1208[5:3]};
assign col_out_1210 = {u_ca_out_1210[2:0], u_ca_out_1209[5:3]};
assign col_out_1211 = {u_ca_out_1211[2:0], u_ca_out_1210[5:3]};
assign col_out_1212 = {u_ca_out_1212[2:0], u_ca_out_1211[5:3]};
assign col_out_1213 = {u_ca_out_1213[2:0], u_ca_out_1212[5:3]};
assign col_out_1214 = {u_ca_out_1214[2:0], u_ca_out_1213[5:3]};
assign col_out_1215 = {u_ca_out_1215[2:0], u_ca_out_1214[5:3]};
assign col_out_1216 = {u_ca_out_1216[2:0], u_ca_out_1215[5:3]};
assign col_out_1217 = {u_ca_out_1217[2:0], u_ca_out_1216[5:3]};
assign col_out_1218 = {u_ca_out_1218[2:0], u_ca_out_1217[5:3]};
assign col_out_1219 = {u_ca_out_1219[2:0], u_ca_out_1218[5:3]};
assign col_out_1220 = {u_ca_out_1220[2:0], u_ca_out_1219[5:3]};
assign col_out_1221 = {u_ca_out_1221[2:0], u_ca_out_1220[5:3]};
assign col_out_1222 = {u_ca_out_1222[2:0], u_ca_out_1221[5:3]};
assign col_out_1223 = {u_ca_out_1223[2:0], u_ca_out_1222[5:3]};
assign col_out_1224 = {u_ca_out_1224[2:0], u_ca_out_1223[5:3]};
assign col_out_1225 = {u_ca_out_1225[2:0], u_ca_out_1224[5:3]};
assign col_out_1226 = {u_ca_out_1226[2:0], u_ca_out_1225[5:3]};
assign col_out_1227 = {u_ca_out_1227[2:0], u_ca_out_1226[5:3]};
assign col_out_1228 = {u_ca_out_1228[2:0], u_ca_out_1227[5:3]};
assign col_out_1229 = {u_ca_out_1229[2:0], u_ca_out_1228[5:3]};
assign col_out_1230 = {u_ca_out_1230[2:0], u_ca_out_1229[5:3]};
assign col_out_1231 = {u_ca_out_1231[2:0], u_ca_out_1230[5:3]};
assign col_out_1232 = {u_ca_out_1232[2:0], u_ca_out_1231[5:3]};
assign col_out_1233 = {u_ca_out_1233[2:0], u_ca_out_1232[5:3]};
assign col_out_1234 = {u_ca_out_1234[2:0], u_ca_out_1233[5:3]};
assign col_out_1235 = {u_ca_out_1235[2:0], u_ca_out_1234[5:3]};
assign col_out_1236 = {u_ca_out_1236[2:0], u_ca_out_1235[5:3]};
assign col_out_1237 = {u_ca_out_1237[2:0], u_ca_out_1236[5:3]};
assign col_out_1238 = {u_ca_out_1238[2:0], u_ca_out_1237[5:3]};
assign col_out_1239 = {u_ca_out_1239[2:0], u_ca_out_1238[5:3]};
assign col_out_1240 = {u_ca_out_1240[2:0], u_ca_out_1239[5:3]};
assign col_out_1241 = {u_ca_out_1241[2:0], u_ca_out_1240[5:3]};
assign col_out_1242 = {u_ca_out_1242[2:0], u_ca_out_1241[5:3]};
assign col_out_1243 = {u_ca_out_1243[2:0], u_ca_out_1242[5:3]};
assign col_out_1244 = {u_ca_out_1244[2:0], u_ca_out_1243[5:3]};
assign col_out_1245 = {u_ca_out_1245[2:0], u_ca_out_1244[5:3]};
assign col_out_1246 = {u_ca_out_1246[2:0], u_ca_out_1245[5:3]};
assign col_out_1247 = {u_ca_out_1247[2:0], u_ca_out_1246[5:3]};
assign col_out_1248 = {u_ca_out_1248[2:0], u_ca_out_1247[5:3]};
assign col_out_1249 = {u_ca_out_1249[2:0], u_ca_out_1248[5:3]};
assign col_out_1250 = {u_ca_out_1250[2:0], u_ca_out_1249[5:3]};
assign col_out_1251 = {u_ca_out_1251[2:0], u_ca_out_1250[5:3]};
assign col_out_1252 = {u_ca_out_1252[2:0], u_ca_out_1251[5:3]};
assign col_out_1253 = {u_ca_out_1253[2:0], u_ca_out_1252[5:3]};
assign col_out_1254 = {u_ca_out_1254[2:0], u_ca_out_1253[5:3]};
assign col_out_1255 = {u_ca_out_1255[2:0], u_ca_out_1254[5:3]};
assign col_out_1256 = {u_ca_out_1256[2:0], u_ca_out_1255[5:3]};
assign col_out_1257 = {u_ca_out_1257[2:0], u_ca_out_1256[5:3]};
assign col_out_1258 = {u_ca_out_1258[2:0], u_ca_out_1257[5:3]};
assign col_out_1259 = {u_ca_out_1259[2:0], u_ca_out_1258[5:3]};
assign col_out_1260 = {u_ca_out_1260[2:0], u_ca_out_1259[5:3]};
assign col_out_1261 = {u_ca_out_1261[2:0], u_ca_out_1260[5:3]};
assign col_out_1262 = {u_ca_out_1262[2:0], u_ca_out_1261[5:3]};
assign col_out_1263 = {u_ca_out_1263[2:0], u_ca_out_1262[5:3]};
assign col_out_1264 = {u_ca_out_1264[2:0], u_ca_out_1263[5:3]};
assign col_out_1265 = {u_ca_out_1265[2:0], u_ca_out_1264[5:3]};
assign col_out_1266 = {u_ca_out_1266[2:0], u_ca_out_1265[5:3]};
assign col_out_1267 = {u_ca_out_1267[2:0], u_ca_out_1266[5:3]};
assign col_out_1268 = {u_ca_out_1268[2:0], u_ca_out_1267[5:3]};
assign col_out_1269 = {u_ca_out_1269[2:0], u_ca_out_1268[5:3]};
assign col_out_1270 = {u_ca_out_1270[2:0], u_ca_out_1269[5:3]};
assign col_out_1271 = {u_ca_out_1271[2:0], u_ca_out_1270[5:3]};
assign col_out_1272 = {u_ca_out_1272[2:0], u_ca_out_1271[5:3]};
assign col_out_1273 = {u_ca_out_1273[2:0], u_ca_out_1272[5:3]};
assign col_out_1274 = {u_ca_out_1274[2:0], u_ca_out_1273[5:3]};
assign col_out_1275 = {u_ca_out_1275[2:0], u_ca_out_1274[5:3]};
assign col_out_1276 = {u_ca_out_1276[2:0], u_ca_out_1275[5:3]};
assign col_out_1277 = {u_ca_out_1277[2:0], u_ca_out_1276[5:3]};
assign col_out_1278 = {u_ca_out_1278[2:0], u_ca_out_1277[5:3]};
assign col_out_1279 = {u_ca_out_1279[2:0], u_ca_out_1278[5:3]};
assign col_out_1280 = {u_ca_out_1280[2:0], u_ca_out_1279[5:3]};
assign col_out_1281 = {u_ca_out_1281[2:0], u_ca_out_1280[5:3]};
assign col_out_1282 = {u_ca_out_1282[2:0], u_ca_out_1281[5:3]};
assign col_out_1283 = {u_ca_out_1283[2:0], u_ca_out_1282[5:3]};
assign col_out_1284 = {u_ca_out_1284[2:0], u_ca_out_1283[5:3]};
assign col_out_1285 = {u_ca_out_1285[2:0], u_ca_out_1284[5:3]};
assign col_out_1286 = {u_ca_out_1286[2:0], u_ca_out_1285[5:3]};
assign col_out_1287 = {u_ca_out_1287[2:0], u_ca_out_1286[5:3]};
assign col_out_1288 = {{3{1'b0}}, u_ca_out_1287[5:3]};

//---------------------------------------------------------


endmodule
module xpb_5_740
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5b3ee2ab8bf542db3a2ec0fc227618aea89cf0804d94391174eabc72a617828e5e2a2e688630c8c2e2cadf2d65d0fabbda7776e42e03e744c1a4d201c73dfb79f76b89b479c1aec0f4438bc2439e27d2ed1a66ceda58e83aaed30fe2f6004091c543df1959131c6fcc121cc53d4aee64e22fbfb619cf48ed008b02496e61349c;
    5'b00010 : xpb = 1024'h5d0800155fc50eda9580a213491ea0bdfc3ddcfc5b0d1ab6bf8bf8f992c5814b90bdf58423b12f726377f13e843e4ad50d4c5e23954fe3dd2aa64a553a982427a87deba43f2603cd5ed14e1ee608b74e62fd405282ba364a8198dcb31d5de915b802c09015d4052116452ab82c5b6a07585a089e35334a9baa6898e53e002cd;
    5'b00011 : xpb = 1024'h610f62ace1f193c8e386cb1d570802ba8860ce5013450abce0e37c023f43daa317360dc0c86bdbba09025e414e14df692b4c3cc66758e582944f36a71ae77dbc71f3686ebdb40efdca30a0a431feb347d34a3ad402848b9f56ec9dae27d61f2320c40b225a705cc1dd766f70c010a50557b5603ffd227d96bb318bd7c2413769;
    5'b00100 : xpb = 1024'hba10002abf8a1db52b014426923d417bf87bb9f8b61a356d7f17f1f3258b0297217beb0847625ee4c6efe27d087c95aa1a98bc472a9fc7ba554c94aa7530484f50fbd7487e4c079abda29c3dcc116e9cc5fa80a505746c950331b9663abbd22b700581202ba80a422c8a557058b6d40eb0b4113c6a66953754d131ca7c0059a;
    5'b00101 : xpb = 1024'h66dfe2ae37ede4b68cded53e8b99ecc66824ac1fd8f5dc684cdc3b91d87032b7d041ed190aa6eeb12f39dd553658c4167c2102a8a0ade3c066f99b4c6e90fffeec7b472901a66f3aa01db586205f3ebcb97a0ed92ab02f03ff062b7959abfdb47c44372b5bcd9d13eedac21c42d65ba5cd3b00c9e075b24075d8156616213a36;
    5'b00110 : xpb = 1024'h1171800401f4f2c8fc081e639db5be239f4b996f5112750243ea3eaecb85083e2b239e08c6b138e572a67d3bb8cbae07f27e51a6abfefab977ff2deffafc86c76f979c2ecbd720b681c73ea5cb21a25eb28f7c0f7882ea2df84ca96195819bb41280841b0417c0f6342cf802885123e16090e19da9f99dfd2ff39caafba00867;
    5'b00111 : xpb = 1024'h6cb062af8dea35a43636df5fc02bd6d247e889ef9ea6ae13b8d4fb21719c8acc894dcc714ce201a855715c691e9ca8c3ccf5c88ada02e1fe39a3fff1c23a8241670325e34598cf77760aca680ebfca319fa9e2de52dbd268a71fb9448b81dc45d7c463345d2add66003f14c7c59c124642c0a153c3c8e6ea307e9ef46a013d03;
    5'b01000 : xpb = 1024'h1742000557f143b6a5602884d247a82f7f0f773f16c346adafe2fe3e64b16052e42f7d6108ec4bdc98ddfc4fa10f92b543531788e553f8f74aa992954ea60909ea1f7ae90fc980f357b45387b9822dd398bf5014a0ae8d92a066372cc7577a456e00b0240575014845914aae0b16da81d61682278d4cd2a6ea9a26394f800b34;
    5'b01001 : xpb = 1024'h7280e2b0e3e68691df8ee980f4bdc0de27ac67bf64577fbf24cdbab10ac8e2e14259abc98f1d149f7ba8db7d06e08d711dca8e6d1357e03c0c4e649715e40483e18b049d898b2fb44bf7df49fd2055a685d9b6e37b0775cd4f39470fbd57bad733448f3d5e881db811a367734861c8e6b84641dda71c1b93eb252882bde13fd0;
    5'b01010 : xpb = 1024'h1d128006aded94a44eb832a606d9923b5ed3550edc7418591bdbbdcdfdddb8679d3b5cb94b275ed3bf157b63895377629427dd6b1ea8f7351d53f73aa24f8b4c64a759a353bbe1302da16869a7e2b9487eef2419c8da30f7487fc4f7f92d58d6c980dc2d06d2419a56f59d598ddc91224b9c22b170a00750a540afc7a3600e01;
    5'b01011 : xpb = 1024'h785162b239e2d77f88e6f3a2294faaea0770458f2a08516a90c67a40a3f53af5fb658b21d1582796a1e05a90ef24721e6e9f544f4cacde79def8c93c698d86c65c12e357cd7d8ff121e4f42beb80e11b6c098ae8a3331931f752d4daef2d99688ec4bb465fe55e0a2307ba1ecb277f872dcbe2678a6f503da5cbb21111c1429d;
    5'b01100 : xpb = 1024'h22e3000803e9e591f8103cc73b6b7c473e9732dea224ea0487d47d5d970a107c56473c118d6271cae54cfa7771975c0fe4fca34d57fdf572effe5bdff5f90d8edf2f385d97ae416d038e7d4b964344bd651ef81ef105d45bf09952c32b03376825010836082f81ec6859f00510a247c2c121c33b53f33bfa5fe73955f74010ce;
    5'b01101 : xpb = 1024'h7e21e2b38fdf286d323efdc35de194f5e734235eefb92315fcbf39d03d21930ab4716a7a13933a8dc817d9a4d76856cbbf741a318601dcb7b1a32de1bd370908d69ac212116ff02df7d2090dd9e16c9052395eedcb5ebc969f6c62a6210377f9ea44e74f61429e5c346c0cca4ded3627a35182f16dc284e760723b9f65a1456a;
    5'b01110 : xpb = 1024'h28b3800959e6367fa16846e86ffd66531e5b10ae67d5bbaff3cd3ced303668910f531b69cf9d84c20b84798b59db40bd35d1692f9152f3b0c2a8c08549a28fd159b71717dba0a1a9d97b922d84a3d0324b4ecc24193177c098b2e08e5cd915f98081343f098cc23e79be42b09367fe6336a763c5374670a41a8dc2e44b20139b;
    5'b01111 : xpb = 1024'h83f262b4e5db795adb9707e492737f01c6f8012eb569f4c168b7f95fd64deb1f6d7d49d255ce4d84ee4f58b8bfac3b791048e013bf56daf5844d928710e08b4b5122a0cc5562506acdbf1defc841f805386932f2f38a5ffb4785f07152d9568b45c51358629fdeae45d05f75d0b2ecc818d7237b5115b9911b18c52db9814837;
    5'b10000 : xpb = 1024'h2e84000aafe2876d4ac05109a48f505efe1eee7e2d868d5b5fc5fc7cc962c0a5c85efac211d897b931bbf89f421f256a86a62f11caa7f1ee9553252a9d4c1213d43ef5d21f9301e6af68a70f73045ba7317ea029415d1b2540cc6e598eaef48adc0160480aea02908b22955c162db503ac2d044f1a99a54dd5344c729f001668;
    5'b10001 : xpb = 1024'h89c2e2b63bd7ca4884ef1205c705690da6bbdefe7b1ac66cd4b0b8ef6f7a43342689292a9809607c1486d7cca7f02026611da5f5f8abd93356f7f72c648a0d8dcbaa7f869954b0a7a3ac32d1b6a2837a1e9906f81bb6035fef9f7e3c84af351ca1453f6163fd1f005734b2215378a3688e5cc4053468ee3ad5bf4ebc0d614b04;
    5'b10010 : xpb = 1024'h3454800c05ded85af4185b2ad9213a6adde2cc4df3375f06cbbebc0c628f18ba816ada1a5413aab057f377b32a630a17d77af4f403fcf02c67fd89cff0f594564ec6d48c638562238555bbf16164e71c17ae742e6988be89e8e5fc24c084d31c37818c510c4742e29c86e80798f36ba421b2a4d8fdecd9f78fdad600f2e01935;
    5'b10011 : xpb = 1024'h8f9362b791d41b362e471c26fb975319867fbcce40cb981840a9787f08a69b48df950882da4473733abe56e0903404d3b1f26bd83200d77129a25bd1b8338fd046325e40dd4710e4799947b3a5030eef04c8dafd43e1a6c497b90c07b68513adfcc56b6a655a5f52689904ccd63e5a0903e2648f17bc22e49065d84a61414dd1;
    5'b10100 : xpb = 1024'h3a25000d5bdb29489d70654c0db32476bda6aa1db8e830b237b77b9bfbbb70cf3a76b972964ebda77e2af6c712a6eec5284fbad63d51ee6a3aa7ee75449f1698c94eb346a777c2605b42d0d34fc57290fdde483391b461ee90ff89eff25ab1ad9301b85a0da48334adeb3ab31bb9224497384562e1400ea14a815f8f46c01c02;
    5'b10101 : xpb = 1024'h9563e2b8e7d06c23d79f264830293d2566439a9e067c69c3aca2380ea1d2f35d98a0e7db1c7f866a60f5d5f47877e98102c731ba6b55d5aefc4cc0770bdd1212c0ba3cfb213971214f865c9593639a63eaf8af026c0d4a293fd299d2e85af23f5845977366b79fa479fd5778590410a979680518fb0f578e4b0c61d8b521509e;
    5'b10110 : xpb = 1024'h3ff5800eb1d77a3646c86f6d42450e829d6a87ed7e99025da3b03b2b94e7c8e3f38298cad889d09ea46275dafaead372792480b876a6eca80d52531a984898db43d69200eb6a229d312fe5b53e25fe05e40e1c38b9e00553391917bb2430903eee81e4630f01c386bf4f8d5e9e7ed8e50cbde5ecc493434b0527e91d9aa01ecf;
    5'b10111 : xpb = 1024'h9b3462ba3dccbd1180f7306964bb27314607786dcc2d3b6f189af79e3aff4b7251acc7335eba9961872d550860bbce2e539bf79ca4aad3eccef7251c5f8694553b421bb5652bd15e2573717781c425d8d12883079438ed8de7ec279e1a30d0d0b3c5c37c6814dff68b61aa23dbc9c749eeeda5a2de628c3805b2eb670901536b;
    5'b11000 : xpb = 1024'h45c6001007d3cb23f020798e76d6f88e7d2e65bd4449d4090fa8fabb2e1420f8ac8e78231ac4e395ca99f4eee32eb81fc9f9469aaffbeae5dffcb7bfebf21b1dbe5e70bb2f5c82da071cfa972c86897aca3df03de20ba8b7e132a58656066ed04a02106c105f03d8d0b3e00a21448f8582438676a7e677f4bfce72abee80219c;
    5'b11001 : xpb = 1024'ha104e2bb93c90dff2a4f3a8a994d113d25cb563d91de0d1a8493b72dd42ba3870ab8a68ba0f5ac58ad64d41c48ffb2dba470bd7eddffd22aa1a189c1b3301697b5c9fa6fa91e319afb6086597024b14db758570cbc6490f29005b5694c06af620f45ef85697220489cc5fccf5e8f7dea6473462cc1b5c0e1c05974f55ce15638;
    5'b11010 : xpb = 1024'h4b9680115dd01c11997883afab68e29a5cf2438d09faa5b47ba1ba4ac740790d659a577b5cfff68cf0d17402cb729ccd1ace0c7ce950e923b2a71c653f9b9d6038e64f75734ee316dd0a0f791ae714efb06dc4430a374c1c894c335187dc4d61a5823c7511bc442ae21832b5a40a4625f7c927008b39ac9e7a74fc3a42602469;
    5'b11011 : xpb = 1024'ha6d562bce9c55eecd3a744abcddefb49058f340d578edec5f08c76bd6d57fb9bc3c485e3e330bf4fd39c533031439788f54583611754d068744bee6706d998da3051d929ed1091d7d14d9b3b5e853cc29d882b11e4903457381f43347ddc8df36ac61b8e6acf609aae2a4f7ae155348ad9f8e6b6a508f58b7afffe83b0c15905;
    5'b11100 : xpb = 1024'h51670012b3cc6cff42d08dd0dffacca63cb6215ccfab775fe79a79da606cd1221ea636d39f3b09841708f316b3b6817a6ba2d25f22a5e7618551810a93451fa2b36e2e2fb7414353b2f7245b0947a064969d98483262ef813165c11cb9b22bf30102687e1319847cf37c856126cffcc66d4ec78a6e8ce148351b85c896402736;
    5'b11101 : xpb = 1024'haca5e2be3fc1afda7cff4ecd0270e554e55311dd1d3fb0715c85364d068453b07cd0653c256bd246f9d3d24419877c36461a494350a9cea646f6530c5a831b1caad9b7e43102f214a73ab01d4ce5c83783b7ff170cbbd7bbe038d0ffafb26c84c64647976c2ca0ecbf8ea226641aeb2b4f7e8740885c2a3535a6881204a15bd2;
    5'b11110 : xpb = 1024'h5737801409c8bdecec2897f2148cb6b21c79ff2c955c490b53933969f9992936d7b2162be1761c7b3d40722a9bfa6627bc7798415bfae59f57fbe5afe6eea1e52df60ce9fb33a39088e4393cf7a82bd97ccd6c4d5a8e92e5d97f4ee7eb880a845c8294871476c4cf04e0d80ca995b366e2d4681451e015f1efc20f56ea202a03;
    5'b11111 : xpb = 1024'h1c91d69d3cfcbff5b51e11726a8880f53a0ec7c0d78e1a54aa13c86ecadfebd3293c71b9d8066af80ad12111e6d501932d4e73f674bfc9869017853735a28adb11261efc564550c6a8dc25ca26a8f7b75e2d983a8614e0fd2c5ccd0275da883f2bee176bcc0e8b14a330df2ef107ba2762a48e81b6401aea9dd969bcf9ef834;
    endcase
end

endmodule

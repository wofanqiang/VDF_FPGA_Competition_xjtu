module xpb_5_370
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h76924e4de078bf74252ef23221bd98503f2cfeb451f94f2da618fd0f0fd83dd441274a45348e1778811bfb2fd5ef09a3f51f36426d1dade54f93133edce913265ba9429ee780e5cbf033f3fb6fb2fd8d4cc5dcd69aa152f6126706f6bc8e240f2951e9d3e52a7fc5e8fb9c76fefe3743fdfb3a4ff0a84783984b9714e9fa35b8;
    5'b00010 : xpb = 1024'h3c775745ff034a1f7f586c8d3320e94f0ce3fa37ce7afde3ce5540c86cadcea07f0617119ef5b06262d9b718c880027d8624449eb7888b7eee86e71f7effb19b4303508f1f70ce52cdcde554468a36e9a586c014a8bc78db6f417bf2bef1a58c239c417e198c06fe4b37520f062c485ead1c95bd910531d6ea27b3254b120505;
    5'b00011 : xpb = 1024'h25c603e1d8dd4cad981e6e844843a4dda9af5bb4afcac99f6918481c9835f6cbce4e3de095d494c44977301bb10fb57172952fb01f369188d7abb00211650102a5d5e7f5760b6d9ab67d6ad1d617045fe47a352b6d79ec0cc1bf0eec15527091de699284ded8e36ad7307a70d5a59795c3df12b31621c2a3c03cf35ac29d452;
    5'b00100 : xpb = 1024'h78eeae8bfe06943efeb0d91a6641d29e19c7f46f9cf5fbc79caa8190d95b9d40fe0c2e233deb60c4c5b36e31910004fb0c48893d6f1116fddd0dce3efdff63368606a11e3ee19ca59b9bcaa88d146dd34b0d80295178f1b6de82f7e57de34b18473882fc33180dfc966ea41e0c5890bd5a392b7b220a63add44f664a96240a0a;
    5'b00101 : xpb = 1024'h3ed3b7841c911eea58da537577a5239ce77eeff31977aa7dc4e6c54a36312e0d3beafaefa852f9aea7712a1a8390fdd49d4d9799b97bf4977c01a21fa01601ab6d60af0e76d1852c7935bc0163eba72fa3ce63675f94179c3b5d6ce18046cc954182daa667799534f8aa59b61386a1d8095a86e8c2674e01262b825af73bd957;
    5'b00110 : xpb = 1024'h4b8c07c3b1ba995b303cdd08908749bb535eb7695f95933ed2309039306bed979c9c7bc12ba9298892ee6037621f6ae2e52a5f603e6d2311af57600422ca02054babcfeaec16db356cfad5a3ac2e08bfc8f46a56daf3d819837e1dd82aa4e123bcd32509bdb1c6d5ae60f4e1ab4b2f2b87be25662c4385478079e6b5853a8a4;
    5'b00111 : xpb = 1024'h7b4b0eca1b946909d832c002aac60cebf462ea2ae7f2a861933c0612a2defcadbaf112014748aa110a4ae1334c1100522371dc38710480166a88893f1f15b346b063ff9d9642537f4703a155aa75de194955237c08509077aa9ee8d43f387221651f1c2481059c3343e1abc519b2ea36b6771ca6536c7fd810533580424dde5c;
    5'b01000 : xpb = 1024'h413017c23a1ef3b5325c3a5dbc295deac219e5ae64745717bb7849cbffb48d79f8cfdecdb1b042faec089d1c3ea1f92bb476ea94bb6f5db0097c5d1fc12c51bb97be0d8dce323c06249d92ae814d1775a21606ba166bb65d07795dd0419bf39e5f6973ceb567236ba61d615d20e0fb5165987813f3c96a2b622f5190a365ada9;
    5'b01001 : xpb = 1024'h71520ba58a97e608c85b4b8cd8caee98fd0e131e0f605cde3b48d855c8a1e4636aeab9a1c17dbe4cdc659053132f205457bf8f105da3b49a87031006342f0307f181b7e0622248d02378407582450d1fad6e9f82486dc426453d2cc43ff751b59b3cb78e9c8aaa4085916f5280f0c6c14b9d3819426547eb40b6da1047d7cf6;
    5'b01010 : xpb = 1024'h7da76f0839223dd4b1b4a6eaef4a4739cefddfe632ef54fb89cd8a946c625c1a77d5f5df50a5f35d4ee254350721fba93a9b2f3372f7e92ef803443f402c0356dac15e1ceda30a58f26b7802c7d74e5f479cc6cebf282f3876bad9c3008d992a8305b54ccef32a69f154b36c270d43b012b50dd184ce9c024c5704b5ee77b2ae;
    5'b01011 : xpb = 1024'h438c780057acc8800bde214600ad98389cb4db69af7103b1b209ce4dc937ece6b5b4c2abbb0d8c4730a0101df9b2f482cba03d8fbd62c6c896f7181fe242a1cbc21b6c0d2592f2dfd005695b9eae87bba05daa0ccd43551dd3954ebf02f11aa77d500cf70354b1a2539069042e3b54cac1d6693f252b86559e3320c64f8f81fb;
    5'b01100 : xpb = 1024'h97180f87637532b66079ba11210e9376a6bd6ed2bf2b267da461207260d7db2f3938f7825752531125dcc06ec43ed5c5ca54bec07cda46235eaec0084594040a97579fd5d82db66ad9f5ab47585c117f91e8d4adb5e7b03306fc3bb05549c24779a64a137b638dab5cc1e9c356965e570f7c4acc58870a8f00f3cd6b0a75148;
    5'b01101 : xpb = 1024'h8003cf4656b0129f8b368dd333ce8187a998d5a17dec0195805f0f1635e5bb8734bad9bd5a033ca99379c736c232f70051c4822e74eb5247857dff3f61425367051ebc9c4503c1329dd34eafe538bea545e46a2175ffcdf942d6cab1c1e2c033a0ec4e751ce0b8a09ec7bb1334679d296ef2fefcb630b82c885ad3eb9aa18700;
    5'b01110 : xpb = 1024'h45e8d83e753a9d4ae560082e4531d286774fd124fa6db04ba89b52cf92bb4c537299a689c46ad5937537831fb4c3efd9e2c9908abf562fe12471d3200358f1dbec78ca8c7cf3a9b97b6d4008bc0ff8019ea54d5f841af3de9fb13fadc44641b09b36a61f51423fd9010370ab3b95ae441e145a6a568da27fda36effbfbb9564d;
    5'b01111 : xpb = 1024'hbcde13693c527f63f898289569523854506cca876ef5f01d0d79688ef90dd1fb07873562ed26e7d56f53f08a754e8b373ce9ee709c10d7ac365a700a56f9050d3d2d87cb4e392405907316192e7315df766309d923619c3fc8bb4a9c6a9c32d9580fdc985a3c711633f264342c3bf5ecd35b5d7f6ea8cd32c130c0c5cd1259a;
    5'b10000 : xpb = 1024'h82602f84743de76a64b874bb7852bbd58433cb5cc8e8ae2f76f09397ff691af3f19fbd9b636085f5d8113a387d43f25768edd52976debb6012f8ba3f8258a3772f7c1b1b9c64780c493b255d029a2eeb442c0d742cd76cba0ef2bba08337e73cbed2e79d6ace46d74c3ac2ba41c1f6a2cb30f027e792d456c45ea32146cb5b52;
    5'b10001 : xpb = 1024'h4845387c92c87215bee1ef1689b60cd451eac6e0456a5ce59f2cd7515c3eabc02f7e8a67cdc81edfb9cef6216fd4eb30f9f2e385c14998f9b1ec8e20246f41ec16d6290bd454609326d516b5d97168479cecf0b23af2929f6bcd309c859b68b9b91d3f479f2fce0fae76785248f007bd7a524b9587efbeaa163abf31a7e32a9f;
    5'b10010 : xpb = 1024'he2a4174b152fcc1190b69719b195dd31fa1c263c1ec0b9bc7691b0ab9143c8c6d5d5734382fb7c99b8cb20a6265e40a8af7f1e20bb4769350e06200c685e060fe3036fc0c44491a046f080eb048a1a3f5add3f0490db884c8a7a59887feea36b36796f1d391554810b22dea501e18d82973a703284ca8fd6816db4208faf9ec;
    5'b10011 : xpb = 1024'h84bc8fc291cbbc353e3a5ba3bcd6f6235ecec11813e55ac96d821819c8ec7a60ae84a1796cbdcf421ca8ad3a3854edae8017282478d22478a073753fa36ef38759d9799af3c52ee5f4a2fc0a1ffb9f314273b0c6e3af0b7adb0eac8f448d0e45dcb980c5b8bbd50df9adca614f1c501c276ee15318f4f08100627256f2f52fa4;
    5'b10100 : xpb = 1024'h4aa198bab05646e09863d5fece3a47222c85bc9b9067097f95be5bd325c20b2cec636e45d725682bfe6669232ae5e688111c3680c33d02123f674920458591fc4133878b2bb5176cd23ced62f6d2d88d9b349404f1ca316037e9218b46f08fc2d703d86fed1d5c465be97ff9564a6136d6903cc0b951dad4523e8e67540cfef1;
    5'b10101 : xpb = 1024'h1086a1b2cee0d18bf28d5059df9d9820fa3cb81f0ce8b835bdfa9f8c82979bf92a423b12418d0115e024250c1d76df61a22144dd0da7dfabde5b1d00e79c3071288d957b63a4fff3afd6debbcdaa11e9f3f57742ffe5574594c396874954113fd14e301a217ee37ebe2535915d78725185b1982e59aec527a41aaa77b524ce3e;
    5'b10110 : xpb = 1024'h8718f000af59910017bc428c015b30713969b6d35ee2076364139c9b926fd9cd6b698557761b188e6140203bf365e90597407b1f7ac58d912dee303fc48543978436d81a4b25e5bfa00ad2b73d5d0f7740bb54199a86aa3ba72a9d7e05e2354efaa019ee06a96344a720d2085c76a99583acd27e4a570cab3c66418c9f1f03f6;
    5'b10111 : xpb = 1024'h4cfdf8f8cde41bab71e5bce712be81700720b256db63b6198c4fe054ef456a99a9485223e082b17842fddc24e5f6e1df2845897bc5306b2acce20420669be20c6b90e60a8315ce467da4c410143448d3997c3757a8a1d0210405127a0845b6cbf4ea71983b0aea7d095c87a063a4bab032ce2debeab3f6fe8e425d9d0036d343;
    5'b11000 : xpb = 1024'h12e301f0ec6ea656cc0f37422421d26ed4d7adda57e564cfb48c240e4c1afb65e7271ef04aea4a6224bb980dd887dab8b94a97d80f9b48c46bd5d80108b2808152eaf3fabb05b6cd5b3eb568eb0b822ff23d1a95b6bcf60660df87760aa93848ef34c9426f6c71b56b983d386ad2cbcae1ef89598b10e151e01e79ad614ea290;
    5'b11001 : xpb = 1024'h8975503ecce765caf13e297445df6abf1404ac8ea9deb3fd5aa5211d5bf3393a284e69357f7861daa5d7933dae76e45cae69ce1a7cb8f6a9bb68eb3fe59b93a7ae943699a2869c994b72a9645abe7fbd3f02f76c515e48fc73468e6cc7375c581886b3165496f17b5493d9af69d1030edfeac3a97bb928d5786a10c24b48d848;
    5'b11010 : xpb = 1024'h4f5a5936eb71f0764b67a3cf5742bbbde1bba812266062b382e164d6b8c8ca06662d3601e9dffac487954f26a107dd363f6edc76c723d4435a5cbf2087b2321c95ee4489da768520290c9abd3195b91997c3daaa5f796ee1d0210368c99addd512d10ac088f878b3b6cf8f4770ff14298f0c1f171c161328ca462cd2ac60a795;
    5'b11011 : xpb = 1024'h153f622f09fc7b21a5911e2a68a60cbcaf72a395a2e21169ab1da890159e5ad2a40c02ce544793ae69530b0f9398d60fd073ead3118eb1dcf950930129c8d0917d48527a12666da706a68c16086cf275f084bde86d9494c72cfb7864cbfe5f520d1b626abd59ffec190b44df782d25443e2d7a84bc72fd7c1c2248e30d7876e2;
    5'b11100 : xpb = 1024'h8bd1b07cea753a95cac0105c8a63a50cee9fa249f4db60975136a59f257698a6e5334d1388d5ab26ea6f063f6987dfb3c59321157eac5fc248e3a64006b1e3b7d8f19518f9e75372f6da8011781ff0033d4a9abf0835e7bd3f627f5b888c8361366d4c3ea2847fb20206e156772b5c883c28b4d4ad1b44ffb46ddff7f772ac9a;
    5'b11101 : xpb = 1024'h51b6b97508ffc54124e98ab79bc6f60bbc569dcd715d0f4d7972e958824c2973231219dff33d4410cc2cc2285c18d88d56982f71c9173d5be7d77a20a8c8822cc04ba30931d73bf9d474716a4ef7295f960b7dfd16510da29c3cf4578af004de30b7a3e8d6e606ea644296ee7e596da2eb4a10424d782f530649fc08588a7be7;
    5'b11110 : xpb = 1024'h179bc26d278a4fec7f130512ad2a470a8a0d9950eddebe03a1af2d11df21ba3f60f0e6ac5da4dcfaadea7e114ea9d166e79d3dce13821af586cb4e014adf20a1a7a5b0f969c72480b20e62c325ce62bbeecc613b246c3387f91769538d53865b2b01fb930b478e22c67e4c8685877ebd9a6b6bafedd519a658261818b9a24b34;
    5'b11111 : xpb = 1024'h8e2e10bb08030f60a441f744cee7df5ac93a98053fd80d3147c82a20eef9f813a21830f19232f4732f0679412498db0adcbc7410809fc8dad65e614027c833c8034ef39851480a4ca24256be958160493b923e11bf0d867e0b7e704a49e1aa6a5453e566f0720de8af79e8fd8485b6019866a5ffde7d6129f071af2da39c80ec;
    endcase
end

endmodule

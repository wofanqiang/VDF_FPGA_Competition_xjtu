module compressor_array_236_2_1280_row
(
    input [235:0] col_in_0,
    input [235:0] col_in_1,
    input [235:0] col_in_2,
    input [235:0] col_in_3,
    input [235:0] col_in_4,
    input [235:0] col_in_5,
    input [235:0] col_in_6,
    input [235:0] col_in_7,
    input [235:0] col_in_8,
    input [235:0] col_in_9,
    input [235:0] col_in_10,
    input [235:0] col_in_11,
    input [235:0] col_in_12,
    input [235:0] col_in_13,
    input [235:0] col_in_14,
    input [235:0] col_in_15,
    input [235:0] col_in_16,
    input [235:0] col_in_17,
    input [235:0] col_in_18,
    input [235:0] col_in_19,
    input [235:0] col_in_20,
    input [235:0] col_in_21,
    input [235:0] col_in_22,
    input [235:0] col_in_23,
    input [235:0] col_in_24,
    input [235:0] col_in_25,
    input [235:0] col_in_26,
    input [235:0] col_in_27,
    input [235:0] col_in_28,
    input [235:0] col_in_29,
    input [235:0] col_in_30,
    input [235:0] col_in_31,
    input [235:0] col_in_32,
    input [235:0] col_in_33,
    input [235:0] col_in_34,
    input [235:0] col_in_35,
    input [235:0] col_in_36,
    input [235:0] col_in_37,
    input [235:0] col_in_38,
    input [235:0] col_in_39,
    input [235:0] col_in_40,
    input [235:0] col_in_41,
    input [235:0] col_in_42,
    input [235:0] col_in_43,
    input [235:0] col_in_44,
    input [235:0] col_in_45,
    input [235:0] col_in_46,
    input [235:0] col_in_47,
    input [235:0] col_in_48,
    input [235:0] col_in_49,
    input [235:0] col_in_50,
    input [235:0] col_in_51,
    input [235:0] col_in_52,
    input [235:0] col_in_53,
    input [235:0] col_in_54,
    input [235:0] col_in_55,
    input [235:0] col_in_56,
    input [235:0] col_in_57,
    input [235:0] col_in_58,
    input [235:0] col_in_59,
    input [235:0] col_in_60,
    input [235:0] col_in_61,
    input [235:0] col_in_62,
    input [235:0] col_in_63,
    input [235:0] col_in_64,
    input [235:0] col_in_65,
    input [235:0] col_in_66,
    input [235:0] col_in_67,
    input [235:0] col_in_68,
    input [235:0] col_in_69,
    input [235:0] col_in_70,
    input [235:0] col_in_71,
    input [235:0] col_in_72,
    input [235:0] col_in_73,
    input [235:0] col_in_74,
    input [235:0] col_in_75,
    input [235:0] col_in_76,
    input [235:0] col_in_77,
    input [235:0] col_in_78,
    input [235:0] col_in_79,
    input [235:0] col_in_80,
    input [235:0] col_in_81,
    input [235:0] col_in_82,
    input [235:0] col_in_83,
    input [235:0] col_in_84,
    input [235:0] col_in_85,
    input [235:0] col_in_86,
    input [235:0] col_in_87,
    input [235:0] col_in_88,
    input [235:0] col_in_89,
    input [235:0] col_in_90,
    input [235:0] col_in_91,
    input [235:0] col_in_92,
    input [235:0] col_in_93,
    input [235:0] col_in_94,
    input [235:0] col_in_95,
    input [235:0] col_in_96,
    input [235:0] col_in_97,
    input [235:0] col_in_98,
    input [235:0] col_in_99,
    input [235:0] col_in_100,
    input [235:0] col_in_101,
    input [235:0] col_in_102,
    input [235:0] col_in_103,
    input [235:0] col_in_104,
    input [235:0] col_in_105,
    input [235:0] col_in_106,
    input [235:0] col_in_107,
    input [235:0] col_in_108,
    input [235:0] col_in_109,
    input [235:0] col_in_110,
    input [235:0] col_in_111,
    input [235:0] col_in_112,
    input [235:0] col_in_113,
    input [235:0] col_in_114,
    input [235:0] col_in_115,
    input [235:0] col_in_116,
    input [235:0] col_in_117,
    input [235:0] col_in_118,
    input [235:0] col_in_119,
    input [235:0] col_in_120,
    input [235:0] col_in_121,
    input [235:0] col_in_122,
    input [235:0] col_in_123,
    input [235:0] col_in_124,
    input [235:0] col_in_125,
    input [235:0] col_in_126,
    input [235:0] col_in_127,
    input [235:0] col_in_128,
    input [235:0] col_in_129,
    input [235:0] col_in_130,
    input [235:0] col_in_131,
    input [235:0] col_in_132,
    input [235:0] col_in_133,
    input [235:0] col_in_134,
    input [235:0] col_in_135,
    input [235:0] col_in_136,
    input [235:0] col_in_137,
    input [235:0] col_in_138,
    input [235:0] col_in_139,
    input [235:0] col_in_140,
    input [235:0] col_in_141,
    input [235:0] col_in_142,
    input [235:0] col_in_143,
    input [235:0] col_in_144,
    input [235:0] col_in_145,
    input [235:0] col_in_146,
    input [235:0] col_in_147,
    input [235:0] col_in_148,
    input [235:0] col_in_149,
    input [235:0] col_in_150,
    input [235:0] col_in_151,
    input [235:0] col_in_152,
    input [235:0] col_in_153,
    input [235:0] col_in_154,
    input [235:0] col_in_155,
    input [235:0] col_in_156,
    input [235:0] col_in_157,
    input [235:0] col_in_158,
    input [235:0] col_in_159,
    input [235:0] col_in_160,
    input [235:0] col_in_161,
    input [235:0] col_in_162,
    input [235:0] col_in_163,
    input [235:0] col_in_164,
    input [235:0] col_in_165,
    input [235:0] col_in_166,
    input [235:0] col_in_167,
    input [235:0] col_in_168,
    input [235:0] col_in_169,
    input [235:0] col_in_170,
    input [235:0] col_in_171,
    input [235:0] col_in_172,
    input [235:0] col_in_173,
    input [235:0] col_in_174,
    input [235:0] col_in_175,
    input [235:0] col_in_176,
    input [235:0] col_in_177,
    input [235:0] col_in_178,
    input [235:0] col_in_179,
    input [235:0] col_in_180,
    input [235:0] col_in_181,
    input [235:0] col_in_182,
    input [235:0] col_in_183,
    input [235:0] col_in_184,
    input [235:0] col_in_185,
    input [235:0] col_in_186,
    input [235:0] col_in_187,
    input [235:0] col_in_188,
    input [235:0] col_in_189,
    input [235:0] col_in_190,
    input [235:0] col_in_191,
    input [235:0] col_in_192,
    input [235:0] col_in_193,
    input [235:0] col_in_194,
    input [235:0] col_in_195,
    input [235:0] col_in_196,
    input [235:0] col_in_197,
    input [235:0] col_in_198,
    input [235:0] col_in_199,
    input [235:0] col_in_200,
    input [235:0] col_in_201,
    input [235:0] col_in_202,
    input [235:0] col_in_203,
    input [235:0] col_in_204,
    input [235:0] col_in_205,
    input [235:0] col_in_206,
    input [235:0] col_in_207,
    input [235:0] col_in_208,
    input [235:0] col_in_209,
    input [235:0] col_in_210,
    input [235:0] col_in_211,
    input [235:0] col_in_212,
    input [235:0] col_in_213,
    input [235:0] col_in_214,
    input [235:0] col_in_215,
    input [235:0] col_in_216,
    input [235:0] col_in_217,
    input [235:0] col_in_218,
    input [235:0] col_in_219,
    input [235:0] col_in_220,
    input [235:0] col_in_221,
    input [235:0] col_in_222,
    input [235:0] col_in_223,
    input [235:0] col_in_224,
    input [235:0] col_in_225,
    input [235:0] col_in_226,
    input [235:0] col_in_227,
    input [235:0] col_in_228,
    input [235:0] col_in_229,
    input [235:0] col_in_230,
    input [235:0] col_in_231,
    input [235:0] col_in_232,
    input [235:0] col_in_233,
    input [235:0] col_in_234,
    input [235:0] col_in_235,
    input [235:0] col_in_236,
    input [235:0] col_in_237,
    input [235:0] col_in_238,
    input [235:0] col_in_239,
    input [235:0] col_in_240,
    input [235:0] col_in_241,
    input [235:0] col_in_242,
    input [235:0] col_in_243,
    input [235:0] col_in_244,
    input [235:0] col_in_245,
    input [235:0] col_in_246,
    input [235:0] col_in_247,
    input [235:0] col_in_248,
    input [235:0] col_in_249,
    input [235:0] col_in_250,
    input [235:0] col_in_251,
    input [235:0] col_in_252,
    input [235:0] col_in_253,
    input [235:0] col_in_254,
    input [235:0] col_in_255,
    input [235:0] col_in_256,
    input [235:0] col_in_257,
    input [235:0] col_in_258,
    input [235:0] col_in_259,
    input [235:0] col_in_260,
    input [235:0] col_in_261,
    input [235:0] col_in_262,
    input [235:0] col_in_263,
    input [235:0] col_in_264,
    input [235:0] col_in_265,
    input [235:0] col_in_266,
    input [235:0] col_in_267,
    input [235:0] col_in_268,
    input [235:0] col_in_269,
    input [235:0] col_in_270,
    input [235:0] col_in_271,
    input [235:0] col_in_272,
    input [235:0] col_in_273,
    input [235:0] col_in_274,
    input [235:0] col_in_275,
    input [235:0] col_in_276,
    input [235:0] col_in_277,
    input [235:0] col_in_278,
    input [235:0] col_in_279,
    input [235:0] col_in_280,
    input [235:0] col_in_281,
    input [235:0] col_in_282,
    input [235:0] col_in_283,
    input [235:0] col_in_284,
    input [235:0] col_in_285,
    input [235:0] col_in_286,
    input [235:0] col_in_287,
    input [235:0] col_in_288,
    input [235:0] col_in_289,
    input [235:0] col_in_290,
    input [235:0] col_in_291,
    input [235:0] col_in_292,
    input [235:0] col_in_293,
    input [235:0] col_in_294,
    input [235:0] col_in_295,
    input [235:0] col_in_296,
    input [235:0] col_in_297,
    input [235:0] col_in_298,
    input [235:0] col_in_299,
    input [235:0] col_in_300,
    input [235:0] col_in_301,
    input [235:0] col_in_302,
    input [235:0] col_in_303,
    input [235:0] col_in_304,
    input [235:0] col_in_305,
    input [235:0] col_in_306,
    input [235:0] col_in_307,
    input [235:0] col_in_308,
    input [235:0] col_in_309,
    input [235:0] col_in_310,
    input [235:0] col_in_311,
    input [235:0] col_in_312,
    input [235:0] col_in_313,
    input [235:0] col_in_314,
    input [235:0] col_in_315,
    input [235:0] col_in_316,
    input [235:0] col_in_317,
    input [235:0] col_in_318,
    input [235:0] col_in_319,
    input [235:0] col_in_320,
    input [235:0] col_in_321,
    input [235:0] col_in_322,
    input [235:0] col_in_323,
    input [235:0] col_in_324,
    input [235:0] col_in_325,
    input [235:0] col_in_326,
    input [235:0] col_in_327,
    input [235:0] col_in_328,
    input [235:0] col_in_329,
    input [235:0] col_in_330,
    input [235:0] col_in_331,
    input [235:0] col_in_332,
    input [235:0] col_in_333,
    input [235:0] col_in_334,
    input [235:0] col_in_335,
    input [235:0] col_in_336,
    input [235:0] col_in_337,
    input [235:0] col_in_338,
    input [235:0] col_in_339,
    input [235:0] col_in_340,
    input [235:0] col_in_341,
    input [235:0] col_in_342,
    input [235:0] col_in_343,
    input [235:0] col_in_344,
    input [235:0] col_in_345,
    input [235:0] col_in_346,
    input [235:0] col_in_347,
    input [235:0] col_in_348,
    input [235:0] col_in_349,
    input [235:0] col_in_350,
    input [235:0] col_in_351,
    input [235:0] col_in_352,
    input [235:0] col_in_353,
    input [235:0] col_in_354,
    input [235:0] col_in_355,
    input [235:0] col_in_356,
    input [235:0] col_in_357,
    input [235:0] col_in_358,
    input [235:0] col_in_359,
    input [235:0] col_in_360,
    input [235:0] col_in_361,
    input [235:0] col_in_362,
    input [235:0] col_in_363,
    input [235:0] col_in_364,
    input [235:0] col_in_365,
    input [235:0] col_in_366,
    input [235:0] col_in_367,
    input [235:0] col_in_368,
    input [235:0] col_in_369,
    input [235:0] col_in_370,
    input [235:0] col_in_371,
    input [235:0] col_in_372,
    input [235:0] col_in_373,
    input [235:0] col_in_374,
    input [235:0] col_in_375,
    input [235:0] col_in_376,
    input [235:0] col_in_377,
    input [235:0] col_in_378,
    input [235:0] col_in_379,
    input [235:0] col_in_380,
    input [235:0] col_in_381,
    input [235:0] col_in_382,
    input [235:0] col_in_383,
    input [235:0] col_in_384,
    input [235:0] col_in_385,
    input [235:0] col_in_386,
    input [235:0] col_in_387,
    input [235:0] col_in_388,
    input [235:0] col_in_389,
    input [235:0] col_in_390,
    input [235:0] col_in_391,
    input [235:0] col_in_392,
    input [235:0] col_in_393,
    input [235:0] col_in_394,
    input [235:0] col_in_395,
    input [235:0] col_in_396,
    input [235:0] col_in_397,
    input [235:0] col_in_398,
    input [235:0] col_in_399,
    input [235:0] col_in_400,
    input [235:0] col_in_401,
    input [235:0] col_in_402,
    input [235:0] col_in_403,
    input [235:0] col_in_404,
    input [235:0] col_in_405,
    input [235:0] col_in_406,
    input [235:0] col_in_407,
    input [235:0] col_in_408,
    input [235:0] col_in_409,
    input [235:0] col_in_410,
    input [235:0] col_in_411,
    input [235:0] col_in_412,
    input [235:0] col_in_413,
    input [235:0] col_in_414,
    input [235:0] col_in_415,
    input [235:0] col_in_416,
    input [235:0] col_in_417,
    input [235:0] col_in_418,
    input [235:0] col_in_419,
    input [235:0] col_in_420,
    input [235:0] col_in_421,
    input [235:0] col_in_422,
    input [235:0] col_in_423,
    input [235:0] col_in_424,
    input [235:0] col_in_425,
    input [235:0] col_in_426,
    input [235:0] col_in_427,
    input [235:0] col_in_428,
    input [235:0] col_in_429,
    input [235:0] col_in_430,
    input [235:0] col_in_431,
    input [235:0] col_in_432,
    input [235:0] col_in_433,
    input [235:0] col_in_434,
    input [235:0] col_in_435,
    input [235:0] col_in_436,
    input [235:0] col_in_437,
    input [235:0] col_in_438,
    input [235:0] col_in_439,
    input [235:0] col_in_440,
    input [235:0] col_in_441,
    input [235:0] col_in_442,
    input [235:0] col_in_443,
    input [235:0] col_in_444,
    input [235:0] col_in_445,
    input [235:0] col_in_446,
    input [235:0] col_in_447,
    input [235:0] col_in_448,
    input [235:0] col_in_449,
    input [235:0] col_in_450,
    input [235:0] col_in_451,
    input [235:0] col_in_452,
    input [235:0] col_in_453,
    input [235:0] col_in_454,
    input [235:0] col_in_455,
    input [235:0] col_in_456,
    input [235:0] col_in_457,
    input [235:0] col_in_458,
    input [235:0] col_in_459,
    input [235:0] col_in_460,
    input [235:0] col_in_461,
    input [235:0] col_in_462,
    input [235:0] col_in_463,
    input [235:0] col_in_464,
    input [235:0] col_in_465,
    input [235:0] col_in_466,
    input [235:0] col_in_467,
    input [235:0] col_in_468,
    input [235:0] col_in_469,
    input [235:0] col_in_470,
    input [235:0] col_in_471,
    input [235:0] col_in_472,
    input [235:0] col_in_473,
    input [235:0] col_in_474,
    input [235:0] col_in_475,
    input [235:0] col_in_476,
    input [235:0] col_in_477,
    input [235:0] col_in_478,
    input [235:0] col_in_479,
    input [235:0] col_in_480,
    input [235:0] col_in_481,
    input [235:0] col_in_482,
    input [235:0] col_in_483,
    input [235:0] col_in_484,
    input [235:0] col_in_485,
    input [235:0] col_in_486,
    input [235:0] col_in_487,
    input [235:0] col_in_488,
    input [235:0] col_in_489,
    input [235:0] col_in_490,
    input [235:0] col_in_491,
    input [235:0] col_in_492,
    input [235:0] col_in_493,
    input [235:0] col_in_494,
    input [235:0] col_in_495,
    input [235:0] col_in_496,
    input [235:0] col_in_497,
    input [235:0] col_in_498,
    input [235:0] col_in_499,
    input [235:0] col_in_500,
    input [235:0] col_in_501,
    input [235:0] col_in_502,
    input [235:0] col_in_503,
    input [235:0] col_in_504,
    input [235:0] col_in_505,
    input [235:0] col_in_506,
    input [235:0] col_in_507,
    input [235:0] col_in_508,
    input [235:0] col_in_509,
    input [235:0] col_in_510,
    input [235:0] col_in_511,
    input [235:0] col_in_512,
    input [235:0] col_in_513,
    input [235:0] col_in_514,
    input [235:0] col_in_515,
    input [235:0] col_in_516,
    input [235:0] col_in_517,
    input [235:0] col_in_518,
    input [235:0] col_in_519,
    input [235:0] col_in_520,
    input [235:0] col_in_521,
    input [235:0] col_in_522,
    input [235:0] col_in_523,
    input [235:0] col_in_524,
    input [235:0] col_in_525,
    input [235:0] col_in_526,
    input [235:0] col_in_527,
    input [235:0] col_in_528,
    input [235:0] col_in_529,
    input [235:0] col_in_530,
    input [235:0] col_in_531,
    input [235:0] col_in_532,
    input [235:0] col_in_533,
    input [235:0] col_in_534,
    input [235:0] col_in_535,
    input [235:0] col_in_536,
    input [235:0] col_in_537,
    input [235:0] col_in_538,
    input [235:0] col_in_539,
    input [235:0] col_in_540,
    input [235:0] col_in_541,
    input [235:0] col_in_542,
    input [235:0] col_in_543,
    input [235:0] col_in_544,
    input [235:0] col_in_545,
    input [235:0] col_in_546,
    input [235:0] col_in_547,
    input [235:0] col_in_548,
    input [235:0] col_in_549,
    input [235:0] col_in_550,
    input [235:0] col_in_551,
    input [235:0] col_in_552,
    input [235:0] col_in_553,
    input [235:0] col_in_554,
    input [235:0] col_in_555,
    input [235:0] col_in_556,
    input [235:0] col_in_557,
    input [235:0] col_in_558,
    input [235:0] col_in_559,
    input [235:0] col_in_560,
    input [235:0] col_in_561,
    input [235:0] col_in_562,
    input [235:0] col_in_563,
    input [235:0] col_in_564,
    input [235:0] col_in_565,
    input [235:0] col_in_566,
    input [235:0] col_in_567,
    input [235:0] col_in_568,
    input [235:0] col_in_569,
    input [235:0] col_in_570,
    input [235:0] col_in_571,
    input [235:0] col_in_572,
    input [235:0] col_in_573,
    input [235:0] col_in_574,
    input [235:0] col_in_575,
    input [235:0] col_in_576,
    input [235:0] col_in_577,
    input [235:0] col_in_578,
    input [235:0] col_in_579,
    input [235:0] col_in_580,
    input [235:0] col_in_581,
    input [235:0] col_in_582,
    input [235:0] col_in_583,
    input [235:0] col_in_584,
    input [235:0] col_in_585,
    input [235:0] col_in_586,
    input [235:0] col_in_587,
    input [235:0] col_in_588,
    input [235:0] col_in_589,
    input [235:0] col_in_590,
    input [235:0] col_in_591,
    input [235:0] col_in_592,
    input [235:0] col_in_593,
    input [235:0] col_in_594,
    input [235:0] col_in_595,
    input [235:0] col_in_596,
    input [235:0] col_in_597,
    input [235:0] col_in_598,
    input [235:0] col_in_599,
    input [235:0] col_in_600,
    input [235:0] col_in_601,
    input [235:0] col_in_602,
    input [235:0] col_in_603,
    input [235:0] col_in_604,
    input [235:0] col_in_605,
    input [235:0] col_in_606,
    input [235:0] col_in_607,
    input [235:0] col_in_608,
    input [235:0] col_in_609,
    input [235:0] col_in_610,
    input [235:0] col_in_611,
    input [235:0] col_in_612,
    input [235:0] col_in_613,
    input [235:0] col_in_614,
    input [235:0] col_in_615,
    input [235:0] col_in_616,
    input [235:0] col_in_617,
    input [235:0] col_in_618,
    input [235:0] col_in_619,
    input [235:0] col_in_620,
    input [235:0] col_in_621,
    input [235:0] col_in_622,
    input [235:0] col_in_623,
    input [235:0] col_in_624,
    input [235:0] col_in_625,
    input [235:0] col_in_626,
    input [235:0] col_in_627,
    input [235:0] col_in_628,
    input [235:0] col_in_629,
    input [235:0] col_in_630,
    input [235:0] col_in_631,
    input [235:0] col_in_632,
    input [235:0] col_in_633,
    input [235:0] col_in_634,
    input [235:0] col_in_635,
    input [235:0] col_in_636,
    input [235:0] col_in_637,
    input [235:0] col_in_638,
    input [235:0] col_in_639,
    input [235:0] col_in_640,
    input [235:0] col_in_641,
    input [235:0] col_in_642,
    input [235:0] col_in_643,
    input [235:0] col_in_644,
    input [235:0] col_in_645,
    input [235:0] col_in_646,
    input [235:0] col_in_647,
    input [235:0] col_in_648,
    input [235:0] col_in_649,
    input [235:0] col_in_650,
    input [235:0] col_in_651,
    input [235:0] col_in_652,
    input [235:0] col_in_653,
    input [235:0] col_in_654,
    input [235:0] col_in_655,
    input [235:0] col_in_656,
    input [235:0] col_in_657,
    input [235:0] col_in_658,
    input [235:0] col_in_659,
    input [235:0] col_in_660,
    input [235:0] col_in_661,
    input [235:0] col_in_662,
    input [235:0] col_in_663,
    input [235:0] col_in_664,
    input [235:0] col_in_665,
    input [235:0] col_in_666,
    input [235:0] col_in_667,
    input [235:0] col_in_668,
    input [235:0] col_in_669,
    input [235:0] col_in_670,
    input [235:0] col_in_671,
    input [235:0] col_in_672,
    input [235:0] col_in_673,
    input [235:0] col_in_674,
    input [235:0] col_in_675,
    input [235:0] col_in_676,
    input [235:0] col_in_677,
    input [235:0] col_in_678,
    input [235:0] col_in_679,
    input [235:0] col_in_680,
    input [235:0] col_in_681,
    input [235:0] col_in_682,
    input [235:0] col_in_683,
    input [235:0] col_in_684,
    input [235:0] col_in_685,
    input [235:0] col_in_686,
    input [235:0] col_in_687,
    input [235:0] col_in_688,
    input [235:0] col_in_689,
    input [235:0] col_in_690,
    input [235:0] col_in_691,
    input [235:0] col_in_692,
    input [235:0] col_in_693,
    input [235:0] col_in_694,
    input [235:0] col_in_695,
    input [235:0] col_in_696,
    input [235:0] col_in_697,
    input [235:0] col_in_698,
    input [235:0] col_in_699,
    input [235:0] col_in_700,
    input [235:0] col_in_701,
    input [235:0] col_in_702,
    input [235:0] col_in_703,
    input [235:0] col_in_704,
    input [235:0] col_in_705,
    input [235:0] col_in_706,
    input [235:0] col_in_707,
    input [235:0] col_in_708,
    input [235:0] col_in_709,
    input [235:0] col_in_710,
    input [235:0] col_in_711,
    input [235:0] col_in_712,
    input [235:0] col_in_713,
    input [235:0] col_in_714,
    input [235:0] col_in_715,
    input [235:0] col_in_716,
    input [235:0] col_in_717,
    input [235:0] col_in_718,
    input [235:0] col_in_719,
    input [235:0] col_in_720,
    input [235:0] col_in_721,
    input [235:0] col_in_722,
    input [235:0] col_in_723,
    input [235:0] col_in_724,
    input [235:0] col_in_725,
    input [235:0] col_in_726,
    input [235:0] col_in_727,
    input [235:0] col_in_728,
    input [235:0] col_in_729,
    input [235:0] col_in_730,
    input [235:0] col_in_731,
    input [235:0] col_in_732,
    input [235:0] col_in_733,
    input [235:0] col_in_734,
    input [235:0] col_in_735,
    input [235:0] col_in_736,
    input [235:0] col_in_737,
    input [235:0] col_in_738,
    input [235:0] col_in_739,
    input [235:0] col_in_740,
    input [235:0] col_in_741,
    input [235:0] col_in_742,
    input [235:0] col_in_743,
    input [235:0] col_in_744,
    input [235:0] col_in_745,
    input [235:0] col_in_746,
    input [235:0] col_in_747,
    input [235:0] col_in_748,
    input [235:0] col_in_749,
    input [235:0] col_in_750,
    input [235:0] col_in_751,
    input [235:0] col_in_752,
    input [235:0] col_in_753,
    input [235:0] col_in_754,
    input [235:0] col_in_755,
    input [235:0] col_in_756,
    input [235:0] col_in_757,
    input [235:0] col_in_758,
    input [235:0] col_in_759,
    input [235:0] col_in_760,
    input [235:0] col_in_761,
    input [235:0] col_in_762,
    input [235:0] col_in_763,
    input [235:0] col_in_764,
    input [235:0] col_in_765,
    input [235:0] col_in_766,
    input [235:0] col_in_767,
    input [235:0] col_in_768,
    input [235:0] col_in_769,
    input [235:0] col_in_770,
    input [235:0] col_in_771,
    input [235:0] col_in_772,
    input [235:0] col_in_773,
    input [235:0] col_in_774,
    input [235:0] col_in_775,
    input [235:0] col_in_776,
    input [235:0] col_in_777,
    input [235:0] col_in_778,
    input [235:0] col_in_779,
    input [235:0] col_in_780,
    input [235:0] col_in_781,
    input [235:0] col_in_782,
    input [235:0] col_in_783,
    input [235:0] col_in_784,
    input [235:0] col_in_785,
    input [235:0] col_in_786,
    input [235:0] col_in_787,
    input [235:0] col_in_788,
    input [235:0] col_in_789,
    input [235:0] col_in_790,
    input [235:0] col_in_791,
    input [235:0] col_in_792,
    input [235:0] col_in_793,
    input [235:0] col_in_794,
    input [235:0] col_in_795,
    input [235:0] col_in_796,
    input [235:0] col_in_797,
    input [235:0] col_in_798,
    input [235:0] col_in_799,
    input [235:0] col_in_800,
    input [235:0] col_in_801,
    input [235:0] col_in_802,
    input [235:0] col_in_803,
    input [235:0] col_in_804,
    input [235:0] col_in_805,
    input [235:0] col_in_806,
    input [235:0] col_in_807,
    input [235:0] col_in_808,
    input [235:0] col_in_809,
    input [235:0] col_in_810,
    input [235:0] col_in_811,
    input [235:0] col_in_812,
    input [235:0] col_in_813,
    input [235:0] col_in_814,
    input [235:0] col_in_815,
    input [235:0] col_in_816,
    input [235:0] col_in_817,
    input [235:0] col_in_818,
    input [235:0] col_in_819,
    input [235:0] col_in_820,
    input [235:0] col_in_821,
    input [235:0] col_in_822,
    input [235:0] col_in_823,
    input [235:0] col_in_824,
    input [235:0] col_in_825,
    input [235:0] col_in_826,
    input [235:0] col_in_827,
    input [235:0] col_in_828,
    input [235:0] col_in_829,
    input [235:0] col_in_830,
    input [235:0] col_in_831,
    input [235:0] col_in_832,
    input [235:0] col_in_833,
    input [235:0] col_in_834,
    input [235:0] col_in_835,
    input [235:0] col_in_836,
    input [235:0] col_in_837,
    input [235:0] col_in_838,
    input [235:0] col_in_839,
    input [235:0] col_in_840,
    input [235:0] col_in_841,
    input [235:0] col_in_842,
    input [235:0] col_in_843,
    input [235:0] col_in_844,
    input [235:0] col_in_845,
    input [235:0] col_in_846,
    input [235:0] col_in_847,
    input [235:0] col_in_848,
    input [235:0] col_in_849,
    input [235:0] col_in_850,
    input [235:0] col_in_851,
    input [235:0] col_in_852,
    input [235:0] col_in_853,
    input [235:0] col_in_854,
    input [235:0] col_in_855,
    input [235:0] col_in_856,
    input [235:0] col_in_857,
    input [235:0] col_in_858,
    input [235:0] col_in_859,
    input [235:0] col_in_860,
    input [235:0] col_in_861,
    input [235:0] col_in_862,
    input [235:0] col_in_863,
    input [235:0] col_in_864,
    input [235:0] col_in_865,
    input [235:0] col_in_866,
    input [235:0] col_in_867,
    input [235:0] col_in_868,
    input [235:0] col_in_869,
    input [235:0] col_in_870,
    input [235:0] col_in_871,
    input [235:0] col_in_872,
    input [235:0] col_in_873,
    input [235:0] col_in_874,
    input [235:0] col_in_875,
    input [235:0] col_in_876,
    input [235:0] col_in_877,
    input [235:0] col_in_878,
    input [235:0] col_in_879,
    input [235:0] col_in_880,
    input [235:0] col_in_881,
    input [235:0] col_in_882,
    input [235:0] col_in_883,
    input [235:0] col_in_884,
    input [235:0] col_in_885,
    input [235:0] col_in_886,
    input [235:0] col_in_887,
    input [235:0] col_in_888,
    input [235:0] col_in_889,
    input [235:0] col_in_890,
    input [235:0] col_in_891,
    input [235:0] col_in_892,
    input [235:0] col_in_893,
    input [235:0] col_in_894,
    input [235:0] col_in_895,
    input [235:0] col_in_896,
    input [235:0] col_in_897,
    input [235:0] col_in_898,
    input [235:0] col_in_899,
    input [235:0] col_in_900,
    input [235:0] col_in_901,
    input [235:0] col_in_902,
    input [235:0] col_in_903,
    input [235:0] col_in_904,
    input [235:0] col_in_905,
    input [235:0] col_in_906,
    input [235:0] col_in_907,
    input [235:0] col_in_908,
    input [235:0] col_in_909,
    input [235:0] col_in_910,
    input [235:0] col_in_911,
    input [235:0] col_in_912,
    input [235:0] col_in_913,
    input [235:0] col_in_914,
    input [235:0] col_in_915,
    input [235:0] col_in_916,
    input [235:0] col_in_917,
    input [235:0] col_in_918,
    input [235:0] col_in_919,
    input [235:0] col_in_920,
    input [235:0] col_in_921,
    input [235:0] col_in_922,
    input [235:0] col_in_923,
    input [235:0] col_in_924,
    input [235:0] col_in_925,
    input [235:0] col_in_926,
    input [235:0] col_in_927,
    input [235:0] col_in_928,
    input [235:0] col_in_929,
    input [235:0] col_in_930,
    input [235:0] col_in_931,
    input [235:0] col_in_932,
    input [235:0] col_in_933,
    input [235:0] col_in_934,
    input [235:0] col_in_935,
    input [235:0] col_in_936,
    input [235:0] col_in_937,
    input [235:0] col_in_938,
    input [235:0] col_in_939,
    input [235:0] col_in_940,
    input [235:0] col_in_941,
    input [235:0] col_in_942,
    input [235:0] col_in_943,
    input [235:0] col_in_944,
    input [235:0] col_in_945,
    input [235:0] col_in_946,
    input [235:0] col_in_947,
    input [235:0] col_in_948,
    input [235:0] col_in_949,
    input [235:0] col_in_950,
    input [235:0] col_in_951,
    input [235:0] col_in_952,
    input [235:0] col_in_953,
    input [235:0] col_in_954,
    input [235:0] col_in_955,
    input [235:0] col_in_956,
    input [235:0] col_in_957,
    input [235:0] col_in_958,
    input [235:0] col_in_959,
    input [235:0] col_in_960,
    input [235:0] col_in_961,
    input [235:0] col_in_962,
    input [235:0] col_in_963,
    input [235:0] col_in_964,
    input [235:0] col_in_965,
    input [235:0] col_in_966,
    input [235:0] col_in_967,
    input [235:0] col_in_968,
    input [235:0] col_in_969,
    input [235:0] col_in_970,
    input [235:0] col_in_971,
    input [235:0] col_in_972,
    input [235:0] col_in_973,
    input [235:0] col_in_974,
    input [235:0] col_in_975,
    input [235:0] col_in_976,
    input [235:0] col_in_977,
    input [235:0] col_in_978,
    input [235:0] col_in_979,
    input [235:0] col_in_980,
    input [235:0] col_in_981,
    input [235:0] col_in_982,
    input [235:0] col_in_983,
    input [235:0] col_in_984,
    input [235:0] col_in_985,
    input [235:0] col_in_986,
    input [235:0] col_in_987,
    input [235:0] col_in_988,
    input [235:0] col_in_989,
    input [235:0] col_in_990,
    input [235:0] col_in_991,
    input [235:0] col_in_992,
    input [235:0] col_in_993,
    input [235:0] col_in_994,
    input [235:0] col_in_995,
    input [235:0] col_in_996,
    input [235:0] col_in_997,
    input [235:0] col_in_998,
    input [235:0] col_in_999,
    input [235:0] col_in_1000,
    input [235:0] col_in_1001,
    input [235:0] col_in_1002,
    input [235:0] col_in_1003,
    input [235:0] col_in_1004,
    input [235:0] col_in_1005,
    input [235:0] col_in_1006,
    input [235:0] col_in_1007,
    input [235:0] col_in_1008,
    input [235:0] col_in_1009,
    input [235:0] col_in_1010,
    input [235:0] col_in_1011,
    input [235:0] col_in_1012,
    input [235:0] col_in_1013,
    input [235:0] col_in_1014,
    input [235:0] col_in_1015,
    input [235:0] col_in_1016,
    input [235:0] col_in_1017,
    input [235:0] col_in_1018,
    input [235:0] col_in_1019,
    input [235:0] col_in_1020,
    input [235:0] col_in_1021,
    input [235:0] col_in_1022,
    input [235:0] col_in_1023,
    input [235:0] col_in_1024,
    input [235:0] col_in_1025,
    input [235:0] col_in_1026,
    input [235:0] col_in_1027,
    input [235:0] col_in_1028,
    input [235:0] col_in_1029,
    input [235:0] col_in_1030,
    input [235:0] col_in_1031,
    input [235:0] col_in_1032,
    input [235:0] col_in_1033,
    input [235:0] col_in_1034,
    input [235:0] col_in_1035,
    input [235:0] col_in_1036,
    input [235:0] col_in_1037,
    input [235:0] col_in_1038,
    input [235:0] col_in_1039,
    input [235:0] col_in_1040,
    input [235:0] col_in_1041,
    input [235:0] col_in_1042,
    input [235:0] col_in_1043,
    input [235:0] col_in_1044,
    input [235:0] col_in_1045,
    input [235:0] col_in_1046,
    input [235:0] col_in_1047,
    input [235:0] col_in_1048,
    input [235:0] col_in_1049,
    input [235:0] col_in_1050,
    input [235:0] col_in_1051,
    input [235:0] col_in_1052,
    input [235:0] col_in_1053,
    input [235:0] col_in_1054,
    input [235:0] col_in_1055,
    input [235:0] col_in_1056,
    input [235:0] col_in_1057,
    input [235:0] col_in_1058,
    input [235:0] col_in_1059,
    input [235:0] col_in_1060,
    input [235:0] col_in_1061,
    input [235:0] col_in_1062,
    input [235:0] col_in_1063,
    input [235:0] col_in_1064,
    input [235:0] col_in_1065,
    input [235:0] col_in_1066,
    input [235:0] col_in_1067,
    input [235:0] col_in_1068,
    input [235:0] col_in_1069,
    input [235:0] col_in_1070,
    input [235:0] col_in_1071,
    input [235:0] col_in_1072,
    input [235:0] col_in_1073,
    input [235:0] col_in_1074,
    input [235:0] col_in_1075,
    input [235:0] col_in_1076,
    input [235:0] col_in_1077,
    input [235:0] col_in_1078,
    input [235:0] col_in_1079,
    input [235:0] col_in_1080,
    input [235:0] col_in_1081,
    input [235:0] col_in_1082,
    input [235:0] col_in_1083,
    input [235:0] col_in_1084,
    input [235:0] col_in_1085,
    input [235:0] col_in_1086,
    input [235:0] col_in_1087,
    input [235:0] col_in_1088,
    input [235:0] col_in_1089,
    input [235:0] col_in_1090,
    input [235:0] col_in_1091,
    input [235:0] col_in_1092,
    input [235:0] col_in_1093,
    input [235:0] col_in_1094,
    input [235:0] col_in_1095,
    input [235:0] col_in_1096,
    input [235:0] col_in_1097,
    input [235:0] col_in_1098,
    input [235:0] col_in_1099,
    input [235:0] col_in_1100,
    input [235:0] col_in_1101,
    input [235:0] col_in_1102,
    input [235:0] col_in_1103,
    input [235:0] col_in_1104,
    input [235:0] col_in_1105,
    input [235:0] col_in_1106,
    input [235:0] col_in_1107,
    input [235:0] col_in_1108,
    input [235:0] col_in_1109,
    input [235:0] col_in_1110,
    input [235:0] col_in_1111,
    input [235:0] col_in_1112,
    input [235:0] col_in_1113,
    input [235:0] col_in_1114,
    input [235:0] col_in_1115,
    input [235:0] col_in_1116,
    input [235:0] col_in_1117,
    input [235:0] col_in_1118,
    input [235:0] col_in_1119,
    input [235:0] col_in_1120,
    input [235:0] col_in_1121,
    input [235:0] col_in_1122,
    input [235:0] col_in_1123,
    input [235:0] col_in_1124,
    input [235:0] col_in_1125,
    input [235:0] col_in_1126,
    input [235:0] col_in_1127,
    input [235:0] col_in_1128,
    input [235:0] col_in_1129,
    input [235:0] col_in_1130,
    input [235:0] col_in_1131,
    input [235:0] col_in_1132,
    input [235:0] col_in_1133,
    input [235:0] col_in_1134,
    input [235:0] col_in_1135,
    input [235:0] col_in_1136,
    input [235:0] col_in_1137,
    input [235:0] col_in_1138,
    input [235:0] col_in_1139,
    input [235:0] col_in_1140,
    input [235:0] col_in_1141,
    input [235:0] col_in_1142,
    input [235:0] col_in_1143,
    input [235:0] col_in_1144,
    input [235:0] col_in_1145,
    input [235:0] col_in_1146,
    input [235:0] col_in_1147,
    input [235:0] col_in_1148,
    input [235:0] col_in_1149,
    input [235:0] col_in_1150,
    input [235:0] col_in_1151,
    input [235:0] col_in_1152,
    input [235:0] col_in_1153,
    input [235:0] col_in_1154,
    input [235:0] col_in_1155,
    input [235:0] col_in_1156,
    input [235:0] col_in_1157,
    input [235:0] col_in_1158,
    input [235:0] col_in_1159,
    input [235:0] col_in_1160,
    input [235:0] col_in_1161,
    input [235:0] col_in_1162,
    input [235:0] col_in_1163,
    input [235:0] col_in_1164,
    input [235:0] col_in_1165,
    input [235:0] col_in_1166,
    input [235:0] col_in_1167,
    input [235:0] col_in_1168,
    input [235:0] col_in_1169,
    input [235:0] col_in_1170,
    input [235:0] col_in_1171,
    input [235:0] col_in_1172,
    input [235:0] col_in_1173,
    input [235:0] col_in_1174,
    input [235:0] col_in_1175,
    input [235:0] col_in_1176,
    input [235:0] col_in_1177,
    input [235:0] col_in_1178,
    input [235:0] col_in_1179,
    input [235:0] col_in_1180,
    input [235:0] col_in_1181,
    input [235:0] col_in_1182,
    input [235:0] col_in_1183,
    input [235:0] col_in_1184,
    input [235:0] col_in_1185,
    input [235:0] col_in_1186,
    input [235:0] col_in_1187,
    input [235:0] col_in_1188,
    input [235:0] col_in_1189,
    input [235:0] col_in_1190,
    input [235:0] col_in_1191,
    input [235:0] col_in_1192,
    input [235:0] col_in_1193,
    input [235:0] col_in_1194,
    input [235:0] col_in_1195,
    input [235:0] col_in_1196,
    input [235:0] col_in_1197,
    input [235:0] col_in_1198,
    input [235:0] col_in_1199,
    input [235:0] col_in_1200,
    input [235:0] col_in_1201,
    input [235:0] col_in_1202,
    input [235:0] col_in_1203,
    input [235:0] col_in_1204,
    input [235:0] col_in_1205,
    input [235:0] col_in_1206,
    input [235:0] col_in_1207,
    input [235:0] col_in_1208,
    input [235:0] col_in_1209,
    input [235:0] col_in_1210,
    input [235:0] col_in_1211,
    input [235:0] col_in_1212,
    input [235:0] col_in_1213,
    input [235:0] col_in_1214,
    input [235:0] col_in_1215,
    input [235:0] col_in_1216,
    input [235:0] col_in_1217,
    input [235:0] col_in_1218,
    input [235:0] col_in_1219,
    input [235:0] col_in_1220,
    input [235:0] col_in_1221,
    input [235:0] col_in_1222,
    input [235:0] col_in_1223,
    input [235:0] col_in_1224,
    input [235:0] col_in_1225,
    input [235:0] col_in_1226,
    input [235:0] col_in_1227,
    input [235:0] col_in_1228,
    input [235:0] col_in_1229,
    input [235:0] col_in_1230,
    input [235:0] col_in_1231,
    input [235:0] col_in_1232,
    input [235:0] col_in_1233,
    input [235:0] col_in_1234,
    input [235:0] col_in_1235,
    input [235:0] col_in_1236,
    input [235:0] col_in_1237,
    input [235:0] col_in_1238,
    input [235:0] col_in_1239,
    input [235:0] col_in_1240,
    input [235:0] col_in_1241,
    input [235:0] col_in_1242,
    input [235:0] col_in_1243,
    input [235:0] col_in_1244,
    input [235:0] col_in_1245,
    input [235:0] col_in_1246,
    input [235:0] col_in_1247,
    input [235:0] col_in_1248,
    input [235:0] col_in_1249,
    input [235:0] col_in_1250,
    input [235:0] col_in_1251,
    input [235:0] col_in_1252,
    input [235:0] col_in_1253,
    input [235:0] col_in_1254,
    input [235:0] col_in_1255,
    input [235:0] col_in_1256,
    input [235:0] col_in_1257,
    input [235:0] col_in_1258,
    input [235:0] col_in_1259,
    input [235:0] col_in_1260,
    input [235:0] col_in_1261,
    input [235:0] col_in_1262,
    input [235:0] col_in_1263,
    input [235:0] col_in_1264,
    input [235:0] col_in_1265,
    input [235:0] col_in_1266,
    input [235:0] col_in_1267,
    input [235:0] col_in_1268,
    input [235:0] col_in_1269,
    input [235:0] col_in_1270,
    input [235:0] col_in_1271,
    input [235:0] col_in_1272,
    input [235:0] col_in_1273,
    input [235:0] col_in_1274,
    input [235:0] col_in_1275,
    input [235:0] col_in_1276,
    input [235:0] col_in_1277,
    input [235:0] col_in_1278,
    input [235:0] col_in_1279,


    output [1287:0] row_out_0,
    output [1287:0] row_out_1
);


wire [1:0] u_col_out_0;
wire [1:0] u_col_out_1;
wire [1:0] u_col_out_2;
wire [1:0] u_col_out_3;
wire [1:0] u_col_out_4;
wire [1:0] u_col_out_5;
wire [1:0] u_col_out_6;
wire [1:0] u_col_out_7;
wire [1:0] u_col_out_8;
wire [1:0] u_col_out_9;
wire [1:0] u_col_out_10;
wire [1:0] u_col_out_11;
wire [1:0] u_col_out_12;
wire [1:0] u_col_out_13;
wire [1:0] u_col_out_14;
wire [1:0] u_col_out_15;
wire [1:0] u_col_out_16;
wire [1:0] u_col_out_17;
wire [1:0] u_col_out_18;
wire [1:0] u_col_out_19;
wire [1:0] u_col_out_20;
wire [1:0] u_col_out_21;
wire [1:0] u_col_out_22;
wire [1:0] u_col_out_23;
wire [1:0] u_col_out_24;
wire [1:0] u_col_out_25;
wire [1:0] u_col_out_26;
wire [1:0] u_col_out_27;
wire [1:0] u_col_out_28;
wire [1:0] u_col_out_29;
wire [1:0] u_col_out_30;
wire [1:0] u_col_out_31;
wire [1:0] u_col_out_32;
wire [1:0] u_col_out_33;
wire [1:0] u_col_out_34;
wire [1:0] u_col_out_35;
wire [1:0] u_col_out_36;
wire [1:0] u_col_out_37;
wire [1:0] u_col_out_38;
wire [1:0] u_col_out_39;
wire [1:0] u_col_out_40;
wire [1:0] u_col_out_41;
wire [1:0] u_col_out_42;
wire [1:0] u_col_out_43;
wire [1:0] u_col_out_44;
wire [1:0] u_col_out_45;
wire [1:0] u_col_out_46;
wire [1:0] u_col_out_47;
wire [1:0] u_col_out_48;
wire [1:0] u_col_out_49;
wire [1:0] u_col_out_50;
wire [1:0] u_col_out_51;
wire [1:0] u_col_out_52;
wire [1:0] u_col_out_53;
wire [1:0] u_col_out_54;
wire [1:0] u_col_out_55;
wire [1:0] u_col_out_56;
wire [1:0] u_col_out_57;
wire [1:0] u_col_out_58;
wire [1:0] u_col_out_59;
wire [1:0] u_col_out_60;
wire [1:0] u_col_out_61;
wire [1:0] u_col_out_62;
wire [1:0] u_col_out_63;
wire [1:0] u_col_out_64;
wire [1:0] u_col_out_65;
wire [1:0] u_col_out_66;
wire [1:0] u_col_out_67;
wire [1:0] u_col_out_68;
wire [1:0] u_col_out_69;
wire [1:0] u_col_out_70;
wire [1:0] u_col_out_71;
wire [1:0] u_col_out_72;
wire [1:0] u_col_out_73;
wire [1:0] u_col_out_74;
wire [1:0] u_col_out_75;
wire [1:0] u_col_out_76;
wire [1:0] u_col_out_77;
wire [1:0] u_col_out_78;
wire [1:0] u_col_out_79;
wire [1:0] u_col_out_80;
wire [1:0] u_col_out_81;
wire [1:0] u_col_out_82;
wire [1:0] u_col_out_83;
wire [1:0] u_col_out_84;
wire [1:0] u_col_out_85;
wire [1:0] u_col_out_86;
wire [1:0] u_col_out_87;
wire [1:0] u_col_out_88;
wire [1:0] u_col_out_89;
wire [1:0] u_col_out_90;
wire [1:0] u_col_out_91;
wire [1:0] u_col_out_92;
wire [1:0] u_col_out_93;
wire [1:0] u_col_out_94;
wire [1:0] u_col_out_95;
wire [1:0] u_col_out_96;
wire [1:0] u_col_out_97;
wire [1:0] u_col_out_98;
wire [1:0] u_col_out_99;
wire [1:0] u_col_out_100;
wire [1:0] u_col_out_101;
wire [1:0] u_col_out_102;
wire [1:0] u_col_out_103;
wire [1:0] u_col_out_104;
wire [1:0] u_col_out_105;
wire [1:0] u_col_out_106;
wire [1:0] u_col_out_107;
wire [1:0] u_col_out_108;
wire [1:0] u_col_out_109;
wire [1:0] u_col_out_110;
wire [1:0] u_col_out_111;
wire [1:0] u_col_out_112;
wire [1:0] u_col_out_113;
wire [1:0] u_col_out_114;
wire [1:0] u_col_out_115;
wire [1:0] u_col_out_116;
wire [1:0] u_col_out_117;
wire [1:0] u_col_out_118;
wire [1:0] u_col_out_119;
wire [1:0] u_col_out_120;
wire [1:0] u_col_out_121;
wire [1:0] u_col_out_122;
wire [1:0] u_col_out_123;
wire [1:0] u_col_out_124;
wire [1:0] u_col_out_125;
wire [1:0] u_col_out_126;
wire [1:0] u_col_out_127;
wire [1:0] u_col_out_128;
wire [1:0] u_col_out_129;
wire [1:0] u_col_out_130;
wire [1:0] u_col_out_131;
wire [1:0] u_col_out_132;
wire [1:0] u_col_out_133;
wire [1:0] u_col_out_134;
wire [1:0] u_col_out_135;
wire [1:0] u_col_out_136;
wire [1:0] u_col_out_137;
wire [1:0] u_col_out_138;
wire [1:0] u_col_out_139;
wire [1:0] u_col_out_140;
wire [1:0] u_col_out_141;
wire [1:0] u_col_out_142;
wire [1:0] u_col_out_143;
wire [1:0] u_col_out_144;
wire [1:0] u_col_out_145;
wire [1:0] u_col_out_146;
wire [1:0] u_col_out_147;
wire [1:0] u_col_out_148;
wire [1:0] u_col_out_149;
wire [1:0] u_col_out_150;
wire [1:0] u_col_out_151;
wire [1:0] u_col_out_152;
wire [1:0] u_col_out_153;
wire [1:0] u_col_out_154;
wire [1:0] u_col_out_155;
wire [1:0] u_col_out_156;
wire [1:0] u_col_out_157;
wire [1:0] u_col_out_158;
wire [1:0] u_col_out_159;
wire [1:0] u_col_out_160;
wire [1:0] u_col_out_161;
wire [1:0] u_col_out_162;
wire [1:0] u_col_out_163;
wire [1:0] u_col_out_164;
wire [1:0] u_col_out_165;
wire [1:0] u_col_out_166;
wire [1:0] u_col_out_167;
wire [1:0] u_col_out_168;
wire [1:0] u_col_out_169;
wire [1:0] u_col_out_170;
wire [1:0] u_col_out_171;
wire [1:0] u_col_out_172;
wire [1:0] u_col_out_173;
wire [1:0] u_col_out_174;
wire [1:0] u_col_out_175;
wire [1:0] u_col_out_176;
wire [1:0] u_col_out_177;
wire [1:0] u_col_out_178;
wire [1:0] u_col_out_179;
wire [1:0] u_col_out_180;
wire [1:0] u_col_out_181;
wire [1:0] u_col_out_182;
wire [1:0] u_col_out_183;
wire [1:0] u_col_out_184;
wire [1:0] u_col_out_185;
wire [1:0] u_col_out_186;
wire [1:0] u_col_out_187;
wire [1:0] u_col_out_188;
wire [1:0] u_col_out_189;
wire [1:0] u_col_out_190;
wire [1:0] u_col_out_191;
wire [1:0] u_col_out_192;
wire [1:0] u_col_out_193;
wire [1:0] u_col_out_194;
wire [1:0] u_col_out_195;
wire [1:0] u_col_out_196;
wire [1:0] u_col_out_197;
wire [1:0] u_col_out_198;
wire [1:0] u_col_out_199;
wire [1:0] u_col_out_200;
wire [1:0] u_col_out_201;
wire [1:0] u_col_out_202;
wire [1:0] u_col_out_203;
wire [1:0] u_col_out_204;
wire [1:0] u_col_out_205;
wire [1:0] u_col_out_206;
wire [1:0] u_col_out_207;
wire [1:0] u_col_out_208;
wire [1:0] u_col_out_209;
wire [1:0] u_col_out_210;
wire [1:0] u_col_out_211;
wire [1:0] u_col_out_212;
wire [1:0] u_col_out_213;
wire [1:0] u_col_out_214;
wire [1:0] u_col_out_215;
wire [1:0] u_col_out_216;
wire [1:0] u_col_out_217;
wire [1:0] u_col_out_218;
wire [1:0] u_col_out_219;
wire [1:0] u_col_out_220;
wire [1:0] u_col_out_221;
wire [1:0] u_col_out_222;
wire [1:0] u_col_out_223;
wire [1:0] u_col_out_224;
wire [1:0] u_col_out_225;
wire [1:0] u_col_out_226;
wire [1:0] u_col_out_227;
wire [1:0] u_col_out_228;
wire [1:0] u_col_out_229;
wire [1:0] u_col_out_230;
wire [1:0] u_col_out_231;
wire [1:0] u_col_out_232;
wire [1:0] u_col_out_233;
wire [1:0] u_col_out_234;
wire [1:0] u_col_out_235;
wire [1:0] u_col_out_236;
wire [1:0] u_col_out_237;
wire [1:0] u_col_out_238;
wire [1:0] u_col_out_239;
wire [1:0] u_col_out_240;
wire [1:0] u_col_out_241;
wire [1:0] u_col_out_242;
wire [1:0] u_col_out_243;
wire [1:0] u_col_out_244;
wire [1:0] u_col_out_245;
wire [1:0] u_col_out_246;
wire [1:0] u_col_out_247;
wire [1:0] u_col_out_248;
wire [1:0] u_col_out_249;
wire [1:0] u_col_out_250;
wire [1:0] u_col_out_251;
wire [1:0] u_col_out_252;
wire [1:0] u_col_out_253;
wire [1:0] u_col_out_254;
wire [1:0] u_col_out_255;
wire [1:0] u_col_out_256;
wire [1:0] u_col_out_257;
wire [1:0] u_col_out_258;
wire [1:0] u_col_out_259;
wire [1:0] u_col_out_260;
wire [1:0] u_col_out_261;
wire [1:0] u_col_out_262;
wire [1:0] u_col_out_263;
wire [1:0] u_col_out_264;
wire [1:0] u_col_out_265;
wire [1:0] u_col_out_266;
wire [1:0] u_col_out_267;
wire [1:0] u_col_out_268;
wire [1:0] u_col_out_269;
wire [1:0] u_col_out_270;
wire [1:0] u_col_out_271;
wire [1:0] u_col_out_272;
wire [1:0] u_col_out_273;
wire [1:0] u_col_out_274;
wire [1:0] u_col_out_275;
wire [1:0] u_col_out_276;
wire [1:0] u_col_out_277;
wire [1:0] u_col_out_278;
wire [1:0] u_col_out_279;
wire [1:0] u_col_out_280;
wire [1:0] u_col_out_281;
wire [1:0] u_col_out_282;
wire [1:0] u_col_out_283;
wire [1:0] u_col_out_284;
wire [1:0] u_col_out_285;
wire [1:0] u_col_out_286;
wire [1:0] u_col_out_287;
wire [1:0] u_col_out_288;
wire [1:0] u_col_out_289;
wire [1:0] u_col_out_290;
wire [1:0] u_col_out_291;
wire [1:0] u_col_out_292;
wire [1:0] u_col_out_293;
wire [1:0] u_col_out_294;
wire [1:0] u_col_out_295;
wire [1:0] u_col_out_296;
wire [1:0] u_col_out_297;
wire [1:0] u_col_out_298;
wire [1:0] u_col_out_299;
wire [1:0] u_col_out_300;
wire [1:0] u_col_out_301;
wire [1:0] u_col_out_302;
wire [1:0] u_col_out_303;
wire [1:0] u_col_out_304;
wire [1:0] u_col_out_305;
wire [1:0] u_col_out_306;
wire [1:0] u_col_out_307;
wire [1:0] u_col_out_308;
wire [1:0] u_col_out_309;
wire [1:0] u_col_out_310;
wire [1:0] u_col_out_311;
wire [1:0] u_col_out_312;
wire [1:0] u_col_out_313;
wire [1:0] u_col_out_314;
wire [1:0] u_col_out_315;
wire [1:0] u_col_out_316;
wire [1:0] u_col_out_317;
wire [1:0] u_col_out_318;
wire [1:0] u_col_out_319;
wire [1:0] u_col_out_320;
wire [1:0] u_col_out_321;
wire [1:0] u_col_out_322;
wire [1:0] u_col_out_323;
wire [1:0] u_col_out_324;
wire [1:0] u_col_out_325;
wire [1:0] u_col_out_326;
wire [1:0] u_col_out_327;
wire [1:0] u_col_out_328;
wire [1:0] u_col_out_329;
wire [1:0] u_col_out_330;
wire [1:0] u_col_out_331;
wire [1:0] u_col_out_332;
wire [1:0] u_col_out_333;
wire [1:0] u_col_out_334;
wire [1:0] u_col_out_335;
wire [1:0] u_col_out_336;
wire [1:0] u_col_out_337;
wire [1:0] u_col_out_338;
wire [1:0] u_col_out_339;
wire [1:0] u_col_out_340;
wire [1:0] u_col_out_341;
wire [1:0] u_col_out_342;
wire [1:0] u_col_out_343;
wire [1:0] u_col_out_344;
wire [1:0] u_col_out_345;
wire [1:0] u_col_out_346;
wire [1:0] u_col_out_347;
wire [1:0] u_col_out_348;
wire [1:0] u_col_out_349;
wire [1:0] u_col_out_350;
wire [1:0] u_col_out_351;
wire [1:0] u_col_out_352;
wire [1:0] u_col_out_353;
wire [1:0] u_col_out_354;
wire [1:0] u_col_out_355;
wire [1:0] u_col_out_356;
wire [1:0] u_col_out_357;
wire [1:0] u_col_out_358;
wire [1:0] u_col_out_359;
wire [1:0] u_col_out_360;
wire [1:0] u_col_out_361;
wire [1:0] u_col_out_362;
wire [1:0] u_col_out_363;
wire [1:0] u_col_out_364;
wire [1:0] u_col_out_365;
wire [1:0] u_col_out_366;
wire [1:0] u_col_out_367;
wire [1:0] u_col_out_368;
wire [1:0] u_col_out_369;
wire [1:0] u_col_out_370;
wire [1:0] u_col_out_371;
wire [1:0] u_col_out_372;
wire [1:0] u_col_out_373;
wire [1:0] u_col_out_374;
wire [1:0] u_col_out_375;
wire [1:0] u_col_out_376;
wire [1:0] u_col_out_377;
wire [1:0] u_col_out_378;
wire [1:0] u_col_out_379;
wire [1:0] u_col_out_380;
wire [1:0] u_col_out_381;
wire [1:0] u_col_out_382;
wire [1:0] u_col_out_383;
wire [1:0] u_col_out_384;
wire [1:0] u_col_out_385;
wire [1:0] u_col_out_386;
wire [1:0] u_col_out_387;
wire [1:0] u_col_out_388;
wire [1:0] u_col_out_389;
wire [1:0] u_col_out_390;
wire [1:0] u_col_out_391;
wire [1:0] u_col_out_392;
wire [1:0] u_col_out_393;
wire [1:0] u_col_out_394;
wire [1:0] u_col_out_395;
wire [1:0] u_col_out_396;
wire [1:0] u_col_out_397;
wire [1:0] u_col_out_398;
wire [1:0] u_col_out_399;
wire [1:0] u_col_out_400;
wire [1:0] u_col_out_401;
wire [1:0] u_col_out_402;
wire [1:0] u_col_out_403;
wire [1:0] u_col_out_404;
wire [1:0] u_col_out_405;
wire [1:0] u_col_out_406;
wire [1:0] u_col_out_407;
wire [1:0] u_col_out_408;
wire [1:0] u_col_out_409;
wire [1:0] u_col_out_410;
wire [1:0] u_col_out_411;
wire [1:0] u_col_out_412;
wire [1:0] u_col_out_413;
wire [1:0] u_col_out_414;
wire [1:0] u_col_out_415;
wire [1:0] u_col_out_416;
wire [1:0] u_col_out_417;
wire [1:0] u_col_out_418;
wire [1:0] u_col_out_419;
wire [1:0] u_col_out_420;
wire [1:0] u_col_out_421;
wire [1:0] u_col_out_422;
wire [1:0] u_col_out_423;
wire [1:0] u_col_out_424;
wire [1:0] u_col_out_425;
wire [1:0] u_col_out_426;
wire [1:0] u_col_out_427;
wire [1:0] u_col_out_428;
wire [1:0] u_col_out_429;
wire [1:0] u_col_out_430;
wire [1:0] u_col_out_431;
wire [1:0] u_col_out_432;
wire [1:0] u_col_out_433;
wire [1:0] u_col_out_434;
wire [1:0] u_col_out_435;
wire [1:0] u_col_out_436;
wire [1:0] u_col_out_437;
wire [1:0] u_col_out_438;
wire [1:0] u_col_out_439;
wire [1:0] u_col_out_440;
wire [1:0] u_col_out_441;
wire [1:0] u_col_out_442;
wire [1:0] u_col_out_443;
wire [1:0] u_col_out_444;
wire [1:0] u_col_out_445;
wire [1:0] u_col_out_446;
wire [1:0] u_col_out_447;
wire [1:0] u_col_out_448;
wire [1:0] u_col_out_449;
wire [1:0] u_col_out_450;
wire [1:0] u_col_out_451;
wire [1:0] u_col_out_452;
wire [1:0] u_col_out_453;
wire [1:0] u_col_out_454;
wire [1:0] u_col_out_455;
wire [1:0] u_col_out_456;
wire [1:0] u_col_out_457;
wire [1:0] u_col_out_458;
wire [1:0] u_col_out_459;
wire [1:0] u_col_out_460;
wire [1:0] u_col_out_461;
wire [1:0] u_col_out_462;
wire [1:0] u_col_out_463;
wire [1:0] u_col_out_464;
wire [1:0] u_col_out_465;
wire [1:0] u_col_out_466;
wire [1:0] u_col_out_467;
wire [1:0] u_col_out_468;
wire [1:0] u_col_out_469;
wire [1:0] u_col_out_470;
wire [1:0] u_col_out_471;
wire [1:0] u_col_out_472;
wire [1:0] u_col_out_473;
wire [1:0] u_col_out_474;
wire [1:0] u_col_out_475;
wire [1:0] u_col_out_476;
wire [1:0] u_col_out_477;
wire [1:0] u_col_out_478;
wire [1:0] u_col_out_479;
wire [1:0] u_col_out_480;
wire [1:0] u_col_out_481;
wire [1:0] u_col_out_482;
wire [1:0] u_col_out_483;
wire [1:0] u_col_out_484;
wire [1:0] u_col_out_485;
wire [1:0] u_col_out_486;
wire [1:0] u_col_out_487;
wire [1:0] u_col_out_488;
wire [1:0] u_col_out_489;
wire [1:0] u_col_out_490;
wire [1:0] u_col_out_491;
wire [1:0] u_col_out_492;
wire [1:0] u_col_out_493;
wire [1:0] u_col_out_494;
wire [1:0] u_col_out_495;
wire [1:0] u_col_out_496;
wire [1:0] u_col_out_497;
wire [1:0] u_col_out_498;
wire [1:0] u_col_out_499;
wire [1:0] u_col_out_500;
wire [1:0] u_col_out_501;
wire [1:0] u_col_out_502;
wire [1:0] u_col_out_503;
wire [1:0] u_col_out_504;
wire [1:0] u_col_out_505;
wire [1:0] u_col_out_506;
wire [1:0] u_col_out_507;
wire [1:0] u_col_out_508;
wire [1:0] u_col_out_509;
wire [1:0] u_col_out_510;
wire [1:0] u_col_out_511;
wire [1:0] u_col_out_512;
wire [1:0] u_col_out_513;
wire [1:0] u_col_out_514;
wire [1:0] u_col_out_515;
wire [1:0] u_col_out_516;
wire [1:0] u_col_out_517;
wire [1:0] u_col_out_518;
wire [1:0] u_col_out_519;
wire [1:0] u_col_out_520;
wire [1:0] u_col_out_521;
wire [1:0] u_col_out_522;
wire [1:0] u_col_out_523;
wire [1:0] u_col_out_524;
wire [1:0] u_col_out_525;
wire [1:0] u_col_out_526;
wire [1:0] u_col_out_527;
wire [1:0] u_col_out_528;
wire [1:0] u_col_out_529;
wire [1:0] u_col_out_530;
wire [1:0] u_col_out_531;
wire [1:0] u_col_out_532;
wire [1:0] u_col_out_533;
wire [1:0] u_col_out_534;
wire [1:0] u_col_out_535;
wire [1:0] u_col_out_536;
wire [1:0] u_col_out_537;
wire [1:0] u_col_out_538;
wire [1:0] u_col_out_539;
wire [1:0] u_col_out_540;
wire [1:0] u_col_out_541;
wire [1:0] u_col_out_542;
wire [1:0] u_col_out_543;
wire [1:0] u_col_out_544;
wire [1:0] u_col_out_545;
wire [1:0] u_col_out_546;
wire [1:0] u_col_out_547;
wire [1:0] u_col_out_548;
wire [1:0] u_col_out_549;
wire [1:0] u_col_out_550;
wire [1:0] u_col_out_551;
wire [1:0] u_col_out_552;
wire [1:0] u_col_out_553;
wire [1:0] u_col_out_554;
wire [1:0] u_col_out_555;
wire [1:0] u_col_out_556;
wire [1:0] u_col_out_557;
wire [1:0] u_col_out_558;
wire [1:0] u_col_out_559;
wire [1:0] u_col_out_560;
wire [1:0] u_col_out_561;
wire [1:0] u_col_out_562;
wire [1:0] u_col_out_563;
wire [1:0] u_col_out_564;
wire [1:0] u_col_out_565;
wire [1:0] u_col_out_566;
wire [1:0] u_col_out_567;
wire [1:0] u_col_out_568;
wire [1:0] u_col_out_569;
wire [1:0] u_col_out_570;
wire [1:0] u_col_out_571;
wire [1:0] u_col_out_572;
wire [1:0] u_col_out_573;
wire [1:0] u_col_out_574;
wire [1:0] u_col_out_575;
wire [1:0] u_col_out_576;
wire [1:0] u_col_out_577;
wire [1:0] u_col_out_578;
wire [1:0] u_col_out_579;
wire [1:0] u_col_out_580;
wire [1:0] u_col_out_581;
wire [1:0] u_col_out_582;
wire [1:0] u_col_out_583;
wire [1:0] u_col_out_584;
wire [1:0] u_col_out_585;
wire [1:0] u_col_out_586;
wire [1:0] u_col_out_587;
wire [1:0] u_col_out_588;
wire [1:0] u_col_out_589;
wire [1:0] u_col_out_590;
wire [1:0] u_col_out_591;
wire [1:0] u_col_out_592;
wire [1:0] u_col_out_593;
wire [1:0] u_col_out_594;
wire [1:0] u_col_out_595;
wire [1:0] u_col_out_596;
wire [1:0] u_col_out_597;
wire [1:0] u_col_out_598;
wire [1:0] u_col_out_599;
wire [1:0] u_col_out_600;
wire [1:0] u_col_out_601;
wire [1:0] u_col_out_602;
wire [1:0] u_col_out_603;
wire [1:0] u_col_out_604;
wire [1:0] u_col_out_605;
wire [1:0] u_col_out_606;
wire [1:0] u_col_out_607;
wire [1:0] u_col_out_608;
wire [1:0] u_col_out_609;
wire [1:0] u_col_out_610;
wire [1:0] u_col_out_611;
wire [1:0] u_col_out_612;
wire [1:0] u_col_out_613;
wire [1:0] u_col_out_614;
wire [1:0] u_col_out_615;
wire [1:0] u_col_out_616;
wire [1:0] u_col_out_617;
wire [1:0] u_col_out_618;
wire [1:0] u_col_out_619;
wire [1:0] u_col_out_620;
wire [1:0] u_col_out_621;
wire [1:0] u_col_out_622;
wire [1:0] u_col_out_623;
wire [1:0] u_col_out_624;
wire [1:0] u_col_out_625;
wire [1:0] u_col_out_626;
wire [1:0] u_col_out_627;
wire [1:0] u_col_out_628;
wire [1:0] u_col_out_629;
wire [1:0] u_col_out_630;
wire [1:0] u_col_out_631;
wire [1:0] u_col_out_632;
wire [1:0] u_col_out_633;
wire [1:0] u_col_out_634;
wire [1:0] u_col_out_635;
wire [1:0] u_col_out_636;
wire [1:0] u_col_out_637;
wire [1:0] u_col_out_638;
wire [1:0] u_col_out_639;
wire [1:0] u_col_out_640;
wire [1:0] u_col_out_641;
wire [1:0] u_col_out_642;
wire [1:0] u_col_out_643;
wire [1:0] u_col_out_644;
wire [1:0] u_col_out_645;
wire [1:0] u_col_out_646;
wire [1:0] u_col_out_647;
wire [1:0] u_col_out_648;
wire [1:0] u_col_out_649;
wire [1:0] u_col_out_650;
wire [1:0] u_col_out_651;
wire [1:0] u_col_out_652;
wire [1:0] u_col_out_653;
wire [1:0] u_col_out_654;
wire [1:0] u_col_out_655;
wire [1:0] u_col_out_656;
wire [1:0] u_col_out_657;
wire [1:0] u_col_out_658;
wire [1:0] u_col_out_659;
wire [1:0] u_col_out_660;
wire [1:0] u_col_out_661;
wire [1:0] u_col_out_662;
wire [1:0] u_col_out_663;
wire [1:0] u_col_out_664;
wire [1:0] u_col_out_665;
wire [1:0] u_col_out_666;
wire [1:0] u_col_out_667;
wire [1:0] u_col_out_668;
wire [1:0] u_col_out_669;
wire [1:0] u_col_out_670;
wire [1:0] u_col_out_671;
wire [1:0] u_col_out_672;
wire [1:0] u_col_out_673;
wire [1:0] u_col_out_674;
wire [1:0] u_col_out_675;
wire [1:0] u_col_out_676;
wire [1:0] u_col_out_677;
wire [1:0] u_col_out_678;
wire [1:0] u_col_out_679;
wire [1:0] u_col_out_680;
wire [1:0] u_col_out_681;
wire [1:0] u_col_out_682;
wire [1:0] u_col_out_683;
wire [1:0] u_col_out_684;
wire [1:0] u_col_out_685;
wire [1:0] u_col_out_686;
wire [1:0] u_col_out_687;
wire [1:0] u_col_out_688;
wire [1:0] u_col_out_689;
wire [1:0] u_col_out_690;
wire [1:0] u_col_out_691;
wire [1:0] u_col_out_692;
wire [1:0] u_col_out_693;
wire [1:0] u_col_out_694;
wire [1:0] u_col_out_695;
wire [1:0] u_col_out_696;
wire [1:0] u_col_out_697;
wire [1:0] u_col_out_698;
wire [1:0] u_col_out_699;
wire [1:0] u_col_out_700;
wire [1:0] u_col_out_701;
wire [1:0] u_col_out_702;
wire [1:0] u_col_out_703;
wire [1:0] u_col_out_704;
wire [1:0] u_col_out_705;
wire [1:0] u_col_out_706;
wire [1:0] u_col_out_707;
wire [1:0] u_col_out_708;
wire [1:0] u_col_out_709;
wire [1:0] u_col_out_710;
wire [1:0] u_col_out_711;
wire [1:0] u_col_out_712;
wire [1:0] u_col_out_713;
wire [1:0] u_col_out_714;
wire [1:0] u_col_out_715;
wire [1:0] u_col_out_716;
wire [1:0] u_col_out_717;
wire [1:0] u_col_out_718;
wire [1:0] u_col_out_719;
wire [1:0] u_col_out_720;
wire [1:0] u_col_out_721;
wire [1:0] u_col_out_722;
wire [1:0] u_col_out_723;
wire [1:0] u_col_out_724;
wire [1:0] u_col_out_725;
wire [1:0] u_col_out_726;
wire [1:0] u_col_out_727;
wire [1:0] u_col_out_728;
wire [1:0] u_col_out_729;
wire [1:0] u_col_out_730;
wire [1:0] u_col_out_731;
wire [1:0] u_col_out_732;
wire [1:0] u_col_out_733;
wire [1:0] u_col_out_734;
wire [1:0] u_col_out_735;
wire [1:0] u_col_out_736;
wire [1:0] u_col_out_737;
wire [1:0] u_col_out_738;
wire [1:0] u_col_out_739;
wire [1:0] u_col_out_740;
wire [1:0] u_col_out_741;
wire [1:0] u_col_out_742;
wire [1:0] u_col_out_743;
wire [1:0] u_col_out_744;
wire [1:0] u_col_out_745;
wire [1:0] u_col_out_746;
wire [1:0] u_col_out_747;
wire [1:0] u_col_out_748;
wire [1:0] u_col_out_749;
wire [1:0] u_col_out_750;
wire [1:0] u_col_out_751;
wire [1:0] u_col_out_752;
wire [1:0] u_col_out_753;
wire [1:0] u_col_out_754;
wire [1:0] u_col_out_755;
wire [1:0] u_col_out_756;
wire [1:0] u_col_out_757;
wire [1:0] u_col_out_758;
wire [1:0] u_col_out_759;
wire [1:0] u_col_out_760;
wire [1:0] u_col_out_761;
wire [1:0] u_col_out_762;
wire [1:0] u_col_out_763;
wire [1:0] u_col_out_764;
wire [1:0] u_col_out_765;
wire [1:0] u_col_out_766;
wire [1:0] u_col_out_767;
wire [1:0] u_col_out_768;
wire [1:0] u_col_out_769;
wire [1:0] u_col_out_770;
wire [1:0] u_col_out_771;
wire [1:0] u_col_out_772;
wire [1:0] u_col_out_773;
wire [1:0] u_col_out_774;
wire [1:0] u_col_out_775;
wire [1:0] u_col_out_776;
wire [1:0] u_col_out_777;
wire [1:0] u_col_out_778;
wire [1:0] u_col_out_779;
wire [1:0] u_col_out_780;
wire [1:0] u_col_out_781;
wire [1:0] u_col_out_782;
wire [1:0] u_col_out_783;
wire [1:0] u_col_out_784;
wire [1:0] u_col_out_785;
wire [1:0] u_col_out_786;
wire [1:0] u_col_out_787;
wire [1:0] u_col_out_788;
wire [1:0] u_col_out_789;
wire [1:0] u_col_out_790;
wire [1:0] u_col_out_791;
wire [1:0] u_col_out_792;
wire [1:0] u_col_out_793;
wire [1:0] u_col_out_794;
wire [1:0] u_col_out_795;
wire [1:0] u_col_out_796;
wire [1:0] u_col_out_797;
wire [1:0] u_col_out_798;
wire [1:0] u_col_out_799;
wire [1:0] u_col_out_800;
wire [1:0] u_col_out_801;
wire [1:0] u_col_out_802;
wire [1:0] u_col_out_803;
wire [1:0] u_col_out_804;
wire [1:0] u_col_out_805;
wire [1:0] u_col_out_806;
wire [1:0] u_col_out_807;
wire [1:0] u_col_out_808;
wire [1:0] u_col_out_809;
wire [1:0] u_col_out_810;
wire [1:0] u_col_out_811;
wire [1:0] u_col_out_812;
wire [1:0] u_col_out_813;
wire [1:0] u_col_out_814;
wire [1:0] u_col_out_815;
wire [1:0] u_col_out_816;
wire [1:0] u_col_out_817;
wire [1:0] u_col_out_818;
wire [1:0] u_col_out_819;
wire [1:0] u_col_out_820;
wire [1:0] u_col_out_821;
wire [1:0] u_col_out_822;
wire [1:0] u_col_out_823;
wire [1:0] u_col_out_824;
wire [1:0] u_col_out_825;
wire [1:0] u_col_out_826;
wire [1:0] u_col_out_827;
wire [1:0] u_col_out_828;
wire [1:0] u_col_out_829;
wire [1:0] u_col_out_830;
wire [1:0] u_col_out_831;
wire [1:0] u_col_out_832;
wire [1:0] u_col_out_833;
wire [1:0] u_col_out_834;
wire [1:0] u_col_out_835;
wire [1:0] u_col_out_836;
wire [1:0] u_col_out_837;
wire [1:0] u_col_out_838;
wire [1:0] u_col_out_839;
wire [1:0] u_col_out_840;
wire [1:0] u_col_out_841;
wire [1:0] u_col_out_842;
wire [1:0] u_col_out_843;
wire [1:0] u_col_out_844;
wire [1:0] u_col_out_845;
wire [1:0] u_col_out_846;
wire [1:0] u_col_out_847;
wire [1:0] u_col_out_848;
wire [1:0] u_col_out_849;
wire [1:0] u_col_out_850;
wire [1:0] u_col_out_851;
wire [1:0] u_col_out_852;
wire [1:0] u_col_out_853;
wire [1:0] u_col_out_854;
wire [1:0] u_col_out_855;
wire [1:0] u_col_out_856;
wire [1:0] u_col_out_857;
wire [1:0] u_col_out_858;
wire [1:0] u_col_out_859;
wire [1:0] u_col_out_860;
wire [1:0] u_col_out_861;
wire [1:0] u_col_out_862;
wire [1:0] u_col_out_863;
wire [1:0] u_col_out_864;
wire [1:0] u_col_out_865;
wire [1:0] u_col_out_866;
wire [1:0] u_col_out_867;
wire [1:0] u_col_out_868;
wire [1:0] u_col_out_869;
wire [1:0] u_col_out_870;
wire [1:0] u_col_out_871;
wire [1:0] u_col_out_872;
wire [1:0] u_col_out_873;
wire [1:0] u_col_out_874;
wire [1:0] u_col_out_875;
wire [1:0] u_col_out_876;
wire [1:0] u_col_out_877;
wire [1:0] u_col_out_878;
wire [1:0] u_col_out_879;
wire [1:0] u_col_out_880;
wire [1:0] u_col_out_881;
wire [1:0] u_col_out_882;
wire [1:0] u_col_out_883;
wire [1:0] u_col_out_884;
wire [1:0] u_col_out_885;
wire [1:0] u_col_out_886;
wire [1:0] u_col_out_887;
wire [1:0] u_col_out_888;
wire [1:0] u_col_out_889;
wire [1:0] u_col_out_890;
wire [1:0] u_col_out_891;
wire [1:0] u_col_out_892;
wire [1:0] u_col_out_893;
wire [1:0] u_col_out_894;
wire [1:0] u_col_out_895;
wire [1:0] u_col_out_896;
wire [1:0] u_col_out_897;
wire [1:0] u_col_out_898;
wire [1:0] u_col_out_899;
wire [1:0] u_col_out_900;
wire [1:0] u_col_out_901;
wire [1:0] u_col_out_902;
wire [1:0] u_col_out_903;
wire [1:0] u_col_out_904;
wire [1:0] u_col_out_905;
wire [1:0] u_col_out_906;
wire [1:0] u_col_out_907;
wire [1:0] u_col_out_908;
wire [1:0] u_col_out_909;
wire [1:0] u_col_out_910;
wire [1:0] u_col_out_911;
wire [1:0] u_col_out_912;
wire [1:0] u_col_out_913;
wire [1:0] u_col_out_914;
wire [1:0] u_col_out_915;
wire [1:0] u_col_out_916;
wire [1:0] u_col_out_917;
wire [1:0] u_col_out_918;
wire [1:0] u_col_out_919;
wire [1:0] u_col_out_920;
wire [1:0] u_col_out_921;
wire [1:0] u_col_out_922;
wire [1:0] u_col_out_923;
wire [1:0] u_col_out_924;
wire [1:0] u_col_out_925;
wire [1:0] u_col_out_926;
wire [1:0] u_col_out_927;
wire [1:0] u_col_out_928;
wire [1:0] u_col_out_929;
wire [1:0] u_col_out_930;
wire [1:0] u_col_out_931;
wire [1:0] u_col_out_932;
wire [1:0] u_col_out_933;
wire [1:0] u_col_out_934;
wire [1:0] u_col_out_935;
wire [1:0] u_col_out_936;
wire [1:0] u_col_out_937;
wire [1:0] u_col_out_938;
wire [1:0] u_col_out_939;
wire [1:0] u_col_out_940;
wire [1:0] u_col_out_941;
wire [1:0] u_col_out_942;
wire [1:0] u_col_out_943;
wire [1:0] u_col_out_944;
wire [1:0] u_col_out_945;
wire [1:0] u_col_out_946;
wire [1:0] u_col_out_947;
wire [1:0] u_col_out_948;
wire [1:0] u_col_out_949;
wire [1:0] u_col_out_950;
wire [1:0] u_col_out_951;
wire [1:0] u_col_out_952;
wire [1:0] u_col_out_953;
wire [1:0] u_col_out_954;
wire [1:0] u_col_out_955;
wire [1:0] u_col_out_956;
wire [1:0] u_col_out_957;
wire [1:0] u_col_out_958;
wire [1:0] u_col_out_959;
wire [1:0] u_col_out_960;
wire [1:0] u_col_out_961;
wire [1:0] u_col_out_962;
wire [1:0] u_col_out_963;
wire [1:0] u_col_out_964;
wire [1:0] u_col_out_965;
wire [1:0] u_col_out_966;
wire [1:0] u_col_out_967;
wire [1:0] u_col_out_968;
wire [1:0] u_col_out_969;
wire [1:0] u_col_out_970;
wire [1:0] u_col_out_971;
wire [1:0] u_col_out_972;
wire [1:0] u_col_out_973;
wire [1:0] u_col_out_974;
wire [1:0] u_col_out_975;
wire [1:0] u_col_out_976;
wire [1:0] u_col_out_977;
wire [1:0] u_col_out_978;
wire [1:0] u_col_out_979;
wire [1:0] u_col_out_980;
wire [1:0] u_col_out_981;
wire [1:0] u_col_out_982;
wire [1:0] u_col_out_983;
wire [1:0] u_col_out_984;
wire [1:0] u_col_out_985;
wire [1:0] u_col_out_986;
wire [1:0] u_col_out_987;
wire [1:0] u_col_out_988;
wire [1:0] u_col_out_989;
wire [1:0] u_col_out_990;
wire [1:0] u_col_out_991;
wire [1:0] u_col_out_992;
wire [1:0] u_col_out_993;
wire [1:0] u_col_out_994;
wire [1:0] u_col_out_995;
wire [1:0] u_col_out_996;
wire [1:0] u_col_out_997;
wire [1:0] u_col_out_998;
wire [1:0] u_col_out_999;
wire [1:0] u_col_out_1000;
wire [1:0] u_col_out_1001;
wire [1:0] u_col_out_1002;
wire [1:0] u_col_out_1003;
wire [1:0] u_col_out_1004;
wire [1:0] u_col_out_1005;
wire [1:0] u_col_out_1006;
wire [1:0] u_col_out_1007;
wire [1:0] u_col_out_1008;
wire [1:0] u_col_out_1009;
wire [1:0] u_col_out_1010;
wire [1:0] u_col_out_1011;
wire [1:0] u_col_out_1012;
wire [1:0] u_col_out_1013;
wire [1:0] u_col_out_1014;
wire [1:0] u_col_out_1015;
wire [1:0] u_col_out_1016;
wire [1:0] u_col_out_1017;
wire [1:0] u_col_out_1018;
wire [1:0] u_col_out_1019;
wire [1:0] u_col_out_1020;
wire [1:0] u_col_out_1021;
wire [1:0] u_col_out_1022;
wire [1:0] u_col_out_1023;
wire [1:0] u_col_out_1024;
wire [1:0] u_col_out_1025;
wire [1:0] u_col_out_1026;
wire [1:0] u_col_out_1027;
wire [1:0] u_col_out_1028;
wire [1:0] u_col_out_1029;
wire [1:0] u_col_out_1030;
wire [1:0] u_col_out_1031;
wire [1:0] u_col_out_1032;
wire [1:0] u_col_out_1033;
wire [1:0] u_col_out_1034;
wire [1:0] u_col_out_1035;
wire [1:0] u_col_out_1036;
wire [1:0] u_col_out_1037;
wire [1:0] u_col_out_1038;
wire [1:0] u_col_out_1039;
wire [1:0] u_col_out_1040;
wire [1:0] u_col_out_1041;
wire [1:0] u_col_out_1042;
wire [1:0] u_col_out_1043;
wire [1:0] u_col_out_1044;
wire [1:0] u_col_out_1045;
wire [1:0] u_col_out_1046;
wire [1:0] u_col_out_1047;
wire [1:0] u_col_out_1048;
wire [1:0] u_col_out_1049;
wire [1:0] u_col_out_1050;
wire [1:0] u_col_out_1051;
wire [1:0] u_col_out_1052;
wire [1:0] u_col_out_1053;
wire [1:0] u_col_out_1054;
wire [1:0] u_col_out_1055;
wire [1:0] u_col_out_1056;
wire [1:0] u_col_out_1057;
wire [1:0] u_col_out_1058;
wire [1:0] u_col_out_1059;
wire [1:0] u_col_out_1060;
wire [1:0] u_col_out_1061;
wire [1:0] u_col_out_1062;
wire [1:0] u_col_out_1063;
wire [1:0] u_col_out_1064;
wire [1:0] u_col_out_1065;
wire [1:0] u_col_out_1066;
wire [1:0] u_col_out_1067;
wire [1:0] u_col_out_1068;
wire [1:0] u_col_out_1069;
wire [1:0] u_col_out_1070;
wire [1:0] u_col_out_1071;
wire [1:0] u_col_out_1072;
wire [1:0] u_col_out_1073;
wire [1:0] u_col_out_1074;
wire [1:0] u_col_out_1075;
wire [1:0] u_col_out_1076;
wire [1:0] u_col_out_1077;
wire [1:0] u_col_out_1078;
wire [1:0] u_col_out_1079;
wire [1:0] u_col_out_1080;
wire [1:0] u_col_out_1081;
wire [1:0] u_col_out_1082;
wire [1:0] u_col_out_1083;
wire [1:0] u_col_out_1084;
wire [1:0] u_col_out_1085;
wire [1:0] u_col_out_1086;
wire [1:0] u_col_out_1087;
wire [1:0] u_col_out_1088;
wire [1:0] u_col_out_1089;
wire [1:0] u_col_out_1090;
wire [1:0] u_col_out_1091;
wire [1:0] u_col_out_1092;
wire [1:0] u_col_out_1093;
wire [1:0] u_col_out_1094;
wire [1:0] u_col_out_1095;
wire [1:0] u_col_out_1096;
wire [1:0] u_col_out_1097;
wire [1:0] u_col_out_1098;
wire [1:0] u_col_out_1099;
wire [1:0] u_col_out_1100;
wire [1:0] u_col_out_1101;
wire [1:0] u_col_out_1102;
wire [1:0] u_col_out_1103;
wire [1:0] u_col_out_1104;
wire [1:0] u_col_out_1105;
wire [1:0] u_col_out_1106;
wire [1:0] u_col_out_1107;
wire [1:0] u_col_out_1108;
wire [1:0] u_col_out_1109;
wire [1:0] u_col_out_1110;
wire [1:0] u_col_out_1111;
wire [1:0] u_col_out_1112;
wire [1:0] u_col_out_1113;
wire [1:0] u_col_out_1114;
wire [1:0] u_col_out_1115;
wire [1:0] u_col_out_1116;
wire [1:0] u_col_out_1117;
wire [1:0] u_col_out_1118;
wire [1:0] u_col_out_1119;
wire [1:0] u_col_out_1120;
wire [1:0] u_col_out_1121;
wire [1:0] u_col_out_1122;
wire [1:0] u_col_out_1123;
wire [1:0] u_col_out_1124;
wire [1:0] u_col_out_1125;
wire [1:0] u_col_out_1126;
wire [1:0] u_col_out_1127;
wire [1:0] u_col_out_1128;
wire [1:0] u_col_out_1129;
wire [1:0] u_col_out_1130;
wire [1:0] u_col_out_1131;
wire [1:0] u_col_out_1132;
wire [1:0] u_col_out_1133;
wire [1:0] u_col_out_1134;
wire [1:0] u_col_out_1135;
wire [1:0] u_col_out_1136;
wire [1:0] u_col_out_1137;
wire [1:0] u_col_out_1138;
wire [1:0] u_col_out_1139;
wire [1:0] u_col_out_1140;
wire [1:0] u_col_out_1141;
wire [1:0] u_col_out_1142;
wire [1:0] u_col_out_1143;
wire [1:0] u_col_out_1144;
wire [1:0] u_col_out_1145;
wire [1:0] u_col_out_1146;
wire [1:0] u_col_out_1147;
wire [1:0] u_col_out_1148;
wire [1:0] u_col_out_1149;
wire [1:0] u_col_out_1150;
wire [1:0] u_col_out_1151;
wire [1:0] u_col_out_1152;
wire [1:0] u_col_out_1153;
wire [1:0] u_col_out_1154;
wire [1:0] u_col_out_1155;
wire [1:0] u_col_out_1156;
wire [1:0] u_col_out_1157;
wire [1:0] u_col_out_1158;
wire [1:0] u_col_out_1159;
wire [1:0] u_col_out_1160;
wire [1:0] u_col_out_1161;
wire [1:0] u_col_out_1162;
wire [1:0] u_col_out_1163;
wire [1:0] u_col_out_1164;
wire [1:0] u_col_out_1165;
wire [1:0] u_col_out_1166;
wire [1:0] u_col_out_1167;
wire [1:0] u_col_out_1168;
wire [1:0] u_col_out_1169;
wire [1:0] u_col_out_1170;
wire [1:0] u_col_out_1171;
wire [1:0] u_col_out_1172;
wire [1:0] u_col_out_1173;
wire [1:0] u_col_out_1174;
wire [1:0] u_col_out_1175;
wire [1:0] u_col_out_1176;
wire [1:0] u_col_out_1177;
wire [1:0] u_col_out_1178;
wire [1:0] u_col_out_1179;
wire [1:0] u_col_out_1180;
wire [1:0] u_col_out_1181;
wire [1:0] u_col_out_1182;
wire [1:0] u_col_out_1183;
wire [1:0] u_col_out_1184;
wire [1:0] u_col_out_1185;
wire [1:0] u_col_out_1186;
wire [1:0] u_col_out_1187;
wire [1:0] u_col_out_1188;
wire [1:0] u_col_out_1189;
wire [1:0] u_col_out_1190;
wire [1:0] u_col_out_1191;
wire [1:0] u_col_out_1192;
wire [1:0] u_col_out_1193;
wire [1:0] u_col_out_1194;
wire [1:0] u_col_out_1195;
wire [1:0] u_col_out_1196;
wire [1:0] u_col_out_1197;
wire [1:0] u_col_out_1198;
wire [1:0] u_col_out_1199;
wire [1:0] u_col_out_1200;
wire [1:0] u_col_out_1201;
wire [1:0] u_col_out_1202;
wire [1:0] u_col_out_1203;
wire [1:0] u_col_out_1204;
wire [1:0] u_col_out_1205;
wire [1:0] u_col_out_1206;
wire [1:0] u_col_out_1207;
wire [1:0] u_col_out_1208;
wire [1:0] u_col_out_1209;
wire [1:0] u_col_out_1210;
wire [1:0] u_col_out_1211;
wire [1:0] u_col_out_1212;
wire [1:0] u_col_out_1213;
wire [1:0] u_col_out_1214;
wire [1:0] u_col_out_1215;
wire [1:0] u_col_out_1216;
wire [1:0] u_col_out_1217;
wire [1:0] u_col_out_1218;
wire [1:0] u_col_out_1219;
wire [1:0] u_col_out_1220;
wire [1:0] u_col_out_1221;
wire [1:0] u_col_out_1222;
wire [1:0] u_col_out_1223;
wire [1:0] u_col_out_1224;
wire [1:0] u_col_out_1225;
wire [1:0] u_col_out_1226;
wire [1:0] u_col_out_1227;
wire [1:0] u_col_out_1228;
wire [1:0] u_col_out_1229;
wire [1:0] u_col_out_1230;
wire [1:0] u_col_out_1231;
wire [1:0] u_col_out_1232;
wire [1:0] u_col_out_1233;
wire [1:0] u_col_out_1234;
wire [1:0] u_col_out_1235;
wire [1:0] u_col_out_1236;
wire [1:0] u_col_out_1237;
wire [1:0] u_col_out_1238;
wire [1:0] u_col_out_1239;
wire [1:0] u_col_out_1240;
wire [1:0] u_col_out_1241;
wire [1:0] u_col_out_1242;
wire [1:0] u_col_out_1243;
wire [1:0] u_col_out_1244;
wire [1:0] u_col_out_1245;
wire [1:0] u_col_out_1246;
wire [1:0] u_col_out_1247;
wire [1:0] u_col_out_1248;
wire [1:0] u_col_out_1249;
wire [1:0] u_col_out_1250;
wire [1:0] u_col_out_1251;
wire [1:0] u_col_out_1252;
wire [1:0] u_col_out_1253;
wire [1:0] u_col_out_1254;
wire [1:0] u_col_out_1255;
wire [1:0] u_col_out_1256;
wire [1:0] u_col_out_1257;
wire [1:0] u_col_out_1258;
wire [1:0] u_col_out_1259;
wire [1:0] u_col_out_1260;
wire [1:0] u_col_out_1261;
wire [1:0] u_col_out_1262;
wire [1:0] u_col_out_1263;
wire [1:0] u_col_out_1264;
wire [1:0] u_col_out_1265;
wire [1:0] u_col_out_1266;
wire [1:0] u_col_out_1267;
wire [1:0] u_col_out_1268;
wire [1:0] u_col_out_1269;
wire [1:0] u_col_out_1270;
wire [1:0] u_col_out_1271;
wire [1:0] u_col_out_1272;
wire [1:0] u_col_out_1273;
wire [1:0] u_col_out_1274;
wire [1:0] u_col_out_1275;
wire [1:0] u_col_out_1276;
wire [1:0] u_col_out_1277;
wire [1:0] u_col_out_1278;
wire [1:0] u_col_out_1279;
wire [1:0] u_col_out_1280;
wire [1:0] u_col_out_1281;
wire [1:0] u_col_out_1282;
wire [1:0] u_col_out_1283;
wire [1:0] u_col_out_1284;
wire [1:0] u_col_out_1285;
wire [1:0] u_col_out_1286;
wire [1:0] u_col_out_1287;


compressor_array_236_2_1280 u_compressor_array_236_2_1280
(
    .col_in_0(col_in_0),
    .col_in_1(col_in_1),
    .col_in_2(col_in_2),
    .col_in_3(col_in_3),
    .col_in_4(col_in_4),
    .col_in_5(col_in_5),
    .col_in_6(col_in_6),
    .col_in_7(col_in_7),
    .col_in_8(col_in_8),
    .col_in_9(col_in_9),
    .col_in_10(col_in_10),
    .col_in_11(col_in_11),
    .col_in_12(col_in_12),
    .col_in_13(col_in_13),
    .col_in_14(col_in_14),
    .col_in_15(col_in_15),
    .col_in_16(col_in_16),
    .col_in_17(col_in_17),
    .col_in_18(col_in_18),
    .col_in_19(col_in_19),
    .col_in_20(col_in_20),
    .col_in_21(col_in_21),
    .col_in_22(col_in_22),
    .col_in_23(col_in_23),
    .col_in_24(col_in_24),
    .col_in_25(col_in_25),
    .col_in_26(col_in_26),
    .col_in_27(col_in_27),
    .col_in_28(col_in_28),
    .col_in_29(col_in_29),
    .col_in_30(col_in_30),
    .col_in_31(col_in_31),
    .col_in_32(col_in_32),
    .col_in_33(col_in_33),
    .col_in_34(col_in_34),
    .col_in_35(col_in_35),
    .col_in_36(col_in_36),
    .col_in_37(col_in_37),
    .col_in_38(col_in_38),
    .col_in_39(col_in_39),
    .col_in_40(col_in_40),
    .col_in_41(col_in_41),
    .col_in_42(col_in_42),
    .col_in_43(col_in_43),
    .col_in_44(col_in_44),
    .col_in_45(col_in_45),
    .col_in_46(col_in_46),
    .col_in_47(col_in_47),
    .col_in_48(col_in_48),
    .col_in_49(col_in_49),
    .col_in_50(col_in_50),
    .col_in_51(col_in_51),
    .col_in_52(col_in_52),
    .col_in_53(col_in_53),
    .col_in_54(col_in_54),
    .col_in_55(col_in_55),
    .col_in_56(col_in_56),
    .col_in_57(col_in_57),
    .col_in_58(col_in_58),
    .col_in_59(col_in_59),
    .col_in_60(col_in_60),
    .col_in_61(col_in_61),
    .col_in_62(col_in_62),
    .col_in_63(col_in_63),
    .col_in_64(col_in_64),
    .col_in_65(col_in_65),
    .col_in_66(col_in_66),
    .col_in_67(col_in_67),
    .col_in_68(col_in_68),
    .col_in_69(col_in_69),
    .col_in_70(col_in_70),
    .col_in_71(col_in_71),
    .col_in_72(col_in_72),
    .col_in_73(col_in_73),
    .col_in_74(col_in_74),
    .col_in_75(col_in_75),
    .col_in_76(col_in_76),
    .col_in_77(col_in_77),
    .col_in_78(col_in_78),
    .col_in_79(col_in_79),
    .col_in_80(col_in_80),
    .col_in_81(col_in_81),
    .col_in_82(col_in_82),
    .col_in_83(col_in_83),
    .col_in_84(col_in_84),
    .col_in_85(col_in_85),
    .col_in_86(col_in_86),
    .col_in_87(col_in_87),
    .col_in_88(col_in_88),
    .col_in_89(col_in_89),
    .col_in_90(col_in_90),
    .col_in_91(col_in_91),
    .col_in_92(col_in_92),
    .col_in_93(col_in_93),
    .col_in_94(col_in_94),
    .col_in_95(col_in_95),
    .col_in_96(col_in_96),
    .col_in_97(col_in_97),
    .col_in_98(col_in_98),
    .col_in_99(col_in_99),
    .col_in_100(col_in_100),
    .col_in_101(col_in_101),
    .col_in_102(col_in_102),
    .col_in_103(col_in_103),
    .col_in_104(col_in_104),
    .col_in_105(col_in_105),
    .col_in_106(col_in_106),
    .col_in_107(col_in_107),
    .col_in_108(col_in_108),
    .col_in_109(col_in_109),
    .col_in_110(col_in_110),
    .col_in_111(col_in_111),
    .col_in_112(col_in_112),
    .col_in_113(col_in_113),
    .col_in_114(col_in_114),
    .col_in_115(col_in_115),
    .col_in_116(col_in_116),
    .col_in_117(col_in_117),
    .col_in_118(col_in_118),
    .col_in_119(col_in_119),
    .col_in_120(col_in_120),
    .col_in_121(col_in_121),
    .col_in_122(col_in_122),
    .col_in_123(col_in_123),
    .col_in_124(col_in_124),
    .col_in_125(col_in_125),
    .col_in_126(col_in_126),
    .col_in_127(col_in_127),
    .col_in_128(col_in_128),
    .col_in_129(col_in_129),
    .col_in_130(col_in_130),
    .col_in_131(col_in_131),
    .col_in_132(col_in_132),
    .col_in_133(col_in_133),
    .col_in_134(col_in_134),
    .col_in_135(col_in_135),
    .col_in_136(col_in_136),
    .col_in_137(col_in_137),
    .col_in_138(col_in_138),
    .col_in_139(col_in_139),
    .col_in_140(col_in_140),
    .col_in_141(col_in_141),
    .col_in_142(col_in_142),
    .col_in_143(col_in_143),
    .col_in_144(col_in_144),
    .col_in_145(col_in_145),
    .col_in_146(col_in_146),
    .col_in_147(col_in_147),
    .col_in_148(col_in_148),
    .col_in_149(col_in_149),
    .col_in_150(col_in_150),
    .col_in_151(col_in_151),
    .col_in_152(col_in_152),
    .col_in_153(col_in_153),
    .col_in_154(col_in_154),
    .col_in_155(col_in_155),
    .col_in_156(col_in_156),
    .col_in_157(col_in_157),
    .col_in_158(col_in_158),
    .col_in_159(col_in_159),
    .col_in_160(col_in_160),
    .col_in_161(col_in_161),
    .col_in_162(col_in_162),
    .col_in_163(col_in_163),
    .col_in_164(col_in_164),
    .col_in_165(col_in_165),
    .col_in_166(col_in_166),
    .col_in_167(col_in_167),
    .col_in_168(col_in_168),
    .col_in_169(col_in_169),
    .col_in_170(col_in_170),
    .col_in_171(col_in_171),
    .col_in_172(col_in_172),
    .col_in_173(col_in_173),
    .col_in_174(col_in_174),
    .col_in_175(col_in_175),
    .col_in_176(col_in_176),
    .col_in_177(col_in_177),
    .col_in_178(col_in_178),
    .col_in_179(col_in_179),
    .col_in_180(col_in_180),
    .col_in_181(col_in_181),
    .col_in_182(col_in_182),
    .col_in_183(col_in_183),
    .col_in_184(col_in_184),
    .col_in_185(col_in_185),
    .col_in_186(col_in_186),
    .col_in_187(col_in_187),
    .col_in_188(col_in_188),
    .col_in_189(col_in_189),
    .col_in_190(col_in_190),
    .col_in_191(col_in_191),
    .col_in_192(col_in_192),
    .col_in_193(col_in_193),
    .col_in_194(col_in_194),
    .col_in_195(col_in_195),
    .col_in_196(col_in_196),
    .col_in_197(col_in_197),
    .col_in_198(col_in_198),
    .col_in_199(col_in_199),
    .col_in_200(col_in_200),
    .col_in_201(col_in_201),
    .col_in_202(col_in_202),
    .col_in_203(col_in_203),
    .col_in_204(col_in_204),
    .col_in_205(col_in_205),
    .col_in_206(col_in_206),
    .col_in_207(col_in_207),
    .col_in_208(col_in_208),
    .col_in_209(col_in_209),
    .col_in_210(col_in_210),
    .col_in_211(col_in_211),
    .col_in_212(col_in_212),
    .col_in_213(col_in_213),
    .col_in_214(col_in_214),
    .col_in_215(col_in_215),
    .col_in_216(col_in_216),
    .col_in_217(col_in_217),
    .col_in_218(col_in_218),
    .col_in_219(col_in_219),
    .col_in_220(col_in_220),
    .col_in_221(col_in_221),
    .col_in_222(col_in_222),
    .col_in_223(col_in_223),
    .col_in_224(col_in_224),
    .col_in_225(col_in_225),
    .col_in_226(col_in_226),
    .col_in_227(col_in_227),
    .col_in_228(col_in_228),
    .col_in_229(col_in_229),
    .col_in_230(col_in_230),
    .col_in_231(col_in_231),
    .col_in_232(col_in_232),
    .col_in_233(col_in_233),
    .col_in_234(col_in_234),
    .col_in_235(col_in_235),
    .col_in_236(col_in_236),
    .col_in_237(col_in_237),
    .col_in_238(col_in_238),
    .col_in_239(col_in_239),
    .col_in_240(col_in_240),
    .col_in_241(col_in_241),
    .col_in_242(col_in_242),
    .col_in_243(col_in_243),
    .col_in_244(col_in_244),
    .col_in_245(col_in_245),
    .col_in_246(col_in_246),
    .col_in_247(col_in_247),
    .col_in_248(col_in_248),
    .col_in_249(col_in_249),
    .col_in_250(col_in_250),
    .col_in_251(col_in_251),
    .col_in_252(col_in_252),
    .col_in_253(col_in_253),
    .col_in_254(col_in_254),
    .col_in_255(col_in_255),
    .col_in_256(col_in_256),
    .col_in_257(col_in_257),
    .col_in_258(col_in_258),
    .col_in_259(col_in_259),
    .col_in_260(col_in_260),
    .col_in_261(col_in_261),
    .col_in_262(col_in_262),
    .col_in_263(col_in_263),
    .col_in_264(col_in_264),
    .col_in_265(col_in_265),
    .col_in_266(col_in_266),
    .col_in_267(col_in_267),
    .col_in_268(col_in_268),
    .col_in_269(col_in_269),
    .col_in_270(col_in_270),
    .col_in_271(col_in_271),
    .col_in_272(col_in_272),
    .col_in_273(col_in_273),
    .col_in_274(col_in_274),
    .col_in_275(col_in_275),
    .col_in_276(col_in_276),
    .col_in_277(col_in_277),
    .col_in_278(col_in_278),
    .col_in_279(col_in_279),
    .col_in_280(col_in_280),
    .col_in_281(col_in_281),
    .col_in_282(col_in_282),
    .col_in_283(col_in_283),
    .col_in_284(col_in_284),
    .col_in_285(col_in_285),
    .col_in_286(col_in_286),
    .col_in_287(col_in_287),
    .col_in_288(col_in_288),
    .col_in_289(col_in_289),
    .col_in_290(col_in_290),
    .col_in_291(col_in_291),
    .col_in_292(col_in_292),
    .col_in_293(col_in_293),
    .col_in_294(col_in_294),
    .col_in_295(col_in_295),
    .col_in_296(col_in_296),
    .col_in_297(col_in_297),
    .col_in_298(col_in_298),
    .col_in_299(col_in_299),
    .col_in_300(col_in_300),
    .col_in_301(col_in_301),
    .col_in_302(col_in_302),
    .col_in_303(col_in_303),
    .col_in_304(col_in_304),
    .col_in_305(col_in_305),
    .col_in_306(col_in_306),
    .col_in_307(col_in_307),
    .col_in_308(col_in_308),
    .col_in_309(col_in_309),
    .col_in_310(col_in_310),
    .col_in_311(col_in_311),
    .col_in_312(col_in_312),
    .col_in_313(col_in_313),
    .col_in_314(col_in_314),
    .col_in_315(col_in_315),
    .col_in_316(col_in_316),
    .col_in_317(col_in_317),
    .col_in_318(col_in_318),
    .col_in_319(col_in_319),
    .col_in_320(col_in_320),
    .col_in_321(col_in_321),
    .col_in_322(col_in_322),
    .col_in_323(col_in_323),
    .col_in_324(col_in_324),
    .col_in_325(col_in_325),
    .col_in_326(col_in_326),
    .col_in_327(col_in_327),
    .col_in_328(col_in_328),
    .col_in_329(col_in_329),
    .col_in_330(col_in_330),
    .col_in_331(col_in_331),
    .col_in_332(col_in_332),
    .col_in_333(col_in_333),
    .col_in_334(col_in_334),
    .col_in_335(col_in_335),
    .col_in_336(col_in_336),
    .col_in_337(col_in_337),
    .col_in_338(col_in_338),
    .col_in_339(col_in_339),
    .col_in_340(col_in_340),
    .col_in_341(col_in_341),
    .col_in_342(col_in_342),
    .col_in_343(col_in_343),
    .col_in_344(col_in_344),
    .col_in_345(col_in_345),
    .col_in_346(col_in_346),
    .col_in_347(col_in_347),
    .col_in_348(col_in_348),
    .col_in_349(col_in_349),
    .col_in_350(col_in_350),
    .col_in_351(col_in_351),
    .col_in_352(col_in_352),
    .col_in_353(col_in_353),
    .col_in_354(col_in_354),
    .col_in_355(col_in_355),
    .col_in_356(col_in_356),
    .col_in_357(col_in_357),
    .col_in_358(col_in_358),
    .col_in_359(col_in_359),
    .col_in_360(col_in_360),
    .col_in_361(col_in_361),
    .col_in_362(col_in_362),
    .col_in_363(col_in_363),
    .col_in_364(col_in_364),
    .col_in_365(col_in_365),
    .col_in_366(col_in_366),
    .col_in_367(col_in_367),
    .col_in_368(col_in_368),
    .col_in_369(col_in_369),
    .col_in_370(col_in_370),
    .col_in_371(col_in_371),
    .col_in_372(col_in_372),
    .col_in_373(col_in_373),
    .col_in_374(col_in_374),
    .col_in_375(col_in_375),
    .col_in_376(col_in_376),
    .col_in_377(col_in_377),
    .col_in_378(col_in_378),
    .col_in_379(col_in_379),
    .col_in_380(col_in_380),
    .col_in_381(col_in_381),
    .col_in_382(col_in_382),
    .col_in_383(col_in_383),
    .col_in_384(col_in_384),
    .col_in_385(col_in_385),
    .col_in_386(col_in_386),
    .col_in_387(col_in_387),
    .col_in_388(col_in_388),
    .col_in_389(col_in_389),
    .col_in_390(col_in_390),
    .col_in_391(col_in_391),
    .col_in_392(col_in_392),
    .col_in_393(col_in_393),
    .col_in_394(col_in_394),
    .col_in_395(col_in_395),
    .col_in_396(col_in_396),
    .col_in_397(col_in_397),
    .col_in_398(col_in_398),
    .col_in_399(col_in_399),
    .col_in_400(col_in_400),
    .col_in_401(col_in_401),
    .col_in_402(col_in_402),
    .col_in_403(col_in_403),
    .col_in_404(col_in_404),
    .col_in_405(col_in_405),
    .col_in_406(col_in_406),
    .col_in_407(col_in_407),
    .col_in_408(col_in_408),
    .col_in_409(col_in_409),
    .col_in_410(col_in_410),
    .col_in_411(col_in_411),
    .col_in_412(col_in_412),
    .col_in_413(col_in_413),
    .col_in_414(col_in_414),
    .col_in_415(col_in_415),
    .col_in_416(col_in_416),
    .col_in_417(col_in_417),
    .col_in_418(col_in_418),
    .col_in_419(col_in_419),
    .col_in_420(col_in_420),
    .col_in_421(col_in_421),
    .col_in_422(col_in_422),
    .col_in_423(col_in_423),
    .col_in_424(col_in_424),
    .col_in_425(col_in_425),
    .col_in_426(col_in_426),
    .col_in_427(col_in_427),
    .col_in_428(col_in_428),
    .col_in_429(col_in_429),
    .col_in_430(col_in_430),
    .col_in_431(col_in_431),
    .col_in_432(col_in_432),
    .col_in_433(col_in_433),
    .col_in_434(col_in_434),
    .col_in_435(col_in_435),
    .col_in_436(col_in_436),
    .col_in_437(col_in_437),
    .col_in_438(col_in_438),
    .col_in_439(col_in_439),
    .col_in_440(col_in_440),
    .col_in_441(col_in_441),
    .col_in_442(col_in_442),
    .col_in_443(col_in_443),
    .col_in_444(col_in_444),
    .col_in_445(col_in_445),
    .col_in_446(col_in_446),
    .col_in_447(col_in_447),
    .col_in_448(col_in_448),
    .col_in_449(col_in_449),
    .col_in_450(col_in_450),
    .col_in_451(col_in_451),
    .col_in_452(col_in_452),
    .col_in_453(col_in_453),
    .col_in_454(col_in_454),
    .col_in_455(col_in_455),
    .col_in_456(col_in_456),
    .col_in_457(col_in_457),
    .col_in_458(col_in_458),
    .col_in_459(col_in_459),
    .col_in_460(col_in_460),
    .col_in_461(col_in_461),
    .col_in_462(col_in_462),
    .col_in_463(col_in_463),
    .col_in_464(col_in_464),
    .col_in_465(col_in_465),
    .col_in_466(col_in_466),
    .col_in_467(col_in_467),
    .col_in_468(col_in_468),
    .col_in_469(col_in_469),
    .col_in_470(col_in_470),
    .col_in_471(col_in_471),
    .col_in_472(col_in_472),
    .col_in_473(col_in_473),
    .col_in_474(col_in_474),
    .col_in_475(col_in_475),
    .col_in_476(col_in_476),
    .col_in_477(col_in_477),
    .col_in_478(col_in_478),
    .col_in_479(col_in_479),
    .col_in_480(col_in_480),
    .col_in_481(col_in_481),
    .col_in_482(col_in_482),
    .col_in_483(col_in_483),
    .col_in_484(col_in_484),
    .col_in_485(col_in_485),
    .col_in_486(col_in_486),
    .col_in_487(col_in_487),
    .col_in_488(col_in_488),
    .col_in_489(col_in_489),
    .col_in_490(col_in_490),
    .col_in_491(col_in_491),
    .col_in_492(col_in_492),
    .col_in_493(col_in_493),
    .col_in_494(col_in_494),
    .col_in_495(col_in_495),
    .col_in_496(col_in_496),
    .col_in_497(col_in_497),
    .col_in_498(col_in_498),
    .col_in_499(col_in_499),
    .col_in_500(col_in_500),
    .col_in_501(col_in_501),
    .col_in_502(col_in_502),
    .col_in_503(col_in_503),
    .col_in_504(col_in_504),
    .col_in_505(col_in_505),
    .col_in_506(col_in_506),
    .col_in_507(col_in_507),
    .col_in_508(col_in_508),
    .col_in_509(col_in_509),
    .col_in_510(col_in_510),
    .col_in_511(col_in_511),
    .col_in_512(col_in_512),
    .col_in_513(col_in_513),
    .col_in_514(col_in_514),
    .col_in_515(col_in_515),
    .col_in_516(col_in_516),
    .col_in_517(col_in_517),
    .col_in_518(col_in_518),
    .col_in_519(col_in_519),
    .col_in_520(col_in_520),
    .col_in_521(col_in_521),
    .col_in_522(col_in_522),
    .col_in_523(col_in_523),
    .col_in_524(col_in_524),
    .col_in_525(col_in_525),
    .col_in_526(col_in_526),
    .col_in_527(col_in_527),
    .col_in_528(col_in_528),
    .col_in_529(col_in_529),
    .col_in_530(col_in_530),
    .col_in_531(col_in_531),
    .col_in_532(col_in_532),
    .col_in_533(col_in_533),
    .col_in_534(col_in_534),
    .col_in_535(col_in_535),
    .col_in_536(col_in_536),
    .col_in_537(col_in_537),
    .col_in_538(col_in_538),
    .col_in_539(col_in_539),
    .col_in_540(col_in_540),
    .col_in_541(col_in_541),
    .col_in_542(col_in_542),
    .col_in_543(col_in_543),
    .col_in_544(col_in_544),
    .col_in_545(col_in_545),
    .col_in_546(col_in_546),
    .col_in_547(col_in_547),
    .col_in_548(col_in_548),
    .col_in_549(col_in_549),
    .col_in_550(col_in_550),
    .col_in_551(col_in_551),
    .col_in_552(col_in_552),
    .col_in_553(col_in_553),
    .col_in_554(col_in_554),
    .col_in_555(col_in_555),
    .col_in_556(col_in_556),
    .col_in_557(col_in_557),
    .col_in_558(col_in_558),
    .col_in_559(col_in_559),
    .col_in_560(col_in_560),
    .col_in_561(col_in_561),
    .col_in_562(col_in_562),
    .col_in_563(col_in_563),
    .col_in_564(col_in_564),
    .col_in_565(col_in_565),
    .col_in_566(col_in_566),
    .col_in_567(col_in_567),
    .col_in_568(col_in_568),
    .col_in_569(col_in_569),
    .col_in_570(col_in_570),
    .col_in_571(col_in_571),
    .col_in_572(col_in_572),
    .col_in_573(col_in_573),
    .col_in_574(col_in_574),
    .col_in_575(col_in_575),
    .col_in_576(col_in_576),
    .col_in_577(col_in_577),
    .col_in_578(col_in_578),
    .col_in_579(col_in_579),
    .col_in_580(col_in_580),
    .col_in_581(col_in_581),
    .col_in_582(col_in_582),
    .col_in_583(col_in_583),
    .col_in_584(col_in_584),
    .col_in_585(col_in_585),
    .col_in_586(col_in_586),
    .col_in_587(col_in_587),
    .col_in_588(col_in_588),
    .col_in_589(col_in_589),
    .col_in_590(col_in_590),
    .col_in_591(col_in_591),
    .col_in_592(col_in_592),
    .col_in_593(col_in_593),
    .col_in_594(col_in_594),
    .col_in_595(col_in_595),
    .col_in_596(col_in_596),
    .col_in_597(col_in_597),
    .col_in_598(col_in_598),
    .col_in_599(col_in_599),
    .col_in_600(col_in_600),
    .col_in_601(col_in_601),
    .col_in_602(col_in_602),
    .col_in_603(col_in_603),
    .col_in_604(col_in_604),
    .col_in_605(col_in_605),
    .col_in_606(col_in_606),
    .col_in_607(col_in_607),
    .col_in_608(col_in_608),
    .col_in_609(col_in_609),
    .col_in_610(col_in_610),
    .col_in_611(col_in_611),
    .col_in_612(col_in_612),
    .col_in_613(col_in_613),
    .col_in_614(col_in_614),
    .col_in_615(col_in_615),
    .col_in_616(col_in_616),
    .col_in_617(col_in_617),
    .col_in_618(col_in_618),
    .col_in_619(col_in_619),
    .col_in_620(col_in_620),
    .col_in_621(col_in_621),
    .col_in_622(col_in_622),
    .col_in_623(col_in_623),
    .col_in_624(col_in_624),
    .col_in_625(col_in_625),
    .col_in_626(col_in_626),
    .col_in_627(col_in_627),
    .col_in_628(col_in_628),
    .col_in_629(col_in_629),
    .col_in_630(col_in_630),
    .col_in_631(col_in_631),
    .col_in_632(col_in_632),
    .col_in_633(col_in_633),
    .col_in_634(col_in_634),
    .col_in_635(col_in_635),
    .col_in_636(col_in_636),
    .col_in_637(col_in_637),
    .col_in_638(col_in_638),
    .col_in_639(col_in_639),
    .col_in_640(col_in_640),
    .col_in_641(col_in_641),
    .col_in_642(col_in_642),
    .col_in_643(col_in_643),
    .col_in_644(col_in_644),
    .col_in_645(col_in_645),
    .col_in_646(col_in_646),
    .col_in_647(col_in_647),
    .col_in_648(col_in_648),
    .col_in_649(col_in_649),
    .col_in_650(col_in_650),
    .col_in_651(col_in_651),
    .col_in_652(col_in_652),
    .col_in_653(col_in_653),
    .col_in_654(col_in_654),
    .col_in_655(col_in_655),
    .col_in_656(col_in_656),
    .col_in_657(col_in_657),
    .col_in_658(col_in_658),
    .col_in_659(col_in_659),
    .col_in_660(col_in_660),
    .col_in_661(col_in_661),
    .col_in_662(col_in_662),
    .col_in_663(col_in_663),
    .col_in_664(col_in_664),
    .col_in_665(col_in_665),
    .col_in_666(col_in_666),
    .col_in_667(col_in_667),
    .col_in_668(col_in_668),
    .col_in_669(col_in_669),
    .col_in_670(col_in_670),
    .col_in_671(col_in_671),
    .col_in_672(col_in_672),
    .col_in_673(col_in_673),
    .col_in_674(col_in_674),
    .col_in_675(col_in_675),
    .col_in_676(col_in_676),
    .col_in_677(col_in_677),
    .col_in_678(col_in_678),
    .col_in_679(col_in_679),
    .col_in_680(col_in_680),
    .col_in_681(col_in_681),
    .col_in_682(col_in_682),
    .col_in_683(col_in_683),
    .col_in_684(col_in_684),
    .col_in_685(col_in_685),
    .col_in_686(col_in_686),
    .col_in_687(col_in_687),
    .col_in_688(col_in_688),
    .col_in_689(col_in_689),
    .col_in_690(col_in_690),
    .col_in_691(col_in_691),
    .col_in_692(col_in_692),
    .col_in_693(col_in_693),
    .col_in_694(col_in_694),
    .col_in_695(col_in_695),
    .col_in_696(col_in_696),
    .col_in_697(col_in_697),
    .col_in_698(col_in_698),
    .col_in_699(col_in_699),
    .col_in_700(col_in_700),
    .col_in_701(col_in_701),
    .col_in_702(col_in_702),
    .col_in_703(col_in_703),
    .col_in_704(col_in_704),
    .col_in_705(col_in_705),
    .col_in_706(col_in_706),
    .col_in_707(col_in_707),
    .col_in_708(col_in_708),
    .col_in_709(col_in_709),
    .col_in_710(col_in_710),
    .col_in_711(col_in_711),
    .col_in_712(col_in_712),
    .col_in_713(col_in_713),
    .col_in_714(col_in_714),
    .col_in_715(col_in_715),
    .col_in_716(col_in_716),
    .col_in_717(col_in_717),
    .col_in_718(col_in_718),
    .col_in_719(col_in_719),
    .col_in_720(col_in_720),
    .col_in_721(col_in_721),
    .col_in_722(col_in_722),
    .col_in_723(col_in_723),
    .col_in_724(col_in_724),
    .col_in_725(col_in_725),
    .col_in_726(col_in_726),
    .col_in_727(col_in_727),
    .col_in_728(col_in_728),
    .col_in_729(col_in_729),
    .col_in_730(col_in_730),
    .col_in_731(col_in_731),
    .col_in_732(col_in_732),
    .col_in_733(col_in_733),
    .col_in_734(col_in_734),
    .col_in_735(col_in_735),
    .col_in_736(col_in_736),
    .col_in_737(col_in_737),
    .col_in_738(col_in_738),
    .col_in_739(col_in_739),
    .col_in_740(col_in_740),
    .col_in_741(col_in_741),
    .col_in_742(col_in_742),
    .col_in_743(col_in_743),
    .col_in_744(col_in_744),
    .col_in_745(col_in_745),
    .col_in_746(col_in_746),
    .col_in_747(col_in_747),
    .col_in_748(col_in_748),
    .col_in_749(col_in_749),
    .col_in_750(col_in_750),
    .col_in_751(col_in_751),
    .col_in_752(col_in_752),
    .col_in_753(col_in_753),
    .col_in_754(col_in_754),
    .col_in_755(col_in_755),
    .col_in_756(col_in_756),
    .col_in_757(col_in_757),
    .col_in_758(col_in_758),
    .col_in_759(col_in_759),
    .col_in_760(col_in_760),
    .col_in_761(col_in_761),
    .col_in_762(col_in_762),
    .col_in_763(col_in_763),
    .col_in_764(col_in_764),
    .col_in_765(col_in_765),
    .col_in_766(col_in_766),
    .col_in_767(col_in_767),
    .col_in_768(col_in_768),
    .col_in_769(col_in_769),
    .col_in_770(col_in_770),
    .col_in_771(col_in_771),
    .col_in_772(col_in_772),
    .col_in_773(col_in_773),
    .col_in_774(col_in_774),
    .col_in_775(col_in_775),
    .col_in_776(col_in_776),
    .col_in_777(col_in_777),
    .col_in_778(col_in_778),
    .col_in_779(col_in_779),
    .col_in_780(col_in_780),
    .col_in_781(col_in_781),
    .col_in_782(col_in_782),
    .col_in_783(col_in_783),
    .col_in_784(col_in_784),
    .col_in_785(col_in_785),
    .col_in_786(col_in_786),
    .col_in_787(col_in_787),
    .col_in_788(col_in_788),
    .col_in_789(col_in_789),
    .col_in_790(col_in_790),
    .col_in_791(col_in_791),
    .col_in_792(col_in_792),
    .col_in_793(col_in_793),
    .col_in_794(col_in_794),
    .col_in_795(col_in_795),
    .col_in_796(col_in_796),
    .col_in_797(col_in_797),
    .col_in_798(col_in_798),
    .col_in_799(col_in_799),
    .col_in_800(col_in_800),
    .col_in_801(col_in_801),
    .col_in_802(col_in_802),
    .col_in_803(col_in_803),
    .col_in_804(col_in_804),
    .col_in_805(col_in_805),
    .col_in_806(col_in_806),
    .col_in_807(col_in_807),
    .col_in_808(col_in_808),
    .col_in_809(col_in_809),
    .col_in_810(col_in_810),
    .col_in_811(col_in_811),
    .col_in_812(col_in_812),
    .col_in_813(col_in_813),
    .col_in_814(col_in_814),
    .col_in_815(col_in_815),
    .col_in_816(col_in_816),
    .col_in_817(col_in_817),
    .col_in_818(col_in_818),
    .col_in_819(col_in_819),
    .col_in_820(col_in_820),
    .col_in_821(col_in_821),
    .col_in_822(col_in_822),
    .col_in_823(col_in_823),
    .col_in_824(col_in_824),
    .col_in_825(col_in_825),
    .col_in_826(col_in_826),
    .col_in_827(col_in_827),
    .col_in_828(col_in_828),
    .col_in_829(col_in_829),
    .col_in_830(col_in_830),
    .col_in_831(col_in_831),
    .col_in_832(col_in_832),
    .col_in_833(col_in_833),
    .col_in_834(col_in_834),
    .col_in_835(col_in_835),
    .col_in_836(col_in_836),
    .col_in_837(col_in_837),
    .col_in_838(col_in_838),
    .col_in_839(col_in_839),
    .col_in_840(col_in_840),
    .col_in_841(col_in_841),
    .col_in_842(col_in_842),
    .col_in_843(col_in_843),
    .col_in_844(col_in_844),
    .col_in_845(col_in_845),
    .col_in_846(col_in_846),
    .col_in_847(col_in_847),
    .col_in_848(col_in_848),
    .col_in_849(col_in_849),
    .col_in_850(col_in_850),
    .col_in_851(col_in_851),
    .col_in_852(col_in_852),
    .col_in_853(col_in_853),
    .col_in_854(col_in_854),
    .col_in_855(col_in_855),
    .col_in_856(col_in_856),
    .col_in_857(col_in_857),
    .col_in_858(col_in_858),
    .col_in_859(col_in_859),
    .col_in_860(col_in_860),
    .col_in_861(col_in_861),
    .col_in_862(col_in_862),
    .col_in_863(col_in_863),
    .col_in_864(col_in_864),
    .col_in_865(col_in_865),
    .col_in_866(col_in_866),
    .col_in_867(col_in_867),
    .col_in_868(col_in_868),
    .col_in_869(col_in_869),
    .col_in_870(col_in_870),
    .col_in_871(col_in_871),
    .col_in_872(col_in_872),
    .col_in_873(col_in_873),
    .col_in_874(col_in_874),
    .col_in_875(col_in_875),
    .col_in_876(col_in_876),
    .col_in_877(col_in_877),
    .col_in_878(col_in_878),
    .col_in_879(col_in_879),
    .col_in_880(col_in_880),
    .col_in_881(col_in_881),
    .col_in_882(col_in_882),
    .col_in_883(col_in_883),
    .col_in_884(col_in_884),
    .col_in_885(col_in_885),
    .col_in_886(col_in_886),
    .col_in_887(col_in_887),
    .col_in_888(col_in_888),
    .col_in_889(col_in_889),
    .col_in_890(col_in_890),
    .col_in_891(col_in_891),
    .col_in_892(col_in_892),
    .col_in_893(col_in_893),
    .col_in_894(col_in_894),
    .col_in_895(col_in_895),
    .col_in_896(col_in_896),
    .col_in_897(col_in_897),
    .col_in_898(col_in_898),
    .col_in_899(col_in_899),
    .col_in_900(col_in_900),
    .col_in_901(col_in_901),
    .col_in_902(col_in_902),
    .col_in_903(col_in_903),
    .col_in_904(col_in_904),
    .col_in_905(col_in_905),
    .col_in_906(col_in_906),
    .col_in_907(col_in_907),
    .col_in_908(col_in_908),
    .col_in_909(col_in_909),
    .col_in_910(col_in_910),
    .col_in_911(col_in_911),
    .col_in_912(col_in_912),
    .col_in_913(col_in_913),
    .col_in_914(col_in_914),
    .col_in_915(col_in_915),
    .col_in_916(col_in_916),
    .col_in_917(col_in_917),
    .col_in_918(col_in_918),
    .col_in_919(col_in_919),
    .col_in_920(col_in_920),
    .col_in_921(col_in_921),
    .col_in_922(col_in_922),
    .col_in_923(col_in_923),
    .col_in_924(col_in_924),
    .col_in_925(col_in_925),
    .col_in_926(col_in_926),
    .col_in_927(col_in_927),
    .col_in_928(col_in_928),
    .col_in_929(col_in_929),
    .col_in_930(col_in_930),
    .col_in_931(col_in_931),
    .col_in_932(col_in_932),
    .col_in_933(col_in_933),
    .col_in_934(col_in_934),
    .col_in_935(col_in_935),
    .col_in_936(col_in_936),
    .col_in_937(col_in_937),
    .col_in_938(col_in_938),
    .col_in_939(col_in_939),
    .col_in_940(col_in_940),
    .col_in_941(col_in_941),
    .col_in_942(col_in_942),
    .col_in_943(col_in_943),
    .col_in_944(col_in_944),
    .col_in_945(col_in_945),
    .col_in_946(col_in_946),
    .col_in_947(col_in_947),
    .col_in_948(col_in_948),
    .col_in_949(col_in_949),
    .col_in_950(col_in_950),
    .col_in_951(col_in_951),
    .col_in_952(col_in_952),
    .col_in_953(col_in_953),
    .col_in_954(col_in_954),
    .col_in_955(col_in_955),
    .col_in_956(col_in_956),
    .col_in_957(col_in_957),
    .col_in_958(col_in_958),
    .col_in_959(col_in_959),
    .col_in_960(col_in_960),
    .col_in_961(col_in_961),
    .col_in_962(col_in_962),
    .col_in_963(col_in_963),
    .col_in_964(col_in_964),
    .col_in_965(col_in_965),
    .col_in_966(col_in_966),
    .col_in_967(col_in_967),
    .col_in_968(col_in_968),
    .col_in_969(col_in_969),
    .col_in_970(col_in_970),
    .col_in_971(col_in_971),
    .col_in_972(col_in_972),
    .col_in_973(col_in_973),
    .col_in_974(col_in_974),
    .col_in_975(col_in_975),
    .col_in_976(col_in_976),
    .col_in_977(col_in_977),
    .col_in_978(col_in_978),
    .col_in_979(col_in_979),
    .col_in_980(col_in_980),
    .col_in_981(col_in_981),
    .col_in_982(col_in_982),
    .col_in_983(col_in_983),
    .col_in_984(col_in_984),
    .col_in_985(col_in_985),
    .col_in_986(col_in_986),
    .col_in_987(col_in_987),
    .col_in_988(col_in_988),
    .col_in_989(col_in_989),
    .col_in_990(col_in_990),
    .col_in_991(col_in_991),
    .col_in_992(col_in_992),
    .col_in_993(col_in_993),
    .col_in_994(col_in_994),
    .col_in_995(col_in_995),
    .col_in_996(col_in_996),
    .col_in_997(col_in_997),
    .col_in_998(col_in_998),
    .col_in_999(col_in_999),
    .col_in_1000(col_in_1000),
    .col_in_1001(col_in_1001),
    .col_in_1002(col_in_1002),
    .col_in_1003(col_in_1003),
    .col_in_1004(col_in_1004),
    .col_in_1005(col_in_1005),
    .col_in_1006(col_in_1006),
    .col_in_1007(col_in_1007),
    .col_in_1008(col_in_1008),
    .col_in_1009(col_in_1009),
    .col_in_1010(col_in_1010),
    .col_in_1011(col_in_1011),
    .col_in_1012(col_in_1012),
    .col_in_1013(col_in_1013),
    .col_in_1014(col_in_1014),
    .col_in_1015(col_in_1015),
    .col_in_1016(col_in_1016),
    .col_in_1017(col_in_1017),
    .col_in_1018(col_in_1018),
    .col_in_1019(col_in_1019),
    .col_in_1020(col_in_1020),
    .col_in_1021(col_in_1021),
    .col_in_1022(col_in_1022),
    .col_in_1023(col_in_1023),
    .col_in_1024(col_in_1024),
    .col_in_1025(col_in_1025),
    .col_in_1026(col_in_1026),
    .col_in_1027(col_in_1027),
    .col_in_1028(col_in_1028),
    .col_in_1029(col_in_1029),
    .col_in_1030(col_in_1030),
    .col_in_1031(col_in_1031),
    .col_in_1032(col_in_1032),
    .col_in_1033(col_in_1033),
    .col_in_1034(col_in_1034),
    .col_in_1035(col_in_1035),
    .col_in_1036(col_in_1036),
    .col_in_1037(col_in_1037),
    .col_in_1038(col_in_1038),
    .col_in_1039(col_in_1039),
    .col_in_1040(col_in_1040),
    .col_in_1041(col_in_1041),
    .col_in_1042(col_in_1042),
    .col_in_1043(col_in_1043),
    .col_in_1044(col_in_1044),
    .col_in_1045(col_in_1045),
    .col_in_1046(col_in_1046),
    .col_in_1047(col_in_1047),
    .col_in_1048(col_in_1048),
    .col_in_1049(col_in_1049),
    .col_in_1050(col_in_1050),
    .col_in_1051(col_in_1051),
    .col_in_1052(col_in_1052),
    .col_in_1053(col_in_1053),
    .col_in_1054(col_in_1054),
    .col_in_1055(col_in_1055),
    .col_in_1056(col_in_1056),
    .col_in_1057(col_in_1057),
    .col_in_1058(col_in_1058),
    .col_in_1059(col_in_1059),
    .col_in_1060(col_in_1060),
    .col_in_1061(col_in_1061),
    .col_in_1062(col_in_1062),
    .col_in_1063(col_in_1063),
    .col_in_1064(col_in_1064),
    .col_in_1065(col_in_1065),
    .col_in_1066(col_in_1066),
    .col_in_1067(col_in_1067),
    .col_in_1068(col_in_1068),
    .col_in_1069(col_in_1069),
    .col_in_1070(col_in_1070),
    .col_in_1071(col_in_1071),
    .col_in_1072(col_in_1072),
    .col_in_1073(col_in_1073),
    .col_in_1074(col_in_1074),
    .col_in_1075(col_in_1075),
    .col_in_1076(col_in_1076),
    .col_in_1077(col_in_1077),
    .col_in_1078(col_in_1078),
    .col_in_1079(col_in_1079),
    .col_in_1080(col_in_1080),
    .col_in_1081(col_in_1081),
    .col_in_1082(col_in_1082),
    .col_in_1083(col_in_1083),
    .col_in_1084(col_in_1084),
    .col_in_1085(col_in_1085),
    .col_in_1086(col_in_1086),
    .col_in_1087(col_in_1087),
    .col_in_1088(col_in_1088),
    .col_in_1089(col_in_1089),
    .col_in_1090(col_in_1090),
    .col_in_1091(col_in_1091),
    .col_in_1092(col_in_1092),
    .col_in_1093(col_in_1093),
    .col_in_1094(col_in_1094),
    .col_in_1095(col_in_1095),
    .col_in_1096(col_in_1096),
    .col_in_1097(col_in_1097),
    .col_in_1098(col_in_1098),
    .col_in_1099(col_in_1099),
    .col_in_1100(col_in_1100),
    .col_in_1101(col_in_1101),
    .col_in_1102(col_in_1102),
    .col_in_1103(col_in_1103),
    .col_in_1104(col_in_1104),
    .col_in_1105(col_in_1105),
    .col_in_1106(col_in_1106),
    .col_in_1107(col_in_1107),
    .col_in_1108(col_in_1108),
    .col_in_1109(col_in_1109),
    .col_in_1110(col_in_1110),
    .col_in_1111(col_in_1111),
    .col_in_1112(col_in_1112),
    .col_in_1113(col_in_1113),
    .col_in_1114(col_in_1114),
    .col_in_1115(col_in_1115),
    .col_in_1116(col_in_1116),
    .col_in_1117(col_in_1117),
    .col_in_1118(col_in_1118),
    .col_in_1119(col_in_1119),
    .col_in_1120(col_in_1120),
    .col_in_1121(col_in_1121),
    .col_in_1122(col_in_1122),
    .col_in_1123(col_in_1123),
    .col_in_1124(col_in_1124),
    .col_in_1125(col_in_1125),
    .col_in_1126(col_in_1126),
    .col_in_1127(col_in_1127),
    .col_in_1128(col_in_1128),
    .col_in_1129(col_in_1129),
    .col_in_1130(col_in_1130),
    .col_in_1131(col_in_1131),
    .col_in_1132(col_in_1132),
    .col_in_1133(col_in_1133),
    .col_in_1134(col_in_1134),
    .col_in_1135(col_in_1135),
    .col_in_1136(col_in_1136),
    .col_in_1137(col_in_1137),
    .col_in_1138(col_in_1138),
    .col_in_1139(col_in_1139),
    .col_in_1140(col_in_1140),
    .col_in_1141(col_in_1141),
    .col_in_1142(col_in_1142),
    .col_in_1143(col_in_1143),
    .col_in_1144(col_in_1144),
    .col_in_1145(col_in_1145),
    .col_in_1146(col_in_1146),
    .col_in_1147(col_in_1147),
    .col_in_1148(col_in_1148),
    .col_in_1149(col_in_1149),
    .col_in_1150(col_in_1150),
    .col_in_1151(col_in_1151),
    .col_in_1152(col_in_1152),
    .col_in_1153(col_in_1153),
    .col_in_1154(col_in_1154),
    .col_in_1155(col_in_1155),
    .col_in_1156(col_in_1156),
    .col_in_1157(col_in_1157),
    .col_in_1158(col_in_1158),
    .col_in_1159(col_in_1159),
    .col_in_1160(col_in_1160),
    .col_in_1161(col_in_1161),
    .col_in_1162(col_in_1162),
    .col_in_1163(col_in_1163),
    .col_in_1164(col_in_1164),
    .col_in_1165(col_in_1165),
    .col_in_1166(col_in_1166),
    .col_in_1167(col_in_1167),
    .col_in_1168(col_in_1168),
    .col_in_1169(col_in_1169),
    .col_in_1170(col_in_1170),
    .col_in_1171(col_in_1171),
    .col_in_1172(col_in_1172),
    .col_in_1173(col_in_1173),
    .col_in_1174(col_in_1174),
    .col_in_1175(col_in_1175),
    .col_in_1176(col_in_1176),
    .col_in_1177(col_in_1177),
    .col_in_1178(col_in_1178),
    .col_in_1179(col_in_1179),
    .col_in_1180(col_in_1180),
    .col_in_1181(col_in_1181),
    .col_in_1182(col_in_1182),
    .col_in_1183(col_in_1183),
    .col_in_1184(col_in_1184),
    .col_in_1185(col_in_1185),
    .col_in_1186(col_in_1186),
    .col_in_1187(col_in_1187),
    .col_in_1188(col_in_1188),
    .col_in_1189(col_in_1189),
    .col_in_1190(col_in_1190),
    .col_in_1191(col_in_1191),
    .col_in_1192(col_in_1192),
    .col_in_1193(col_in_1193),
    .col_in_1194(col_in_1194),
    .col_in_1195(col_in_1195),
    .col_in_1196(col_in_1196),
    .col_in_1197(col_in_1197),
    .col_in_1198(col_in_1198),
    .col_in_1199(col_in_1199),
    .col_in_1200(col_in_1200),
    .col_in_1201(col_in_1201),
    .col_in_1202(col_in_1202),
    .col_in_1203(col_in_1203),
    .col_in_1204(col_in_1204),
    .col_in_1205(col_in_1205),
    .col_in_1206(col_in_1206),
    .col_in_1207(col_in_1207),
    .col_in_1208(col_in_1208),
    .col_in_1209(col_in_1209),
    .col_in_1210(col_in_1210),
    .col_in_1211(col_in_1211),
    .col_in_1212(col_in_1212),
    .col_in_1213(col_in_1213),
    .col_in_1214(col_in_1214),
    .col_in_1215(col_in_1215),
    .col_in_1216(col_in_1216),
    .col_in_1217(col_in_1217),
    .col_in_1218(col_in_1218),
    .col_in_1219(col_in_1219),
    .col_in_1220(col_in_1220),
    .col_in_1221(col_in_1221),
    .col_in_1222(col_in_1222),
    .col_in_1223(col_in_1223),
    .col_in_1224(col_in_1224),
    .col_in_1225(col_in_1225),
    .col_in_1226(col_in_1226),
    .col_in_1227(col_in_1227),
    .col_in_1228(col_in_1228),
    .col_in_1229(col_in_1229),
    .col_in_1230(col_in_1230),
    .col_in_1231(col_in_1231),
    .col_in_1232(col_in_1232),
    .col_in_1233(col_in_1233),
    .col_in_1234(col_in_1234),
    .col_in_1235(col_in_1235),
    .col_in_1236(col_in_1236),
    .col_in_1237(col_in_1237),
    .col_in_1238(col_in_1238),
    .col_in_1239(col_in_1239),
    .col_in_1240(col_in_1240),
    .col_in_1241(col_in_1241),
    .col_in_1242(col_in_1242),
    .col_in_1243(col_in_1243),
    .col_in_1244(col_in_1244),
    .col_in_1245(col_in_1245),
    .col_in_1246(col_in_1246),
    .col_in_1247(col_in_1247),
    .col_in_1248(col_in_1248),
    .col_in_1249(col_in_1249),
    .col_in_1250(col_in_1250),
    .col_in_1251(col_in_1251),
    .col_in_1252(col_in_1252),
    .col_in_1253(col_in_1253),
    .col_in_1254(col_in_1254),
    .col_in_1255(col_in_1255),
    .col_in_1256(col_in_1256),
    .col_in_1257(col_in_1257),
    .col_in_1258(col_in_1258),
    .col_in_1259(col_in_1259),
    .col_in_1260(col_in_1260),
    .col_in_1261(col_in_1261),
    .col_in_1262(col_in_1262),
    .col_in_1263(col_in_1263),
    .col_in_1264(col_in_1264),
    .col_in_1265(col_in_1265),
    .col_in_1266(col_in_1266),
    .col_in_1267(col_in_1267),
    .col_in_1268(col_in_1268),
    .col_in_1269(col_in_1269),
    .col_in_1270(col_in_1270),
    .col_in_1271(col_in_1271),
    .col_in_1272(col_in_1272),
    .col_in_1273(col_in_1273),
    .col_in_1274(col_in_1274),
    .col_in_1275(col_in_1275),
    .col_in_1276(col_in_1276),
    .col_in_1277(col_in_1277),
    .col_in_1278(col_in_1278),
    .col_in_1279(col_in_1279),


    .col_out_0(u_col_out_0),
    .col_out_1(u_col_out_1),
    .col_out_2(u_col_out_2),
    .col_out_3(u_col_out_3),
    .col_out_4(u_col_out_4),
    .col_out_5(u_col_out_5),
    .col_out_6(u_col_out_6),
    .col_out_7(u_col_out_7),
    .col_out_8(u_col_out_8),
    .col_out_9(u_col_out_9),
    .col_out_10(u_col_out_10),
    .col_out_11(u_col_out_11),
    .col_out_12(u_col_out_12),
    .col_out_13(u_col_out_13),
    .col_out_14(u_col_out_14),
    .col_out_15(u_col_out_15),
    .col_out_16(u_col_out_16),
    .col_out_17(u_col_out_17),
    .col_out_18(u_col_out_18),
    .col_out_19(u_col_out_19),
    .col_out_20(u_col_out_20),
    .col_out_21(u_col_out_21),
    .col_out_22(u_col_out_22),
    .col_out_23(u_col_out_23),
    .col_out_24(u_col_out_24),
    .col_out_25(u_col_out_25),
    .col_out_26(u_col_out_26),
    .col_out_27(u_col_out_27),
    .col_out_28(u_col_out_28),
    .col_out_29(u_col_out_29),
    .col_out_30(u_col_out_30),
    .col_out_31(u_col_out_31),
    .col_out_32(u_col_out_32),
    .col_out_33(u_col_out_33),
    .col_out_34(u_col_out_34),
    .col_out_35(u_col_out_35),
    .col_out_36(u_col_out_36),
    .col_out_37(u_col_out_37),
    .col_out_38(u_col_out_38),
    .col_out_39(u_col_out_39),
    .col_out_40(u_col_out_40),
    .col_out_41(u_col_out_41),
    .col_out_42(u_col_out_42),
    .col_out_43(u_col_out_43),
    .col_out_44(u_col_out_44),
    .col_out_45(u_col_out_45),
    .col_out_46(u_col_out_46),
    .col_out_47(u_col_out_47),
    .col_out_48(u_col_out_48),
    .col_out_49(u_col_out_49),
    .col_out_50(u_col_out_50),
    .col_out_51(u_col_out_51),
    .col_out_52(u_col_out_52),
    .col_out_53(u_col_out_53),
    .col_out_54(u_col_out_54),
    .col_out_55(u_col_out_55),
    .col_out_56(u_col_out_56),
    .col_out_57(u_col_out_57),
    .col_out_58(u_col_out_58),
    .col_out_59(u_col_out_59),
    .col_out_60(u_col_out_60),
    .col_out_61(u_col_out_61),
    .col_out_62(u_col_out_62),
    .col_out_63(u_col_out_63),
    .col_out_64(u_col_out_64),
    .col_out_65(u_col_out_65),
    .col_out_66(u_col_out_66),
    .col_out_67(u_col_out_67),
    .col_out_68(u_col_out_68),
    .col_out_69(u_col_out_69),
    .col_out_70(u_col_out_70),
    .col_out_71(u_col_out_71),
    .col_out_72(u_col_out_72),
    .col_out_73(u_col_out_73),
    .col_out_74(u_col_out_74),
    .col_out_75(u_col_out_75),
    .col_out_76(u_col_out_76),
    .col_out_77(u_col_out_77),
    .col_out_78(u_col_out_78),
    .col_out_79(u_col_out_79),
    .col_out_80(u_col_out_80),
    .col_out_81(u_col_out_81),
    .col_out_82(u_col_out_82),
    .col_out_83(u_col_out_83),
    .col_out_84(u_col_out_84),
    .col_out_85(u_col_out_85),
    .col_out_86(u_col_out_86),
    .col_out_87(u_col_out_87),
    .col_out_88(u_col_out_88),
    .col_out_89(u_col_out_89),
    .col_out_90(u_col_out_90),
    .col_out_91(u_col_out_91),
    .col_out_92(u_col_out_92),
    .col_out_93(u_col_out_93),
    .col_out_94(u_col_out_94),
    .col_out_95(u_col_out_95),
    .col_out_96(u_col_out_96),
    .col_out_97(u_col_out_97),
    .col_out_98(u_col_out_98),
    .col_out_99(u_col_out_99),
    .col_out_100(u_col_out_100),
    .col_out_101(u_col_out_101),
    .col_out_102(u_col_out_102),
    .col_out_103(u_col_out_103),
    .col_out_104(u_col_out_104),
    .col_out_105(u_col_out_105),
    .col_out_106(u_col_out_106),
    .col_out_107(u_col_out_107),
    .col_out_108(u_col_out_108),
    .col_out_109(u_col_out_109),
    .col_out_110(u_col_out_110),
    .col_out_111(u_col_out_111),
    .col_out_112(u_col_out_112),
    .col_out_113(u_col_out_113),
    .col_out_114(u_col_out_114),
    .col_out_115(u_col_out_115),
    .col_out_116(u_col_out_116),
    .col_out_117(u_col_out_117),
    .col_out_118(u_col_out_118),
    .col_out_119(u_col_out_119),
    .col_out_120(u_col_out_120),
    .col_out_121(u_col_out_121),
    .col_out_122(u_col_out_122),
    .col_out_123(u_col_out_123),
    .col_out_124(u_col_out_124),
    .col_out_125(u_col_out_125),
    .col_out_126(u_col_out_126),
    .col_out_127(u_col_out_127),
    .col_out_128(u_col_out_128),
    .col_out_129(u_col_out_129),
    .col_out_130(u_col_out_130),
    .col_out_131(u_col_out_131),
    .col_out_132(u_col_out_132),
    .col_out_133(u_col_out_133),
    .col_out_134(u_col_out_134),
    .col_out_135(u_col_out_135),
    .col_out_136(u_col_out_136),
    .col_out_137(u_col_out_137),
    .col_out_138(u_col_out_138),
    .col_out_139(u_col_out_139),
    .col_out_140(u_col_out_140),
    .col_out_141(u_col_out_141),
    .col_out_142(u_col_out_142),
    .col_out_143(u_col_out_143),
    .col_out_144(u_col_out_144),
    .col_out_145(u_col_out_145),
    .col_out_146(u_col_out_146),
    .col_out_147(u_col_out_147),
    .col_out_148(u_col_out_148),
    .col_out_149(u_col_out_149),
    .col_out_150(u_col_out_150),
    .col_out_151(u_col_out_151),
    .col_out_152(u_col_out_152),
    .col_out_153(u_col_out_153),
    .col_out_154(u_col_out_154),
    .col_out_155(u_col_out_155),
    .col_out_156(u_col_out_156),
    .col_out_157(u_col_out_157),
    .col_out_158(u_col_out_158),
    .col_out_159(u_col_out_159),
    .col_out_160(u_col_out_160),
    .col_out_161(u_col_out_161),
    .col_out_162(u_col_out_162),
    .col_out_163(u_col_out_163),
    .col_out_164(u_col_out_164),
    .col_out_165(u_col_out_165),
    .col_out_166(u_col_out_166),
    .col_out_167(u_col_out_167),
    .col_out_168(u_col_out_168),
    .col_out_169(u_col_out_169),
    .col_out_170(u_col_out_170),
    .col_out_171(u_col_out_171),
    .col_out_172(u_col_out_172),
    .col_out_173(u_col_out_173),
    .col_out_174(u_col_out_174),
    .col_out_175(u_col_out_175),
    .col_out_176(u_col_out_176),
    .col_out_177(u_col_out_177),
    .col_out_178(u_col_out_178),
    .col_out_179(u_col_out_179),
    .col_out_180(u_col_out_180),
    .col_out_181(u_col_out_181),
    .col_out_182(u_col_out_182),
    .col_out_183(u_col_out_183),
    .col_out_184(u_col_out_184),
    .col_out_185(u_col_out_185),
    .col_out_186(u_col_out_186),
    .col_out_187(u_col_out_187),
    .col_out_188(u_col_out_188),
    .col_out_189(u_col_out_189),
    .col_out_190(u_col_out_190),
    .col_out_191(u_col_out_191),
    .col_out_192(u_col_out_192),
    .col_out_193(u_col_out_193),
    .col_out_194(u_col_out_194),
    .col_out_195(u_col_out_195),
    .col_out_196(u_col_out_196),
    .col_out_197(u_col_out_197),
    .col_out_198(u_col_out_198),
    .col_out_199(u_col_out_199),
    .col_out_200(u_col_out_200),
    .col_out_201(u_col_out_201),
    .col_out_202(u_col_out_202),
    .col_out_203(u_col_out_203),
    .col_out_204(u_col_out_204),
    .col_out_205(u_col_out_205),
    .col_out_206(u_col_out_206),
    .col_out_207(u_col_out_207),
    .col_out_208(u_col_out_208),
    .col_out_209(u_col_out_209),
    .col_out_210(u_col_out_210),
    .col_out_211(u_col_out_211),
    .col_out_212(u_col_out_212),
    .col_out_213(u_col_out_213),
    .col_out_214(u_col_out_214),
    .col_out_215(u_col_out_215),
    .col_out_216(u_col_out_216),
    .col_out_217(u_col_out_217),
    .col_out_218(u_col_out_218),
    .col_out_219(u_col_out_219),
    .col_out_220(u_col_out_220),
    .col_out_221(u_col_out_221),
    .col_out_222(u_col_out_222),
    .col_out_223(u_col_out_223),
    .col_out_224(u_col_out_224),
    .col_out_225(u_col_out_225),
    .col_out_226(u_col_out_226),
    .col_out_227(u_col_out_227),
    .col_out_228(u_col_out_228),
    .col_out_229(u_col_out_229),
    .col_out_230(u_col_out_230),
    .col_out_231(u_col_out_231),
    .col_out_232(u_col_out_232),
    .col_out_233(u_col_out_233),
    .col_out_234(u_col_out_234),
    .col_out_235(u_col_out_235),
    .col_out_236(u_col_out_236),
    .col_out_237(u_col_out_237),
    .col_out_238(u_col_out_238),
    .col_out_239(u_col_out_239),
    .col_out_240(u_col_out_240),
    .col_out_241(u_col_out_241),
    .col_out_242(u_col_out_242),
    .col_out_243(u_col_out_243),
    .col_out_244(u_col_out_244),
    .col_out_245(u_col_out_245),
    .col_out_246(u_col_out_246),
    .col_out_247(u_col_out_247),
    .col_out_248(u_col_out_248),
    .col_out_249(u_col_out_249),
    .col_out_250(u_col_out_250),
    .col_out_251(u_col_out_251),
    .col_out_252(u_col_out_252),
    .col_out_253(u_col_out_253),
    .col_out_254(u_col_out_254),
    .col_out_255(u_col_out_255),
    .col_out_256(u_col_out_256),
    .col_out_257(u_col_out_257),
    .col_out_258(u_col_out_258),
    .col_out_259(u_col_out_259),
    .col_out_260(u_col_out_260),
    .col_out_261(u_col_out_261),
    .col_out_262(u_col_out_262),
    .col_out_263(u_col_out_263),
    .col_out_264(u_col_out_264),
    .col_out_265(u_col_out_265),
    .col_out_266(u_col_out_266),
    .col_out_267(u_col_out_267),
    .col_out_268(u_col_out_268),
    .col_out_269(u_col_out_269),
    .col_out_270(u_col_out_270),
    .col_out_271(u_col_out_271),
    .col_out_272(u_col_out_272),
    .col_out_273(u_col_out_273),
    .col_out_274(u_col_out_274),
    .col_out_275(u_col_out_275),
    .col_out_276(u_col_out_276),
    .col_out_277(u_col_out_277),
    .col_out_278(u_col_out_278),
    .col_out_279(u_col_out_279),
    .col_out_280(u_col_out_280),
    .col_out_281(u_col_out_281),
    .col_out_282(u_col_out_282),
    .col_out_283(u_col_out_283),
    .col_out_284(u_col_out_284),
    .col_out_285(u_col_out_285),
    .col_out_286(u_col_out_286),
    .col_out_287(u_col_out_287),
    .col_out_288(u_col_out_288),
    .col_out_289(u_col_out_289),
    .col_out_290(u_col_out_290),
    .col_out_291(u_col_out_291),
    .col_out_292(u_col_out_292),
    .col_out_293(u_col_out_293),
    .col_out_294(u_col_out_294),
    .col_out_295(u_col_out_295),
    .col_out_296(u_col_out_296),
    .col_out_297(u_col_out_297),
    .col_out_298(u_col_out_298),
    .col_out_299(u_col_out_299),
    .col_out_300(u_col_out_300),
    .col_out_301(u_col_out_301),
    .col_out_302(u_col_out_302),
    .col_out_303(u_col_out_303),
    .col_out_304(u_col_out_304),
    .col_out_305(u_col_out_305),
    .col_out_306(u_col_out_306),
    .col_out_307(u_col_out_307),
    .col_out_308(u_col_out_308),
    .col_out_309(u_col_out_309),
    .col_out_310(u_col_out_310),
    .col_out_311(u_col_out_311),
    .col_out_312(u_col_out_312),
    .col_out_313(u_col_out_313),
    .col_out_314(u_col_out_314),
    .col_out_315(u_col_out_315),
    .col_out_316(u_col_out_316),
    .col_out_317(u_col_out_317),
    .col_out_318(u_col_out_318),
    .col_out_319(u_col_out_319),
    .col_out_320(u_col_out_320),
    .col_out_321(u_col_out_321),
    .col_out_322(u_col_out_322),
    .col_out_323(u_col_out_323),
    .col_out_324(u_col_out_324),
    .col_out_325(u_col_out_325),
    .col_out_326(u_col_out_326),
    .col_out_327(u_col_out_327),
    .col_out_328(u_col_out_328),
    .col_out_329(u_col_out_329),
    .col_out_330(u_col_out_330),
    .col_out_331(u_col_out_331),
    .col_out_332(u_col_out_332),
    .col_out_333(u_col_out_333),
    .col_out_334(u_col_out_334),
    .col_out_335(u_col_out_335),
    .col_out_336(u_col_out_336),
    .col_out_337(u_col_out_337),
    .col_out_338(u_col_out_338),
    .col_out_339(u_col_out_339),
    .col_out_340(u_col_out_340),
    .col_out_341(u_col_out_341),
    .col_out_342(u_col_out_342),
    .col_out_343(u_col_out_343),
    .col_out_344(u_col_out_344),
    .col_out_345(u_col_out_345),
    .col_out_346(u_col_out_346),
    .col_out_347(u_col_out_347),
    .col_out_348(u_col_out_348),
    .col_out_349(u_col_out_349),
    .col_out_350(u_col_out_350),
    .col_out_351(u_col_out_351),
    .col_out_352(u_col_out_352),
    .col_out_353(u_col_out_353),
    .col_out_354(u_col_out_354),
    .col_out_355(u_col_out_355),
    .col_out_356(u_col_out_356),
    .col_out_357(u_col_out_357),
    .col_out_358(u_col_out_358),
    .col_out_359(u_col_out_359),
    .col_out_360(u_col_out_360),
    .col_out_361(u_col_out_361),
    .col_out_362(u_col_out_362),
    .col_out_363(u_col_out_363),
    .col_out_364(u_col_out_364),
    .col_out_365(u_col_out_365),
    .col_out_366(u_col_out_366),
    .col_out_367(u_col_out_367),
    .col_out_368(u_col_out_368),
    .col_out_369(u_col_out_369),
    .col_out_370(u_col_out_370),
    .col_out_371(u_col_out_371),
    .col_out_372(u_col_out_372),
    .col_out_373(u_col_out_373),
    .col_out_374(u_col_out_374),
    .col_out_375(u_col_out_375),
    .col_out_376(u_col_out_376),
    .col_out_377(u_col_out_377),
    .col_out_378(u_col_out_378),
    .col_out_379(u_col_out_379),
    .col_out_380(u_col_out_380),
    .col_out_381(u_col_out_381),
    .col_out_382(u_col_out_382),
    .col_out_383(u_col_out_383),
    .col_out_384(u_col_out_384),
    .col_out_385(u_col_out_385),
    .col_out_386(u_col_out_386),
    .col_out_387(u_col_out_387),
    .col_out_388(u_col_out_388),
    .col_out_389(u_col_out_389),
    .col_out_390(u_col_out_390),
    .col_out_391(u_col_out_391),
    .col_out_392(u_col_out_392),
    .col_out_393(u_col_out_393),
    .col_out_394(u_col_out_394),
    .col_out_395(u_col_out_395),
    .col_out_396(u_col_out_396),
    .col_out_397(u_col_out_397),
    .col_out_398(u_col_out_398),
    .col_out_399(u_col_out_399),
    .col_out_400(u_col_out_400),
    .col_out_401(u_col_out_401),
    .col_out_402(u_col_out_402),
    .col_out_403(u_col_out_403),
    .col_out_404(u_col_out_404),
    .col_out_405(u_col_out_405),
    .col_out_406(u_col_out_406),
    .col_out_407(u_col_out_407),
    .col_out_408(u_col_out_408),
    .col_out_409(u_col_out_409),
    .col_out_410(u_col_out_410),
    .col_out_411(u_col_out_411),
    .col_out_412(u_col_out_412),
    .col_out_413(u_col_out_413),
    .col_out_414(u_col_out_414),
    .col_out_415(u_col_out_415),
    .col_out_416(u_col_out_416),
    .col_out_417(u_col_out_417),
    .col_out_418(u_col_out_418),
    .col_out_419(u_col_out_419),
    .col_out_420(u_col_out_420),
    .col_out_421(u_col_out_421),
    .col_out_422(u_col_out_422),
    .col_out_423(u_col_out_423),
    .col_out_424(u_col_out_424),
    .col_out_425(u_col_out_425),
    .col_out_426(u_col_out_426),
    .col_out_427(u_col_out_427),
    .col_out_428(u_col_out_428),
    .col_out_429(u_col_out_429),
    .col_out_430(u_col_out_430),
    .col_out_431(u_col_out_431),
    .col_out_432(u_col_out_432),
    .col_out_433(u_col_out_433),
    .col_out_434(u_col_out_434),
    .col_out_435(u_col_out_435),
    .col_out_436(u_col_out_436),
    .col_out_437(u_col_out_437),
    .col_out_438(u_col_out_438),
    .col_out_439(u_col_out_439),
    .col_out_440(u_col_out_440),
    .col_out_441(u_col_out_441),
    .col_out_442(u_col_out_442),
    .col_out_443(u_col_out_443),
    .col_out_444(u_col_out_444),
    .col_out_445(u_col_out_445),
    .col_out_446(u_col_out_446),
    .col_out_447(u_col_out_447),
    .col_out_448(u_col_out_448),
    .col_out_449(u_col_out_449),
    .col_out_450(u_col_out_450),
    .col_out_451(u_col_out_451),
    .col_out_452(u_col_out_452),
    .col_out_453(u_col_out_453),
    .col_out_454(u_col_out_454),
    .col_out_455(u_col_out_455),
    .col_out_456(u_col_out_456),
    .col_out_457(u_col_out_457),
    .col_out_458(u_col_out_458),
    .col_out_459(u_col_out_459),
    .col_out_460(u_col_out_460),
    .col_out_461(u_col_out_461),
    .col_out_462(u_col_out_462),
    .col_out_463(u_col_out_463),
    .col_out_464(u_col_out_464),
    .col_out_465(u_col_out_465),
    .col_out_466(u_col_out_466),
    .col_out_467(u_col_out_467),
    .col_out_468(u_col_out_468),
    .col_out_469(u_col_out_469),
    .col_out_470(u_col_out_470),
    .col_out_471(u_col_out_471),
    .col_out_472(u_col_out_472),
    .col_out_473(u_col_out_473),
    .col_out_474(u_col_out_474),
    .col_out_475(u_col_out_475),
    .col_out_476(u_col_out_476),
    .col_out_477(u_col_out_477),
    .col_out_478(u_col_out_478),
    .col_out_479(u_col_out_479),
    .col_out_480(u_col_out_480),
    .col_out_481(u_col_out_481),
    .col_out_482(u_col_out_482),
    .col_out_483(u_col_out_483),
    .col_out_484(u_col_out_484),
    .col_out_485(u_col_out_485),
    .col_out_486(u_col_out_486),
    .col_out_487(u_col_out_487),
    .col_out_488(u_col_out_488),
    .col_out_489(u_col_out_489),
    .col_out_490(u_col_out_490),
    .col_out_491(u_col_out_491),
    .col_out_492(u_col_out_492),
    .col_out_493(u_col_out_493),
    .col_out_494(u_col_out_494),
    .col_out_495(u_col_out_495),
    .col_out_496(u_col_out_496),
    .col_out_497(u_col_out_497),
    .col_out_498(u_col_out_498),
    .col_out_499(u_col_out_499),
    .col_out_500(u_col_out_500),
    .col_out_501(u_col_out_501),
    .col_out_502(u_col_out_502),
    .col_out_503(u_col_out_503),
    .col_out_504(u_col_out_504),
    .col_out_505(u_col_out_505),
    .col_out_506(u_col_out_506),
    .col_out_507(u_col_out_507),
    .col_out_508(u_col_out_508),
    .col_out_509(u_col_out_509),
    .col_out_510(u_col_out_510),
    .col_out_511(u_col_out_511),
    .col_out_512(u_col_out_512),
    .col_out_513(u_col_out_513),
    .col_out_514(u_col_out_514),
    .col_out_515(u_col_out_515),
    .col_out_516(u_col_out_516),
    .col_out_517(u_col_out_517),
    .col_out_518(u_col_out_518),
    .col_out_519(u_col_out_519),
    .col_out_520(u_col_out_520),
    .col_out_521(u_col_out_521),
    .col_out_522(u_col_out_522),
    .col_out_523(u_col_out_523),
    .col_out_524(u_col_out_524),
    .col_out_525(u_col_out_525),
    .col_out_526(u_col_out_526),
    .col_out_527(u_col_out_527),
    .col_out_528(u_col_out_528),
    .col_out_529(u_col_out_529),
    .col_out_530(u_col_out_530),
    .col_out_531(u_col_out_531),
    .col_out_532(u_col_out_532),
    .col_out_533(u_col_out_533),
    .col_out_534(u_col_out_534),
    .col_out_535(u_col_out_535),
    .col_out_536(u_col_out_536),
    .col_out_537(u_col_out_537),
    .col_out_538(u_col_out_538),
    .col_out_539(u_col_out_539),
    .col_out_540(u_col_out_540),
    .col_out_541(u_col_out_541),
    .col_out_542(u_col_out_542),
    .col_out_543(u_col_out_543),
    .col_out_544(u_col_out_544),
    .col_out_545(u_col_out_545),
    .col_out_546(u_col_out_546),
    .col_out_547(u_col_out_547),
    .col_out_548(u_col_out_548),
    .col_out_549(u_col_out_549),
    .col_out_550(u_col_out_550),
    .col_out_551(u_col_out_551),
    .col_out_552(u_col_out_552),
    .col_out_553(u_col_out_553),
    .col_out_554(u_col_out_554),
    .col_out_555(u_col_out_555),
    .col_out_556(u_col_out_556),
    .col_out_557(u_col_out_557),
    .col_out_558(u_col_out_558),
    .col_out_559(u_col_out_559),
    .col_out_560(u_col_out_560),
    .col_out_561(u_col_out_561),
    .col_out_562(u_col_out_562),
    .col_out_563(u_col_out_563),
    .col_out_564(u_col_out_564),
    .col_out_565(u_col_out_565),
    .col_out_566(u_col_out_566),
    .col_out_567(u_col_out_567),
    .col_out_568(u_col_out_568),
    .col_out_569(u_col_out_569),
    .col_out_570(u_col_out_570),
    .col_out_571(u_col_out_571),
    .col_out_572(u_col_out_572),
    .col_out_573(u_col_out_573),
    .col_out_574(u_col_out_574),
    .col_out_575(u_col_out_575),
    .col_out_576(u_col_out_576),
    .col_out_577(u_col_out_577),
    .col_out_578(u_col_out_578),
    .col_out_579(u_col_out_579),
    .col_out_580(u_col_out_580),
    .col_out_581(u_col_out_581),
    .col_out_582(u_col_out_582),
    .col_out_583(u_col_out_583),
    .col_out_584(u_col_out_584),
    .col_out_585(u_col_out_585),
    .col_out_586(u_col_out_586),
    .col_out_587(u_col_out_587),
    .col_out_588(u_col_out_588),
    .col_out_589(u_col_out_589),
    .col_out_590(u_col_out_590),
    .col_out_591(u_col_out_591),
    .col_out_592(u_col_out_592),
    .col_out_593(u_col_out_593),
    .col_out_594(u_col_out_594),
    .col_out_595(u_col_out_595),
    .col_out_596(u_col_out_596),
    .col_out_597(u_col_out_597),
    .col_out_598(u_col_out_598),
    .col_out_599(u_col_out_599),
    .col_out_600(u_col_out_600),
    .col_out_601(u_col_out_601),
    .col_out_602(u_col_out_602),
    .col_out_603(u_col_out_603),
    .col_out_604(u_col_out_604),
    .col_out_605(u_col_out_605),
    .col_out_606(u_col_out_606),
    .col_out_607(u_col_out_607),
    .col_out_608(u_col_out_608),
    .col_out_609(u_col_out_609),
    .col_out_610(u_col_out_610),
    .col_out_611(u_col_out_611),
    .col_out_612(u_col_out_612),
    .col_out_613(u_col_out_613),
    .col_out_614(u_col_out_614),
    .col_out_615(u_col_out_615),
    .col_out_616(u_col_out_616),
    .col_out_617(u_col_out_617),
    .col_out_618(u_col_out_618),
    .col_out_619(u_col_out_619),
    .col_out_620(u_col_out_620),
    .col_out_621(u_col_out_621),
    .col_out_622(u_col_out_622),
    .col_out_623(u_col_out_623),
    .col_out_624(u_col_out_624),
    .col_out_625(u_col_out_625),
    .col_out_626(u_col_out_626),
    .col_out_627(u_col_out_627),
    .col_out_628(u_col_out_628),
    .col_out_629(u_col_out_629),
    .col_out_630(u_col_out_630),
    .col_out_631(u_col_out_631),
    .col_out_632(u_col_out_632),
    .col_out_633(u_col_out_633),
    .col_out_634(u_col_out_634),
    .col_out_635(u_col_out_635),
    .col_out_636(u_col_out_636),
    .col_out_637(u_col_out_637),
    .col_out_638(u_col_out_638),
    .col_out_639(u_col_out_639),
    .col_out_640(u_col_out_640),
    .col_out_641(u_col_out_641),
    .col_out_642(u_col_out_642),
    .col_out_643(u_col_out_643),
    .col_out_644(u_col_out_644),
    .col_out_645(u_col_out_645),
    .col_out_646(u_col_out_646),
    .col_out_647(u_col_out_647),
    .col_out_648(u_col_out_648),
    .col_out_649(u_col_out_649),
    .col_out_650(u_col_out_650),
    .col_out_651(u_col_out_651),
    .col_out_652(u_col_out_652),
    .col_out_653(u_col_out_653),
    .col_out_654(u_col_out_654),
    .col_out_655(u_col_out_655),
    .col_out_656(u_col_out_656),
    .col_out_657(u_col_out_657),
    .col_out_658(u_col_out_658),
    .col_out_659(u_col_out_659),
    .col_out_660(u_col_out_660),
    .col_out_661(u_col_out_661),
    .col_out_662(u_col_out_662),
    .col_out_663(u_col_out_663),
    .col_out_664(u_col_out_664),
    .col_out_665(u_col_out_665),
    .col_out_666(u_col_out_666),
    .col_out_667(u_col_out_667),
    .col_out_668(u_col_out_668),
    .col_out_669(u_col_out_669),
    .col_out_670(u_col_out_670),
    .col_out_671(u_col_out_671),
    .col_out_672(u_col_out_672),
    .col_out_673(u_col_out_673),
    .col_out_674(u_col_out_674),
    .col_out_675(u_col_out_675),
    .col_out_676(u_col_out_676),
    .col_out_677(u_col_out_677),
    .col_out_678(u_col_out_678),
    .col_out_679(u_col_out_679),
    .col_out_680(u_col_out_680),
    .col_out_681(u_col_out_681),
    .col_out_682(u_col_out_682),
    .col_out_683(u_col_out_683),
    .col_out_684(u_col_out_684),
    .col_out_685(u_col_out_685),
    .col_out_686(u_col_out_686),
    .col_out_687(u_col_out_687),
    .col_out_688(u_col_out_688),
    .col_out_689(u_col_out_689),
    .col_out_690(u_col_out_690),
    .col_out_691(u_col_out_691),
    .col_out_692(u_col_out_692),
    .col_out_693(u_col_out_693),
    .col_out_694(u_col_out_694),
    .col_out_695(u_col_out_695),
    .col_out_696(u_col_out_696),
    .col_out_697(u_col_out_697),
    .col_out_698(u_col_out_698),
    .col_out_699(u_col_out_699),
    .col_out_700(u_col_out_700),
    .col_out_701(u_col_out_701),
    .col_out_702(u_col_out_702),
    .col_out_703(u_col_out_703),
    .col_out_704(u_col_out_704),
    .col_out_705(u_col_out_705),
    .col_out_706(u_col_out_706),
    .col_out_707(u_col_out_707),
    .col_out_708(u_col_out_708),
    .col_out_709(u_col_out_709),
    .col_out_710(u_col_out_710),
    .col_out_711(u_col_out_711),
    .col_out_712(u_col_out_712),
    .col_out_713(u_col_out_713),
    .col_out_714(u_col_out_714),
    .col_out_715(u_col_out_715),
    .col_out_716(u_col_out_716),
    .col_out_717(u_col_out_717),
    .col_out_718(u_col_out_718),
    .col_out_719(u_col_out_719),
    .col_out_720(u_col_out_720),
    .col_out_721(u_col_out_721),
    .col_out_722(u_col_out_722),
    .col_out_723(u_col_out_723),
    .col_out_724(u_col_out_724),
    .col_out_725(u_col_out_725),
    .col_out_726(u_col_out_726),
    .col_out_727(u_col_out_727),
    .col_out_728(u_col_out_728),
    .col_out_729(u_col_out_729),
    .col_out_730(u_col_out_730),
    .col_out_731(u_col_out_731),
    .col_out_732(u_col_out_732),
    .col_out_733(u_col_out_733),
    .col_out_734(u_col_out_734),
    .col_out_735(u_col_out_735),
    .col_out_736(u_col_out_736),
    .col_out_737(u_col_out_737),
    .col_out_738(u_col_out_738),
    .col_out_739(u_col_out_739),
    .col_out_740(u_col_out_740),
    .col_out_741(u_col_out_741),
    .col_out_742(u_col_out_742),
    .col_out_743(u_col_out_743),
    .col_out_744(u_col_out_744),
    .col_out_745(u_col_out_745),
    .col_out_746(u_col_out_746),
    .col_out_747(u_col_out_747),
    .col_out_748(u_col_out_748),
    .col_out_749(u_col_out_749),
    .col_out_750(u_col_out_750),
    .col_out_751(u_col_out_751),
    .col_out_752(u_col_out_752),
    .col_out_753(u_col_out_753),
    .col_out_754(u_col_out_754),
    .col_out_755(u_col_out_755),
    .col_out_756(u_col_out_756),
    .col_out_757(u_col_out_757),
    .col_out_758(u_col_out_758),
    .col_out_759(u_col_out_759),
    .col_out_760(u_col_out_760),
    .col_out_761(u_col_out_761),
    .col_out_762(u_col_out_762),
    .col_out_763(u_col_out_763),
    .col_out_764(u_col_out_764),
    .col_out_765(u_col_out_765),
    .col_out_766(u_col_out_766),
    .col_out_767(u_col_out_767),
    .col_out_768(u_col_out_768),
    .col_out_769(u_col_out_769),
    .col_out_770(u_col_out_770),
    .col_out_771(u_col_out_771),
    .col_out_772(u_col_out_772),
    .col_out_773(u_col_out_773),
    .col_out_774(u_col_out_774),
    .col_out_775(u_col_out_775),
    .col_out_776(u_col_out_776),
    .col_out_777(u_col_out_777),
    .col_out_778(u_col_out_778),
    .col_out_779(u_col_out_779),
    .col_out_780(u_col_out_780),
    .col_out_781(u_col_out_781),
    .col_out_782(u_col_out_782),
    .col_out_783(u_col_out_783),
    .col_out_784(u_col_out_784),
    .col_out_785(u_col_out_785),
    .col_out_786(u_col_out_786),
    .col_out_787(u_col_out_787),
    .col_out_788(u_col_out_788),
    .col_out_789(u_col_out_789),
    .col_out_790(u_col_out_790),
    .col_out_791(u_col_out_791),
    .col_out_792(u_col_out_792),
    .col_out_793(u_col_out_793),
    .col_out_794(u_col_out_794),
    .col_out_795(u_col_out_795),
    .col_out_796(u_col_out_796),
    .col_out_797(u_col_out_797),
    .col_out_798(u_col_out_798),
    .col_out_799(u_col_out_799),
    .col_out_800(u_col_out_800),
    .col_out_801(u_col_out_801),
    .col_out_802(u_col_out_802),
    .col_out_803(u_col_out_803),
    .col_out_804(u_col_out_804),
    .col_out_805(u_col_out_805),
    .col_out_806(u_col_out_806),
    .col_out_807(u_col_out_807),
    .col_out_808(u_col_out_808),
    .col_out_809(u_col_out_809),
    .col_out_810(u_col_out_810),
    .col_out_811(u_col_out_811),
    .col_out_812(u_col_out_812),
    .col_out_813(u_col_out_813),
    .col_out_814(u_col_out_814),
    .col_out_815(u_col_out_815),
    .col_out_816(u_col_out_816),
    .col_out_817(u_col_out_817),
    .col_out_818(u_col_out_818),
    .col_out_819(u_col_out_819),
    .col_out_820(u_col_out_820),
    .col_out_821(u_col_out_821),
    .col_out_822(u_col_out_822),
    .col_out_823(u_col_out_823),
    .col_out_824(u_col_out_824),
    .col_out_825(u_col_out_825),
    .col_out_826(u_col_out_826),
    .col_out_827(u_col_out_827),
    .col_out_828(u_col_out_828),
    .col_out_829(u_col_out_829),
    .col_out_830(u_col_out_830),
    .col_out_831(u_col_out_831),
    .col_out_832(u_col_out_832),
    .col_out_833(u_col_out_833),
    .col_out_834(u_col_out_834),
    .col_out_835(u_col_out_835),
    .col_out_836(u_col_out_836),
    .col_out_837(u_col_out_837),
    .col_out_838(u_col_out_838),
    .col_out_839(u_col_out_839),
    .col_out_840(u_col_out_840),
    .col_out_841(u_col_out_841),
    .col_out_842(u_col_out_842),
    .col_out_843(u_col_out_843),
    .col_out_844(u_col_out_844),
    .col_out_845(u_col_out_845),
    .col_out_846(u_col_out_846),
    .col_out_847(u_col_out_847),
    .col_out_848(u_col_out_848),
    .col_out_849(u_col_out_849),
    .col_out_850(u_col_out_850),
    .col_out_851(u_col_out_851),
    .col_out_852(u_col_out_852),
    .col_out_853(u_col_out_853),
    .col_out_854(u_col_out_854),
    .col_out_855(u_col_out_855),
    .col_out_856(u_col_out_856),
    .col_out_857(u_col_out_857),
    .col_out_858(u_col_out_858),
    .col_out_859(u_col_out_859),
    .col_out_860(u_col_out_860),
    .col_out_861(u_col_out_861),
    .col_out_862(u_col_out_862),
    .col_out_863(u_col_out_863),
    .col_out_864(u_col_out_864),
    .col_out_865(u_col_out_865),
    .col_out_866(u_col_out_866),
    .col_out_867(u_col_out_867),
    .col_out_868(u_col_out_868),
    .col_out_869(u_col_out_869),
    .col_out_870(u_col_out_870),
    .col_out_871(u_col_out_871),
    .col_out_872(u_col_out_872),
    .col_out_873(u_col_out_873),
    .col_out_874(u_col_out_874),
    .col_out_875(u_col_out_875),
    .col_out_876(u_col_out_876),
    .col_out_877(u_col_out_877),
    .col_out_878(u_col_out_878),
    .col_out_879(u_col_out_879),
    .col_out_880(u_col_out_880),
    .col_out_881(u_col_out_881),
    .col_out_882(u_col_out_882),
    .col_out_883(u_col_out_883),
    .col_out_884(u_col_out_884),
    .col_out_885(u_col_out_885),
    .col_out_886(u_col_out_886),
    .col_out_887(u_col_out_887),
    .col_out_888(u_col_out_888),
    .col_out_889(u_col_out_889),
    .col_out_890(u_col_out_890),
    .col_out_891(u_col_out_891),
    .col_out_892(u_col_out_892),
    .col_out_893(u_col_out_893),
    .col_out_894(u_col_out_894),
    .col_out_895(u_col_out_895),
    .col_out_896(u_col_out_896),
    .col_out_897(u_col_out_897),
    .col_out_898(u_col_out_898),
    .col_out_899(u_col_out_899),
    .col_out_900(u_col_out_900),
    .col_out_901(u_col_out_901),
    .col_out_902(u_col_out_902),
    .col_out_903(u_col_out_903),
    .col_out_904(u_col_out_904),
    .col_out_905(u_col_out_905),
    .col_out_906(u_col_out_906),
    .col_out_907(u_col_out_907),
    .col_out_908(u_col_out_908),
    .col_out_909(u_col_out_909),
    .col_out_910(u_col_out_910),
    .col_out_911(u_col_out_911),
    .col_out_912(u_col_out_912),
    .col_out_913(u_col_out_913),
    .col_out_914(u_col_out_914),
    .col_out_915(u_col_out_915),
    .col_out_916(u_col_out_916),
    .col_out_917(u_col_out_917),
    .col_out_918(u_col_out_918),
    .col_out_919(u_col_out_919),
    .col_out_920(u_col_out_920),
    .col_out_921(u_col_out_921),
    .col_out_922(u_col_out_922),
    .col_out_923(u_col_out_923),
    .col_out_924(u_col_out_924),
    .col_out_925(u_col_out_925),
    .col_out_926(u_col_out_926),
    .col_out_927(u_col_out_927),
    .col_out_928(u_col_out_928),
    .col_out_929(u_col_out_929),
    .col_out_930(u_col_out_930),
    .col_out_931(u_col_out_931),
    .col_out_932(u_col_out_932),
    .col_out_933(u_col_out_933),
    .col_out_934(u_col_out_934),
    .col_out_935(u_col_out_935),
    .col_out_936(u_col_out_936),
    .col_out_937(u_col_out_937),
    .col_out_938(u_col_out_938),
    .col_out_939(u_col_out_939),
    .col_out_940(u_col_out_940),
    .col_out_941(u_col_out_941),
    .col_out_942(u_col_out_942),
    .col_out_943(u_col_out_943),
    .col_out_944(u_col_out_944),
    .col_out_945(u_col_out_945),
    .col_out_946(u_col_out_946),
    .col_out_947(u_col_out_947),
    .col_out_948(u_col_out_948),
    .col_out_949(u_col_out_949),
    .col_out_950(u_col_out_950),
    .col_out_951(u_col_out_951),
    .col_out_952(u_col_out_952),
    .col_out_953(u_col_out_953),
    .col_out_954(u_col_out_954),
    .col_out_955(u_col_out_955),
    .col_out_956(u_col_out_956),
    .col_out_957(u_col_out_957),
    .col_out_958(u_col_out_958),
    .col_out_959(u_col_out_959),
    .col_out_960(u_col_out_960),
    .col_out_961(u_col_out_961),
    .col_out_962(u_col_out_962),
    .col_out_963(u_col_out_963),
    .col_out_964(u_col_out_964),
    .col_out_965(u_col_out_965),
    .col_out_966(u_col_out_966),
    .col_out_967(u_col_out_967),
    .col_out_968(u_col_out_968),
    .col_out_969(u_col_out_969),
    .col_out_970(u_col_out_970),
    .col_out_971(u_col_out_971),
    .col_out_972(u_col_out_972),
    .col_out_973(u_col_out_973),
    .col_out_974(u_col_out_974),
    .col_out_975(u_col_out_975),
    .col_out_976(u_col_out_976),
    .col_out_977(u_col_out_977),
    .col_out_978(u_col_out_978),
    .col_out_979(u_col_out_979),
    .col_out_980(u_col_out_980),
    .col_out_981(u_col_out_981),
    .col_out_982(u_col_out_982),
    .col_out_983(u_col_out_983),
    .col_out_984(u_col_out_984),
    .col_out_985(u_col_out_985),
    .col_out_986(u_col_out_986),
    .col_out_987(u_col_out_987),
    .col_out_988(u_col_out_988),
    .col_out_989(u_col_out_989),
    .col_out_990(u_col_out_990),
    .col_out_991(u_col_out_991),
    .col_out_992(u_col_out_992),
    .col_out_993(u_col_out_993),
    .col_out_994(u_col_out_994),
    .col_out_995(u_col_out_995),
    .col_out_996(u_col_out_996),
    .col_out_997(u_col_out_997),
    .col_out_998(u_col_out_998),
    .col_out_999(u_col_out_999),
    .col_out_1000(u_col_out_1000),
    .col_out_1001(u_col_out_1001),
    .col_out_1002(u_col_out_1002),
    .col_out_1003(u_col_out_1003),
    .col_out_1004(u_col_out_1004),
    .col_out_1005(u_col_out_1005),
    .col_out_1006(u_col_out_1006),
    .col_out_1007(u_col_out_1007),
    .col_out_1008(u_col_out_1008),
    .col_out_1009(u_col_out_1009),
    .col_out_1010(u_col_out_1010),
    .col_out_1011(u_col_out_1011),
    .col_out_1012(u_col_out_1012),
    .col_out_1013(u_col_out_1013),
    .col_out_1014(u_col_out_1014),
    .col_out_1015(u_col_out_1015),
    .col_out_1016(u_col_out_1016),
    .col_out_1017(u_col_out_1017),
    .col_out_1018(u_col_out_1018),
    .col_out_1019(u_col_out_1019),
    .col_out_1020(u_col_out_1020),
    .col_out_1021(u_col_out_1021),
    .col_out_1022(u_col_out_1022),
    .col_out_1023(u_col_out_1023),
    .col_out_1024(u_col_out_1024),
    .col_out_1025(u_col_out_1025),
    .col_out_1026(u_col_out_1026),
    .col_out_1027(u_col_out_1027),
    .col_out_1028(u_col_out_1028),
    .col_out_1029(u_col_out_1029),
    .col_out_1030(u_col_out_1030),
    .col_out_1031(u_col_out_1031),
    .col_out_1032(u_col_out_1032),
    .col_out_1033(u_col_out_1033),
    .col_out_1034(u_col_out_1034),
    .col_out_1035(u_col_out_1035),
    .col_out_1036(u_col_out_1036),
    .col_out_1037(u_col_out_1037),
    .col_out_1038(u_col_out_1038),
    .col_out_1039(u_col_out_1039),
    .col_out_1040(u_col_out_1040),
    .col_out_1041(u_col_out_1041),
    .col_out_1042(u_col_out_1042),
    .col_out_1043(u_col_out_1043),
    .col_out_1044(u_col_out_1044),
    .col_out_1045(u_col_out_1045),
    .col_out_1046(u_col_out_1046),
    .col_out_1047(u_col_out_1047),
    .col_out_1048(u_col_out_1048),
    .col_out_1049(u_col_out_1049),
    .col_out_1050(u_col_out_1050),
    .col_out_1051(u_col_out_1051),
    .col_out_1052(u_col_out_1052),
    .col_out_1053(u_col_out_1053),
    .col_out_1054(u_col_out_1054),
    .col_out_1055(u_col_out_1055),
    .col_out_1056(u_col_out_1056),
    .col_out_1057(u_col_out_1057),
    .col_out_1058(u_col_out_1058),
    .col_out_1059(u_col_out_1059),
    .col_out_1060(u_col_out_1060),
    .col_out_1061(u_col_out_1061),
    .col_out_1062(u_col_out_1062),
    .col_out_1063(u_col_out_1063),
    .col_out_1064(u_col_out_1064),
    .col_out_1065(u_col_out_1065),
    .col_out_1066(u_col_out_1066),
    .col_out_1067(u_col_out_1067),
    .col_out_1068(u_col_out_1068),
    .col_out_1069(u_col_out_1069),
    .col_out_1070(u_col_out_1070),
    .col_out_1071(u_col_out_1071),
    .col_out_1072(u_col_out_1072),
    .col_out_1073(u_col_out_1073),
    .col_out_1074(u_col_out_1074),
    .col_out_1075(u_col_out_1075),
    .col_out_1076(u_col_out_1076),
    .col_out_1077(u_col_out_1077),
    .col_out_1078(u_col_out_1078),
    .col_out_1079(u_col_out_1079),
    .col_out_1080(u_col_out_1080),
    .col_out_1081(u_col_out_1081),
    .col_out_1082(u_col_out_1082),
    .col_out_1083(u_col_out_1083),
    .col_out_1084(u_col_out_1084),
    .col_out_1085(u_col_out_1085),
    .col_out_1086(u_col_out_1086),
    .col_out_1087(u_col_out_1087),
    .col_out_1088(u_col_out_1088),
    .col_out_1089(u_col_out_1089),
    .col_out_1090(u_col_out_1090),
    .col_out_1091(u_col_out_1091),
    .col_out_1092(u_col_out_1092),
    .col_out_1093(u_col_out_1093),
    .col_out_1094(u_col_out_1094),
    .col_out_1095(u_col_out_1095),
    .col_out_1096(u_col_out_1096),
    .col_out_1097(u_col_out_1097),
    .col_out_1098(u_col_out_1098),
    .col_out_1099(u_col_out_1099),
    .col_out_1100(u_col_out_1100),
    .col_out_1101(u_col_out_1101),
    .col_out_1102(u_col_out_1102),
    .col_out_1103(u_col_out_1103),
    .col_out_1104(u_col_out_1104),
    .col_out_1105(u_col_out_1105),
    .col_out_1106(u_col_out_1106),
    .col_out_1107(u_col_out_1107),
    .col_out_1108(u_col_out_1108),
    .col_out_1109(u_col_out_1109),
    .col_out_1110(u_col_out_1110),
    .col_out_1111(u_col_out_1111),
    .col_out_1112(u_col_out_1112),
    .col_out_1113(u_col_out_1113),
    .col_out_1114(u_col_out_1114),
    .col_out_1115(u_col_out_1115),
    .col_out_1116(u_col_out_1116),
    .col_out_1117(u_col_out_1117),
    .col_out_1118(u_col_out_1118),
    .col_out_1119(u_col_out_1119),
    .col_out_1120(u_col_out_1120),
    .col_out_1121(u_col_out_1121),
    .col_out_1122(u_col_out_1122),
    .col_out_1123(u_col_out_1123),
    .col_out_1124(u_col_out_1124),
    .col_out_1125(u_col_out_1125),
    .col_out_1126(u_col_out_1126),
    .col_out_1127(u_col_out_1127),
    .col_out_1128(u_col_out_1128),
    .col_out_1129(u_col_out_1129),
    .col_out_1130(u_col_out_1130),
    .col_out_1131(u_col_out_1131),
    .col_out_1132(u_col_out_1132),
    .col_out_1133(u_col_out_1133),
    .col_out_1134(u_col_out_1134),
    .col_out_1135(u_col_out_1135),
    .col_out_1136(u_col_out_1136),
    .col_out_1137(u_col_out_1137),
    .col_out_1138(u_col_out_1138),
    .col_out_1139(u_col_out_1139),
    .col_out_1140(u_col_out_1140),
    .col_out_1141(u_col_out_1141),
    .col_out_1142(u_col_out_1142),
    .col_out_1143(u_col_out_1143),
    .col_out_1144(u_col_out_1144),
    .col_out_1145(u_col_out_1145),
    .col_out_1146(u_col_out_1146),
    .col_out_1147(u_col_out_1147),
    .col_out_1148(u_col_out_1148),
    .col_out_1149(u_col_out_1149),
    .col_out_1150(u_col_out_1150),
    .col_out_1151(u_col_out_1151),
    .col_out_1152(u_col_out_1152),
    .col_out_1153(u_col_out_1153),
    .col_out_1154(u_col_out_1154),
    .col_out_1155(u_col_out_1155),
    .col_out_1156(u_col_out_1156),
    .col_out_1157(u_col_out_1157),
    .col_out_1158(u_col_out_1158),
    .col_out_1159(u_col_out_1159),
    .col_out_1160(u_col_out_1160),
    .col_out_1161(u_col_out_1161),
    .col_out_1162(u_col_out_1162),
    .col_out_1163(u_col_out_1163),
    .col_out_1164(u_col_out_1164),
    .col_out_1165(u_col_out_1165),
    .col_out_1166(u_col_out_1166),
    .col_out_1167(u_col_out_1167),
    .col_out_1168(u_col_out_1168),
    .col_out_1169(u_col_out_1169),
    .col_out_1170(u_col_out_1170),
    .col_out_1171(u_col_out_1171),
    .col_out_1172(u_col_out_1172),
    .col_out_1173(u_col_out_1173),
    .col_out_1174(u_col_out_1174),
    .col_out_1175(u_col_out_1175),
    .col_out_1176(u_col_out_1176),
    .col_out_1177(u_col_out_1177),
    .col_out_1178(u_col_out_1178),
    .col_out_1179(u_col_out_1179),
    .col_out_1180(u_col_out_1180),
    .col_out_1181(u_col_out_1181),
    .col_out_1182(u_col_out_1182),
    .col_out_1183(u_col_out_1183),
    .col_out_1184(u_col_out_1184),
    .col_out_1185(u_col_out_1185),
    .col_out_1186(u_col_out_1186),
    .col_out_1187(u_col_out_1187),
    .col_out_1188(u_col_out_1188),
    .col_out_1189(u_col_out_1189),
    .col_out_1190(u_col_out_1190),
    .col_out_1191(u_col_out_1191),
    .col_out_1192(u_col_out_1192),
    .col_out_1193(u_col_out_1193),
    .col_out_1194(u_col_out_1194),
    .col_out_1195(u_col_out_1195),
    .col_out_1196(u_col_out_1196),
    .col_out_1197(u_col_out_1197),
    .col_out_1198(u_col_out_1198),
    .col_out_1199(u_col_out_1199),
    .col_out_1200(u_col_out_1200),
    .col_out_1201(u_col_out_1201),
    .col_out_1202(u_col_out_1202),
    .col_out_1203(u_col_out_1203),
    .col_out_1204(u_col_out_1204),
    .col_out_1205(u_col_out_1205),
    .col_out_1206(u_col_out_1206),
    .col_out_1207(u_col_out_1207),
    .col_out_1208(u_col_out_1208),
    .col_out_1209(u_col_out_1209),
    .col_out_1210(u_col_out_1210),
    .col_out_1211(u_col_out_1211),
    .col_out_1212(u_col_out_1212),
    .col_out_1213(u_col_out_1213),
    .col_out_1214(u_col_out_1214),
    .col_out_1215(u_col_out_1215),
    .col_out_1216(u_col_out_1216),
    .col_out_1217(u_col_out_1217),
    .col_out_1218(u_col_out_1218),
    .col_out_1219(u_col_out_1219),
    .col_out_1220(u_col_out_1220),
    .col_out_1221(u_col_out_1221),
    .col_out_1222(u_col_out_1222),
    .col_out_1223(u_col_out_1223),
    .col_out_1224(u_col_out_1224),
    .col_out_1225(u_col_out_1225),
    .col_out_1226(u_col_out_1226),
    .col_out_1227(u_col_out_1227),
    .col_out_1228(u_col_out_1228),
    .col_out_1229(u_col_out_1229),
    .col_out_1230(u_col_out_1230),
    .col_out_1231(u_col_out_1231),
    .col_out_1232(u_col_out_1232),
    .col_out_1233(u_col_out_1233),
    .col_out_1234(u_col_out_1234),
    .col_out_1235(u_col_out_1235),
    .col_out_1236(u_col_out_1236),
    .col_out_1237(u_col_out_1237),
    .col_out_1238(u_col_out_1238),
    .col_out_1239(u_col_out_1239),
    .col_out_1240(u_col_out_1240),
    .col_out_1241(u_col_out_1241),
    .col_out_1242(u_col_out_1242),
    .col_out_1243(u_col_out_1243),
    .col_out_1244(u_col_out_1244),
    .col_out_1245(u_col_out_1245),
    .col_out_1246(u_col_out_1246),
    .col_out_1247(u_col_out_1247),
    .col_out_1248(u_col_out_1248),
    .col_out_1249(u_col_out_1249),
    .col_out_1250(u_col_out_1250),
    .col_out_1251(u_col_out_1251),
    .col_out_1252(u_col_out_1252),
    .col_out_1253(u_col_out_1253),
    .col_out_1254(u_col_out_1254),
    .col_out_1255(u_col_out_1255),
    .col_out_1256(u_col_out_1256),
    .col_out_1257(u_col_out_1257),
    .col_out_1258(u_col_out_1258),
    .col_out_1259(u_col_out_1259),
    .col_out_1260(u_col_out_1260),
    .col_out_1261(u_col_out_1261),
    .col_out_1262(u_col_out_1262),
    .col_out_1263(u_col_out_1263),
    .col_out_1264(u_col_out_1264),
    .col_out_1265(u_col_out_1265),
    .col_out_1266(u_col_out_1266),
    .col_out_1267(u_col_out_1267),
    .col_out_1268(u_col_out_1268),
    .col_out_1269(u_col_out_1269),
    .col_out_1270(u_col_out_1270),
    .col_out_1271(u_col_out_1271),
    .col_out_1272(u_col_out_1272),
    .col_out_1273(u_col_out_1273),
    .col_out_1274(u_col_out_1274),
    .col_out_1275(u_col_out_1275),
    .col_out_1276(u_col_out_1276),
    .col_out_1277(u_col_out_1277),
    .col_out_1278(u_col_out_1278),
    .col_out_1279(u_col_out_1279),
    .col_out_1280(u_col_out_1280),
    .col_out_1281(u_col_out_1281),
    .col_out_1282(u_col_out_1282),
    .col_out_1283(u_col_out_1283),
    .col_out_1284(u_col_out_1284),
    .col_out_1285(u_col_out_1285),
    .col_out_1286(u_col_out_1286),
    .col_out_1287(u_col_out_1287)
);


assign row_out_0 = {u_col_out_1287[0], u_col_out_1286[0], u_col_out_1285[0], u_col_out_1284[0], u_col_out_1283[0], u_col_out_1282[0], u_col_out_1281[0], u_col_out_1280[0], u_col_out_1279[0], u_col_out_1278[0], u_col_out_1277[0], u_col_out_1276[0], u_col_out_1275[0], u_col_out_1274[0], u_col_out_1273[0], u_col_out_1272[0], u_col_out_1271[0], u_col_out_1270[0], u_col_out_1269[0], u_col_out_1268[0], u_col_out_1267[0], u_col_out_1266[0], u_col_out_1265[0], u_col_out_1264[0], u_col_out_1263[0], u_col_out_1262[0], u_col_out_1261[0], u_col_out_1260[0], u_col_out_1259[0], u_col_out_1258[0], u_col_out_1257[0], u_col_out_1256[0], u_col_out_1255[0], u_col_out_1254[0], u_col_out_1253[0], u_col_out_1252[0], u_col_out_1251[0], u_col_out_1250[0], u_col_out_1249[0], u_col_out_1248[0], u_col_out_1247[0], u_col_out_1246[0], u_col_out_1245[0], u_col_out_1244[0], u_col_out_1243[0], u_col_out_1242[0], u_col_out_1241[0], u_col_out_1240[0], u_col_out_1239[0], u_col_out_1238[0], u_col_out_1237[0], u_col_out_1236[0], u_col_out_1235[0], u_col_out_1234[0], u_col_out_1233[0], u_col_out_1232[0], u_col_out_1231[0], u_col_out_1230[0], u_col_out_1229[0], u_col_out_1228[0], u_col_out_1227[0], u_col_out_1226[0], u_col_out_1225[0], u_col_out_1224[0], u_col_out_1223[0], u_col_out_1222[0], u_col_out_1221[0], u_col_out_1220[0], u_col_out_1219[0], u_col_out_1218[0], u_col_out_1217[0], u_col_out_1216[0], u_col_out_1215[0], u_col_out_1214[0], u_col_out_1213[0], u_col_out_1212[0], u_col_out_1211[0], u_col_out_1210[0], u_col_out_1209[0], u_col_out_1208[0], u_col_out_1207[0], u_col_out_1206[0], u_col_out_1205[0], u_col_out_1204[0], u_col_out_1203[0], u_col_out_1202[0], u_col_out_1201[0], u_col_out_1200[0], u_col_out_1199[0], u_col_out_1198[0], u_col_out_1197[0], u_col_out_1196[0], u_col_out_1195[0], u_col_out_1194[0], u_col_out_1193[0], u_col_out_1192[0], u_col_out_1191[0], u_col_out_1190[0], u_col_out_1189[0], u_col_out_1188[0], u_col_out_1187[0], u_col_out_1186[0], u_col_out_1185[0], u_col_out_1184[0], u_col_out_1183[0], u_col_out_1182[0], u_col_out_1181[0], u_col_out_1180[0], u_col_out_1179[0], u_col_out_1178[0], u_col_out_1177[0], u_col_out_1176[0], u_col_out_1175[0], u_col_out_1174[0], u_col_out_1173[0], u_col_out_1172[0], u_col_out_1171[0], u_col_out_1170[0], u_col_out_1169[0], u_col_out_1168[0], u_col_out_1167[0], u_col_out_1166[0], u_col_out_1165[0], u_col_out_1164[0], u_col_out_1163[0], u_col_out_1162[0], u_col_out_1161[0], u_col_out_1160[0], u_col_out_1159[0], u_col_out_1158[0], u_col_out_1157[0], u_col_out_1156[0], u_col_out_1155[0], u_col_out_1154[0], u_col_out_1153[0], u_col_out_1152[0], u_col_out_1151[0], u_col_out_1150[0], u_col_out_1149[0], u_col_out_1148[0], u_col_out_1147[0], u_col_out_1146[0], u_col_out_1145[0], u_col_out_1144[0], u_col_out_1143[0], u_col_out_1142[0], u_col_out_1141[0], u_col_out_1140[0], u_col_out_1139[0], u_col_out_1138[0], u_col_out_1137[0], u_col_out_1136[0], u_col_out_1135[0], u_col_out_1134[0], u_col_out_1133[0], u_col_out_1132[0], u_col_out_1131[0], u_col_out_1130[0], u_col_out_1129[0], u_col_out_1128[0], u_col_out_1127[0], u_col_out_1126[0], u_col_out_1125[0], u_col_out_1124[0], u_col_out_1123[0], u_col_out_1122[0], u_col_out_1121[0], u_col_out_1120[0], u_col_out_1119[0], u_col_out_1118[0], u_col_out_1117[0], u_col_out_1116[0], u_col_out_1115[0], u_col_out_1114[0], u_col_out_1113[0], u_col_out_1112[0], u_col_out_1111[0], u_col_out_1110[0], u_col_out_1109[0], u_col_out_1108[0], u_col_out_1107[0], u_col_out_1106[0], u_col_out_1105[0], u_col_out_1104[0], u_col_out_1103[0], u_col_out_1102[0], u_col_out_1101[0], u_col_out_1100[0], u_col_out_1099[0], u_col_out_1098[0], u_col_out_1097[0], u_col_out_1096[0], u_col_out_1095[0], u_col_out_1094[0], u_col_out_1093[0], u_col_out_1092[0], u_col_out_1091[0], u_col_out_1090[0], u_col_out_1089[0], u_col_out_1088[0], u_col_out_1087[0], u_col_out_1086[0], u_col_out_1085[0], u_col_out_1084[0], u_col_out_1083[0], u_col_out_1082[0], u_col_out_1081[0], u_col_out_1080[0], u_col_out_1079[0], u_col_out_1078[0], u_col_out_1077[0], u_col_out_1076[0], u_col_out_1075[0], u_col_out_1074[0], u_col_out_1073[0], u_col_out_1072[0], u_col_out_1071[0], u_col_out_1070[0], u_col_out_1069[0], u_col_out_1068[0], u_col_out_1067[0], u_col_out_1066[0], u_col_out_1065[0], u_col_out_1064[0], u_col_out_1063[0], u_col_out_1062[0], u_col_out_1061[0], u_col_out_1060[0], u_col_out_1059[0], u_col_out_1058[0], u_col_out_1057[0], u_col_out_1056[0], u_col_out_1055[0], u_col_out_1054[0], u_col_out_1053[0], u_col_out_1052[0], u_col_out_1051[0], u_col_out_1050[0], u_col_out_1049[0], u_col_out_1048[0], u_col_out_1047[0], u_col_out_1046[0], u_col_out_1045[0], u_col_out_1044[0], u_col_out_1043[0], u_col_out_1042[0], u_col_out_1041[0], u_col_out_1040[0], u_col_out_1039[0], u_col_out_1038[0], u_col_out_1037[0], u_col_out_1036[0], u_col_out_1035[0], u_col_out_1034[0], u_col_out_1033[0], u_col_out_1032[0], u_col_out_1031[0], u_col_out_1030[0], u_col_out_1029[0], u_col_out_1028[0], u_col_out_1027[0], u_col_out_1026[0], u_col_out_1025[0], u_col_out_1024[0], u_col_out_1023[0], u_col_out_1022[0], u_col_out_1021[0], u_col_out_1020[0], u_col_out_1019[0], u_col_out_1018[0], u_col_out_1017[0], u_col_out_1016[0], u_col_out_1015[0], u_col_out_1014[0], u_col_out_1013[0], u_col_out_1012[0], u_col_out_1011[0], u_col_out_1010[0], u_col_out_1009[0], u_col_out_1008[0], u_col_out_1007[0], u_col_out_1006[0], u_col_out_1005[0], u_col_out_1004[0], u_col_out_1003[0], u_col_out_1002[0], u_col_out_1001[0], u_col_out_1000[0], u_col_out_999[0], u_col_out_998[0], u_col_out_997[0], u_col_out_996[0], u_col_out_995[0], u_col_out_994[0], u_col_out_993[0], u_col_out_992[0], u_col_out_991[0], u_col_out_990[0], u_col_out_989[0], u_col_out_988[0], u_col_out_987[0], u_col_out_986[0], u_col_out_985[0], u_col_out_984[0], u_col_out_983[0], u_col_out_982[0], u_col_out_981[0], u_col_out_980[0], u_col_out_979[0], u_col_out_978[0], u_col_out_977[0], u_col_out_976[0], u_col_out_975[0], u_col_out_974[0], u_col_out_973[0], u_col_out_972[0], u_col_out_971[0], u_col_out_970[0], u_col_out_969[0], u_col_out_968[0], u_col_out_967[0], u_col_out_966[0], u_col_out_965[0], u_col_out_964[0], u_col_out_963[0], u_col_out_962[0], u_col_out_961[0], u_col_out_960[0], u_col_out_959[0], u_col_out_958[0], u_col_out_957[0], u_col_out_956[0], u_col_out_955[0], u_col_out_954[0], u_col_out_953[0], u_col_out_952[0], u_col_out_951[0], u_col_out_950[0], u_col_out_949[0], u_col_out_948[0], u_col_out_947[0], u_col_out_946[0], u_col_out_945[0], u_col_out_944[0], u_col_out_943[0], u_col_out_942[0], u_col_out_941[0], u_col_out_940[0], u_col_out_939[0], u_col_out_938[0], u_col_out_937[0], u_col_out_936[0], u_col_out_935[0], u_col_out_934[0], u_col_out_933[0], u_col_out_932[0], u_col_out_931[0], u_col_out_930[0], u_col_out_929[0], u_col_out_928[0], u_col_out_927[0], u_col_out_926[0], u_col_out_925[0], u_col_out_924[0], u_col_out_923[0], u_col_out_922[0], u_col_out_921[0], u_col_out_920[0], u_col_out_919[0], u_col_out_918[0], u_col_out_917[0], u_col_out_916[0], u_col_out_915[0], u_col_out_914[0], u_col_out_913[0], u_col_out_912[0], u_col_out_911[0], u_col_out_910[0], u_col_out_909[0], u_col_out_908[0], u_col_out_907[0], u_col_out_906[0], u_col_out_905[0], u_col_out_904[0], u_col_out_903[0], u_col_out_902[0], u_col_out_901[0], u_col_out_900[0], u_col_out_899[0], u_col_out_898[0], u_col_out_897[0], u_col_out_896[0], u_col_out_895[0], u_col_out_894[0], u_col_out_893[0], u_col_out_892[0], u_col_out_891[0], u_col_out_890[0], u_col_out_889[0], u_col_out_888[0], u_col_out_887[0], u_col_out_886[0], u_col_out_885[0], u_col_out_884[0], u_col_out_883[0], u_col_out_882[0], u_col_out_881[0], u_col_out_880[0], u_col_out_879[0], u_col_out_878[0], u_col_out_877[0], u_col_out_876[0], u_col_out_875[0], u_col_out_874[0], u_col_out_873[0], u_col_out_872[0], u_col_out_871[0], u_col_out_870[0], u_col_out_869[0], u_col_out_868[0], u_col_out_867[0], u_col_out_866[0], u_col_out_865[0], u_col_out_864[0], u_col_out_863[0], u_col_out_862[0], u_col_out_861[0], u_col_out_860[0], u_col_out_859[0], u_col_out_858[0], u_col_out_857[0], u_col_out_856[0], u_col_out_855[0], u_col_out_854[0], u_col_out_853[0], u_col_out_852[0], u_col_out_851[0], u_col_out_850[0], u_col_out_849[0], u_col_out_848[0], u_col_out_847[0], u_col_out_846[0], u_col_out_845[0], u_col_out_844[0], u_col_out_843[0], u_col_out_842[0], u_col_out_841[0], u_col_out_840[0], u_col_out_839[0], u_col_out_838[0], u_col_out_837[0], u_col_out_836[0], u_col_out_835[0], u_col_out_834[0], u_col_out_833[0], u_col_out_832[0], u_col_out_831[0], u_col_out_830[0], u_col_out_829[0], u_col_out_828[0], u_col_out_827[0], u_col_out_826[0], u_col_out_825[0], u_col_out_824[0], u_col_out_823[0], u_col_out_822[0], u_col_out_821[0], u_col_out_820[0], u_col_out_819[0], u_col_out_818[0], u_col_out_817[0], u_col_out_816[0], u_col_out_815[0], u_col_out_814[0], u_col_out_813[0], u_col_out_812[0], u_col_out_811[0], u_col_out_810[0], u_col_out_809[0], u_col_out_808[0], u_col_out_807[0], u_col_out_806[0], u_col_out_805[0], u_col_out_804[0], u_col_out_803[0], u_col_out_802[0], u_col_out_801[0], u_col_out_800[0], u_col_out_799[0], u_col_out_798[0], u_col_out_797[0], u_col_out_796[0], u_col_out_795[0], u_col_out_794[0], u_col_out_793[0], u_col_out_792[0], u_col_out_791[0], u_col_out_790[0], u_col_out_789[0], u_col_out_788[0], u_col_out_787[0], u_col_out_786[0], u_col_out_785[0], u_col_out_784[0], u_col_out_783[0], u_col_out_782[0], u_col_out_781[0], u_col_out_780[0], u_col_out_779[0], u_col_out_778[0], u_col_out_777[0], u_col_out_776[0], u_col_out_775[0], u_col_out_774[0], u_col_out_773[0], u_col_out_772[0], u_col_out_771[0], u_col_out_770[0], u_col_out_769[0], u_col_out_768[0], u_col_out_767[0], u_col_out_766[0], u_col_out_765[0], u_col_out_764[0], u_col_out_763[0], u_col_out_762[0], u_col_out_761[0], u_col_out_760[0], u_col_out_759[0], u_col_out_758[0], u_col_out_757[0], u_col_out_756[0], u_col_out_755[0], u_col_out_754[0], u_col_out_753[0], u_col_out_752[0], u_col_out_751[0], u_col_out_750[0], u_col_out_749[0], u_col_out_748[0], u_col_out_747[0], u_col_out_746[0], u_col_out_745[0], u_col_out_744[0], u_col_out_743[0], u_col_out_742[0], u_col_out_741[0], u_col_out_740[0], u_col_out_739[0], u_col_out_738[0], u_col_out_737[0], u_col_out_736[0], u_col_out_735[0], u_col_out_734[0], u_col_out_733[0], u_col_out_732[0], u_col_out_731[0], u_col_out_730[0], u_col_out_729[0], u_col_out_728[0], u_col_out_727[0], u_col_out_726[0], u_col_out_725[0], u_col_out_724[0], u_col_out_723[0], u_col_out_722[0], u_col_out_721[0], u_col_out_720[0], u_col_out_719[0], u_col_out_718[0], u_col_out_717[0], u_col_out_716[0], u_col_out_715[0], u_col_out_714[0], u_col_out_713[0], u_col_out_712[0], u_col_out_711[0], u_col_out_710[0], u_col_out_709[0], u_col_out_708[0], u_col_out_707[0], u_col_out_706[0], u_col_out_705[0], u_col_out_704[0], u_col_out_703[0], u_col_out_702[0], u_col_out_701[0], u_col_out_700[0], u_col_out_699[0], u_col_out_698[0], u_col_out_697[0], u_col_out_696[0], u_col_out_695[0], u_col_out_694[0], u_col_out_693[0], u_col_out_692[0], u_col_out_691[0], u_col_out_690[0], u_col_out_689[0], u_col_out_688[0], u_col_out_687[0], u_col_out_686[0], u_col_out_685[0], u_col_out_684[0], u_col_out_683[0], u_col_out_682[0], u_col_out_681[0], u_col_out_680[0], u_col_out_679[0], u_col_out_678[0], u_col_out_677[0], u_col_out_676[0], u_col_out_675[0], u_col_out_674[0], u_col_out_673[0], u_col_out_672[0], u_col_out_671[0], u_col_out_670[0], u_col_out_669[0], u_col_out_668[0], u_col_out_667[0], u_col_out_666[0], u_col_out_665[0], u_col_out_664[0], u_col_out_663[0], u_col_out_662[0], u_col_out_661[0], u_col_out_660[0], u_col_out_659[0], u_col_out_658[0], u_col_out_657[0], u_col_out_656[0], u_col_out_655[0], u_col_out_654[0], u_col_out_653[0], u_col_out_652[0], u_col_out_651[0], u_col_out_650[0], u_col_out_649[0], u_col_out_648[0], u_col_out_647[0], u_col_out_646[0], u_col_out_645[0], u_col_out_644[0], u_col_out_643[0], u_col_out_642[0], u_col_out_641[0], u_col_out_640[0], u_col_out_639[0], u_col_out_638[0], u_col_out_637[0], u_col_out_636[0], u_col_out_635[0], u_col_out_634[0], u_col_out_633[0], u_col_out_632[0], u_col_out_631[0], u_col_out_630[0], u_col_out_629[0], u_col_out_628[0], u_col_out_627[0], u_col_out_626[0], u_col_out_625[0], u_col_out_624[0], u_col_out_623[0], u_col_out_622[0], u_col_out_621[0], u_col_out_620[0], u_col_out_619[0], u_col_out_618[0], u_col_out_617[0], u_col_out_616[0], u_col_out_615[0], u_col_out_614[0], u_col_out_613[0], u_col_out_612[0], u_col_out_611[0], u_col_out_610[0], u_col_out_609[0], u_col_out_608[0], u_col_out_607[0], u_col_out_606[0], u_col_out_605[0], u_col_out_604[0], u_col_out_603[0], u_col_out_602[0], u_col_out_601[0], u_col_out_600[0], u_col_out_599[0], u_col_out_598[0], u_col_out_597[0], u_col_out_596[0], u_col_out_595[0], u_col_out_594[0], u_col_out_593[0], u_col_out_592[0], u_col_out_591[0], u_col_out_590[0], u_col_out_589[0], u_col_out_588[0], u_col_out_587[0], u_col_out_586[0], u_col_out_585[0], u_col_out_584[0], u_col_out_583[0], u_col_out_582[0], u_col_out_581[0], u_col_out_580[0], u_col_out_579[0], u_col_out_578[0], u_col_out_577[0], u_col_out_576[0], u_col_out_575[0], u_col_out_574[0], u_col_out_573[0], u_col_out_572[0], u_col_out_571[0], u_col_out_570[0], u_col_out_569[0], u_col_out_568[0], u_col_out_567[0], u_col_out_566[0], u_col_out_565[0], u_col_out_564[0], u_col_out_563[0], u_col_out_562[0], u_col_out_561[0], u_col_out_560[0], u_col_out_559[0], u_col_out_558[0], u_col_out_557[0], u_col_out_556[0], u_col_out_555[0], u_col_out_554[0], u_col_out_553[0], u_col_out_552[0], u_col_out_551[0], u_col_out_550[0], u_col_out_549[0], u_col_out_548[0], u_col_out_547[0], u_col_out_546[0], u_col_out_545[0], u_col_out_544[0], u_col_out_543[0], u_col_out_542[0], u_col_out_541[0], u_col_out_540[0], u_col_out_539[0], u_col_out_538[0], u_col_out_537[0], u_col_out_536[0], u_col_out_535[0], u_col_out_534[0], u_col_out_533[0], u_col_out_532[0], u_col_out_531[0], u_col_out_530[0], u_col_out_529[0], u_col_out_528[0], u_col_out_527[0], u_col_out_526[0], u_col_out_525[0], u_col_out_524[0], u_col_out_523[0], u_col_out_522[0], u_col_out_521[0], u_col_out_520[0], u_col_out_519[0], u_col_out_518[0], u_col_out_517[0], u_col_out_516[0], u_col_out_515[0], u_col_out_514[0], u_col_out_513[0], u_col_out_512[0], u_col_out_511[0], u_col_out_510[0], u_col_out_509[0], u_col_out_508[0], u_col_out_507[0], u_col_out_506[0], u_col_out_505[0], u_col_out_504[0], u_col_out_503[0], u_col_out_502[0], u_col_out_501[0], u_col_out_500[0], u_col_out_499[0], u_col_out_498[0], u_col_out_497[0], u_col_out_496[0], u_col_out_495[0], u_col_out_494[0], u_col_out_493[0], u_col_out_492[0], u_col_out_491[0], u_col_out_490[0], u_col_out_489[0], u_col_out_488[0], u_col_out_487[0], u_col_out_486[0], u_col_out_485[0], u_col_out_484[0], u_col_out_483[0], u_col_out_482[0], u_col_out_481[0], u_col_out_480[0], u_col_out_479[0], u_col_out_478[0], u_col_out_477[0], u_col_out_476[0], u_col_out_475[0], u_col_out_474[0], u_col_out_473[0], u_col_out_472[0], u_col_out_471[0], u_col_out_470[0], u_col_out_469[0], u_col_out_468[0], u_col_out_467[0], u_col_out_466[0], u_col_out_465[0], u_col_out_464[0], u_col_out_463[0], u_col_out_462[0], u_col_out_461[0], u_col_out_460[0], u_col_out_459[0], u_col_out_458[0], u_col_out_457[0], u_col_out_456[0], u_col_out_455[0], u_col_out_454[0], u_col_out_453[0], u_col_out_452[0], u_col_out_451[0], u_col_out_450[0], u_col_out_449[0], u_col_out_448[0], u_col_out_447[0], u_col_out_446[0], u_col_out_445[0], u_col_out_444[0], u_col_out_443[0], u_col_out_442[0], u_col_out_441[0], u_col_out_440[0], u_col_out_439[0], u_col_out_438[0], u_col_out_437[0], u_col_out_436[0], u_col_out_435[0], u_col_out_434[0], u_col_out_433[0], u_col_out_432[0], u_col_out_431[0], u_col_out_430[0], u_col_out_429[0], u_col_out_428[0], u_col_out_427[0], u_col_out_426[0], u_col_out_425[0], u_col_out_424[0], u_col_out_423[0], u_col_out_422[0], u_col_out_421[0], u_col_out_420[0], u_col_out_419[0], u_col_out_418[0], u_col_out_417[0], u_col_out_416[0], u_col_out_415[0], u_col_out_414[0], u_col_out_413[0], u_col_out_412[0], u_col_out_411[0], u_col_out_410[0], u_col_out_409[0], u_col_out_408[0], u_col_out_407[0], u_col_out_406[0], u_col_out_405[0], u_col_out_404[0], u_col_out_403[0], u_col_out_402[0], u_col_out_401[0], u_col_out_400[0], u_col_out_399[0], u_col_out_398[0], u_col_out_397[0], u_col_out_396[0], u_col_out_395[0], u_col_out_394[0], u_col_out_393[0], u_col_out_392[0], u_col_out_391[0], u_col_out_390[0], u_col_out_389[0], u_col_out_388[0], u_col_out_387[0], u_col_out_386[0], u_col_out_385[0], u_col_out_384[0], u_col_out_383[0], u_col_out_382[0], u_col_out_381[0], u_col_out_380[0], u_col_out_379[0], u_col_out_378[0], u_col_out_377[0], u_col_out_376[0], u_col_out_375[0], u_col_out_374[0], u_col_out_373[0], u_col_out_372[0], u_col_out_371[0], u_col_out_370[0], u_col_out_369[0], u_col_out_368[0], u_col_out_367[0], u_col_out_366[0], u_col_out_365[0], u_col_out_364[0], u_col_out_363[0], u_col_out_362[0], u_col_out_361[0], u_col_out_360[0], u_col_out_359[0], u_col_out_358[0], u_col_out_357[0], u_col_out_356[0], u_col_out_355[0], u_col_out_354[0], u_col_out_353[0], u_col_out_352[0], u_col_out_351[0], u_col_out_350[0], u_col_out_349[0], u_col_out_348[0], u_col_out_347[0], u_col_out_346[0], u_col_out_345[0], u_col_out_344[0], u_col_out_343[0], u_col_out_342[0], u_col_out_341[0], u_col_out_340[0], u_col_out_339[0], u_col_out_338[0], u_col_out_337[0], u_col_out_336[0], u_col_out_335[0], u_col_out_334[0], u_col_out_333[0], u_col_out_332[0], u_col_out_331[0], u_col_out_330[0], u_col_out_329[0], u_col_out_328[0], u_col_out_327[0], u_col_out_326[0], u_col_out_325[0], u_col_out_324[0], u_col_out_323[0], u_col_out_322[0], u_col_out_321[0], u_col_out_320[0], u_col_out_319[0], u_col_out_318[0], u_col_out_317[0], u_col_out_316[0], u_col_out_315[0], u_col_out_314[0], u_col_out_313[0], u_col_out_312[0], u_col_out_311[0], u_col_out_310[0], u_col_out_309[0], u_col_out_308[0], u_col_out_307[0], u_col_out_306[0], u_col_out_305[0], u_col_out_304[0], u_col_out_303[0], u_col_out_302[0], u_col_out_301[0], u_col_out_300[0], u_col_out_299[0], u_col_out_298[0], u_col_out_297[0], u_col_out_296[0], u_col_out_295[0], u_col_out_294[0], u_col_out_293[0], u_col_out_292[0], u_col_out_291[0], u_col_out_290[0], u_col_out_289[0], u_col_out_288[0], u_col_out_287[0], u_col_out_286[0], u_col_out_285[0], u_col_out_284[0], u_col_out_283[0], u_col_out_282[0], u_col_out_281[0], u_col_out_280[0], u_col_out_279[0], u_col_out_278[0], u_col_out_277[0], u_col_out_276[0], u_col_out_275[0], u_col_out_274[0], u_col_out_273[0], u_col_out_272[0], u_col_out_271[0], u_col_out_270[0], u_col_out_269[0], u_col_out_268[0], u_col_out_267[0], u_col_out_266[0], u_col_out_265[0], u_col_out_264[0], u_col_out_263[0], u_col_out_262[0], u_col_out_261[0], u_col_out_260[0], u_col_out_259[0], u_col_out_258[0], u_col_out_257[0], u_col_out_256[0], u_col_out_255[0], u_col_out_254[0], u_col_out_253[0], u_col_out_252[0], u_col_out_251[0], u_col_out_250[0], u_col_out_249[0], u_col_out_248[0], u_col_out_247[0], u_col_out_246[0], u_col_out_245[0], u_col_out_244[0], u_col_out_243[0], u_col_out_242[0], u_col_out_241[0], u_col_out_240[0], u_col_out_239[0], u_col_out_238[0], u_col_out_237[0], u_col_out_236[0], u_col_out_235[0], u_col_out_234[0], u_col_out_233[0], u_col_out_232[0], u_col_out_231[0], u_col_out_230[0], u_col_out_229[0], u_col_out_228[0], u_col_out_227[0], u_col_out_226[0], u_col_out_225[0], u_col_out_224[0], u_col_out_223[0], u_col_out_222[0], u_col_out_221[0], u_col_out_220[0], u_col_out_219[0], u_col_out_218[0], u_col_out_217[0], u_col_out_216[0], u_col_out_215[0], u_col_out_214[0], u_col_out_213[0], u_col_out_212[0], u_col_out_211[0], u_col_out_210[0], u_col_out_209[0], u_col_out_208[0], u_col_out_207[0], u_col_out_206[0], u_col_out_205[0], u_col_out_204[0], u_col_out_203[0], u_col_out_202[0], u_col_out_201[0], u_col_out_200[0], u_col_out_199[0], u_col_out_198[0], u_col_out_197[0], u_col_out_196[0], u_col_out_195[0], u_col_out_194[0], u_col_out_193[0], u_col_out_192[0], u_col_out_191[0], u_col_out_190[0], u_col_out_189[0], u_col_out_188[0], u_col_out_187[0], u_col_out_186[0], u_col_out_185[0], u_col_out_184[0], u_col_out_183[0], u_col_out_182[0], u_col_out_181[0], u_col_out_180[0], u_col_out_179[0], u_col_out_178[0], u_col_out_177[0], u_col_out_176[0], u_col_out_175[0], u_col_out_174[0], u_col_out_173[0], u_col_out_172[0], u_col_out_171[0], u_col_out_170[0], u_col_out_169[0], u_col_out_168[0], u_col_out_167[0], u_col_out_166[0], u_col_out_165[0], u_col_out_164[0], u_col_out_163[0], u_col_out_162[0], u_col_out_161[0], u_col_out_160[0], u_col_out_159[0], u_col_out_158[0], u_col_out_157[0], u_col_out_156[0], u_col_out_155[0], u_col_out_154[0], u_col_out_153[0], u_col_out_152[0], u_col_out_151[0], u_col_out_150[0], u_col_out_149[0], u_col_out_148[0], u_col_out_147[0], u_col_out_146[0], u_col_out_145[0], u_col_out_144[0], u_col_out_143[0], u_col_out_142[0], u_col_out_141[0], u_col_out_140[0], u_col_out_139[0], u_col_out_138[0], u_col_out_137[0], u_col_out_136[0], u_col_out_135[0], u_col_out_134[0], u_col_out_133[0], u_col_out_132[0], u_col_out_131[0], u_col_out_130[0], u_col_out_129[0], u_col_out_128[0], u_col_out_127[0], u_col_out_126[0], u_col_out_125[0], u_col_out_124[0], u_col_out_123[0], u_col_out_122[0], u_col_out_121[0], u_col_out_120[0], u_col_out_119[0], u_col_out_118[0], u_col_out_117[0], u_col_out_116[0], u_col_out_115[0], u_col_out_114[0], u_col_out_113[0], u_col_out_112[0], u_col_out_111[0], u_col_out_110[0], u_col_out_109[0], u_col_out_108[0], u_col_out_107[0], u_col_out_106[0], u_col_out_105[0], u_col_out_104[0], u_col_out_103[0], u_col_out_102[0], u_col_out_101[0], u_col_out_100[0], u_col_out_99[0], u_col_out_98[0], u_col_out_97[0], u_col_out_96[0], u_col_out_95[0], u_col_out_94[0], u_col_out_93[0], u_col_out_92[0], u_col_out_91[0], u_col_out_90[0], u_col_out_89[0], u_col_out_88[0], u_col_out_87[0], u_col_out_86[0], u_col_out_85[0], u_col_out_84[0], u_col_out_83[0], u_col_out_82[0], u_col_out_81[0], u_col_out_80[0], u_col_out_79[0], u_col_out_78[0], u_col_out_77[0], u_col_out_76[0], u_col_out_75[0], u_col_out_74[0], u_col_out_73[0], u_col_out_72[0], u_col_out_71[0], u_col_out_70[0], u_col_out_69[0], u_col_out_68[0], u_col_out_67[0], u_col_out_66[0], u_col_out_65[0], u_col_out_64[0], u_col_out_63[0], u_col_out_62[0], u_col_out_61[0], u_col_out_60[0], u_col_out_59[0], u_col_out_58[0], u_col_out_57[0], u_col_out_56[0], u_col_out_55[0], u_col_out_54[0], u_col_out_53[0], u_col_out_52[0], u_col_out_51[0], u_col_out_50[0], u_col_out_49[0], u_col_out_48[0], u_col_out_47[0], u_col_out_46[0], u_col_out_45[0], u_col_out_44[0], u_col_out_43[0], u_col_out_42[0], u_col_out_41[0], u_col_out_40[0], u_col_out_39[0], u_col_out_38[0], u_col_out_37[0], u_col_out_36[0], u_col_out_35[0], u_col_out_34[0], u_col_out_33[0], u_col_out_32[0], u_col_out_31[0], u_col_out_30[0], u_col_out_29[0], u_col_out_28[0], u_col_out_27[0], u_col_out_26[0], u_col_out_25[0], u_col_out_24[0], u_col_out_23[0], u_col_out_22[0], u_col_out_21[0], u_col_out_20[0], u_col_out_19[0], u_col_out_18[0], u_col_out_17[0], u_col_out_16[0], u_col_out_15[0], u_col_out_14[0], u_col_out_13[0], u_col_out_12[0], u_col_out_11[0], u_col_out_10[0], u_col_out_9[0], u_col_out_8[0], u_col_out_7[0], u_col_out_6[0], u_col_out_5[0], u_col_out_4[0], u_col_out_3[0], u_col_out_2[0], u_col_out_1[0], u_col_out_0[0]};


assign row_out_1 = {u_col_out_1287[1], u_col_out_1286[1], u_col_out_1285[1], u_col_out_1284[1], u_col_out_1283[1], u_col_out_1282[1], u_col_out_1281[1], u_col_out_1280[1], u_col_out_1279[1], u_col_out_1278[1], u_col_out_1277[1], u_col_out_1276[1], u_col_out_1275[1], u_col_out_1274[1], u_col_out_1273[1], u_col_out_1272[1], u_col_out_1271[1], u_col_out_1270[1], u_col_out_1269[1], u_col_out_1268[1], u_col_out_1267[1], u_col_out_1266[1], u_col_out_1265[1], u_col_out_1264[1], u_col_out_1263[1], u_col_out_1262[1], u_col_out_1261[1], u_col_out_1260[1], u_col_out_1259[1], u_col_out_1258[1], u_col_out_1257[1], u_col_out_1256[1], u_col_out_1255[1], u_col_out_1254[1], u_col_out_1253[1], u_col_out_1252[1], u_col_out_1251[1], u_col_out_1250[1], u_col_out_1249[1], u_col_out_1248[1], u_col_out_1247[1], u_col_out_1246[1], u_col_out_1245[1], u_col_out_1244[1], u_col_out_1243[1], u_col_out_1242[1], u_col_out_1241[1], u_col_out_1240[1], u_col_out_1239[1], u_col_out_1238[1], u_col_out_1237[1], u_col_out_1236[1], u_col_out_1235[1], u_col_out_1234[1], u_col_out_1233[1], u_col_out_1232[1], u_col_out_1231[1], u_col_out_1230[1], u_col_out_1229[1], u_col_out_1228[1], u_col_out_1227[1], u_col_out_1226[1], u_col_out_1225[1], u_col_out_1224[1], u_col_out_1223[1], u_col_out_1222[1], u_col_out_1221[1], u_col_out_1220[1], u_col_out_1219[1], u_col_out_1218[1], u_col_out_1217[1], u_col_out_1216[1], u_col_out_1215[1], u_col_out_1214[1], u_col_out_1213[1], u_col_out_1212[1], u_col_out_1211[1], u_col_out_1210[1], u_col_out_1209[1], u_col_out_1208[1], u_col_out_1207[1], u_col_out_1206[1], u_col_out_1205[1], u_col_out_1204[1], u_col_out_1203[1], u_col_out_1202[1], u_col_out_1201[1], u_col_out_1200[1], u_col_out_1199[1], u_col_out_1198[1], u_col_out_1197[1], u_col_out_1196[1], u_col_out_1195[1], u_col_out_1194[1], u_col_out_1193[1], u_col_out_1192[1], u_col_out_1191[1], u_col_out_1190[1], u_col_out_1189[1], u_col_out_1188[1], u_col_out_1187[1], u_col_out_1186[1], u_col_out_1185[1], u_col_out_1184[1], u_col_out_1183[1], u_col_out_1182[1], u_col_out_1181[1], u_col_out_1180[1], u_col_out_1179[1], u_col_out_1178[1], u_col_out_1177[1], u_col_out_1176[1], u_col_out_1175[1], u_col_out_1174[1], u_col_out_1173[1], u_col_out_1172[1], u_col_out_1171[1], u_col_out_1170[1], u_col_out_1169[1], u_col_out_1168[1], u_col_out_1167[1], u_col_out_1166[1], u_col_out_1165[1], u_col_out_1164[1], u_col_out_1163[1], u_col_out_1162[1], u_col_out_1161[1], u_col_out_1160[1], u_col_out_1159[1], u_col_out_1158[1], u_col_out_1157[1], u_col_out_1156[1], u_col_out_1155[1], u_col_out_1154[1], u_col_out_1153[1], u_col_out_1152[1], u_col_out_1151[1], u_col_out_1150[1], u_col_out_1149[1], u_col_out_1148[1], u_col_out_1147[1], u_col_out_1146[1], u_col_out_1145[1], u_col_out_1144[1], u_col_out_1143[1], u_col_out_1142[1], u_col_out_1141[1], u_col_out_1140[1], u_col_out_1139[1], u_col_out_1138[1], u_col_out_1137[1], u_col_out_1136[1], u_col_out_1135[1], u_col_out_1134[1], u_col_out_1133[1], u_col_out_1132[1], u_col_out_1131[1], u_col_out_1130[1], u_col_out_1129[1], u_col_out_1128[1], u_col_out_1127[1], u_col_out_1126[1], u_col_out_1125[1], u_col_out_1124[1], u_col_out_1123[1], u_col_out_1122[1], u_col_out_1121[1], u_col_out_1120[1], u_col_out_1119[1], u_col_out_1118[1], u_col_out_1117[1], u_col_out_1116[1], u_col_out_1115[1], u_col_out_1114[1], u_col_out_1113[1], u_col_out_1112[1], u_col_out_1111[1], u_col_out_1110[1], u_col_out_1109[1], u_col_out_1108[1], u_col_out_1107[1], u_col_out_1106[1], u_col_out_1105[1], u_col_out_1104[1], u_col_out_1103[1], u_col_out_1102[1], u_col_out_1101[1], u_col_out_1100[1], u_col_out_1099[1], u_col_out_1098[1], u_col_out_1097[1], u_col_out_1096[1], u_col_out_1095[1], u_col_out_1094[1], u_col_out_1093[1], u_col_out_1092[1], u_col_out_1091[1], u_col_out_1090[1], u_col_out_1089[1], u_col_out_1088[1], u_col_out_1087[1], u_col_out_1086[1], u_col_out_1085[1], u_col_out_1084[1], u_col_out_1083[1], u_col_out_1082[1], u_col_out_1081[1], u_col_out_1080[1], u_col_out_1079[1], u_col_out_1078[1], u_col_out_1077[1], u_col_out_1076[1], u_col_out_1075[1], u_col_out_1074[1], u_col_out_1073[1], u_col_out_1072[1], u_col_out_1071[1], u_col_out_1070[1], u_col_out_1069[1], u_col_out_1068[1], u_col_out_1067[1], u_col_out_1066[1], u_col_out_1065[1], u_col_out_1064[1], u_col_out_1063[1], u_col_out_1062[1], u_col_out_1061[1], u_col_out_1060[1], u_col_out_1059[1], u_col_out_1058[1], u_col_out_1057[1], u_col_out_1056[1], u_col_out_1055[1], u_col_out_1054[1], u_col_out_1053[1], u_col_out_1052[1], u_col_out_1051[1], u_col_out_1050[1], u_col_out_1049[1], u_col_out_1048[1], u_col_out_1047[1], u_col_out_1046[1], u_col_out_1045[1], u_col_out_1044[1], u_col_out_1043[1], u_col_out_1042[1], u_col_out_1041[1], u_col_out_1040[1], u_col_out_1039[1], u_col_out_1038[1], u_col_out_1037[1], u_col_out_1036[1], u_col_out_1035[1], u_col_out_1034[1], u_col_out_1033[1], u_col_out_1032[1], u_col_out_1031[1], u_col_out_1030[1], u_col_out_1029[1], u_col_out_1028[1], u_col_out_1027[1], u_col_out_1026[1], u_col_out_1025[1], u_col_out_1024[1], u_col_out_1023[1], u_col_out_1022[1], u_col_out_1021[1], u_col_out_1020[1], u_col_out_1019[1], u_col_out_1018[1], u_col_out_1017[1], u_col_out_1016[1], u_col_out_1015[1], u_col_out_1014[1], u_col_out_1013[1], u_col_out_1012[1], u_col_out_1011[1], u_col_out_1010[1], u_col_out_1009[1], u_col_out_1008[1], u_col_out_1007[1], u_col_out_1006[1], u_col_out_1005[1], u_col_out_1004[1], u_col_out_1003[1], u_col_out_1002[1], u_col_out_1001[1], u_col_out_1000[1], u_col_out_999[1], u_col_out_998[1], u_col_out_997[1], u_col_out_996[1], u_col_out_995[1], u_col_out_994[1], u_col_out_993[1], u_col_out_992[1], u_col_out_991[1], u_col_out_990[1], u_col_out_989[1], u_col_out_988[1], u_col_out_987[1], u_col_out_986[1], u_col_out_985[1], u_col_out_984[1], u_col_out_983[1], u_col_out_982[1], u_col_out_981[1], u_col_out_980[1], u_col_out_979[1], u_col_out_978[1], u_col_out_977[1], u_col_out_976[1], u_col_out_975[1], u_col_out_974[1], u_col_out_973[1], u_col_out_972[1], u_col_out_971[1], u_col_out_970[1], u_col_out_969[1], u_col_out_968[1], u_col_out_967[1], u_col_out_966[1], u_col_out_965[1], u_col_out_964[1], u_col_out_963[1], u_col_out_962[1], u_col_out_961[1], u_col_out_960[1], u_col_out_959[1], u_col_out_958[1], u_col_out_957[1], u_col_out_956[1], u_col_out_955[1], u_col_out_954[1], u_col_out_953[1], u_col_out_952[1], u_col_out_951[1], u_col_out_950[1], u_col_out_949[1], u_col_out_948[1], u_col_out_947[1], u_col_out_946[1], u_col_out_945[1], u_col_out_944[1], u_col_out_943[1], u_col_out_942[1], u_col_out_941[1], u_col_out_940[1], u_col_out_939[1], u_col_out_938[1], u_col_out_937[1], u_col_out_936[1], u_col_out_935[1], u_col_out_934[1], u_col_out_933[1], u_col_out_932[1], u_col_out_931[1], u_col_out_930[1], u_col_out_929[1], u_col_out_928[1], u_col_out_927[1], u_col_out_926[1], u_col_out_925[1], u_col_out_924[1], u_col_out_923[1], u_col_out_922[1], u_col_out_921[1], u_col_out_920[1], u_col_out_919[1], u_col_out_918[1], u_col_out_917[1], u_col_out_916[1], u_col_out_915[1], u_col_out_914[1], u_col_out_913[1], u_col_out_912[1], u_col_out_911[1], u_col_out_910[1], u_col_out_909[1], u_col_out_908[1], u_col_out_907[1], u_col_out_906[1], u_col_out_905[1], u_col_out_904[1], u_col_out_903[1], u_col_out_902[1], u_col_out_901[1], u_col_out_900[1], u_col_out_899[1], u_col_out_898[1], u_col_out_897[1], u_col_out_896[1], u_col_out_895[1], u_col_out_894[1], u_col_out_893[1], u_col_out_892[1], u_col_out_891[1], u_col_out_890[1], u_col_out_889[1], u_col_out_888[1], u_col_out_887[1], u_col_out_886[1], u_col_out_885[1], u_col_out_884[1], u_col_out_883[1], u_col_out_882[1], u_col_out_881[1], u_col_out_880[1], u_col_out_879[1], u_col_out_878[1], u_col_out_877[1], u_col_out_876[1], u_col_out_875[1], u_col_out_874[1], u_col_out_873[1], u_col_out_872[1], u_col_out_871[1], u_col_out_870[1], u_col_out_869[1], u_col_out_868[1], u_col_out_867[1], u_col_out_866[1], u_col_out_865[1], u_col_out_864[1], u_col_out_863[1], u_col_out_862[1], u_col_out_861[1], u_col_out_860[1], u_col_out_859[1], u_col_out_858[1], u_col_out_857[1], u_col_out_856[1], u_col_out_855[1], u_col_out_854[1], u_col_out_853[1], u_col_out_852[1], u_col_out_851[1], u_col_out_850[1], u_col_out_849[1], u_col_out_848[1], u_col_out_847[1], u_col_out_846[1], u_col_out_845[1], u_col_out_844[1], u_col_out_843[1], u_col_out_842[1], u_col_out_841[1], u_col_out_840[1], u_col_out_839[1], u_col_out_838[1], u_col_out_837[1], u_col_out_836[1], u_col_out_835[1], u_col_out_834[1], u_col_out_833[1], u_col_out_832[1], u_col_out_831[1], u_col_out_830[1], u_col_out_829[1], u_col_out_828[1], u_col_out_827[1], u_col_out_826[1], u_col_out_825[1], u_col_out_824[1], u_col_out_823[1], u_col_out_822[1], u_col_out_821[1], u_col_out_820[1], u_col_out_819[1], u_col_out_818[1], u_col_out_817[1], u_col_out_816[1], u_col_out_815[1], u_col_out_814[1], u_col_out_813[1], u_col_out_812[1], u_col_out_811[1], u_col_out_810[1], u_col_out_809[1], u_col_out_808[1], u_col_out_807[1], u_col_out_806[1], u_col_out_805[1], u_col_out_804[1], u_col_out_803[1], u_col_out_802[1], u_col_out_801[1], u_col_out_800[1], u_col_out_799[1], u_col_out_798[1], u_col_out_797[1], u_col_out_796[1], u_col_out_795[1], u_col_out_794[1], u_col_out_793[1], u_col_out_792[1], u_col_out_791[1], u_col_out_790[1], u_col_out_789[1], u_col_out_788[1], u_col_out_787[1], u_col_out_786[1], u_col_out_785[1], u_col_out_784[1], u_col_out_783[1], u_col_out_782[1], u_col_out_781[1], u_col_out_780[1], u_col_out_779[1], u_col_out_778[1], u_col_out_777[1], u_col_out_776[1], u_col_out_775[1], u_col_out_774[1], u_col_out_773[1], u_col_out_772[1], u_col_out_771[1], u_col_out_770[1], u_col_out_769[1], u_col_out_768[1], u_col_out_767[1], u_col_out_766[1], u_col_out_765[1], u_col_out_764[1], u_col_out_763[1], u_col_out_762[1], u_col_out_761[1], u_col_out_760[1], u_col_out_759[1], u_col_out_758[1], u_col_out_757[1], u_col_out_756[1], u_col_out_755[1], u_col_out_754[1], u_col_out_753[1], u_col_out_752[1], u_col_out_751[1], u_col_out_750[1], u_col_out_749[1], u_col_out_748[1], u_col_out_747[1], u_col_out_746[1], u_col_out_745[1], u_col_out_744[1], u_col_out_743[1], u_col_out_742[1], u_col_out_741[1], u_col_out_740[1], u_col_out_739[1], u_col_out_738[1], u_col_out_737[1], u_col_out_736[1], u_col_out_735[1], u_col_out_734[1], u_col_out_733[1], u_col_out_732[1], u_col_out_731[1], u_col_out_730[1], u_col_out_729[1], u_col_out_728[1], u_col_out_727[1], u_col_out_726[1], u_col_out_725[1], u_col_out_724[1], u_col_out_723[1], u_col_out_722[1], u_col_out_721[1], u_col_out_720[1], u_col_out_719[1], u_col_out_718[1], u_col_out_717[1], u_col_out_716[1], u_col_out_715[1], u_col_out_714[1], u_col_out_713[1], u_col_out_712[1], u_col_out_711[1], u_col_out_710[1], u_col_out_709[1], u_col_out_708[1], u_col_out_707[1], u_col_out_706[1], u_col_out_705[1], u_col_out_704[1], u_col_out_703[1], u_col_out_702[1], u_col_out_701[1], u_col_out_700[1], u_col_out_699[1], u_col_out_698[1], u_col_out_697[1], u_col_out_696[1], u_col_out_695[1], u_col_out_694[1], u_col_out_693[1], u_col_out_692[1], u_col_out_691[1], u_col_out_690[1], u_col_out_689[1], u_col_out_688[1], u_col_out_687[1], u_col_out_686[1], u_col_out_685[1], u_col_out_684[1], u_col_out_683[1], u_col_out_682[1], u_col_out_681[1], u_col_out_680[1], u_col_out_679[1], u_col_out_678[1], u_col_out_677[1], u_col_out_676[1], u_col_out_675[1], u_col_out_674[1], u_col_out_673[1], u_col_out_672[1], u_col_out_671[1], u_col_out_670[1], u_col_out_669[1], u_col_out_668[1], u_col_out_667[1], u_col_out_666[1], u_col_out_665[1], u_col_out_664[1], u_col_out_663[1], u_col_out_662[1], u_col_out_661[1], u_col_out_660[1], u_col_out_659[1], u_col_out_658[1], u_col_out_657[1], u_col_out_656[1], u_col_out_655[1], u_col_out_654[1], u_col_out_653[1], u_col_out_652[1], u_col_out_651[1], u_col_out_650[1], u_col_out_649[1], u_col_out_648[1], u_col_out_647[1], u_col_out_646[1], u_col_out_645[1], u_col_out_644[1], u_col_out_643[1], u_col_out_642[1], u_col_out_641[1], u_col_out_640[1], u_col_out_639[1], u_col_out_638[1], u_col_out_637[1], u_col_out_636[1], u_col_out_635[1], u_col_out_634[1], u_col_out_633[1], u_col_out_632[1], u_col_out_631[1], u_col_out_630[1], u_col_out_629[1], u_col_out_628[1], u_col_out_627[1], u_col_out_626[1], u_col_out_625[1], u_col_out_624[1], u_col_out_623[1], u_col_out_622[1], u_col_out_621[1], u_col_out_620[1], u_col_out_619[1], u_col_out_618[1], u_col_out_617[1], u_col_out_616[1], u_col_out_615[1], u_col_out_614[1], u_col_out_613[1], u_col_out_612[1], u_col_out_611[1], u_col_out_610[1], u_col_out_609[1], u_col_out_608[1], u_col_out_607[1], u_col_out_606[1], u_col_out_605[1], u_col_out_604[1], u_col_out_603[1], u_col_out_602[1], u_col_out_601[1], u_col_out_600[1], u_col_out_599[1], u_col_out_598[1], u_col_out_597[1], u_col_out_596[1], u_col_out_595[1], u_col_out_594[1], u_col_out_593[1], u_col_out_592[1], u_col_out_591[1], u_col_out_590[1], u_col_out_589[1], u_col_out_588[1], u_col_out_587[1], u_col_out_586[1], u_col_out_585[1], u_col_out_584[1], u_col_out_583[1], u_col_out_582[1], u_col_out_581[1], u_col_out_580[1], u_col_out_579[1], u_col_out_578[1], u_col_out_577[1], u_col_out_576[1], u_col_out_575[1], u_col_out_574[1], u_col_out_573[1], u_col_out_572[1], u_col_out_571[1], u_col_out_570[1], u_col_out_569[1], u_col_out_568[1], u_col_out_567[1], u_col_out_566[1], u_col_out_565[1], u_col_out_564[1], u_col_out_563[1], u_col_out_562[1], u_col_out_561[1], u_col_out_560[1], u_col_out_559[1], u_col_out_558[1], u_col_out_557[1], u_col_out_556[1], u_col_out_555[1], u_col_out_554[1], u_col_out_553[1], u_col_out_552[1], u_col_out_551[1], u_col_out_550[1], u_col_out_549[1], u_col_out_548[1], u_col_out_547[1], u_col_out_546[1], u_col_out_545[1], u_col_out_544[1], u_col_out_543[1], u_col_out_542[1], u_col_out_541[1], u_col_out_540[1], u_col_out_539[1], u_col_out_538[1], u_col_out_537[1], u_col_out_536[1], u_col_out_535[1], u_col_out_534[1], u_col_out_533[1], u_col_out_532[1], u_col_out_531[1], u_col_out_530[1], u_col_out_529[1], u_col_out_528[1], u_col_out_527[1], u_col_out_526[1], u_col_out_525[1], u_col_out_524[1], u_col_out_523[1], u_col_out_522[1], u_col_out_521[1], u_col_out_520[1], u_col_out_519[1], u_col_out_518[1], u_col_out_517[1], u_col_out_516[1], u_col_out_515[1], u_col_out_514[1], u_col_out_513[1], u_col_out_512[1], u_col_out_511[1], u_col_out_510[1], u_col_out_509[1], u_col_out_508[1], u_col_out_507[1], u_col_out_506[1], u_col_out_505[1], u_col_out_504[1], u_col_out_503[1], u_col_out_502[1], u_col_out_501[1], u_col_out_500[1], u_col_out_499[1], u_col_out_498[1], u_col_out_497[1], u_col_out_496[1], u_col_out_495[1], u_col_out_494[1], u_col_out_493[1], u_col_out_492[1], u_col_out_491[1], u_col_out_490[1], u_col_out_489[1], u_col_out_488[1], u_col_out_487[1], u_col_out_486[1], u_col_out_485[1], u_col_out_484[1], u_col_out_483[1], u_col_out_482[1], u_col_out_481[1], u_col_out_480[1], u_col_out_479[1], u_col_out_478[1], u_col_out_477[1], u_col_out_476[1], u_col_out_475[1], u_col_out_474[1], u_col_out_473[1], u_col_out_472[1], u_col_out_471[1], u_col_out_470[1], u_col_out_469[1], u_col_out_468[1], u_col_out_467[1], u_col_out_466[1], u_col_out_465[1], u_col_out_464[1], u_col_out_463[1], u_col_out_462[1], u_col_out_461[1], u_col_out_460[1], u_col_out_459[1], u_col_out_458[1], u_col_out_457[1], u_col_out_456[1], u_col_out_455[1], u_col_out_454[1], u_col_out_453[1], u_col_out_452[1], u_col_out_451[1], u_col_out_450[1], u_col_out_449[1], u_col_out_448[1], u_col_out_447[1], u_col_out_446[1], u_col_out_445[1], u_col_out_444[1], u_col_out_443[1], u_col_out_442[1], u_col_out_441[1], u_col_out_440[1], u_col_out_439[1], u_col_out_438[1], u_col_out_437[1], u_col_out_436[1], u_col_out_435[1], u_col_out_434[1], u_col_out_433[1], u_col_out_432[1], u_col_out_431[1], u_col_out_430[1], u_col_out_429[1], u_col_out_428[1], u_col_out_427[1], u_col_out_426[1], u_col_out_425[1], u_col_out_424[1], u_col_out_423[1], u_col_out_422[1], u_col_out_421[1], u_col_out_420[1], u_col_out_419[1], u_col_out_418[1], u_col_out_417[1], u_col_out_416[1], u_col_out_415[1], u_col_out_414[1], u_col_out_413[1], u_col_out_412[1], u_col_out_411[1], u_col_out_410[1], u_col_out_409[1], u_col_out_408[1], u_col_out_407[1], u_col_out_406[1], u_col_out_405[1], u_col_out_404[1], u_col_out_403[1], u_col_out_402[1], u_col_out_401[1], u_col_out_400[1], u_col_out_399[1], u_col_out_398[1], u_col_out_397[1], u_col_out_396[1], u_col_out_395[1], u_col_out_394[1], u_col_out_393[1], u_col_out_392[1], u_col_out_391[1], u_col_out_390[1], u_col_out_389[1], u_col_out_388[1], u_col_out_387[1], u_col_out_386[1], u_col_out_385[1], u_col_out_384[1], u_col_out_383[1], u_col_out_382[1], u_col_out_381[1], u_col_out_380[1], u_col_out_379[1], u_col_out_378[1], u_col_out_377[1], u_col_out_376[1], u_col_out_375[1], u_col_out_374[1], u_col_out_373[1], u_col_out_372[1], u_col_out_371[1], u_col_out_370[1], u_col_out_369[1], u_col_out_368[1], u_col_out_367[1], u_col_out_366[1], u_col_out_365[1], u_col_out_364[1], u_col_out_363[1], u_col_out_362[1], u_col_out_361[1], u_col_out_360[1], u_col_out_359[1], u_col_out_358[1], u_col_out_357[1], u_col_out_356[1], u_col_out_355[1], u_col_out_354[1], u_col_out_353[1], u_col_out_352[1], u_col_out_351[1], u_col_out_350[1], u_col_out_349[1], u_col_out_348[1], u_col_out_347[1], u_col_out_346[1], u_col_out_345[1], u_col_out_344[1], u_col_out_343[1], u_col_out_342[1], u_col_out_341[1], u_col_out_340[1], u_col_out_339[1], u_col_out_338[1], u_col_out_337[1], u_col_out_336[1], u_col_out_335[1], u_col_out_334[1], u_col_out_333[1], u_col_out_332[1], u_col_out_331[1], u_col_out_330[1], u_col_out_329[1], u_col_out_328[1], u_col_out_327[1], u_col_out_326[1], u_col_out_325[1], u_col_out_324[1], u_col_out_323[1], u_col_out_322[1], u_col_out_321[1], u_col_out_320[1], u_col_out_319[1], u_col_out_318[1], u_col_out_317[1], u_col_out_316[1], u_col_out_315[1], u_col_out_314[1], u_col_out_313[1], u_col_out_312[1], u_col_out_311[1], u_col_out_310[1], u_col_out_309[1], u_col_out_308[1], u_col_out_307[1], u_col_out_306[1], u_col_out_305[1], u_col_out_304[1], u_col_out_303[1], u_col_out_302[1], u_col_out_301[1], u_col_out_300[1], u_col_out_299[1], u_col_out_298[1], u_col_out_297[1], u_col_out_296[1], u_col_out_295[1], u_col_out_294[1], u_col_out_293[1], u_col_out_292[1], u_col_out_291[1], u_col_out_290[1], u_col_out_289[1], u_col_out_288[1], u_col_out_287[1], u_col_out_286[1], u_col_out_285[1], u_col_out_284[1], u_col_out_283[1], u_col_out_282[1], u_col_out_281[1], u_col_out_280[1], u_col_out_279[1], u_col_out_278[1], u_col_out_277[1], u_col_out_276[1], u_col_out_275[1], u_col_out_274[1], u_col_out_273[1], u_col_out_272[1], u_col_out_271[1], u_col_out_270[1], u_col_out_269[1], u_col_out_268[1], u_col_out_267[1], u_col_out_266[1], u_col_out_265[1], u_col_out_264[1], u_col_out_263[1], u_col_out_262[1], u_col_out_261[1], u_col_out_260[1], u_col_out_259[1], u_col_out_258[1], u_col_out_257[1], u_col_out_256[1], u_col_out_255[1], u_col_out_254[1], u_col_out_253[1], u_col_out_252[1], u_col_out_251[1], u_col_out_250[1], u_col_out_249[1], u_col_out_248[1], u_col_out_247[1], u_col_out_246[1], u_col_out_245[1], u_col_out_244[1], u_col_out_243[1], u_col_out_242[1], u_col_out_241[1], u_col_out_240[1], u_col_out_239[1], u_col_out_238[1], u_col_out_237[1], u_col_out_236[1], u_col_out_235[1], u_col_out_234[1], u_col_out_233[1], u_col_out_232[1], u_col_out_231[1], u_col_out_230[1], u_col_out_229[1], u_col_out_228[1], u_col_out_227[1], u_col_out_226[1], u_col_out_225[1], u_col_out_224[1], u_col_out_223[1], u_col_out_222[1], u_col_out_221[1], u_col_out_220[1], u_col_out_219[1], u_col_out_218[1], u_col_out_217[1], u_col_out_216[1], u_col_out_215[1], u_col_out_214[1], u_col_out_213[1], u_col_out_212[1], u_col_out_211[1], u_col_out_210[1], u_col_out_209[1], u_col_out_208[1], u_col_out_207[1], u_col_out_206[1], u_col_out_205[1], u_col_out_204[1], u_col_out_203[1], u_col_out_202[1], u_col_out_201[1], u_col_out_200[1], u_col_out_199[1], u_col_out_198[1], u_col_out_197[1], u_col_out_196[1], u_col_out_195[1], u_col_out_194[1], u_col_out_193[1], u_col_out_192[1], u_col_out_191[1], u_col_out_190[1], u_col_out_189[1], u_col_out_188[1], u_col_out_187[1], u_col_out_186[1], u_col_out_185[1], u_col_out_184[1], u_col_out_183[1], u_col_out_182[1], u_col_out_181[1], u_col_out_180[1], u_col_out_179[1], u_col_out_178[1], u_col_out_177[1], u_col_out_176[1], u_col_out_175[1], u_col_out_174[1], u_col_out_173[1], u_col_out_172[1], u_col_out_171[1], u_col_out_170[1], u_col_out_169[1], u_col_out_168[1], u_col_out_167[1], u_col_out_166[1], u_col_out_165[1], u_col_out_164[1], u_col_out_163[1], u_col_out_162[1], u_col_out_161[1], u_col_out_160[1], u_col_out_159[1], u_col_out_158[1], u_col_out_157[1], u_col_out_156[1], u_col_out_155[1], u_col_out_154[1], u_col_out_153[1], u_col_out_152[1], u_col_out_151[1], u_col_out_150[1], u_col_out_149[1], u_col_out_148[1], u_col_out_147[1], u_col_out_146[1], u_col_out_145[1], u_col_out_144[1], u_col_out_143[1], u_col_out_142[1], u_col_out_141[1], u_col_out_140[1], u_col_out_139[1], u_col_out_138[1], u_col_out_137[1], u_col_out_136[1], u_col_out_135[1], u_col_out_134[1], u_col_out_133[1], u_col_out_132[1], u_col_out_131[1], u_col_out_130[1], u_col_out_129[1], u_col_out_128[1], u_col_out_127[1], u_col_out_126[1], u_col_out_125[1], u_col_out_124[1], u_col_out_123[1], u_col_out_122[1], u_col_out_121[1], u_col_out_120[1], u_col_out_119[1], u_col_out_118[1], u_col_out_117[1], u_col_out_116[1], u_col_out_115[1], u_col_out_114[1], u_col_out_113[1], u_col_out_112[1], u_col_out_111[1], u_col_out_110[1], u_col_out_109[1], u_col_out_108[1], u_col_out_107[1], u_col_out_106[1], u_col_out_105[1], u_col_out_104[1], u_col_out_103[1], u_col_out_102[1], u_col_out_101[1], u_col_out_100[1], u_col_out_99[1], u_col_out_98[1], u_col_out_97[1], u_col_out_96[1], u_col_out_95[1], u_col_out_94[1], u_col_out_93[1], u_col_out_92[1], u_col_out_91[1], u_col_out_90[1], u_col_out_89[1], u_col_out_88[1], u_col_out_87[1], u_col_out_86[1], u_col_out_85[1], u_col_out_84[1], u_col_out_83[1], u_col_out_82[1], u_col_out_81[1], u_col_out_80[1], u_col_out_79[1], u_col_out_78[1], u_col_out_77[1], u_col_out_76[1], u_col_out_75[1], u_col_out_74[1], u_col_out_73[1], u_col_out_72[1], u_col_out_71[1], u_col_out_70[1], u_col_out_69[1], u_col_out_68[1], u_col_out_67[1], u_col_out_66[1], u_col_out_65[1], u_col_out_64[1], u_col_out_63[1], u_col_out_62[1], u_col_out_61[1], u_col_out_60[1], u_col_out_59[1], u_col_out_58[1], u_col_out_57[1], u_col_out_56[1], u_col_out_55[1], u_col_out_54[1], u_col_out_53[1], u_col_out_52[1], u_col_out_51[1], u_col_out_50[1], u_col_out_49[1], u_col_out_48[1], u_col_out_47[1], u_col_out_46[1], u_col_out_45[1], u_col_out_44[1], u_col_out_43[1], u_col_out_42[1], u_col_out_41[1], u_col_out_40[1], u_col_out_39[1], u_col_out_38[1], u_col_out_37[1], u_col_out_36[1], u_col_out_35[1], u_col_out_34[1], u_col_out_33[1], u_col_out_32[1], u_col_out_31[1], u_col_out_30[1], u_col_out_29[1], u_col_out_28[1], u_col_out_27[1], u_col_out_26[1], u_col_out_25[1], u_col_out_24[1], u_col_out_23[1], u_col_out_22[1], u_col_out_21[1], u_col_out_20[1], u_col_out_19[1], u_col_out_18[1], u_col_out_17[1], u_col_out_16[1], u_col_out_15[1], u_col_out_14[1], u_col_out_13[1], u_col_out_12[1], u_col_out_11[1], u_col_out_10[1], u_col_out_9[1], u_col_out_8[1], u_col_out_7[1], u_col_out_6[1], u_col_out_5[1], u_col_out_4[1], u_col_out_3[1], u_col_out_2[1], u_col_out_1[1], u_col_out_0[1]};


endmodule



module xpb_5_725
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h72cdcd0336923806de61c9f428806e3384eed7dca4358e5516d34de2c06e914db1fede9bd16b7fad8de3ab037627f2daf7f313cbdf643c907d157d1e868c3e7f255f463a754d519537502b2d6e8793ff7eb4f5c3852d040a23ececa0e2ad90132de29de90529c8676ee659d02ae0a2e1c41e25cadd48abf3e81e812d3ee4b8ff;
    5'b00010 : xpb = 1024'h34ee54b0ab363b44f1be1c1140a695159867ac8872f37c32afc9e26fcdda759360b53fbed8b080cc7c6916c008f1d4eb8bcbffb19c15a8d5498bbaded246084cd66f57c63b09a5e55c0653b8443363ce0964f1ee7dd3db03924d47470b307d942cbda9a8598a9841570cccc15df11f9a39626cb36a45fab789cd8755f4e70b93;
    5'b00011 : xpb = 1024'ha7bc21b3e1c8734bd01fe605692703491d56846517290a87c69d30528e4906e112b41e5aaa1c007a0a4cc1c37f19c7c683bf137d7b79e565c6a137fd58d246cbfbce9e00b056f77a93567ee5b2baf7cd8819e7b20300df0db63a33e7edde0da75aa047915eb460a8c5f3269188d1c27bfd80927e478ea6ab71ec088333cbc492;
    5'b00100 : xpb = 1024'h69dca961566c7689e37c3822814d2a2b30cf5910e5e6f8655f93c4df9bb4eb26c16a7f7db1610198f8d22d8011e3a9d71797ff63382b51aa931775bda48c1099acdeaf8c76134bcab80ca7708866c79c12c9e3dcfba7b607249a8e8e1660fb28597b5350b3153082ae199982bbe23f3472c4d966d48bf56f139b0eabe9ce1726;
    5'b00101 : xpb = 1024'h2bfd310ecb1079c7f6d88a3f9973510d44482dbcb4a4e642f88a596ca920cf6c7020e0a0b8a602b7e757993ca4ad8be7ab70eb48f4dcbdef5f8db37df045da675deec1183bcfa01adcc2cffb5e12976a9d79e007f44e8d0092fae9343ee3e8a958565f100776005c96400c73eef2bbece809204f61894432b54a14d49fd069ba;
    5'b00110 : xpb = 1024'h9ecafe1201a2b1ced53a5433c1f3bf40c937059958da74980f5da74f698f60ba221fbf3c8a118265753b44401ad57ec2a363ff14d440fa7fdca3309c76d218e6834e0752b11cf1b01412fb28cc9a2b6a1c2ed5cb797b910ab6e7d5d5219178bc8638fcf90c9fc8c40526664419d35eceac27461a3ed1f0269d689601deb522b9;
    5'b00111 : xpb = 1024'h60eb85bf7646b50ce896a650da19e622dcafda4527986275a8543bdc76fb44ffd0d6205f9156838463c0affcad9f60d3373ceafa90f266c4a9196e5cc28be2b4345e18de76d9460038c923b3a245fb38a6ded1f6722268042548307b4a14663d851408b86100989ded4cd9354ce3db87216b8d02cbcf3eea3f179c2a94b7754d;
    5'b01000 : xpb = 1024'h230c0d6ceaeab84afbf2f86df2400d04f028aef0f6565053414ad069846729457f8c8182989b84a352461bb9406942e3cb15d6e04da3d309758fac1d0e45ac81e56e2a6a3c959a505d7f4c3e77f1cb07318ece216ac93efd93a88b21729753be83ef1477b5616877d5734c267ff4583f96afd3eb58cc8dade0c6a2534ab9c7e1;
    5'b01001 : xpb = 1024'h95d9da70217cf051da54c2621ac07b38751786cd9a8bdea8581e1e4c44d5ba93318b601e6a070450e029c6bcb69135bec308eaac2d080f99f2a5293b94d1eb010acd70a4b1e2ebe594cf776be6795f06b043c3e4eff64307b79577c25544e3d1b1d1b260ba8b30df4459a5f6aad4fb215acdf9b6361539a1c8e52380899e80e0;
    5'b01010 : xpb = 1024'h57fa621d9620f38fedb1147f32e6a21a88905b796949cc85f114b2d952419ed8e041c141714c056fceaf3279495b17cf56e1d691e9b97bdebf1b66fbe08bb4cebbdd8230779f4035b9859ff6bc252ed53af3c00fe89d1a0125f5d2687dc7d152b0acbe200eec00b92c8018e7dde577d9d012409ec31288656a9429a93fa0d374;
    5'b01011 : xpb = 1024'h1a1ae9cb0ac4f6ce010d669c4b0cc8fc9c0930253807ba638a0b47665fad831e8ef822647891068ebd349e35dc24f9dfeabac277a66ae8238b91a4bc2c457e9c6ced93bc3d5b9485de3bc88191d0fea3c5a3bc3ae143f0fa94562d0ea64abed3af87c9df634cd09314a68bd910f5f49245568787500fd7290c432fd1f5a32608;
    5'b01100 : xpb = 1024'h8ce8b6ce41572ed4df6f3090738d373020f80801dc3d48b8a0de9549201c146c40f7010049fc863c4b184939524cecbae2add64385cf24b408a721dab2d1bd1b924cd9f6b2a8e61b158bf3af005892a34458b1fe6670f504b84319af88f84ee6dd6a67c8687698fa838ce5a93bd697740974ad522d58831cf461b0ff3487df07;
    5'b01101 : xpb = 1024'h4f093e7bb5fb3212f2cb82ad8bb35e123470dcadaafb369639d529d62d87f8b1efad62235141875b399db4f5e516cecb7686c229428090f8d51d5f9afe8b86e9435ceb8278653a6b3a421c39d6046271cf08ae295f17cbfe26a37455b17b3c67dc457387bcd768d46bb3589a6ee7142c7eb8f43aba55d1e09610b727ea8a319b;
    5'b01110 : xpb = 1024'h1129c6292a9f35510627d4caa3d984f447e9b15979b92473d2cbbe633af3dcf79e63c3465886887a282320b277e0b0dc0a5fae0eff31fd3da1939d5b4a4550b6f46cfd0e3e218ebb5ef844c4abb0324059b8aa5457bea2f79503cefbd9fe29e8db207f47113838ae53d9cb8ba1f790e4f3fd3b23475320a437bfbd50a08c842f;
    5'b01111 : xpb = 1024'h83f7932c61316d57e4899ebecc59f327ccd889361deeb2c8e99f0c45fb626e455062a1e229f20827b606cbb5ee08a3b70252c1dade9639ce1ea91a79d0d18f3619cc4348b36ee05096486ff21a37c63fd86da017dceba701b8f0bb9cbcabb9fc09031d3016620115c2c0255bccd833c6b81b60ee249bcc981fde3e7ddf713d2e;
    5'b10000 : xpb = 1024'h46181ad9d5d57095f7e5f0dbe4801a09e0515de1ecaca0a68295a0d308ce528aff19030531370946a48c377280d285c7962badc09b47a612eb1f583a1c8b5903cadc54d4792b34a0bafe987cefe3960e631d9c42d5927dfb27511642e52ea77d07de28ef6ac2d0efaae6984cffe8b07f2d5fa7d6b1991b5bc18d44a695738fc2;
    5'b10001 : xpb = 1024'h838a2874a7973d40b4242f8fca640ebf3ca328dbb6a8e841b8c3560163a36d0adcf6428387c0a659311a32f139c67d82a0499a657f91257b79595fa684522d17bec66603ee788f0dfb4c107c58f65dcedcd986dce3954f495b170e90db194fe06b934aebf23a0c9930d0b3e32f92d37a2a3eebf3e966a1f633c4acf4b75e256;
    5'b10010 : xpb = 1024'h7b066f8a810babdae9a40ced2526af1f78b90a6a5fa01cd9325f8342d6a8c81e5fce42c409e78a1320f54e3289c45ab321f7ad72375d4ee834ab1318eed16150a14bac9ab434da861704ec353416f9dc6c828e31536658feb99e5d89f05f2511349bd297c44d693101f3650e5dd9d01966c2148a1bdf16134b5acbfc8a5a9b55;
    5'b10011 : xpb = 1024'h3d26f737f5afaf18fd005f0a3d4cd6018c31df162e5e0ab6cb5617cfe414ac640e84a3e7112c8b320f7ab9ef1c8e3cc3b5d09957f40ebb2d012150d93a8b2b1e525bbe2679f12ed63bbb14c009c2c9aaf7328a5c4c0d2ff827feb83018e212923376de5718ae390aea19d7ff90ea4cd1dc065b72a8dc64d6ed09d225405cede9;
    5'b10100 : xpb = 1024'haff4c43b2c41e71fdb6228fe65cd44351120b6f2d293990be22965b2a4833db1c0838282e2980adf9d5e64f292b62f9eadc3ad23d372f7bd7e36cdf7c117699d77bb0460ef3e806b730b3fed784a5daa75e7801fd13a34024beba4d0fb8fa2a561597c401dd80172590031cfbbcaefb3a024813d862510cad52853527f41a6e8;
    5'b10101 : xpb = 1024'h72154be8a0e5ea5deebe7b1b7df36b1724998b9ea15186e97b1ffa3fb1ef21f76f39e3a5e9dd0bfe8be3d0af258011af419c9909902464024aad0bb80cd1336b28cb15ecb4fad4bb97c168784df62d7900977c4ac9e10afbba4bff7724129026603487ff7238d14c4126a4c0eedb6c6c1568c82613225f8e76d7597b3543f97c;
    5'b10110 : xpb = 1024'h3435d3961589ed9c021acd38961991f93812604a700f74c714168eccbf5b063d1df044c8f1220d1d7a693c6bb849f3bfd57584ef4cd5d04717234978588afd38d9db27787ab7290bbc77910323a1fd478b477875c287e1f528ac5a1d4c957da75f0f93bec699a126294d17b221ebe9248aad0f0ea01fae5218865fa3eb464c10;
    5'b10111 : xpb = 1024'ha703a0994c1c25a2e07c972cbe9a002cbd0138271445031c2ae9dcaf7fc9978acfef2364c28d8ccb084ce76f2e71e69acd6898bb2c3a0cd79438c696df173bb7ff3a6db2f0047aa0f3c7bc309229914709fc6e3947b4e5ff4c9946be2f430dba8cf231a7cbc3698d983371824ccc8c064ecb34d97d685a4600a4e0d12a2b050f;
    5'b11000 : xpb = 1024'h69242846c0c028e0f3d8e949d6c0270ed07a0cd2e302f0f9c3e0713c8d357bd07ea58487c9d28de9f6d2532bc13bc8ab614184a0e8eb791c60af04572ad10585b04a7f3eb5c0cef1187de4bb67d5611594ac6a64405bbcf8baf9a16457c5fb3b8bcd3d67202439678059e4737fdd08bec40f7bc20a65a909a253e6f9e02d57a3;
    5'b11001 : xpb = 1024'h2b44aff435642c1f07353b66eee64df0e3f2e17eb1c0ded75cd705c99aa160162d5be5aad1178f08e557bee85405aabbf51a7086a59ce5612d254217768acf53615a90ca7b7d23413d340d463d8130e41f5c668f390293f22959fc0a8048e8bc8aa849267485094168805764b2ed85773953c2aa9762f7cd4402ed22962faa37;
    5'b11010 : xpb = 1024'h9e127cf76bf66425e597055b1766bc2468e1b95b55f66d2c73aa53ac5b0ff163df5ac446a2830eb6733b69ebca2d9d96ed0d8452850121f1aa3abf35fd170dd286b9d704f0ca74d674843873ac08c4e39e115c52be2f97fc4d46e8ab62f678cfb88ae70f79aed1a8d766b134ddce2858fd71e87574aba3c12c216e4fd5146336;
    5'b11011 : xpb = 1024'h603304a4e09a6763f8f357782f8ce3067c5a8e0724b45b0a0ca0e839687bd5a98e112569a9c80fd561c0d5a85cf77fa780e6703841b28e3676b0fcf648d0d7a037c9e890b686c926993a60fe81b494b228c1587db6d66ef5bba743518b796650b765f2cece0fa182bf8d242610dea51172b62f5e01a8f284cdd074788b16b5ca;
    5'b11100 : xpb = 1024'h22538c52553e6aa20c4fa99547b309e88fd362b2f37248e7a5977cc675e7b9ef3cc7868cb10d10f450464164efc161b814bf5c1dfe63fa7b43273ab6948aa16de8d9fa1c7c431d76bdf0898957606480b37154a8af7d45ef2a079df7b3fc53d1b640fe8e2270715ca7b3971743ef21c9e7fa76468ea641486f7f7aa14119085e;
    5'b11101 : xpb = 1024'h952159558bd0a2a8eab173897033781c14c23a8f97a7d73cbc6acaa936564b3ceec66528827890a1de29ec6865e954930cb26fe9ddc8370bc03cb7d51b16dfed0e394056f1906f0bf540b4b6c5e7f88032264a6c34aa49f94df48a9896a9e3e4e4239c77279a39c41699f0e76ecfc4abac189c116beeed3c579dfbce7ffdc15d;
    5'b11110 : xpb = 1024'h5741e1030074a5e6fe0dc5a688599efe283b0f3b6665c51a55615f3643c22f829d7cc64b89bd91c0ccaf5824f8b336a3a08b5bcf9a79a3508cb2f59566d0a9babf4951e2b74cc35c19f6dd419b93c84ebcd646972d5120f2bc54e53ebf2cd165e2fea8367bfb099dfec063d8a1e04164215ce2f9f8ec3bfff94d01f7360013f1;
    5'b11111 : xpb = 1024'h196268b07518a925116a17c3a07fc5e03bb3e3e73523b2f7ee57f3c3512e13c84c33276e910292dfbb34c3e18b7d18b4346447b5572b0f9559293355b28a73887059636e7d0917ac3ead05cc713f981d478642c225f7f7ec2ab53fe4e7afbee6e1d9b3f5d05bd977e6e6d6c9d4f0be1c96a129e285e98ac39afc081fec026685;
    endcase
end

endmodule

module xpb_5_835
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h83a33ec5ce5ea065a45ff9b7765ef8956a3fedf3c7a72ab3f6708a0a6ca87ad2a33ceb7f87e08956b6e5f8607a48d38cffbd73ccb1b559986cc840ca1f05a0b6be6125f89bafa32df2c953d7b97858ae2a44d945b778d15d54a1544236c4cea8c06f12d9e1fd8ac2ffe746b80ea6aad531f2ce120465e32be561e13da16399cc;
    5'b00010 : xpb = 1024'h56993835dacf0c027dba7b97dc63a9d96309d8b6b9d6b4f06f045abf264e489d43315986459a941ece6db17a1133964f9b60bfb340b7e2e528f142360338ccbc0873174287ce4916d2f8a50cda14ed2b6084b8f2e26b75a9f3b61689b35efabf51d6938a13321cf8790ea691257d2f81150bbd41b880692784544776b9e4cd2d;
    5'b00011 : xpb = 1024'h298f31a5e73f779f5714fd7842685b1d5bd3c379ac063f2ce7982b73dff41667e325c78d03549ee6e5f56a93a81e591237040b99cfba6c31e51a43a1e76bf8c15285088c73eceeffb327f641fab181a896c498a00d5e19f692cad8d12ff926d5e33e143a4466af2df236066a3c53b42cf824ac716c9aef232346adafd266008e;
    5'b00100 : xpb = 1024'had32706bb59e1804fb74f72fb8c753b2c613b16d73ad69e0de08b57e4c9c913a8662b30c8b35283d9cdb62f422672c9f36c17f66816fc5ca51e2846c0671997810e62e850f9c922da5f14a19b429da56c10971e5c4d6eb53e76c2d1366bdf57ea3ad2714266439f0f21d4d224afa5f022a177a837100d24f08a88eed73c99a5a;
    5'b00101 : xpb = 1024'h802869dbc20e83a1d4cf79101ecc04f6bedd9c3065dcf41d569c863306425f052657211348ef3305b4631c0db951ef61d264cb4d10724f170e0b85d7eaa4c57d5af81fcefbbb381686209b4ed4c66ed3f7495192efc98fa08680ef5ae35821953514a7c45798cc266b44acfb61d0e3ae0d3069b3251b584aa79af5268c4acdbb;
    5'b00110 : xpb = 1024'h531e634bce7eef3eae29faf084d0b63ab7a786f3580c7e59cf3056e7bfe82ccfc64b8f1a06a93dcdcbead527503cb2246e0817339f74d863ca348743ced7f182a50a1118e7d9ddff664fec83f56303512d8931401abc33ed2595b1a25ff24dabc67c287488cd5e5be46c0cd478a76859f04958e2d935de46468d5b5fa4cc011c;
    5'b00111 : xpb = 1024'h26145cbbdaef5adb87847cd0ead5677eb07171b64a3c089647c4279c798dfa9a663ffd20c4634895e3728e40e72774e709ab631a2e7761b0865d88afb30b1d87ef1c0262d3f883e8467f3db915ff97ce63c910ed45aed839c4aa73e9dc8c79c257e3a924ba01f0915d936cad8f7ded05d36248128d506441e57fc198bd4d347d;
    5'b01000 : xpb = 1024'ha9b79b81a94dfb412be47688613460141ab15faa11e3334a3e34b1a6e636756d097ce8a04c43d1ec9a5886a1617048740968d6e6e02cbb48f325c979d210be3ead7d285b6fa8271639489190cf77f07c8e0dea32fd27a997194bc82c1351486b1852bbfe9bff7b545d7ab3659e2497db0555162491b6476dcae1a2d65eb0ce49;
    5'b01001 : xpb = 1024'h7cad94f1b5be66de053ef868c7391158137b4a6d0412bd86b6c8825b9fdc4337a97156a709fddcb4b1e03fbaf85b0b36a50c22cd6f2f4495af4ecae5b643ea43f78f19a55bc6ccff1977e2c5f01484f9c44dc9e0281a4de3b8608a738feb7481a9ba3caecd340d89d6a2133eb4fb1c86e86e055445d0cd6969d4090f773201aa;
    5'b01010 : xpb = 1024'h4fa38e61c22ed27ade997a492d3dc29c0c45352ff64247c32f5c5310598211024965c4adc7b7e77cc967f8d48f45cdf940af6eb3fe31cde26b77cc519a77164941a10aef47e572e7f9a733fb10b11976fa8da98d530cf23057754cbb0c85a0983b21bd5efe689fbf4fc97317cbd1a132cb86f483f9eb536508c66f488fb3350b;
    5'b01011 : xpb = 1024'h229987d1ce9f3e17b7f3fc29934273e0050f1ff2e871d1ffa7f023c51327decce95a32b48571f244e0efb1ee263090bbdc52ba9a8d34572f27a0cdbd7eaa424e8bb2fc39340418d0d9d68530314dadf430cd893a7dff967cf68a0f02891fccaecc893e0f2f9d31f4c8f0d2f0e2a825deae9fe3b3ae05d960a7b8d581a834686c;
    5'b01100 : xpb = 1024'ha63cc6979cfdde7d5c53f5e109a16c756f4f0de6b018fcb39e60adcf7fd0599f8c971e340d527b9b97d5aa4ea0796448dc102e673ee9b0c794690e879dafe3054a142231cfb3bbfecc9fd907eac606a25b126280357867da4b2b6344bfe49b578cf850e9119abcb7c8d819a8f14ed0b3e092b1c5b26bbc8c8d1ab6bf49980238;
    5'b01101 : xpb = 1024'h7932c007a96e4a1a35ae77c16fa61db96818f8a9a24886f016f47e843976276a2c8b8c3acb0c8663af5d63683764270b77b37a4dcdec3a1450920ff381e30f0a9426137bbbd261e7accf2a3d0b629b1f9152422d606b0c26ea40258c3c7ec76e1e5fd19942cf4eed41ff79820825555fc3aba0f5668642882c0d1cf862193599;
    5'b01110 : xpb = 1024'h4c28b977b5deb5b70f08f9a1d5aacefd60e2e36c9478112c8f884f38f31bf534cc7ffa4188c6912bc6e51c81ce4ee9ce1356c6345ceec3610cbb115f66163b0fde3804c5a7f107d08cfe7b722bff2f9cc79221da8b5db0738954e7d3b918f384afc752497403e122bb26d95b1efbda0ba6c490251aa0c883caff83317a9a68fa;
    5'b01111 : xpb = 1024'h1f1eb2e7c24f2153e8637b823baf804159acce2f86a79b69081c1fedacc1c2ff6c74684846809bf3de6cd59b6539ac90aefa121aebf14cadc8e412cb4a4967152849f60f940fadb96d2dcca74c9bc419fdd20187b65054c02869aa1b35b31f9b412ed2f9a5387358344e393435d25eb789dd7f54cebb4e7f69f1e96a931b9c5b;
    5'b10000 : xpb = 1024'ha2c1f1ad90adc1b98cc37539b20e78d6c3ecbc234e4ec61cfe8ca9f8196a3dd20fb153c7ce61254a9552cdfbdf82801daeb785e79da6a64635ac5395694f07cbe6ab1c082fbf50e75ff7207f06141cc82816dacd6dc9261d7d0afe5d6c77ee44019de5d38735fe1b34357fec4479098cbbd04d66d32131ab4f53caa8347f3627;
    5'b10001 : xpb = 1024'h75b7eb1d9d1e2d56661df71a18132a1abcb6a6e6407e505977207aacd3100b9cafa5c1ce8c1b3012acda8715766d42e04a5ad1ce2ca92f92f1d555014d8233d130bd0d521bddf6d0402671b426b0b1455e56ba7a98bbca6a1c1fc0a4e9121a5a93056683b86a9050ad5cdfc55b4f8e389ee93c96873bb7a6ee4630e14d006988;
    5'b10010 : xpb = 1024'h48ade48da98e98f33f7878fa7e17db5eb58091a932adda95efb44b618cb5d9674f9a2fd549d53adac462402f0d5805a2e5fe1db4bbabb8dfadfe566d31b55fd67acefe9c07fc9cb92055c2e9474d45c294969a27c3ae6eb6bb3482ec65ac4671246ce733e99f228626843f9e722612e482022bc63b563da28d38971a65819ce9;
    5'b10011 : xpb = 1024'h1ba3ddfdb5ff049018d2fadae41c8ca2ae4a7c6c24dd64d268481c16465ba731ef8e9ddc078f45a2dbe9f948a442c86581a1699b4aae422c6a2757d915e88bdbc4e0efe5f41b42a20085141e67e9da3fcad679d4eea113035a494533e2467287b5d467e41ad3b4bb9fab9f7788fc9790651b1af5ef70c39e2c2afd537e02d04a;
    5'b10100 : xpb = 1024'h9f471cc3845da4f5bd32f4925a7b8538188a6a5fec848f865eb8a620b304220492cb895b8f6fcef992cff1a91e8b9bf2815edd67fc639bc4d6ef98a334ee2c92834215de8fcae5cff34e67f6216232edf51b531aa619e460aeea9976190b413076437abdfcd13f7e9f92e62f97a34265970de907f3d6a6ca118cde911f666a16;
    5'b10101 : xpb = 1024'h723d163390ce1092968d7672c080367c11545522deb419c2d74c76d56ca9efcf32bff7624d29d9c1aa57aac2b5765eb51d02294e8b66251193189a0f19215897cd5407287be98bb8d37db92b41fec76b2b5b32c7d10c88ad4dff5bbd95a56d4707aafb6e2e05d1b418ba4608ae79c7117a26d837a7f12cc5b07f44ca37e79d77;
    5'b10110 : xpb = 1024'h45330fa39d3e7c2f6fe7f8532684e7c00a1e3fe5d0e3a3ff4fe0478a264fbd99d2b465690ae3e489c1df63dc4c612177b8a575351a68ae5e4f419b7afd54849d1765f872680831a1b3ad0a60629b5be8619b1274fbff2cf9ed141e05123f995d99127c1e5f3a63e991e1a5e1c5504bbd5d3fc7675c0bb2c14f71ab035068d0d8;
    5'b10111 : xpb = 1024'h18290913a9aee7cc49427a338c89990402e82aa8c3132e3bc874183edff58b6472a8d36fc89def51d9671cf5e34be43a5448c11ba96b37ab0b6a9ce6e187b0a26177e9bc5426d78a93dc5b958337f06597daf22226f1d1468c28e04c8ed9c5742a79fcce906ef61f0b0905badc26d0694058b697102638bcee64113c68ea0439;
    5'b11000 : xpb = 1024'h9bcc47d9780d8831eda273eb02e891996d28189c8aba58efbee4a2494c9e063715e5beef507e78a8904d15565d94b7c7540634e85b2091437832ddb1008d51591fd90fb4efd67ab886a5af6d3cb04913c21fcb67de6aa2a3e0ca348ec59e941ceae90fa8726c80e20af04c72eacd7b3e724b84a9148c1be8d3c5f27a0a4d9e05;
    5'b11001 : xpb = 1024'h6ec24149847df3cec6fcf5cb68ed42dd65f2035f7ce9e32c377872fe0643d401b5da2cf60e388370a7d4ce6ff47f7a89efa980ceea231a90345bdf1ce4c07d5e69eb00fedbf520a166d500a25d4cdd90f85fab15095d46f07fdef6d64238c0337c509058a3a113178417ac4c01a3ffea556473d8c8a6a1e472b858b322ced166;
    5'b11010 : xpb = 1024'h41b83ab990ee5f6ba05777abcef1f4215ebbee226f196d68b00c43b2bfe9a1cc55ce9afccbf28e38bf5c87898b6a3d4c8b4cccb57925a3dcf084e088c8f3a963b3fcf248c813c68a470451d77de9720e2e9f8ac2344feb3d1ef3b91dbed2ec4a0db81108d4d5a54cfd3f0c25187a8496387d63087cc127e011aabeec3b5004c7;
    5'b11011 : xpb = 1024'h14ae34299d5ecb0879b1f98c34f6a5655785d8e56148f7a528a01467798f6f96f5c3090389ac9900d6e440a32255000f26f0189c08282d29acade1f4ad26d568fe0ee392b4326c732733a30c9e86068b64df6a6f5f428f89be087b653b6d18609f1f91b9060a378276666bfe2f5109421b96523830dbaddbb09d252553d13828;
    5'b11100 : xpb = 1024'h985172ef6bbd6b6e1e11f343ab559dfac1c5c6d928f022591f109e71e637ea6998fff483118d22578dca39039c9dd39c26ad8c68b9dd86c2197622becc2c761fbc70098b4fe20fa119fcf6e457fe5f398f2443b516bb60e712a9cfa77231e7095f8ea492e807c245764db2b63df7b4174d89204a3541910795ff0662f534d1f4;
    5'b11101 : xpb = 1024'h6b476c5f782dd70af76c7524115a4f3eba8fb19c1b1fac9597a46f269fddb83438f46289cf472d1fa551f21d3388965ec250d84f48e0100ed59f242ab05fa2250681fad53c00b589fa2c4819789af3b6c564236241ae0533b1be91eeeecc131ff0f62543193c547aef75128f54ce38c330a20f79e95c170334f16c9c0db60555;
    5'b11110 : xpb = 1024'h3e3d65cf849e42a7d0c6f704775f0082b3599c5f0d4f36d210383fdb598385fed8e8d0908d0137e7bcd9ab36ca7359215df42435d7e2995b91c825969492ce2a5093ec1f281f5b72da5b994e99378833fba4030f6ca0a98050d354366b663f36825da5f34a70e6b0689c72686ba4bd6f13bafea99d769cfed3e3d2d5263738b6;
    5'b11111 : xpb = 1024'h11335f3f910eae44aa2178e4dd63b1c6ac238721ff7ec10e88cc1090132953c978dd3e974abb42afd4616450615e1be3f997701c66e522a84df1270278c5fa2f9aa5dd69143e015bba8aea83b9d41cb131e3e2bc97934dccefe8167de8006b4d13c526a37ba578e5e1c3d241827b421af6d3edd9519122fa72d6390e3eb86c17;
    endcase
end

endmodule

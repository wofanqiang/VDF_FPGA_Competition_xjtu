module xpb_5_815
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha8088772548a740a1d3b18e0e2a93007a938118b5df94f706ff7df0c860e138eed5a890722cca66e1a302c91414ef391267ebf4bc3df875dbe3fefaf58f2e04bcad7ab93311a2957fe74a86bad2a49568b73a8edcf448d0e581c9b7580f8a583e094999e475035a264e32de826307061c6ab61cdbf3a5992c2c40fa02d6adafa;
    5'b00010 : xpb = 1024'h9f63c98ee726b34b6f70b9eab4f818bde0fa1fe5e67afe69621304c359197a15d76c94957b72ce4d950219db9f3fd657e8e356b1650c3e6fcbe0a00077134be621602277b2a3556aea4f4e34c178ce7c22e258431202ed0bfaaca4f047c6a8759221a112ddd772b7430674f15490ba9a3e7ce4b92e2955f53f18a43bd1f34f89;
    5'b00011 : xpb = 1024'h96bf0bab79c2f28cc1a65af48747017418bc2e406efcad62542e2a7a2c24e09cc17ea023d418f62d0fd40725fd30b91eab47ee170638f581d98150519533b78077e8995c342c817dd629f3fdd5c753a1ba51079854c14d099d3cae6b0e94ab6743aea887745eafcc2129bbfa82f104d2b64e67a49d185257bb6d38d7767bc418;
    5'b00100 : xpb = 1024'h8e1a4dc80c5f31ce13dbfbfe5995ea2a507e3c9af77e5c5b46495030ff304723ab90abb22cbf1e0c8aa5f4705b219be56dac857ca765ac93e72200a2b354231ace711040b5b5ad90c20499c6ea15d8c751bfb6ed977fad073fccb7e5d562ae58f53baffc0ae5ece0ff4d0303b1514f0b2e1fea900c074eba37c1cd731b0438a7;
    5'b00101 : xpb = 1024'h85758fe49efb710f66119d082be4d2e088404af580000b54386475e7d23badaa95a2b740856545ec0577e1bab9127eac30111ce2489263a5f4c2b0f3d1748eb524f98725373ed9a3addf3f8ffe645dece92e6642da3e0d04e25cc1609c30b14aa6c8b770a16d29f5dd704a0cdfb19943a5f16d7b7af64b1cb416620ebf8cad36;
    5'b00110 : xpb = 1024'h7cd0d2013197b050b8473e11fe33bb96c00259500881ba4d2a7f9b9ea54714317fb4c2cede0b6dcb8049cf0517036172f275b447e9bf1ab802636144ef94fa4f7b81fe09b8c805b699b9e55912b2e312809d15981cfc6d0284eccadb62feb43c5855bee537f4670abb9391160e11e37c1dc2f066e9e5477f306af6aa641521c5;
    5'b00111 : xpb = 1024'h742c141dc433ef920a7cdf1bd082a44cf7c467aa910369461c9ac15578527ab869c6ce5d36b195aafb1bbc4f74f44439b4da4bad8aebd1ca100411960db565e9d20a74ee3a5131c985948b2227016838180bc4ed5fbacd00277cd45629ccb72e09e2c659ce7ba41f99b6d81f3c722db49594735258d443e1acbf8b46089d9654;
    5'b01000 : xpb = 1024'h6b87563a56d02ed35cb28025a2d18d032f8676051985183f0eb5e70c4b5de13f53d8d9eb8f57bd8a75eda999d2e52700773ee3132c1888dc1da4c1e72bd5d1842892ebd2bbda5ddc716f30eb3b4fed5daf7a7442a2792cfdca0cddd0f09aba1fbb6fcdce6502e13477da1f286ad277ed0d65f63dc7c3404429141fe1ad260ae3;
    5'b01001 : xpb = 1024'h62e29856e96c6e14aee8212f752075b96748845fa206c73800d10cc31e6947c63deae579e7fde569f0bf96e430d609c739a37a78cd453fee2b45723849f63d1e7f1b62b73d6389ef5d49d6b44f9e728346e92397e5378cfb6c9ce74bb768bd116cfcd542fb8a1e4955fd66319932c2258537792936b23ca6a568b47d51ae7f72;
    5'b01010 : xpb = 1024'h5a3dda737c08ad56011dc239476f5e6f9f0a92ba2a887630f2ec3279f174ae4d27fcf10840a40d496b91842e8ec6ec8dfc0811de6e71f70038e622896816a8b8d5a3d99bbeecb60249247c7d63ecf7a8de57d2ed27f5ecf90f2cf0c67e36c0031e89dcb792115b5e3420ad3ac7930c5dfd08fc14a5a1390921bd4918f636f401;
    5'b01011 : xpb = 1024'h51991c900ea4ec975353634319be4725d6cca114b30a2529e5075830c48014d4120efc96994a3528e6637178ecb7cf54be6ca9440f9eae124686d2da863714532c2c50804075e21534ff2246783b7cce75c682426ab44cf6b1bcfa414504c2f4d016e42c289898731243f443f5f3569674da7f001490356b9e11ddb49abf6890;
    5'b01100 : xpb = 1024'h48f45eaca1412bd8a589044cec0d2fdc0e8eaf6f3b8bd422d7227de7978b7b5afc210824f1f05d0861355ec34aa8b21b80d140a9b0cb65245427832ba4577fed82b4c764c1ff0e2820d9c80f8c8a01f40d353197ad72acf4544d03bc0bd2c5e681a3eba0bf1fd587f0673b4d2453a0ceecac01eb837f31ce1a6672503f47dd1f;
    5'b01101 : xpb = 1024'h404fa0c933dd6b19f7bea556be5c18924650bdc9c40d831bc93da39e6a96e1e1e63313b34a9684e7dc074c0da89994e24335d80f51f81c3661c8337cc277eb87d93d3e4943883a3b0cb46dd8a0d88719a4a3e0ecf0310cf1f6dd0d36d2a0c8d83330f31555a7129cce8a825652b3eb07647d84d6f26e2e3096bb06ebe3d051ae;
    5'b01110 : xpb = 1024'h37aae2e5c679aa5b49f4466090ab01487e12cc244c8f3214bb58c9553da24868d0451f41a33cacc756d93958068a77a9059a6f74f324d3486f68e3cde09857222fc5b52dc511664df88f13a1b5270c3f3c12904232ef6cef996d16b1996ecbc9e4bdfa89ec2e4fb1acadc95f8114353fdc4f07c2615d2a93130f9b878858c63d;
    5'b01111 : xpb = 1024'h2f0625025915e99c9c29e76a62f9e9feb5d4da7ed510e10dad73ef0c10adaeefba572acffbe2d4a6d1ab26a2647b5a6fc7ff06da94518a5a7d09941efeb8c2bc864e2c12469a9260e469b96ac9759164d3813f9775adcced3bfd202c603ccebb964b01fe82b58cc68ad11068af747f7854208aadd04c26f58f6430232ce13acc;
    5'b10000 : xpb = 1024'h2661671eebb228ddee5f88743548d2b4ed96e8d95d9290069f8f14c2e3b91576a469365e5488fc864c7d13ecc26c3d368a639e40357e416c8aaa44701cd92e56dcd6a2f6c823be73d0445f33ddc4168a6aefeeecb86c2ceade8d29a7270ad1ad47d80973193cc9db68f45771ddd4c9b0cbf20d993f3b23580bb8c4bed169af5b;
    5'b10001 : xpb = 1024'h1dbca93b7e4e681f4095297e0797bb6b2558f733e6143eff91aa3a79b6c47bfd8e7b41ecad2f2465c74f0137205d1ffd4cc835a5d6aaf87e984af4c13af999f1335f19db49acea86bc1f04fcf2129bb0025e9e41fb2a8ce8811d3321edd8d49ef96510e7afc406f047179e7b0c3513e943c39084ae2a1fba880d595a75f223ea;
    5'b10010 : xpb = 1024'h1517eb5810eaa76092caca87d9e6a4215d1b058e6e95edf883c5603089cfe284788d4d7b05d54c454220ee817e4e02c40f2ccd0b77d7af90a5eba512591a058b89e790bfcb361699a7f9aac6066120d599cd4d973de8ece623ad3c9cb4a6d790aaf2185c464b4405253ae5843a955e21bb9513701d191c1d0461edf61a7a9879;
    5'b10011 : xpb = 1024'hc732d74a386e6a1e5006b91ac358cd794dd13e8f7179cf175e085e75cdb490b629f59095e7b7424bcf2dbcbdc3ee58ad1916471190466a2b38c5563773a7125e07007a44cbf42ac93d4508f1aafa5fb313bfcec80a74ce3c63d46177b74da825c7f1fd0dcd2811a035e2c8d68f5a85a3366965b8c08187f80b68291bf030d08;
    5'b10100 : xpb = 1024'h3ce6f91362325e337360c9b7e84758dcc9f22437f994bea67fbab9e2fe6af924cb16497b7219c0437c4c9163a2fc85193f5fbd6ba311db4c12d05b4955adcc036f87e88ce486ebf7faef6582efe2b20c8aaac41c365ace168cd4f924242dd740e0c27457359be2ee18173969755f292ab381946faf714e1fd0b172d638b8197;
    5'b10101 : xpb = 1024'habd6f7038aad99ed5471257c612da59575d733cedd929b5ad7f38aaab5f4c3213a0bed9ed9ee427251f4f5a77b7ebbe2ba74bb227e10a5127f6cf563ee4dbd0c01d02a1bff6298177e239ec3dc287477541e552f92aa39efc0e9eb07c33b82f7eea0c0e3baa9f3d14664a17ebd8662f471e37b14ba316e74bfcf26cd90f65c91;
    5'b10110 : xpb = 1024'ha33239201d49d92ea6a6c686337c8e4bad99422966144a53ca0eb061890029a8241df92d32946a51ccc6e2f1d96f9ea97cd952881f3d5c248d0da5b50c6e28a65858a10080ebc42a69fe448cf076f99ceb8d0484d56899ed6379f4828a0985e9a02dc858513130e62487e887ebe6ad2ce9b4fe0029206ad73c23bb69357ed120;
    5'b10111 : xpb = 1024'h9a8d7b3cafe6186ff8dc679005cb7701e55b5083ee95f94cbc29d6185c0b902f0e3004bb8b3a92314798d03c376081703f3de9edc06a13369aae56062a8e9440aee117e50274f03d55d8ea5604c57ec282fbb3da1826f9eb0609fdfd50d788db51bacfcce7b86dfb02ab2f911a46f765618680eb980f6739b8785004da0745af;
    5'b11000 : xpb = 1024'h91e8bd59428257b14b120899d81a5fb81d1d5ede7717a845ae44fbcf2f16f6b5f8421049e3e0ba10c26abd869551643701a281536196ca48a84f065748aeffdb05698ec983fe1c5041b3901f191403e81a6a632f5ae559e8a89a077817a58bcd0347d7417e3fab0fe0ce769a48a7419dd95803d706fe639c34cce4a07e8fba3e;
    5'b11001 : xpb = 1024'h8943ff75d51e96f29d47a9a3aa69486e54df6d38ff99573ea060218602225d3ce2541bd83c86e1f03d3caad0f34246fdc40718b902c3815ab5efb6a866cf6b755bf205ae058748632d8e35e82d62890db1d912849da3b9e64b2a10f2de738ebeb4d4deb614c6e824bef1bda377078bd6512986c275ed5ffeb121793c23182ecd;
    5'b11010 : xpb = 1024'h809f419267bad633ef7d4aad7cb831248ca17b93881b0637927b473cd52dc3c3cc662766952d09cfb80e981b513329c4866bb01ea3f0386cc39066f984efd70fb27a7c92871074761968dbb141b10e334947c1d9e06219e3edba1a6da54191b06661e62aab4e25399d1504aca567d60ec8fb09ade4dc5c612d760dd7c7a0a35c;
    5'b11011 : xpb = 1024'h77fa83aefa57157541b2ebb74f0719dac46389ee109cb53084966cf3a8392a4ab67832f4edd331af32e08565af240c8b48d04784451cef7ed131174aa31042aa0902f3770899a0890543817a55ff9358e0b6712f232079e1904a23e86c0f94a217eeed9f41d5624e7b384bb5d3c8204740cc8c9953cb58c3a9caa2736c2917eb;
    5'b11100 : xpb = 1024'h6f55c5cb8cf354b693e88cc121560290fc259848991e642976b192aa7b4490d1a08a3e834679598eadb272b00d14ef520b34dee9e649a690ded1c79bc130ae445f8b6a5b8a22cc9bf11e27436a4e187e7825208465ded9df32da2d6332dd9793c97bf513d85c9f63595b92bf02286a7fb89e0f84c2ba5526261f370f10b18c7a;
    5'b11101 : xpb = 1024'h66b107e81f8f93f7e61e2dcaf3a4eb4733e7a6a321a0132268ccb8614e4ff7588a9c4a119f1f816e28845ffa6b05d218cd99764f87765da2ec7277ecdf5119deb613e1400babf8aedcf8cd0c7e9c9da40f93cfd9a89d39dcd56a36ddf9ab9a857b08fc886ee3dc78377ed9c83088b4b8306f927031a95188a273cbaab53a0109;
    5'b11110 : xpb = 1024'h5e0c4a04b22bd3393853ced4c5f3d3fd6ba9b4fdaa21c21b5ae7de18215b5ddf74ae559ff7c5a94da3564d44c8f6b4df8ffe0db528a314b4fa13283dfd7185790c9c58248d3524c1c8d372d592eb22c9a7027f2eeb5b99da77fa4058c0799d772c9603fd056b198d15a220d15ee8fef0a841155ba0984deb1ec8604659c27598;
    5'b11111 : xpb = 1024'h55678c2144c8127a8a896fde9842bcb3a36bc35832a371144d0303cef466c4665ec0612e506bd12d1e283a8f26e797a65262a51ac9cfcbc707b3d88f1b91f1136324cf090ebe50d4b4ae189ea739a7ef3e712e842e19f9d81a8a49d38747a068de230b719bf256a1f3c567da8d494929201298470f874a4d9b1cf4e1fe4aea27;
    endcase
end

endmodule

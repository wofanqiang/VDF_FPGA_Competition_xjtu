module xpb_5_700
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h32f4d89edacb63b23c5e2a3c2d998058c45308effeeff647a8d235f1ccec365fa80b9c0311bc2d8df6b349c6c391ba389a81dac64c15710064dd65bc996575c0bc8d8e5f4cc7bcd80b3642bc5f9f03f21a5f5500a9efcce67e9c333019410ab82f618c3cb81da7a086df52ba2f811c7cc83f3bf57c60f75d7ce05339092a668e;
    5'b00010 : xpb = 1024'h65e9b13db596c76478bc54785b3300b188a611dffddfec8f51a46be399d86cbf5017380623785b1bed66938d872374713503b58c982ae200c9bacb7932caeb81791b1cbe998f79b0166c8578bf3e07e434beaa0153df99ccfd386660328215705ec31879703b4f410dbea5745f0238f9907e77eaf8c1eebaf9c0a6721254cd1c;
    5'b00011 : xpb = 1024'h98de89dc90622b16b51a7eb488cc810a4cf91acffccfe2d6fa76a1d566c4a31ef822d409353488a9e419dd544ab52ea9cf859052e44053012e983135cc30614235a8ab1de657368821a2c8351edd0bd64f1dff01fdcf66b37bd499904bc320288e24a4b62858f6e1949df82e8e83557658bdb3e07522e61876a0f9ab1b7f33aa;
    5'b00100 : xpb = 1024'h1b261d25a93f5a0026733119a60bba119fd6208f264838a7256c1e7180ae2c769ce5f2937cca37a93b6ee7d42ae8d81805ed43330da2f3b5e2d657942ac362517de704ce838df61b1a3f084ee5a04b9775785a6a1b39068944e43ac5aad9884e8e7e9ec92fada5f494bd6409c6344bc9d22310f3a1388045ad11d1df9bc733cd;
    5'b00101 : xpb = 1024'h4e1af5c4840abdb262d15b55d3a53a6a6429297f25382eeece3e54634d9a62d644f18e968e8665373222319aee7a9250a06f1df959b864b647b3bd50c428d8123a74932dd055b2f325754b0b453f4f898fd7af6ac528d36fc3806df5c41a9306bde02b05e7cb4d951b9cb6c3f5b568469a624ce91d9977a329f22518a4f19a5b;
    5'b00110 : xpb = 1024'h810fce635ed621649f2f8592013ebac3287c326f2428253677108a551a869935ecfd2a99a04292c528d57b61b20c4c893af0f8bfa5cdd5b6ac91230d5d8e4dd2f702218d1d1d6fcb30ab8dc7a4de537baa37046b6f18a056421ca125dd5b9dbeed41b7429fe8f535a27c097e253684c362a188de99fa6f00a6d27851ae1c00e9;
    5'b00111 : xpb = 1024'h35761ac77b3504e108837f71e7df3ca7b59382e4da07b06a20606f13470228d91c04923e7d841c4802a85e1923ff5f77158ab9fcf30766b60cf496bbc214ee23f407b3dba542f5e2947cde16ba1933cd0915fd38c82402c0b2c425b3c7205e4ed9bb155a73da448a29b75595ce77b16dc06e5f1c610092ddd4350862e64010c;
    5'b01000 : xpb = 1024'h364c3a4b527eb4004ce662334c1774233fac411e4c90714e4ad83ce3015c58ed39cbe526f9946f5276ddcfa855d1b0300bda86661b45e76bc5acaf285586c4a2fbce099d071bec36347e109dcb40972eeaf0b4d436720d1289c8758b55b3109d1cfd3d925f5b4be9297ac8138c689793a44621e74271008b5a23a3bf378e679a;
    5'b01001 : xpb = 1024'h694112ea2d4a17b289448c6f79b0f47c03ff4a0e4b806795f3aa72d4ce488f4ce1d7812a0b509ce06d91196f19636a68a65c612c675b586c2a8a14e4eeec3a63b85b97fc53e3a90e3fb4535a2adf9b21055009d4e061d9f90864a8bb6ef41b554c5ec9cf1778f389b05a1acdbbe9b4106c855ddcbed1f7e8d703f6f840b8ce28;
    5'b01010 : xpb = 1024'h9c35eb8908157b64c5a2b6aba74a74d4c85252fe4a705ddd9c7ca8c69b34c5ac89e31d2d1d0cca6e64446335dcf524a140de3bf2b370c96c8f677aa18851b02474e9265ba0ab65e64aea96168a7e9f131faf5ed58a51a6df8700dbeb8835260d7bc0560bcf969b2a37396d87eb6ad08d34c499d23b32ef4653e44a3149e334b6;
    5'b01011 : xpb = 1024'h1e7d7ed220f2aa4e36fb6910c489addc1b2f58bd73e8b3adc7722562b51e4f042ea63bb764a2796dbb996db5bd28ce0f7745eed2dcd36a2143a5a0ffe6e4b133bd27800c3de225794386d6305141ded44609ba3da7bb46b550107d20e74b8e337c1a501ed6eb4a3d3758d963231bc6e0ae29f6e5674889738a552265ca2b34d9;
    5'b01100 : xpb = 1024'h51725770fbbe0e007359934cf2232e34df8261ad72d8a9f570445b54820a8563d6b1d7ba765ea6fbb24cb77c80ba884811c7c99928e8db21a88306bc804a26f479b50e6b8aa9e2514ebd18ecb0e0e2c660690f3e51ab139bceacb051008c98ebab7bdc5b8f08f1ddbe382c1d529ce35d766932dae3a980d10735759ed3559b67;
    5'b01101 : xpb = 1024'h8467300fd68971b2afb7bd891fbcae8da3d56a9d71c8a03d191691464ef6bbc37ebd73bd881ad489a9000143444c4280ac49a45f74fe4c220d606c7919af9cb536429ccad7719f2959f35ba9107fe6b87ac8643efb9ae0824d48e38119cda3a3dadd68984726997e45177ed7821dffda3ea86ed0600a782e8415c8d7dc8001f5;
    5'b01110 : xpb = 1024'h6aec358ef66a09c21106fee3cfbe794f6b2705c9b40f60d440c0de268e0451b23809247cfb0838900550bc3247febeee2b1573f9e60ecd6c19e92d778429dc47e80f67b74a85ebc528f9bc2d7432679a122bfa719048058165884b678e40bc9db3762ab4e7b48914536eab2b9cef62db80dcbe38c20125bba86a10c5cc80218;
    5'b01111 : xpb = 1024'h39a39bf7ca32044e5d6e9a2a6a9567edbb05794c9a30ec54ecde43d435cc7b7acb8c2e4ae16cb116f7085589e811a6277d333205ea765dd7267bf89411a813853b0e84dac1701b945dc5de7f36e22a6bbb8214a7c2f44d3e94f4b7e6922516820a98eee80698f031cc163d6ce95012aa804d07d9088109b93766f44565f268a6;
    5'b10000 : xpb = 1024'h6c987496a4fd680099ccc466982ee8467f58823c9920e29c95b079c602b8b1da7397ca4df328dea4edbb9f50aba3606017b50ccc368bced78b595e50ab0d8945f79c133a0e37d86c68fc213b96812e5dd5e169a86ce41a251390eb16ab66213a39fa7b24beb697d252f5902718d12f27488c43ce84e20116b447477e6f1ccf34;
    5'b10001 : xpb = 1024'h9f8d4d357fc8cbb2d62aeea2c5c8689f43ab8b2c9810d8e43e82afb7cfa4e83a1ba3665104e50c32e46ee9176f351a98b236e79282a13fd7f036c40d4472ff06b429a1995aff9544743263f7f620324ff040bea916d3e70b922d1e46c4a72bf2695c076176d43f72d9d4e2e148524ba410cb7fc40142f87431279ab7784735c2;
    5'b10010 : xpb = 1024'h21d4e07e98a5fa9c4783a107e307a1a6968890ebc1892eb469782c53e98e7191c06684db4c7abb323bc3f3974f68c406e89e9a72ac03e08ca474ea6ba3060015fc67fb49f83654d76ccea411bce37211169b1a11343d86e15b3cbf7c23bd941869b601747e28ee85d9f44ebc800341f78a30dcd72d5892a1679872ebf88f35e5;
    5'b10011 : xpb = 1024'h54c9b91d73715e4e83e1cb4410a121ff5adb99dbc07924fc124a6245b67aa7f1687220de5e36e8c032773d5e12fa7e3f83207538f819518d095250283c6b75d6b8f589a944fe11af7804e6ce1c82760330fa6f11de2d53c7d9d8f2ac3cfe9ed099178db13646962660d3a176af845e74527018cca9b989fee478c62501b99c73;
    5'b10100 : xpb = 1024'h87be91bc4e3cc200c03ff5803e3aa2581f2ea2cbbf691b43bb1c98378366de51107dbce16ff3164e292a8724d68c38781da24fff442ec28d6e2fb5e4d5d0eb977583180891c5ce87833b298a7c2179f54b59c412881d20ae587525dc563fa988c87919edee643dc6e7b2f430df057af11aaf54c2261a815c6159195e0ae40301;
    5'b10101 : xpb = 1024'ha0625056719f0ea3198a7e55b79db5f720ba88ae8e17113e61214d39d5067a8b540db6bb788c54d807f91a4b6bfe1e6540a02df6d916342226ddc433463eca6bdc171b92efc8e1a7bd769a442e4b9b671b41f7aa586c0842184c711b55611aec8d31400f5b8ecd9e7d2600c16b671449414b1d552301b8997c9f1928b2c0324;
    5'b10110 : xpb = 1024'h3cfafda441e5549c6df6d22189135bb8365eb17ae7d1675b8ee44ac56a3c9e085d4c776ec944f2db7732db6b7a519c1eee8bdda5b9a6d442874b41ffcdc962677a4f00187bc44af2870dac60a283bda88c13747b4f768d6aa020fa41ce971c66f834a03dadd6947a6eb1b2c646378dc15c53edcace9112e714aa44cb945669b2;
    5'b10111 : xpb = 1024'h6fefd6431cb0b84eaa54fc5db6acdc10fab1ba6ae6c15da337b680b73728d46805581371db0120696de625323de35657890db86c05bc4542ec28a7bc672ed82836dc8e77c88c07ca9243ef1d0222c19aa672c97bf9665a511ebd2d71e7d8271f27962c7a65f43c1af591058075b8aa3e249329c04af20a44918a98049d80d040;
    5'b11000 : xpb = 1024'ha2e4aee1f77c1c00e6b32699e4465c69bf04c35ae5b153eae088b6a904150ac7ad63af74ecbd4df764996ef901751090238f933251d1b64351060d7900944de8f36a1cd71553c4a29d7a31d961c1c58cc0d21e7ca35627379d5960a2011931d756f7b8b71e11e3bb7c70583aa539c6baecd265b5c75301a20e6aeb3da6ab36ce;
    5'b11001 : xpb = 1024'h252c422b10594aea580bd8ff0185957111e1c91a0f29a9bb0b7e33451dfe941f5226cdff3452fcf6bbee7978e1a8b9fe59f746127b3456f8054433d75f274ef83ba87687b28a8435961671f32885054de72c79e4c0bfc70d666901d7602f99fd5751b2ca256692ce7c8fc415dceabd0e6637c2c8f3689bcf44dbc37226f336f1;
    5'b11010 : xpb = 1024'h58211ac9eb24ae9c946a033b2f1f15c9d634d20a0e19a002b4506936eaeaca7efa326a02460f2a84b2a1c33fa53a7436f47920d8c749c7f86a219993f88cc4b8f83604e6ff52410da14cb4af88240940018bcee56aaf93f3e50535077970a4b586b33f06dd843a6f036f16d00c6bd98b2e76febe6fc9932cc1bc16ab301d9d7f;
    5'b11011 : xpb = 1024'h8b15f368c5f0124ed0c82d775cb896229a87dafa0d09964a5d229f28b7d700dea23e060557cb5812a9550d0668cc2e6f8efafb9f135f38f8cefeff5091f23a79b4c393464c19fde5ac82f76be7c30d321beb23e6149f60da63a1683792b1af6db614cb4395a1e20f8a4e698a3becf607f6b63ab3ec2a8a8a3e9c69e43948040d;
    5'b11100 : xpb = 1024'hd5d86b1decd41384220dfdc79f7cf29ed64e0b93681ec1a88181bc4d1c08a364701248f9f61071200aa178648ffd7ddc562ae7f3cc1d9ad833d25aef0853b88fd01ecf6e950bd78a51f3785ae864cf342457f4e320900b02cb1096cf1c81793b66ec5569cf691228a6dd565739dec5b701b97c7184024b7750d4218b9900430;
    5'b11101 : xpb = 1024'h40525f50b998a4ea7e7f0a18a7914f82b1b7e9a93571e26230ea51b69eacc095ef0cc092b11d349ff75d614d0c9192165fe4894588d74aade81a8b6b89eab149b98f7b5636187a50b0557a420e2550e55ca4d44edbf8cd96ab4d3c9d0b09224be5d05193551438c3114d281fa31f08d8385ad3bc94a11c14f1ed9551c2ba6abe;
    5'b11110 : xpb = 1024'h734737ef9464089cbadd3454d52acfdb760af2993461d8a9d9bc87a86b98f6f597185c95c2d9622dee10ab13d0234c4efa66640bd4ecbbae4cf7f1282350270a761d09b582e03728bb8bbcfe6dc454d77704294f85e89a7d29e96fcd244a2d041531ddd00d31e063982c7ad9d2a02555009a0fb2110213726ecde88acbe4d14c;
    5'b11111 : xpb = 1024'ha63c108e6f2f6c4ef73b5e9102c450343a5dfb893351cef1828ebd9a38852d553f23f898d4958fbbe4c3f4da93b5068794e83ed221022caeb1d556e4bcb59ccb32aa9814cfa7f400c6c1ffbacd6358c991637e502fd86763a885a2fd3d8b37bc44936a0cc54f88041f0bcd94022141d1c8d94ba78d630acfebae3bc3d50f37da;
    endcase
end

endmodule

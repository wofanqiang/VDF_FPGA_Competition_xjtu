module xpb_5_855
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h938a6ca37e01841d4fb007f20e9bf153717ad5e92ebe6b0ed10cf31e8ac46a0b109204c8673cdaeb4fd96616dccdfd389d9e5137c4fc3bdbe0896f4720645df2151433ebd4573ab05889951bc9b0bf8c358fb2759ba1d48c9bf35ff09fb92f63006237671b83744fc0126657be2536390160800184b6d2b120692b1606a5f664;
    5'b00010 : xpb = 1024'h766793f13a14d371d45a980d0cdd9b55717fa8a1880535a6243d2ce76286270e1ddb8c180453374800548ce6d63de9a6d7227a896745a76c10739f3005f64732b5d93328f91d781b9e792794fa85bae7771a6b52aabd7c08825a2de68547bc33d1bcdca4863df011f964e5d0847a4648b3e72120b9224831fa62db278469865d;
    5'b00011 : xpb = 1024'h5944bb3ef62822c6590528280b1f455771847b59e14c003d776d66b03a47e4112b251367a16993a4b0cfb3b6cfadd61510a6a3db098f12fc405dcf18eb883073569e32661de3b586e468ba0e2b5ab642b8a5242fb9d9238468c0fbdc6ad64904a31781e1f0f86bd432b765494acf5658666dc23fed8dbdb2d45c8b39022d1656;
    5'b00100 : xpb = 1024'h3c21e28cb23b721addafb8430960ef5971894e123a92cad4ca9da0791209a114386e9ab73e7ff001614ada86c91dc2834a2acd2cabd87e8c7047ff01d11a19b3f76331a342a9f2f22a584c875c2fb19dfa2fdd0cc8f4cb004f27c9d25064d5d57472271f5bb2e7966c09e4c21124666818f4635f21f93333ae563b4a7ff0a64f;
    5'b00101 : xpb = 1024'h1eff09da6e4ec16f625a485e07a2995b718e20ca93d9956c1dcdda41e9cb5e1745b82206db964c5e11c60156c28daef183aef67e4e21ea1ca0322eeab6ac02f4982830e06770305d7047df008d04acf93bba95e9d810727c358e97c835f362a645cccc5cc66d6358a55c643ad7797677cb7b047e5664a8b4884feb5bfdb43648;
    5'b00110 : xpb = 1024'h1dc31282a6210c3e704d87905e4435d7192f382ed20600370fe140ac18d1b1a5301a95678aca8bac2412826bbfd9b5fbd331fcff06b55acd01c5ed39c3dec3538ed301d8c366dc8b6377179bdd9a8547d454ec6e72c19f81bf565be1b81ef771727719a3127df1adeaee3b39dce86877e01a59d8ad01e3562499b6d7b77c641;
    5'b00111 : xpb = 1024'h95669dcba86394e136b4e06b148034b0e30dc96c1bdecb12420b07294c5185256393ae1edfe983a6121a8e3d98cb98985ad17107b5679188b0a5ce1abca24a274e016409608da8790ec10695878a67e0b2d5013c82cdee84b7e8c5aebb3b1eda1789a9014cab536a9ec14a0b5bf3bcc07f62259f0f86f0e682b2c683821dbca5;
    5'b01000 : xpb = 1024'h7843c5196476e435bb5f708612c1deb2e3129c24752595a9953b40f22413422870dd356e7cffe002c295b50d923b850694559a5957b0fd18e08ffe03a2343367eec663468553e5e454b0990eb85f633bf45fba1991e996009e4f93a4a0c9abaae8e44e3eb765cf2cd813c9842248ccd031e8c6be43f266675cac7694ffe14c9e;
    5'b01001 : xpb = 1024'h5b20ec67208a338a400a00a1110388b4e3176edcce6c6040e86b7abafbd4ff2b7e26bcbe1a163c5f7310dbdd8bab7174cdd9c3aaf9fa68a9107a2dec87c61ca88f8b6283aa1a234f9aa02b87e9345e9735ea72f6a1053d7c84b6619a8658387bba3ef37c22204aef116648fce89ddcdfe46f67dd785ddbe836a626a67da4dc97;
    5'b01010 : xpb = 1024'h3dfe13b4dc9d82dec4b490bc0f4532b6e31c419527b32ad83b9bb483d396bc2e8b70440db72c98bc238c02ad851b5de3075decfc9c43d43940645dd56d5805e9305061c0cee060bae08fbe011a0959f277752bd3b020e4f86b1d2f906be6c54c8b9998b98cdac6b14ab8c875aef2ecef96f608fcacc95169109fd6b7fb686c90;
    5'b01011 : xpb = 1024'h20db3b0298b0d233495f20d70d86dcb8e321144d80f9f56f8ecbee4cab58793198b9cb5d5442f518d407297d7e8b4a5140e2164e3e8d3fc9704e8dbe52e9ef29d11560fdf3a69e26267f507a4ade554db8ffe4b0bf3c8c745183fd865175521d5cf43df6f7954273840b47ee7547fcff497caa1be134c6e9ea9986c9792bfc89;
    5'b01100 : xpb = 1024'h3b8625054c42187ce09b0f20bc886bae325e705da40c006e1fc2815831a3634a60352acf15951758482504d77fb36bf7a663f9fe0d6ab59a038bda7387bd86a71da603b186cdb916c6ee2f37bb350a8fa8a9d8dce5833f037eacb7c3703deee2e4ee334624fbe35bd5dc7673b9d0d0efc034b3b15a03c6ac49336daf6ef8c82;
    5'b01101 : xpb = 1024'h9742cef3d2c5a5a51db9b8e41a64780e54a0bcef08ff2b15b3091b340ddea03fb695577558962c60d45bb66454c933f8180490d7a5d2e73580c22cee58e0365c86ee9426ecc41641c4f8780f45641035301a500369fa087cd3de2b6cd6bd0e512eb11a9b7dd332857d702dbef9c24347fd63cb3c9a570f1be4fc61f0fd9582e6;
    5'b01110 : xpb = 1024'h7a1ff6418ed8f4f9a26448ff18a6221054a58fa76245f5ad063954fce5a05d42c3dedec4f5ac88bd84d6dd344e3920665188ba29481c52c5b0ac5cd73e721f9d27b39364118a53ad0ae80a8876390b9071a508e07915aff8ba44f962bc4b9b22000bbfd8e88dae47b6c2ad37c0175357afea6c5bcec2849cbef612027b5912df;
    5'b01111 : xpb = 1024'h5cfd1d8f4aec444e270ed91a16e7cc1254aa625fbb8cc04459698ec5bd621a45d128661492c2e51a3552040447a90cd48b0ce37aea65be55e0968cc0240408ddc87892a13650911850d79d01a70e06ebb32fc1bd88315774a0abc758a1da27f2d166651653482a09f0152cb0866c636762710d7b032dfa1d98efc213f91ca2d8;
    5'b10000 : xpb = 1024'h3fda44dd06ff93a2abb969351529761454af351814d38adbac99c88e9523d748de71ed642fd94176e5cd2ad44118f942c4910ccc8caf29e61080bca90995f21e693d91de5b16ce8396c72f7ad7e30246f4ba7a9a974cfef08712954e8768b4c3a2c10a53be02a5cc2967ac294cc1737714f7ae9a37996f9e72e9722576e032d1;
    5'b10001 : xpb = 1024'h22b76c2ac312e2f73063f950136b201654b407d06e1a5572ffca02576ce5944bebbb74b3ccef9dd3964851a43a88e5b0fe15361e2ef89576406aec91ef27db5f0a02911b7fdd0beedcb6c1f408b7fda236453377a668a66c6d7963446cf74194741baf9128bd218e62ba2ba213168386c77e4fb96c04e51f4ce32236f4a3c2ca;
    5'b10010 : xpb = 1024'h59493787f26324bb50e896b11acca1854b8da88c761200a52fa3c2044a7514ef904fc036a05fa3046c3787433f8d21f37995f6fd142010670551c7ad4b9c49faac79058a4a3495a22a6546d398cf8fd77cfec54b5844de853e0313a5285ce65457654ce93779d509c0cab1ad96b93967a04f0d8a0705aa026dcd248726752c3;
    5'b10011 : xpb = 1024'h991f001bfd27b66904be915d2048bb6bc633b071f61f8b1924072f3ecf6bbb5a099700cbd142d51b969cde8b10c6cf57d537b0a7963e3ce250de8bc1f51e2291bfdbc44478fa840a7b2fe989033db889ad5f9eca51262274efd3912af23efdc845d88c35aefb11a05c1f11729790c9cf7b6570da25272d514745fd5e790d4927;
    5'b10100 : xpb = 1024'h7bfc2769b93b05bd896921781e8a656dc638832a4f6655b077376907a72d785d16e0881b6e5931784718055b0a36bbc60ebbd9f93887a87280c8bbaadab00bd260a0c3819dc0c175c11f7c023412b3e4eeea57a76041c9f0d63a5f20d7cd8a991733317319b58d62957190eb5de5d9df2dec11f95992a2d2213fad6ff6d0d920;
    5'b10101 : xpb = 1024'h5ed94eb7754e55120e13b1931ccc0f6fc63d55e2a8ad2047ca67a2d07eef3560242a0f6b0b6f8dd4f7932c2b03a6a8344840034adad11402b0b2eb93c041f5130165c2bec286fee1070f0e7b64e7af40307510846f5d716cbca12d16bd5c1769e88dd6b084700924cec41064243ae9eee072b3188dfe1852fb395d8174946919;
    5'b10110 : xpb = 1024'h41b676053161a46692be41ae1b0db971c642289b01f3eadf1d97dc9956b0f263317396baa885ea31a80e52fafd1694a281c42c9c7d1a7f92e09d1b7ca5d3de53a22ac1fbe74d3c4c4cfea0f495bcaa9b71ffc9617e7918e8a307fb0ca2eaa43ab9e87bedef2a84e708168fdcea8ff9fe92f95437c2698dd3d5330d92f257f912;
    5'b10111 : xpb = 1024'h24939d52ed74f3bb1768d1c9194f6373c646fb535b3ab57670c816622e72af663ebd1e0a459c468e588979caf6868110bb4855ee1f63eb2310874b658b65c79442efc1390c1379b792ee336dc691a5f6b38a823e8d94c064896ec9028879310b8b43212b59e500a941690f55b0e50a0e457ff556f6d50354af2cbda4701b890b;
    5'b11000 : xpb = 1024'h770c4a0a988430f9c1361e417910d75c64bce0bb481800dc3f8502b06346c694c06a559e2b2a2eb0904a09aeff66d7ef4cc7f3fc1ad56b340717b4e70f7b0d4e3b4c07630d9b722d8ddc5e6f766a151f5153b1b9cb067e06fd596f86e07bddc5c9dc668c49f7c6b7abb8ece773a1a1df80696762b4078d589266db5eddf1904;
    5'b11001 : xpb = 1024'h9afb31442789c72cebc369d6262cfec937c6a3f4e33feb1c9505434990f8d6745c98aa2249ef7dd658de06b1ccc46ab7926ad07786a9928f20faea95915c0ec6f8c8f4620530f1d331675b02c11760de2aa4ed9138523c6d0bc8f6e90dc0ed3f5cfffdcfe022f0bb3acdf526355f5056f9671677aff74b86a98f98cbf4850f68;
    5'b11010 : xpb = 1024'h7dd85891e39d1681706df9f1246ea8cb37cb76ad3c86b5b3e8357d1268ba937769e23171e705da3309592d81c6345725cbeef9c928f2fe1f50e51a7e76edf807998df39f29f72f3e7756ed7bf1ec5c396c2fa66e476de3e8f22fc4def34f7a102e5aa30d4add6c7d7420749efbb46066abedb796e462c107838948dd72489f61;
    5'b11011 : xpb = 1024'h60b57fdf9fb065d5f5188a0c22b052cd37d0496595cd804b3b65b6db407c507a772bb8c1841c368fb9d45451bfa443940573231acb3c69af80cf4a675c7fe1483a52f2dc4ebd6ca9bd467ff522c15794adba5f4b56898b64d89692d4d8de06e0ffb5484ab597e83fad72f417c20970765e7458b618ce36885d82f8eef00c2f5a;
    5'b11100 : xpb = 1024'h4392a72d5bc3b52a79c31a2720f1fccf37d51c1def144ae28e95f0a4183e0d7d84754011213292ec6a4f7b21b91430023ef74c6c6d85d53fb0b97a504211ca88db17f2197383aa150336126e539652efef45182865a532e0befd60cabe6c93b1d10fed8820526401e6c57390885e808610faf9d54d39ac09377ca9006dcfbf53;
    5'b11101 : xpb = 1024'h266fce7b17d7047efe6daa421f33a6d137d9eed6485b1579e1c62a6cefffca8091bec760be48ef491acaa1f1b2841c70787b75be0fcf40cfe0a3aa3927a3b3c97bdcf1569849e7804925a4e7846b4e4b30cfd10574c0da5ca5642ec0a3fb2082a26a92c58b0cdfc42017f3094eb39095c3819af481a5218a11765911eb934f4c;
    5'b11110 : xpb = 1024'h94cf5c8d3ea53d383183a5d1d7550d337dec18ea1a1e01134f66435c7c187839f084eb05b5f4ba5cb45c8c1abf408deb1ff9f0fb218ac60108dda220d359d0a1ca1f093bd1024eb8f153760b54049a6725a89e283dc81d88bcafcb68989ad5373c53802f5c75b86596a72821508a0a576083c13b610970aeb7009236956df45;
    5'b11111 : xpb = 1024'h9cd7626c51ebd7f0d2c8424f2c114226a9599777d0604b20060357545285f18eaf9a5378c29c26911b1f2ed888c206174f9df0477714e83bf11749692d99fafc31b6247f91675f9be79ecc7c7ef10932a7ea3c581f7e566527be5ca72942dcb674276f6a114acfd6197cd8d9d32dd6de7768bc153ac769bc0bd934396ffcd5a9;
    endcase
end

endmodule

module xpb_5_665
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1e7c66fd1aa407e3e2e164ec92e142500ff57d04b4e1fd691505b105ebd4013a48f5969ee2a702dcfb5c7c003f8e6fdcffb6e1bb1a4b0cfcbaf39cfea0721cc1773b7c5d4ffe074f2e8f18dcf32f9fc047317e70b75305fee9f937605b3e2856c554f6e604f808680b4010a5bd0cf6f3a9ad5fbd37c53d40b5b9b2051ef9c22c;
    5'b00010 : xpb = 1024'h3cf8cdfa35480fc7c5c2c9d925c284a01feafa0969c3fad22a0b620bd7a8027491eb2d3dc54e05b9f6b8f8007f1cdfb9ff6dc376349619f975e739fd40e43982ee76f8ba9ffc0e9e5d1e31b9e65f3f808e62fce16ea60bfdd3f26ec0b67c50ad8aa9edcc09f010d01680214b7a19ede7535abf7a6f8a7a816b73640a3df38458;
    5'b00011 : xpb = 1024'h5b7534f74fec17aba8a42ec5b8a3c6f02fe0770e1ea5f83b3f111311c37c03aedae0c3dca7f50896f2157400beab4f96ff24a5314ee126f630dad6fbe156564465b27517effa15ed8bad4a96d98edf40d5947b5225f911fcbdeba62111ba79044ffee4b20ee8193821c031f13726e4dafd081f37a74fb7c2212d160f5ced4684;
    5'b00100 : xpb = 1024'h79f19bf46a901f8f8b8593b24b8509403fd5f412d387f5a45416c417af5004e923d65a7b8a9c0b73ed71f000fe39bf73fedb86ec692c33f2ebce73fa81c87305dcedf1753ff81d3cba3c6373ccbe7f011cc5f9c2dd4c17fba7e4dd816cf8a15b1553db9813e021a02d004296f433dbcea6b57ef4df14f502d6e6c8147be708b0;
    5'b00101 : xpb = 1024'h986e02f1853427736e66f89ede664b904fcb71178869f30d691c751d9b2406236ccbf11a6d430e50e8ce6c013dc82f50fe9268a7837740efa6c210f9223a8fc754296dd28ff6248be8cb7c50bfee1ec163f77833949f1dfa91de14e1c836c9b1daa8d27e18d82a083840533cb140d2c25062deb216da32438ca07a199ae0cadc;
    5'b00110 : xpb = 1024'h63d2498dde9fa8e8642e5b460ed468eee4aeaeb67d44fff00456ccdd3f55a55b2790a4085c3929f44cca8ba99f88e639a2f227c7b0f7da0b1166e9987da37d75715b58130632e9604c0928b1a41fa50b723fd0bbf6bf6e8c64aba47694a4f7670f6373a6d0739e2bcc07d03767da38cab365f8cfe541253fbeab11a30f8269d;
    5'b00111 : xpb = 1024'h24b98b95f88e027269244aa0f3ce88defe4067f01cb64d68154b1dd3bfc95b8ffb6ea0df686a957c402924bad986fe4099e60437955a8a9d6c0a0b98284c5498ce5131de806135e5334fab680d719a10fe557b7c76befce7b043f1a7c48877cd364b2e2071ff424ac8008da9338a9a8054e3bf4a36194f94b1a4631f4ff1e8c9;
    5'b01000 : xpb = 1024'h4335f29313320a564c05af8d86afcb2f0e35e4f4d1984ad12a50ced9ab9d5cca4464377e4b1198593b85a0bb19156e1d999ce5f2afa5979a26fda896c8be715a458cae3bd05f3d3461dec44500a139d14586f9ed2e1202e69a3d29081fc6a023fba0250676f74ab2d3409e4ef0979173fe911f076dde8cd5675e15246eebaaf5;
    5'b01001 : xpb = 1024'h61b259902dd6123a2ee7147a19910d7f1e2b61f9867a483a3f567fdf97715e048d59ce1d2db89b3636e21cbb58a3ddfa9953c7adc9f0a496e1f1459569308e1bbcc82a99205d4483906ddd21f3d0d9918cb8785de56508e5843660687b04c87ac0f51bec7bef531ade80aef4ada48867a83e7ec4a5a3ca161d17c7298de56d21;
    5'b01010 : xpb = 1024'h802ec08d487a1a1e11c87966ac724fcf2e20defe3b5c45a3545c30e583455f3ed64f64bc105f9e13323e98bb98324dd7990aa968e43bb1939ce4e29409a2aadd3403a6f6705b4bd2befcf5fee7007951d3e9f6ce9cb80ee46e2f97c8d642f0d1864a12d280e75b82e9c0bf9a6ab17f5b51ebde81dd690756d2d1792eacdf2f4d;
    5'b01011 : xpb = 1024'h9eab278a631e2201f4a9de533f53921f3e165c02f03e430c6961e1eb6f1960791f44fb5af306a0f02d9b14bbd7c0bdb498c18b23fe86be9057d87f92aa14c79eab3f2353c0595321ed8c0edbda3019121b1b753f540b14e35828cf29318119284b9f09b885df63eaf500d04027be764efb993e3f152e4497888b2b33cbd8f179;
    5'b01100 : xpb = 1024'hc7a4931bbd3f51d0c85cb68c1da8d1ddc95d5d6cfa89ffe008ad99ba7eab4ab64f214810b87253e8999517533f11cc7345e44f8f61efb41622cdd330fb46faeae2b6b0260c65d2c098125163483f4a16e47fa177ed7edd18c95748ed2949eece1ec6e74da0e73c57980fa06ecfb4719566cbf19fca824a7f7d5623461f04d3a;
    5'b01101 : xpb = 1024'h2af6b02ed677fd00ef67305554bbcf6dec8b52db848a9d6715908aa193beb5e5ade7ab1fee2e281b84f5cd75737f8ca4341526b4106a083e1d207a31b0268c702566e75fb0c4647b38103df327b39461b5797888362af3d0768eabef2dd2c743a741655adf067c2d84c10aacaa083e0d001a1ed7346d61e8ad8f143980ea0f66;
    5'b01110 : xpb = 1024'h4973172bf11c04e4d2489541e79d11bdfc80cfe0396c9ad02a963ba77f92b71ff6dd41bed0d52af880524975b30dfc8133cc086f2ab5153ad81417305098a9319ca263bd00c26bca669f56d01ae33421fcaaf6f8ed7df9cf6087e34f8910ef9a6c965c40e3fe849590011b5267153500a9c77e946c329f296348c63e9fe3d192;
    5'b01111 : xpb = 1024'h67ef7e290bc00cc8b529fa2e7a7e540e0c764ce4ee4e98393f9becad6b66b85a3fd2d85db37c2dd57baec575f29c6c5e3382ea2a450022379307b42ef10ac5f313dde01a50c07319952e6fad0e12d3e243dc7569a4d0ffce4a811aafe44f17f131eb5326e8f68cfd9b412bf824222bf45374de51a3f7dc6a19027843bedd93be;
    5'b10000 : xpb = 1024'h866be526266414ac980b5f1b0d5f965e1c6bc9e9a33095a254a19db3573ab99488c86efc962330b2770b4176322adc3b3339cbe55f4b2f344dfb512d917ce2b48b195c77a0be7a68c3bd888a014273a28b0df3da5c2405cd347a52103f8d4047f7404a0cedee9565a6813c9de12f22e7fd223e0edbbd19aacebc2a48ddd755ea;
    5'b10001 : xpb = 1024'ha4e84c2341081c907aecc407a040d8ae2c6146ee5812930b69a74eb9430ebaced1be059b78ca338f7267bd7671b94c1832f0ada079963c3108eeee2c31eeff760254d8d4f0bc81b7f24ca166f4721362d23f724b13770bcc1e7389709acb689ebc9540f2f2e69dcdb1c14d439e3c19dba6cf9dcc138256eb8475dc4dfcd11816;
    5'b10010 : xpb = 1024'h12b76dca99bdefab92c8b11d22c7d3accae0c0c2377ceffd00d046697be00f01176b1ec1914ab7ddce65fa2fcde9ab2ace8d6775712e78e213434bcc978ea7860541208391298bc20e41b7a14ec5eef2256bf7233e43e4ba52e02ed63bdeee6352e2a5af4715ada83641770a6378eaa601a31ea6fafc36fbf3c0134e92e873d7;
    5'b10011 : xpb = 1024'h3133d4c7b461f78f75aa1609b5a915fcdad63dc6ec5eed6615d5f76f67b4103b6060b56073f1babac9c276300d781b07ce4449308b7985dece36e8cb3800c4477c7c9ce0e12793113cd0d07e41f58eb26c9d7593f596eab93cd96636971d16ba18379c954c0db610418187b02085e199ab507e6432c1743ca979c553b1e23603;
    5'b10100 : xpb = 1024'h4fb03bc4cf05ff73588b7af6488a584ceacbbacba140eacf2adba87553881175a9564bff5698bd97c51ef2304d068ae4cdfb2aeba5c492db892a85c9d872e108f3b8193e31259a606b5fe95b35252e72b3cef404ace9f0b826d29d96f25b3f10dd8c937b5105be784cc19855dd92d88d54fdde216a86b17d5f337758d0dbf82f;
    5'b10101 : xpb = 1024'h6e2ca2c1e9aa07573b6cdfe2db6b9a9cfac137d05622e8383fe1597b3f5c12aff24be29e393fc074c07b6e308c94fac1cdb20ca6c00f9fd8441e22c878e4fdca6af3959b8123a1af99ef02382854ce32fb007275643cf6b710cbd4f74d996767a2e18a6155fdc6e05801a8fb9a9fcf80feab3ddea24beebe14ed295defd5ba5b;
    5'b10110 : xpb = 1024'h8ca909bf044e0f3b1e4e44cf6e4cdced0ab6b4d50b04e5a154e70a812b3013ea3b41793d1be6c351bbd7ea30cc236a9ecd68ee61da5aacd4ff11bfc719571a8be22f11f8d121a8fec87e1b151b846df34231f0e61b8ffcb5fac50c57a8d78fbe683681475af5cf486341b9a157acc674a8589d9bda112bfecaa6db630ecf7c87;
    5'b10111 : xpb = 1024'hab2570bc1ef2171f012fa9bc012e1f3d1aac31d9bfe6e30a69ecbb871704152484370fdbfe8dc62eb73466310bb1da7bcd1fd01cf4a5b9d1ba055cc5b9c9374d596a8e56211fb04df70d33f20eb40db389636f56d2e302b4e4be43b80415b8152d8b782d5fedd7b06e81ca4714b9bd685205fd5911d6693f80608d682dc93eb3;
    5'b11000 : xpb = 1024'h18f4926377a7ea3a190b96d183b51a3bb92babad9f513ffc0115b3374fd56956c9e42902170e4a7d1332a2ea67e2398e68bc89f1ec3df682c459ba661f68df5d5c56d604c18cba5813024a2c6907e942dc8ff42efdafdba3192ae91da5293dd9c3d8dce9b41ce78af301f40dd9f68e32acd97e33f950494fefaac468c3e09a74;
    5'b11001 : xpb = 1024'h3770f960924bf21dfbecfbbe16965c8bc92128b254333d65161b643d3ba96a9112d9bfa0f9b54d5a0e8f1eeaa770a96b68736bad0689037f7f4d5764bfdafc1ed3925262118ac1a7419163095c37890323c1729fb502e1a20324207e00676630892dd3cfb914eff2fe4204b3970385265686ddf131158690a564766de2da5ca0;
    5'b11010 : xpb = 1024'h55ed605daceffa01dece60aaa9779edbd916a5b709153ace2b211543277d6bcb5bcf563fdc5c503709eb9aeae6ff1948682a4d6820d4107c3a40f463604d18e04acdcebf6188c8f670207be64f6728c36af2f1106c55e7a0ed1d57de5ba58e874e82cab5be0cf85b0982155954107c1a00343dae68dac3d15b1e287301d41ecc;
    5'b11011 : xpb = 1024'h7469c75ac79401e5c1afc5973c58e12be90c22bbbdf738374026c64913516d05a4c4ecdebf035314054816eb268d892567e12f233b1f1d78f534916200bf35a1c2094b1cb186d0459eaf94c34296c883b2246f8123a8ed9fd7168f3eb6e3b6de13d7c19bc30500c314c225ff111d730da9e19d6ba0a0011210d7da7820cde0f8;
    5'b11100 : xpb = 1024'h92e62e57e23809c9a4912a83cf3a237bf9019fc072d935a0552c774eff256e3fedba837da1aa55f100a492eb661bf902679810de556a2a75b0282e60a13152633944c77a0184d794cd3eada035c66843f955edf1dafbf39ec10fc69f1221df34d92cb881c7fd092b200236a4ce2a6a01538efd28d8653e52c6918c7d3fc7a324;
    5'b11101 : xpb = 1024'hb54fff3aeddce4bc6d179951c11e7a9781199452439291ec556eff37f6c27233679ca3ba2ada3f5ca2cfa4c24c58150334cab34d026726ba7c8c0106d0fa733c310f28a1f1e19ee933c3da901a43d34c8272ca05c8cc8cf57c6c04b33564f96f7a1d3e1c2c1905a482606b93673acbae627e03bfdf1e6335dbc37dd5defee5;
    5'b11110 : xpb = 1024'h1f31b6fc5591e4c89f4e7c85e4a260caa776969907258ffb015b200523cac3ac7c5d33429cd1dd1c57ff4ba501dac7f202ebac6e674d7423757028ffa7431734b36c8b85f1efe8ee17c2dcb78349e39393b3f13abd1bd28bdf75a3650e738d5034cf14242124216dafc27111507431bf580fddc0f7a45ba3eb957582f4d8c111;
    5'b11111 : xpb = 1024'h3dae1df97035ecac822fe1727783a31ab76c139dbc078d641660d10b0f9ec4e6c552c9e17f78dff9535bc7a5416937cf02a28e29819881203063c5fe47b533f62aa807e341edf03d4651f59476798353dae56fab746ed88ac96edac569b1b5a6fa240b0a261c29d5bb0281b70d8128b301bd3d7e2f6998e4a14f278813d2833d;
    endcase
end

endmodule

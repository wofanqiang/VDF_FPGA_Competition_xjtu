module xpb_5_690
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h24f8f33393bdfae0e2fcbc1600f644479b673e6cf09c3c068ab7d548e55c4a36c499a91fbf037a7e31cbdf0bc2350cf0da1217cd49d363e411827f17a07154c085fdb0e61983fedd2565fd1daa09d5413785a1fea188865e3790878eb1ee393c3adfed6ec5a0075b7bcad2944755e040c12c97e34926d8376e17844a40dd9b01;
    5'b00010 : xpb = 1024'h49f1e667277bf5c1c5f9782c01ec888f36ce7cd9e138780d156faa91cab8946d8933523f7e06f4fc6397be17846a19e1b4242f9a93a6c7c82304fe2f40e2a9810bfb61cc3307fdba4acbfa3b5413aa826f0b43fd43110cbc6f210f1d63dc727875bfdadd8b400eb6f795a5288eabc08182592fc6924db06edc2f089481bb3602;
    5'b00011 : xpb = 1024'h6eead99abb39f0a2a8f6344202e2ccd6d235bb46d1d4b413a0277fdab014dea44dccfb5f3d0a6f7a95639d23469f26d28e364767dd7a2bac34877d46e153fe4191f912b24c8bfc977031f758fe1d7fc3a690e5fbe499931aa6b196ac15caabb4b09fc84c50e01612736077bcd601a0c24385c7a9db7488a64a468cdec298d103;
    5'b00100 : xpb = 1024'h93e3ccce4ef7eb838bf2f05803d9111e6d9cf9b3c270f01a2adf5523957128db1266a47efc0de9f8c72f7c2f08d433c368485f35274d8f904609fc5e81c5530217f6c398660ffb749597f476a8275504de1687fa86221978de421e3ac7b8e4f0eb7fb5bb16801d6def2b4a511d57810304b25f8d249b60ddb85e112903766c04;
    5'b00101 : xpb = 1024'h82f7aac20c7b19ba3ea3496f4750e14978e34efdd958ba937ba7116c7cac609d3b7d025f0eae5e8599d1bf3e7ab2fe9de404f1c4e6e2328a6ed3c17e764331129a53fcfd002fd0ca863eef1b9556615219730609b2472c6604613cebf7c7b9af75811002b572c3be43636066cdd3b1a7705188e1d76dbe4e0061a6ebb71a09a;
    5'b00110 : xpb = 1024'h2d286ddfb485ac7c86e6f0acf56b525c32f5735cce31c7afc272465fad27104098517945afee60668b68faffa9e03cdab85266e99841870cb86fbb2f87d587d1afa2f0b5e986fbe9cdc9ec0f635f3b56591cd25f3cacf92497d69b5d716ab4d73237fe6ef0f733976001089ab4331b5b3831b071669db41c4e1d9eb8fc4f3b9b;
    5'b00111 : xpb = 1024'h522161134843a75d69e3acc2f66196a3ce5cb1c9bece03b64d2a1ba892835a775ceb22656ef1dae4bd34da0b6c1549cb92647eb6e214eaf0c9f23a472846dc9235a0a19c030afac6f32fe92d0d69109790a2745dde357f82cf6722ec2358ee136d17ebddb6973af2dbcbdb2efb88fb9bf95e4854afc48c53bc3523033d2cd69c;
    5'b01000 : xpb = 1024'h771a5446dc01a23e4ce068d8f757daeb69c3f036af6a3fbcd7e1f0f177dfa4ae2184cb852df55562ef00b9172e4a56bc6c7696842be84ed4db74b95ec8b83152bb9e52821c8ef9a41895e64ab772e5d8c828165c7fbe05e106f7aa7ad547274fa7f7d94c7c37424e5796adc342dedbdcba8ae037f8eb648b2a4ca74d7e0a719d;
    5'b01001 : xpb = 1024'h9c13477a6fbf9d1f2fdd24eef84e1f33052b2ea3a0067bc36299c63a5d3beee4e61e74a4ecf8cfe120cc9822f07f63ad4688ae5175bbb2b8ecf7387669298613419c03683612f8813dfbe368617cbb19ffadb85b21468c3f3e8832098735608be2d7c6bb41d749a9d36180578a34bc1d7bb7781b42123cc298642b97bee80c9e;
    5'b01010 : xpb = 1024'h105ef558418f633747d4692de8ea1c292f1c69dfbb2b17526f74e22d8f958c13a76fa04be1d5cbd0b33a37e7cf565fd3bc809e389cdc46514dda782fcec86622534a7f9fa005fa1950c7dde372aacc2a432e60c13648e58cc08c279d7ef8f735eeb0220056ae5877c86c6c0cd9ba7634ee0a311c3aedb7c9c00c34dd76e34134;
    5'b01011 : xpb = 1024'h3557e88bd54d5e182ad12543e9e06070ca83a84cabc75358fa2cb77674f1d64a6c09496ba0d9464ee50616f3918b6cc49692b605e6afaa355f5cf7476f39bae2d9483085b989f8f6762ddb011cb4a16b7ab402bfd7d16beaf81caf2c30e7307229900f6f1c4e5fd344373ea121105675af36c8ff841490012e23b927b7c0dc35;
    5'b01100 : xpb = 1024'h5a50dbbf690b58f90dcde159ead6a4b865eae6b99c638f5f84e48cbf5a4e208130a2f28b5fdcc0cd16d1f5ff53c079b570a4cdd330830e1970df765f0fab0fa35f45e16bd30df7d39b93d81ec6be76acb239a4be7959f2492fad36bae2d569ae646ffcdde1ee672ec0021135686636b6706360e2cd3b68389c3b3d71f89e7736;
    5'b01101 : xpb = 1024'h7f49cef2fcc953d9f0ca9d6febcce900015225268cffcb660f9c62083faa6ab7f53c9bab1ee03b4b489dd50b15f586a64ab6e5a07a5671fd8261f576b01c6463e5439251ec91f6b0c0f9d53c70c84bede9bf46bd1ae278a7673dbe4994c3a2ea9f4fea4ca78e6e8a3bcce3c9afbc16f7318ff8c6166240700a52c1bc397c1237;
    5'b01110 : xpb = 1024'ha442c22690874ebad3c75985ecc32d479cb963937d9c076c9a5437512506b4eeb9d644cadde3b5c97a69b416d82a939724c8fd6dc429d5e193e4748e508db9246b4143380615f58de65fd25a1ad2212f2144e8bbbc6aff059ece45d846b1dc26da2fd7bb6d2e75e5b797b65df711f737f2bc90a95f8918a7786a46067a59ad38;
    5'b01111 : xpb = 1024'h188e7004625714d2ebbe9dc4dd5f2a3dc6aa9ecf98c0a2fba72f53445760521d7b277071d2c0b1b90cd753dbb7018fbd9ac0ed54eb4a6979f4c7b447b62c99337cefbf6f7008f725f92bccd52c00323f64c59121d16d585320d23b6c3e7572d0e6083300820584b3aca2a2134697b14f650f49aa586493aea0124f4c3254e1ce;
    5'b10000 : xpb = 1024'h3d876337f6150fb3cebb59dade556e856211dd3c895cdf0231e7288d3cbc9c543fc1199191c42c373ea332e779369cae74d30522351dcd5e064a335f569dedf402ed7055898cf6031e91c9f2d60a07809c4b332072f5deb15862c2faf063ac0d20e8206f47a58c0f286d74a78ded9190263be18da18b6be60e29d39673327ccf;
    5'b10001 : xpb = 1024'h6280566b89d30a94b1b815f0df4bb2ccfd791ba979f91b08bc9efdd62218e68b045ac2b150c7a6b5706f11f33b6ba99f4ee51cef7ef1314217ccb276f70f42b488eb213ba310f4e043f7c7108013dcc1d3d0d51f147e650f8ff34a89a251e5495bc80dde0d45936aa438473bd54371d0e7687970eab2441d7c4157e0b41017d0;
    5'b10010 : xpb = 1024'h8779499f1d91057594b4d206e041f71498e05a166a95570f4756d31f077530c1c8f46bd10fcb2133a23af0fefda0b69028f734bcc8c49526294f318e978097750ee8d221bc94f3bd695dc42e2a1db2030b56771db606eb6dc783d21854401e8596a7fb4cd2e59ac6200319d01c995211a895115433d91c54ea58dc2af4edb2d1;
    5'b10011 : xpb = 1024'hac723cd2b14f005677b18e1ce1383b5c344798835b319315d20ea867ecd17af88d8e14f0cece9bb1d406d00abfd5c38103094c8a1297f90a3ad1b0a637f1ec3594e68307d618f29a8ec3c14bd427874442dc191c578f71cbff1459a7062e57c1d187e8bb9885a2219bcdec6463ef325269c1a9377cfff48c5870607535cb4dd2;
    5'b10100 : xpb = 1024'h20bdeab0831ec66e8fa8d25bd1d438525e38d3bf76562ea4dee9c45b1f2b18274edf4097c3ab97a166746fcf9eacbfa779013c7139b88ca29bb4f05f9d90cc44a694ff3f400bf432a18fbbc6e5559854865cc1826c91cb1981184f3afdf1ee6bdd604400ad5cb0ef90d8d819b374ec69dc14623875db6f93801869baedc68268;
    5'b10101 : xpb = 1024'h45b6dde416dcc14f72a58e71d2ca7c99f9a0122c66f26aab69a199a40487625e1378e9b782af121f98404edb60e1cc985313543e838bf086ad376f773e0221052c92b025598ff30fc6f5b8e48f5f6d95bde263810e1a5177b8a8d6c9afe027a81840316f72fcb84b0ca3aaadfacaccaa9d40fa1bbf0247caee2fee052ea41d69;
    5'b10110 : xpb = 1024'h6aafd117aa9abc3055a24a87d3c0c0e195075099578ea6b1f4596eece9e3ac94d81292d741b28c9dca0c2de72316d9892d256c0bcd5f546abeb9ee8ede7375c5b290610b7313f1ecec5bb602396942d6f568057fafa2d7d5f0395e5861ce60e453201ede389cbfa6886e7d424220aceb5e6d91ff082920025c47724f6f81b86a;
    5'b10111 : xpb = 1024'h8fa8c44b3e58b711389f069dd4b70529306e8f06482ae2b87f114435cf3ff6cb9cac3bf700b6071bfbd80cf2e54be67a073783d91732b84ed03c6da67ee4ca86388e11f18c97f0ca11c1b31fe37318182ceda77e512b5e3427c9e5e713bc9a208e000c4cfe3cc70204394fd689768d2c1f9a29e2514ff839ca5ef699b05f536b;
    5'b11000 : xpb = 1024'h3f4722910287d2950964adcc553021f5a5fca42634f7e478bec6029019993fa5dfd679df593030b8e45acb7c422e2a07d2f73c03e534be7311fad5fe483aa954a3c8e28f68af262248dad9af4a12928706e4fe4662db781a9cddb7b0b8030ca99d867921313d5cff9443b8bd8fc474391ece2e34a2b7340f206ffdf685a8801;
    5'b11001 : xpb = 1024'h28ed655ca3e6780a339306f2c6494666f5c708af53ebba4e16a43571e6f5de31229710bdb4967d89c0118bc38657ef9157418b8d8826afcb42a22c7784f4ff55d03a3f0f100ef13f49f3aab89eaafe69a7f3f1e307b63ddfe15e6309bd6e6a06d4b85500d8b3dd2b750f0e202052278453197ac693524b78601e8429a9382302;
    5'b11010 : xpb = 1024'h4de6589037a472eb168fc308c73f8aae912e471c4487f654a15c0abacc522867e730b9dd7399f807f1dd6acf488cfc823153a35ad1fa13af5424ab8f256654165637eff52992f01c6f59a7d648b4d3aadf7993e1a93ec43e18eeea986f5ca3430f98426f9e53e486f0d9e0b467a807c5144612a9dc7923afce360873ea15be03;
    5'b11011 : xpb = 1024'h72df4bc3cb626dcbf98c7f1ec835cef62c9585893524325b2c13e003b1ae729eabca62fd329d728623a949db0ac209730b65bb281bcd779365a72aa6c5d7a8d6dc35a0db4316eef994bfa4f3f2bea8ec16ff35e04ac74a9c507f7227214adc7f4a782fde63f3ebe26ca4b348aefde805d572aa8d259ffbe73c4d8cbe2af35904;
    5'b11100 : xpb = 1024'h97d83ef75f2068acdc893b34c92c133dc7fcc3f625c06e61b6cbb54c970abcd570640c1cf1a0ed04557528e6ccf71663e577d2f565a0db777729a9be6648fd97623351c15c9aedd6ba25a2119cc87e2d4e84d7deec4fd0fa880ff9b5d33915bb85581d4d2993f33de86f85dcf653c846969f42706ec6d41eaa6511086bd0f405;
    5'b11101 : xpb = 1024'hc23ecd530f02ec4f4807f73b9c81033f1edff3240e509f0c3a6d13fc9645a0431b537c3e67de8f3e7e2c8ababce128a5b6fc2dc8cc16f0fd80ce977cbe7dda673e1cdf8c68def6eccf19c8cadf68f3d9205804501522a480a13ef49cafcac65913078923e6b020bdd7a719245d9825e08f1fb7167a24f25d20d1a4e23cc289b;
    5'b11110 : xpb = 1024'h311ce008c4ae29a5d77d3b89babe547b8d553d9f318145f74e5ea688aec0a43af64ee0e3a581637219aea7b76e031f7b3581daa9d694d2f3e98f688f6c593266f9df7edee011ee4bf25799aa5800647ec98b2243a2dab0a641a476d87ceae5a1cc106601040b0967594544268d2f629eca1e9354b0c9275d40249e9864a9c39c;
    5'b11111 : xpb = 1024'h5615d33c586c2486ba79f79fbbb498c328bc7c0c221d81fdd9167bd1941cee71bae88a036484ddf04b7a86c330382c6c0f93f277206836d7fb11e7a70cca87277fdd2fc4f995ed2917bd96c8020a39c00110c442446337047934fe672ed91ede06f0536fc9ab10c2d51016bad48542df8b4b2b37f9efff94ae3c22e2a5875e9d;
    endcase
end

endmodule

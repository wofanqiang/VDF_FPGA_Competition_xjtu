module xpb_5_525
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9b5766e03278934267663ba5ecedd8a0ea02bdf28af409072d8b7f39d610d4a72fb153b447305c9f48378c986094199c42df9887efa41668bd21b1ae060fd77a109e326fef5401bc3fde810a71876e30319a69553e3ff411d60b32620f03d34cbe5843d3975e0cb31ce1d62e5bb53a89261178f71a775984f7cd08266face244;
    5'b00010 : xpb = 1024'h8601886aa302f1bc03c6ff74c98169f0628f78b440707196dd3a451df91efc465c1a29efc43a3aaff110d9e9ddca226e21a50929bc955c85c9a423fdd14d3a42aced30312f1706336d22ff724a33182f6f2fd911eff9bb12f689d2c963dd04074da8f57d7df320d8b303c57dbf9a4ee8fd49130be4a355d9a92a954856775e1d;
    5'b00011 : xpb = 1024'h70aba9f5138d5035a027c343a614fb3fdb1c3375f5ecda268ce90b021c2d23e58883002b414418c099ea273b5b002b40006a79cb8986a2a2d626964d9c8a9d0b493c2df26eda0aaa9a677dda22dec22eacc548cea1b3821417087330b8b634c1dcf9a727648834fe4925b4cd237f6348d480ad20aecf522e5a88226a3d41d9f6;
    5'b00100 : xpb = 1024'h5b55cb7f8417aeaf3c88871282a88c8f53a8ee37ab6942b63c97d0e63f3b4b84b4ebd666be4df6d142c3748cd8363411df2fea6d5677e8bfe2a9089d67c7ffd3e58b2bb3ae9d0f21c7abfc41fb8a6c2dea5ab88b536d4915378713980d8f657c6c4a58d14b1d4923df47a41c876477a8abb8473578fb4e830be5af8c240c55cf;
    5'b00101 : xpb = 1024'h45ffed09f4a20d28d8e94ae15f3c1ddecc35a8f960e5ab45ec4696ca62497323e154aca23b57d4e1eb9cc1de556c3ce3bdf55b0f23692edcef2b7aed3305629c81da2974ee601398f4f07aa9d436162d27f02848052710165805b3ff62689636fb9b0a7b31b25d497569936beb498c0882efe14a43274ad7bd433cae0ad6d1a8;
    5'b00110 : xpb = 1024'h30aa0e94652c6ba2754a0eb03bcfaf2e44c263bb166213d59bf55cae85579ac30dbd82ddb861b2f294760f2fd2a245b59cbacbb0f05a74f9fbaded3cfe42c5651e2927362e2318102234f911ace1c02c65859804b6e0d71778845466b741c6f18aebbc251847716f0b8b82bb4f2ea0685a277b5f0d53472c6ea0c9cff1a14d81;
    5'b00111 : xpb = 1024'h1b54301ed5b6ca1c11aad27f1863407dbd4f1e7ccbde7c654ba42292a865c2623a265919356b91033d4f5c814fd84e877b803c52bd4bbb1708305f8cc980282dba7824f76de61c874f797779858d6a2ba31b07c1689a9e189902f4ce0c1af7ac1a3c6dcefedc8594a1ad720ab313b4c8315f1573d77f43811ffe56f1d86bc95a;
    5'b01000 : xpb = 1024'h5fe51a946412895ae0b964df4f6d1cd35dbd93e815ae4f4fb52e876cb73ea01668f2f54b2756f13e628a9d2cd0e57595a45acf48a3d013414b2d1dc94bd8af656c722b8ada920fe7cbdf5e15e39142ae0b0777e1a546519b981953560f42866a98d1f78e57199ba37cf615a16f8c9280896af88a1ab3fd5d15be413bf364533;
    5'b01001 : xpb = 1024'ha155b88978b9bbd81571d1f3e1e4aa6e1fde97310c4eedfc28de67b0a184bea896408308f9a5cbb32e60366b2da270f59d25457c79e1179cd1d4838a9acd6270676555289cfd22babc9c76ebcfc0825b124ae0d35894592b8f8cc7976ff7fbb367e5634c7ccfa66d54b1378872ae03b12ea8287fbc22995ac928ec3a2ee32777;
    5'b01010 : xpb = 1024'h8bffda13e9441a51b1d295c2be783bbd986b51f2c1cb568bd88d2d94c492e647c2a9594476afa9c3d73983bcaad879c77beab61e46d25db9de56f5da660ac53903b452e9dcc02731e9e0f553a86c2c5a4fe050900a4e202cb00b67fec4d12c6df73614f66364ba92ead326d7d693181105dfc294864e95af7a86795c15ada350;
    5'b01011 : xpb = 1024'h76a9fb9e59ce78cb4e3359919b0bcd0d10f80cb47747bf1b883bf378e7a10de6ef122f7ff3b987d48012d10e280e82995ab026c013c3a3d6ead9682a31482801a00350ab1c832ba9172573bb8117d6598d75c04cbc07e72dd08a086619aa5d288686c6a049f9ceb880f516273a782c70dd175ca9507a92042be4067dfc781f29;
    5'b01100 : xpb = 1024'h61541d28ca58d744ea941d60779f5e5c8984c7762cc427ab37eab95d0aaf35861b7b05bb70c365e528ec1e5fa5448b6b39759761e0b4e9f3f75bda79fc858aca3c524e6c5c4630204469f22359c38058cb0b30096dc1ae2ef108a8cd6e838de315d7784a308ee2de171705769e5d40d0b44ef6be1aa68e58dd41939fe3429b02;
    5'b01101 : xpb = 1024'h4bfe3eb33ae335be86f4e12f5432efac02118237e240903ae7997f412dbd5d2547e3dbf6edcd43f5d1c56bb1227a943d183b0803ada6301103de4cc9c7c2ed92d8a14c2d9c09349771ae708b326f2a5808a09fc61f7b753011874934c35cbe9da52829f41723f703ad38f4c6024255308b8690d2e4d28aad8e9f20c1ca0d16db;
    5'b01110 : xpb = 1024'h36a8603dab6d94382355a4fe30c680fb7a9e3cf997bcf8ca9748452550cb84c4744cb2326ad722067a9eb9029fb09d0ef70078a57a97762e1060bf199300505b74f049eedbcc390e9ef2eef30b1ad45746360f82d1353c313205e99c1835ef583478db9dfdb90b29435ae4156627699062be2ae7aefe87023ffcade3b0d792b4;
    5'b01111 : xpb = 1024'h215281c81bf7f2b1bfb668cd0d5a124af32af7bb4d39615a46f70b0973d9ac63a0b5886de7e10017237806541ce6a5e0d5c5e9474788bc4b1ce331695e3db324113f47b01b8f3d85cc376d5ae3c67e5683cb7f3f82ef033252848a036d0f2012c3c98d47e44e1f4ed97cd364ca0c7df039f5c4fc792a8356f15a3b0597a20e8d;
    5'b10000 : xpb = 1024'hbfca3528c82512b5c172c9be9eda39a6bb7b27d02b5c9e9f6a5d0ed96e7d402cd1e5ea964eade27cc5153a59a1caeb2b48b59e9147a02682965a3b9297b15ecad8e45715b5241fcf97bebc2bc722855c160eefc34a8ca3373032a6ac1e850cd531a3ef1cae333746f9ec2b42df19250112d5f1143567faba2b7c8277e6c8a66;
    5'b10001 : xpb = 1024'ha7540a32befae46dc37d6841d6db7c3b55ba706f8da9d2f1243150276cf8a8a9fccfb25dac1b3ac71488e03dfab0c84ef76af271041e18d0e68755672f8aed66be2c77e14aa643b9395a6ccd2df99685f2fb585172e8be45490e5cccd0ec241a117282c5624140278c8098e289a6ccd9373ed8085dcdd9309a84d04dee196caa;
    5'b10010 : xpb = 1024'h91fe2bbd2f8542e75fde2c10b36f0d8ace472b3143263b80d3e0160b9006d04929388899292518d7bd622d8f77e6d120d6306312d10f5eedf309c7b6fac8502f5a7b75a28a694830669eeb3506a540853090c80e24a28546698cfd3425c554d4a0c3346f48d6544d22a28831ed8be1390e76721d27f9d5854be25d6fd4e3e883;
    5'b10011 : xpb = 1024'h7ca84d47a00fa160fc3eefdf90029eda46d3e5f2f8a2a410838edbefb314f7e855a15ed4a62ef6e8663b7ae0f51cd9f2b4f5d3b49e00a50aff8c3a06c605b2f7f6ca7363ca2c4ca793e3699cdf50ea846e2637cad65c4c478a0b9d9b7a9e858f3013e6192f6b6872b8c477815170f598e5ae0c31f225d1d9fd3fea91bbae645c;
    5'b10100 : xpb = 1024'h67526ed21099ffda989fb3ae6c963029bf60a0b4ae1f0ca0333da1d3d6231f87820a35102338d4f90f14c8327252e2c493bb44566af1eb280c0eac56914315c09319712509ef511ec127e804b7fc9483abbba78788161348aa8a3e02cf77b649bf6497c316007c984ee666d0b55609f8bce5a646bc51ce2eae9d77b3a278e035;
    5'b10101 : xpb = 1024'h51fc905c81245e543500777d4929c17937ed5b76639b752fe2ec67b7f9314726ae730b4ba042b309b7ee1583ef88eb967280b4f837e3314518911ea65c8078892f686ee649b25595ee6c666c90a83e82e951174439cfda49cb08de6a2450e7044eb5496cfc9590bde5085620193b1e58941d405b867dca835ffb04d589435c0e;
    5'b10110 : xpb = 1024'h3ca6b1e6f1aebccdd1613b4c25bd52c8b07a16381917ddbf929b2d9c1c3f6ec5dadbe1871d4c911a60c762d56cbef4685146259a04d47762251390f627bddb51cbb76ca789755a0d1bb0e4d46953e88226e68700eb89a14aeb877ed1792a17bede05fb16e32aa4e37b2a456f7d2032b86b54da7050a9c6d8115891f7700dd7e7;
    5'b10111 : xpb = 1024'h2750d37162391b476dc1ff1b0250e4182906d0f9ce94464f4249f3803f4d96650744b7c29a566f2b09a0b026e9f4fd3a300b963bd1c5bd7f31960345f2fb3e1a68066a68c9385e8448f5633c41ff9281647bf6bd9d43684c0c061f38ce0348796d56acc0c9bfb909114c34bee1054718428c74851ad5c32cc2b61f1956d853c0;
    5'b11000 : xpb = 1024'h11faf4fbd2c379c10a22c2e9dee47567a1938bbb8410aedef1f8b964625bbe0433ad8dfe17604d3bb279fd78672b060c0ed106dd9eb7039c3e187595be38a0e30455682a08fb62fb7639e1a41aab3c80a211667a4efd2f4d2c84bfa022dc7933fca75e6ab054cd2ea76e240e44ea5b7819c40e99e501bf817413ac3b3da2cf99;
    5'b11001 : xpb = 1024'had525bdc053c0d037188fe8fcbd24e088b9649ae0f04b7e61f84389e386c92ab635ee1b25e90a9dafab18a10c7bf1fa851b09f658e5b1a04fb3a2743c448785d14f39a99f84f64b7b61862ae8c32aab0d3abcfcf8d3d235f028ff20231e04c80baffa23e47b2d9e1c44ffa3ca09f96013fd58790ff7919066be0b461ad4fb1dd;
    5'b11010 : xpb = 1024'h97fc7d6675c66b7d0de9c25ea865df580423046fc4812075cf32fe825b7aba4a8fc7b7eddb9a87eba38ad76244f5287a307610075b4c602207bc99938f85db25b142985b3812692ee35ce11664de54b011413f8c3ef6ea60230e926986b97d3b4a5053e82e47ee075a71e98c0484aa61170d21a5c9a5155b1d3e4183941a2db6;
    5'b11011 : xpb = 1024'h82a69ef0e650c9f6aa4a862d84f970a77cafbf3179fd89057ee1c4667e88e1e9bc308e2958a465fc4c6424b3c22b314c0f3b80a9283da63f143f0be35ac33dee4d91961c77d56da610a15f7e3d89feaf4ed6af48f0b0b161438d32d0db92adf5d9a1059214dd022cf093d8db6869bec0ee44bbba93d111afce9bcea57ae4a98f;
    5'b11100 : xpb = 1024'h6d50c07b56db287046ab49fc618d01f6f53c79f32f79f1952e908a4aa1970988e8996464d5ae440cf53d72053f613a1dee00f14af52eec5c20c17e332600a0b6e9e093ddb798721d3de5dde61635a8ae8c6c1f05a26a7862640bd338306bdeb068f1b73bfb72165286b5c82acc4ed320c57c55cf5dfd0e047ff95bc761af2568;
    5'b11101 : xpb = 1024'h57fae205c76586e9e30c0dcb3e2093466dc934b4e4f65a24de3f502ec4a5312815023aa052b8221d9e16bf56bc9742efccc661ecc22032792d43f082f13e037f862f919ef75b76946b2a5c4deee152adca018ec254243f63848a739f85450f6af84268e5e2072a781cd7b77a3033e7809cb3efe428290a593156e8e94879a141;
    5'b11110 : xpb = 1024'h42a5039037efe5637f6cd19a1ab42495e655ef769a72c2b48dee1612e7b358c7416b10dbcfc2002e46f00ca839cd4bc1ab8bd28e8f11789639c662d2bc7b6648227e8f60371e7b0b986edab5c78cfcad0796fe7f05de0664a5091406da1e402587931a8fc89c3e9db2f9a6c99418fbe073eb89f8f25506ade2b4760b2f441d1a;
    5'b11111 : xpb = 1024'h2d4f251aa87a43dd1bcd9568f747b5e55ee2aa384fef2b443d9cdbf70ac180666dd3e7174ccbde3eefc959f9b70354938a5143305c02beb34648d52287b8c910becd8d2176e17f82c5b3591da038a6ac452c6e3bb797cd65c587b46e2ef770e016e3cc39af3152c3491b9618f7fe10404b23240dbc8103029412032d160e98f3;
    endcase
end

endmodule

module xpb_5_670
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5c2a84f68ad9f4906511465f0a64e56ac76190a270e98acd2b668210fb72c6210e486080621fe2d64eb843a580f7a7ac02596fe49be38e1ceb5762fce82750b7a1e3844091ebf78c74e10e7169a923142216ee1c2bc1de89b3681225c4efddfdbf7901f02b14323dc642925cca8e1fa6ab6a9d3b672ed6255708d98d32cc4569;
    5'b00010 : xpb = 1024'h7a7c49753c5b457ff1d14e7046f83841d4d1e140c5b7522d8f04acc43e2df3a19484387fa19471dfe1248041e913e8da098b7e315144bee260f869b957c2cbdcf77d3d27446f1d3d7281a403a7681f75028e29fcafd9002b1439250cfb519694fea71b6a55f6bee05c53dda9d4c192407fb5b947e124f1a67a23815dcb62467;
    5'b00011 : xpb = 1024'h63d2498dde9fa8e8642e5b460ed468eee4aeaeb67d44fff00456ccdd3f55a55b2790a4085c3929f44cca8ba99f88e639a2f227c7b0f7da0b1166e9987da37d75715b58130632e9604c0928b1a41fa50b723fd0bbf6bf6e8c64aba47694a4f7670f6373a6d0739e2bcc07d03767da38cab365f8cfe541253fbeab11a30f8269d0;
    5'b00100 : xpb = 1024'hf4f892ea78b68affe3a29ce08df07083a9a3c2818b6ea45b1e0959887c5be743290870ff4328e3bfc2490083d227d1b41316fc62a2897dc4c1f0d372af8597b9eefa7a4e88de3a7ae50348074ed03eea051c53f95fb2005628724a19f6a32d29fd4e36d4abed7dc0b8a7bb53a9832480ff6b728fc249e34cf44702bb96c48ce;
    5'b00101 : xpb = 1024'h6b7a0e2532655d40634b702d1343ec7301fbccca89a07512dd4717a98338849540d8e790565271124adcd3adbe1a24c7438adfaac60c25f937767034131faa3340d32be57a79db34233142f1de962702c268b35bc1bcfe8f15ef36c7645a10d05f4de55d75d30a19d1cd0e12052651eebb6154646353745a264d49b8ec388e37;
    5'b00110 : xpb = 1024'h16f74dc5fb511d07fd573eb50d4e8a8c57e75a3c25125f688ad0e064cba89dae4bd8ca97ee4bd559fa36d80c5bb3bba8e1ca27a93f3ce3ca722e93d2c07486396e677b775cd4d57b85784ec0af6385e5f07aa7df60f8b00813cab6f26f1f4c3befbf5523f01e43ca114fb98fd7e44b6c17f212bd7a36ed4f36e6a84196226d35;
    5'b00111 : xpb = 1024'h7321d2bc862b11986268851417b36ff71f48eade95fbea35b6376275c71b63cf5a212b18506bb83048ef1bb1dcab6354e423978ddb2071e75d85f6cfa89bd6f1104affb7eec0cd07fa595d32190ca8fa129195fb8cba8e91c732c918340f2a39af3857141b327607d7924beca2726b12c35caff8e165c3748def81cec8eeb29e;
    5'b01000 : xpb = 1024'h1e9f125d4f16d15ffc74539c11be0e1075347850316dd48b63c12b310f8b7ce865210e1fe8651c77f84920107a44fa368262df8c54512fb8983e1a6e55f0b2f73ddf4f49d11bc74f5ca06900e9da07dd40a38a7f2bf6400ac50e49433ed465a53fa9c6da957dafb81714f76a753064901fed6e51f8493c699e88e05772d8919c;
    5'b01001 : xpb = 1024'h7ac99753d9f0c5f0618599fb1c22f37b3c9608f2a2575f588f27ad420afe430973696ea04a84ff4e470163b5fb3ca1e284bc4f70f034bdd583957d6b3e1803aedfc2d38a6307bedbd181777253832af162ba789b57b81e9478765b6903c443a2ff22c8cac091e1f5dd5789c73fbe8436cb580b8d5f78128ef591b9e4a5a4d705;
    5'b01010 : xpb = 1024'h2646d6f4a2dc85b7fb916883162d9194928196643dc949ae3cb175fd536e5c227e6951a7e27e6395f65b681498d638c422fb976f69657ba6be4da109eb6cdfb50d57231c4562b92333c88341245089d490cc6d1ef6f3d00d7651db940e897f0e8f9438913add1ba61cda3545127c7db427e8c9e6765b8b84062b186d4f8eb603;
    5'b01011 : xpb = 1024'h82715beb2db67a4860a2aee2209276ff59e32706aeb2d47b6817f80e4ee122438cb1b228449e466c4513abba19cde07025550754054909c3a9a50406d394306caf3aa75cd74eb0afa8a991b28df9ace8b2e35b3b22b5ae9729b9edb9d3795d0c4f0d3a8165f14de3e31cc7a1dd0a9d5ad3536721dd8a61a95d33f1fa825afb6c;
    5'b01100 : xpb = 1024'h2dee9b8bf6a23a0ffaae7d6a1a9d1518afceb4784a24bed115a1c0c997513b5c97b1952fdc97aab3f46db018b7677751c3944f527e79c794e45d27a580e90c72dccef6eeb9a9aaf70af09d815ec70bcbe0f54fbec1f1601027956de4de3e9877df7eaa47e03c8794229f731fafc896d82fe4257af46dda9e6dcd50832c44da6a;
    5'b01101 : xpb = 1024'h8a192082817c2ea05fbfc3c92501fa837730451abb0e499e410842da92c4017da5f9f5b03eb78d8a4325f3be385f1efdc5edbf371a5d55b1cfb48aa269105d2a7eb27b2f4b95a2837fd1abf2c8702ee0030c3ddaedb33e99dafd800aa32e76759ef7ac380b50b9d1e8e2057c7a56b67edb4ec2b65b9cb0c3c4d62a105f111fd3;
    5'b01110 : xpb = 1024'h359660234a67ee67f9cb92511f0c989ccd1bd28c568033f3ee920b95db341a96b0f9d8b7d6b0f1d1f27ff81cd5f8b5df642d0735938e13830a6cae4116653930ac46cac12df09ccae218b7c1993d8dc3311e325e8ceef012d8d90035adf3b1e12f691bfe859bf3822864b0fa4d14affc37df810f728029b8d56f889908fafed1;
    5'b01111 : xpb = 1024'h91c0e519d541e2f85edcd8b029717e07947d632ec769bec119f88da6d6a6e0b7bf42393838d0d4a841383bc256f05d8b6686771a2f71a19ff5c4113dfe8c89e84e2a4f01bfdc945756f9c63302e6b0d75335207ab8b0ce9c8c41125b72e38fdeeee21deeb0b025bfeea7435717a2cfa2e34a1e4ad9aeffde2c7862263bc7443a;
    5'b10000 : xpb = 1024'h3d3e24ba9e2da2bff8e8a738237c1c20ea68f0a062dba916c78256621f16f9d0ca421c3fd0ca38eff0924020f489f46d04c5bf18a8a25f71307c34dcabe165ee7bbe9e93a2378e9eb940d201d3b40fba814714fe57ec80158a1c92867da8cb4a7f538db52afb5f702e29eed4ea60c9203fdadca3f09278d33d11c0aee5b12338;
    5'b10001 : xpb = 1024'h9968a9b1290797505df9ed972de1018bb1ca8142d3c533e3f2e8d8731a89bff1d88a7cc032ea1bc63f4a83c675819c19071f2efd4485ed8e1bd397d99408b6a61da222d43423862b2e21e0733d5d32cea35e031a83ae5e9f3d84a4ac4298a9483ecc8fa5560f91adf46c8131b4eee8c6eb4579df57c14ef8941a9a3c187d68a1;
    5'b10010 : xpb = 1024'h44e5e951f1f35717f805bc1f27eb9fa507b60eb46f371e39a072a12e62f9d90ae38a5fc7cae3800deea48825131b32faa55e76fbbdb6ab5f568bbb78415d92ac4b367266167e80729068ec420e2a91b1d16ff79e22ea10183b6024d74d5de4b3cf3dff6bd05acb5e33ef2caf87ace24447d638386ea4c7eda4b3f8c4c267479f;
    5'b10011 : xpb = 1024'ha1106e487ccd4ba85d17027e3250850fcf179f56e020a906cbd9233f5e6c9f2bf1d2c0482d0362e43d5ccbca9412daa6a7b7e6e0599a397c41e31e752984e363ed19f6a6a86a77ff0549fab377d3b4c5f386e5ba4eabeea1eec836fd124dc2b18eb7015bfb6efd9bfa31bf0c523b01eaf340d573d5d39e12fbbcd251f5338d08;
    5'b10100 : xpb = 1024'h4c8dade945b90b6ff722d1062c5b232925032cc87b92935c7962ebfaa6dcb844fcd2a34fc4fcc72becb6d02931ac718845f72eded2caf74d7c9b4213d6d9bf6a1aae46388ac572466791068248a113a92198da3dede7a01aeca3b7281d12fe1d1f28712275ba374c39b46a8a24f8fb684fd193ccecb717080c5630da9f1d6c06;
    5'b10101 : xpb = 1024'ha8b832dfd09300005c34176536c00893ec64bd6aec7c1e29a4c96e0ba24f7e660b1b03d0271caa023b6f13ceb2a4193448509ec36eae856a67f2a510bf011021bc91ca791cb169d2dc7214f3b24a36bd43afc85a19a97ea4a00bc94de202dc1adea17312a0ce6989fff6fce6ef871b0efb3c310853e5ed2d635f0a67d1e9b16f;
    5'b10110 : xpb = 1024'h54357280997ebfc7f63fe5ed30caa6ad42504adc87ee087f525336c6eabf977f161ae6d7bf160e49eac9182d503db015e68fe6c1e7df433ba2aac8af6c55ec27ea261a0aff0c641a3eb920c2831795a071c1bcddb8e5301d9de74978ecc817866f12e2d91b19a33a3f79a864c245148c57ccef616ac9662273f868f07bd3906d;
    5'b10111 : xpb = 1024'hb05ff7772458b4585b512c4c3b2f8c1809b1db7ef8d7934c7db9b8d7e6325da0246347582135f12039815bd2d13557c1e8e956a683c2d1588e022bac547d3cdf8c099e4b90f85ba6b39a2f33ecc0b8b493d8aaf9e4a70ea7514f5b9eb1b7f5842e8be4c9462dd57805bc3ac18cd3343303378c9cd1f83c47cb01427dae9fd5d6;
    5'b11000 : xpb = 1024'h5bdd3717ed44741ff55cfad4353a2a315f9d68f094497da22b4381932ea276b92f632a5fb92f5567e8db60316eceeea387289ea4fcf38f29c8ba4f4b01d218e5b99deddd735355ee15e13b02bd8e1797c1ea9f7d83e2c0204f2adbc9bc7d30efbefd548fc0790f28453ee63f5f912db05fc84af5e8dbb53cdb9aa1065889b4d4;
    5'b11001 : xpb = 1024'h75a76b8b63033e78f68c95c2f44c84ab588f6622fbb67f7d8cd4a4e77128fd23a630d675128b9af983564900c6885852567e6a376244cfb037272e9af26f4ebe7323d6f55ae5035782846d18e5b767aeffc9401231e71994d065bf4c7426c5b4f6ec4563ac448d884c191bd324f272dbc59094effbf2e31ec33ff8f027393d2;
    5'b11010 : xpb = 1024'h6384fbaf410a2877f47a0fbb39a9adb57cea8704a0a4f2c50433cc5f728555f348ab6de7b3489c85e6eda8358d602d3127c156881207db17eec9d5e6974e45a38915c1afe79a47c1ed095542f804998f1213821d4ee05023006e6e1a8c324a590ee7c64665d87b164b042419fcdd46d467c3a68a66ee0457433cd91c353fd93b;
    5'b11011 : xpb = 1024'hf023b5009f5e83f8e85de4333b44bced2d614763c16dd1ab1bd951abaf56f0c53ab50ef4b4200cd9647ac942af9c412c6009e868b3898e92981f98544a321a9b6aa1141c9f542094f506111c8d1f872402576a0ee1c019bfe49ee4596f785c49f59360ce023b4c68a86cf97cf9b4051c45464e37dd17d4c53d637a4df29b839;
    5'b11100 : xpb = 1024'h6b2cc04694cfdccff39724a23e1931399a37a518ad0067e7dd24172bb668352d61f3b16fad61e3a3e4fff039abf16bbec85a0e6b271c270614d95c822cca7261588d95825be13995c4316f83327b1b86623c64bd19dde025b1b2006b5be763c25ed237fd0b37e70450c961f49a295ff86fbf021ee5005371aadf113211f5fda2;
    5'b11101 : xpb = 1024'h16a9ffe75dbb9c978da2f32a3823cf52f023328a4872523d8aaddfe6fed84e466cf39477455b47eb9459f498498b02a066995669a04ce4d74f918020da1f4e678621e5143e3c33dd26787b5203487a69904e5940b919919eaf8d809666ac9f2def43a7c3858320b4904c0d726ce75975cc4fc077fbe3cc66bb786fbabbdfdca0;
    5'b11110 : xpb = 1024'h72d484dde8959127f2b439894288b4bdb784c32cb95bdd0ab61461f7fa4b14677b3bf4f7a77b2ac1e312383dca82aa4c68f2c64e3c3072f43ae8e31dc2469f1f28056954d0282b699b5989c36cf19d7db265475ce4db702862f592bc2b9c7d2baebca9b3b09752f2568e9fcf3775791c77ba5db36312a28c12814947eeac2209;
    5'b11111 : xpb = 1024'h1e51c47eb18150ef8cc008113c9352d70d70509e54cdc760639e2ab342bb2d80863bd7ff3f748f09926c3c9c681c412e07320e4cb56130c575a106bc6f9b7b255599b8e6b28325b0fda095923dbefc60e0773be0841721a160d112e73661b8973f2e197a2ae28ca296114b4d0a337299d44b1c0c79f61b81231aa7d098960107;
    endcase
end

endmodule

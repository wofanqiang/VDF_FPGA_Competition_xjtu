module xpb_5_875
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h35ed2fc037e91671f84c888d858c0298d9a2dfbda60a5d4a12477f48e0b6181a2ba3977265fbe46e801fe78f0b5b4f71a4df1da6e024a5b4bf27407dc0d8033fadc9353d7d2b2f352c850a7a9d986f99ea52188bc5091c25bed0953eaa30a3e7e2ddd2d194102b73b37e39dbe69c692b6b50172aa2f9af84ca04ec53b8635669;
    5'b00010 : xpb = 1024'h6bda5f806fd22ce3f099111b0b180531b345bf7b4c14ba94248efe91c16c303457472ee4cbf7c8dd003fcf1e16b69ee349be3b4dc0494b697e4e80fb81b0067f5b926a7afa565e6a590a14f53b30df33d4a431178a12384b7da12a7d546147cfc5bba5a3282056e766fc73b7cd38d256d6a02e5545f35f099409d8a770c6acd2;
    5'b00011 : xpb = 1024'ha1c78f40a7bb4355e8e599a890a407ca8ce89f38f21f17de36d67ddaa222484e82eac65731f3ad4b805fb6ad2211ee54ee9d58f4a06df11e3d75c179428809bf095b9fb877818d9f858f1f6fd8c94ecdbef649a34f1b54713c71bfbbfe91ebb7a8997874bc30825b1a7aad93b3d53b8241f0457fe8ed0e8e5e0ec4fb292a033b;
    5'b00100 : xpb = 1024'h270779ab1db624ff162caa5f05d5c311f5157bc5c2b1d4b0cb4143cdcfd5b360ab45e050cdc9132b61215ef54a0f2cfc2f624eb55ddfc6874bfdc298c88d984d42d5a047451bbf8f9f7a2747dd85fa36b5436896879e438645b5c2ffee97ed0d5c6fb91c9f77b54147390090a2a17e845e667dc83b9b60e2e1a4364a58aaf339;
    5'b00101 : xpb = 1024'h5cf4a96b559f3b710e7932ec8b61c5aaceb85b8368bc31fadd88c316b08bcb7ad6e977c333c4f799e1414684556a7c6dd4416c5c3e046c3c0b25031689659b8cf09ed584c246eec4cbff31c27b1e69d09f9581224ca75fac0486583e98c890f53f4d8bee3387e0b4fab73a6c893de7afc9b694f2de951067aba9229e110e49a2;
    5'b00110 : xpb = 1024'h92e1d92b8d8851e306c5bb7a10edc843a85b3b410ec68f44efd0425f9141e395028d0f3599c0dc0861612e1360c5cbdf79208a031e2911f0ca4c43944a3d9ecc9e680ac23f721df9f8843c3d18b6d96a89e799ae11b07bd1c356ed7d42f934dd222b5ebfc7980c28ae3574486fda50db3506ac1d818ebfec75ae0ef1c971a00b;
    5'b00111 : xpb = 1024'h1821c3960383338c340ccc30861f838b108817cddf594c17843b0852bef54ea72ae8292f359641e84222d65b88c30a86b9e57fc3db9ae759d8d444b3d0432d5ad7e20b510d0c4fea126f44151d7384d38034b8a14a336ae6cc9af0c132ff3632d6019f67aadf3f0edaf3c7455ea693dd517ce465d43d1240f9438040f8f29009;
    5'b01000 : xpb = 1024'h4e0ef3563b6c49fe2c5954be0bab8623ea2af78b8563a9619682879b9fab66c1568bc0a19b922656c242bdea941e59f85ec49d6abbbf8d0e97fb8531911b309a85ab408e8a377f1f3ef44e8fbb0bf46d6a86d12d0f3c870c8b6b85ffdd2fda1ab8df72393eef6a828e7201214542fd08bcccfb907736c1c5c3486c94b155e672;
    5'b01001 : xpb = 1024'h83fc23167355607024a5dd4b913788bcc3cdd7492b6e06aba8ca06e480617edb822f5814018e0ac54262a5799f79a96a03a3bb119be432c35722c5af51f333da337475cc0762ae546b79590a58a4640754d8e9b8d445a3324a3c1b3e87607e029bbd450ad2ff95f641f03afd2bdf6634281d12bb1a30714a8d4d58e869b93cdb;
    5'b01010 : xpb = 1024'h93c0d80e950421951ecee02066944042bfab3d5fc00c37e3d34ccd7ae14e9edaa8a720d9d6370a523244dc1c776e8114468b0d25956082c65aac6ced7f8c2686cee765ad4fce044856460e25d610f704b2608ac0cc8924753801e8277667f584f9385b2b646c8dc6eae8dfa1aaba93644934b036cdec39f10e2ca37993a2cd9;
    5'b01011 : xpb = 1024'h3f293d412139588b4a39768f8bf5469d059d9393a20b20c84f7c4c208ecb0207d62e0980035f5513a3443550d2d23782e947ce79397aade124d2074c98d0c5a81ab7ab9852280f79b1e96b5cfaf97f0a35782137d1d1ae6d1250b3c121972340327158844a56f450222cc7d601481261afe3622e0fd87323dae7b68b519d8342;
    5'b01100 : xpb = 1024'h75166d0159226efd4285ff1d11814935df40735148157e1261c3cb696f811a2201d1a0f2695b398223641cdfde2d86f48e26ec20199f5395e3f947ca59a8c8e7c880e0d5cf533eaede6e75d79891eea41fca39c396daca92d12148ffcbc7c728154f2b55de671fc3d5ab01b1e7e47b8d1b337958b2d222a8a4eca2df0a00d9ab;
    5'b01101 : xpb = 1024'hab039cc1910b856f3ad287aa970d4bceb8e3530eee1fdb5c740b4ab25037323c2d753864cf571df0a384046ee988d666330609c6f9c3f94aa32088481a80cc27764a16134c7e6de40af38052362a5e3e0a1c524f5be3e6b88ff1de3e75f86b0ff82cfe2772774b3789293b8dce80e4b88683908355cbd22d6ef18f32c2643014;
    5'b01110 : xpb = 1024'h3043872c07066718681998610c3f071621102f9bbeb2982f087610a57dea9d4e55d0525e6b2c83d08445acb71186150d73caff87b735ceb3b1a88967a0865ab5afc416a21a189fd424de882a3ae709a7006971429466d5cd9935e18265fe6c65ac033ecf55be7e1db5e78e8abd4d27baa2f9c8cba87a2481f2870081f1e52012;
    5'b01111 : xpb = 1024'h6630b6ec3eef7d8a606620ee91cb09aefab30f5964bcf5791abd8fee5ea0b5688173e9d0d128683f046594461ce1647f18aa1d2e975a746870cfc9e5615e5df55d8d4bdf9743cf09516392a4d87f7940eabb89ce596ff1f3580676c1102f104d8ee111a0e9cea9916965c866a3e990e60e49dff64b73d406bc8becd5aa48767b;
    5'b10000 : xpb = 1024'h9c1de6ac76d893fc58b2a97c17570c47d455ef170ac752c32d050f373f56cd82ad17814337244cad84857bd5283cb3f0bd893ad5777f1a1d2ff70a63223661350b56811d146efe3e7de89d1f7617e8dad50da25a1e790e1916d70bffba5fb43571bee4727dded5051ce402428a85fa117999f720ee6d838b8690d92962abcce4;
    5'b10001 : xpb = 1024'h215dd116ecd375a585f9ba328c88c78f3c82cba3db5a0f95c16fd52a6d0a3894d5729b3cd2f9b28d6547241d5039f297fe4e309634f0ef863e7f0b82a83befc344d081abe209302e97d3a4f77ad49443cb5ac14d56fbfd2e201b0f43aa65b58b2595251a612607eb49a2553f79523d1396102f69411bd5e00a264a78922cbce2;
    5'b10010 : xpb = 1024'h574b00d724bc8c177e4642c01214ca281625ab6181646cdfd3b754734dc050af011632af38f596fbe5670bac5b954209a32d4e3d1515953afda64c006913f302f299b6e95f345f63c458af72186d03ddb5acd9d91c051953deeba482549659730872f7ebf536335efd208f1b5feea63f01604693e4158564d42b36cc4a90134b;
    5'b10011 : xpb = 1024'h8d3830975ca5a2897692cb4d97a0ccc0efc88b1f276eca29e5fed3bc2e7668c92cb9ca219ef17b6a6586f33b66f0917b480c6be3f53a3aefbccd8c7e29ebf642a062ec26dc5f8e98f0ddb9ecb60573779ffef264e10e35799dbc39c0fec6fd5aeb50cabd89465ed2b09ec8f7468b0f6a6cb05dbe870f34e99e30232002f369b4;
    5'b10100 : xpb = 1024'h12781b01d2a08432a3d9dc040cd2880857f567abf80186fc7a6999af5c29d3db5514e41b3ac6e14a46489b838eedd02288d161a4b2ac1058cb558d9daff184d0d9dcecb5a9f9c0890ac8c1c4bac21ee0964c11581991248ea7003d04eeccfeb09f270b656c8d91b8dd5d1bf43557526c89269606d9bd873e21c5946f327459b2;
    5'b10101 : xpb = 1024'h48654ac20a899aa49c266491925e8aa1319847699e0be4468cb118f83cdfebf580b87b8da0c2c5b8c66883129a491f942db07f4b92d0b60d8a7cce1b70c9881087a621f32724efbe374dcc3f585a8e7a809e29e3de9a40b465d0d24398fda2988204de37009dbd2c90db55d01bf3bb97f476ad317cb736c2ebca80c2ead7b01b;
    5'b10110 : xpb = 1024'h7e527a824272b1169472ed1f17ea8d3a0b3b2727441641909ef898411d96040fac5c130006beaa2746886aa1a5a46f05d28f9cf272f55bc249a40e9931a18b50356f5730a4501ef363d2d6b9f5f2fe146af0426fa3a35cda24a16782432e468064e2b10894ade8a044598fac029024c35fc6c45c1fb0e647b5cf6d16a33b0684;
    5'b10111 : xpb = 1024'h39264ecb86d92bfc1b9fdd58d1c4881736803b414a8fe6333635e344b496f21d4b72cf9a2941007274a12e9cda1adad135492b33067312b582c0fb8b7a719de6ee957bf71ea50e37dbdde91faafa97d613d6162dc264bef2de56ac6333447d618b8f1b077f51b867117e2a8f15c67c57c3cfca4725f389c3964de65d2bbf682;
    5'b11000 : xpb = 1024'h397f94acf056a931ba06866312a84b1a4d0ae371bab35bad45aadd7d2bff873c005ac46c088ff475a769fa78d8fcfd1eb833b05a108bd6e017535036787f1d1e1cb28cfcef158018aa42e90c984819174b8f79eea12f6814ecb60004dd64ebbdfb96c4820c0546fa24961c84d7f8d0f0e78d13cf1558e8210369cab98b1f4ceb;
    5'b11001 : xpb = 1024'h6f6cc46d283fbfa3b2530ef098344db326adc32f60bdb8f757f25cc60cb59f562bfe5bde6e8bd8e42789e207e4584c905d12ce00f0b07c94d67a90b43957205dca7bc23a6c40af4dd6c7f38735e088b135e1927a6638843aab86954387958fa5de749753a015726dd8145660be953a1c52dd2af9b85297a5cd6eb70d4382a354;
    5'b11010 : xpb = 1024'ha559f42d6028d615aa9f977e1dc0504c0050a2ed06c816416a39dc0eed6bb77057a1f350d487bd52a7a9c996efb39c0201f1eba7d0d5224995a1d131fa2f239d7844f777e96bde83034cfe01d378f84b2033ab062b41a0606a572a8231c6338dc1526a2534259de18b92903ca531a347be2d42245b4c472a9773a360fbe5f9bd;
    5'b11011 : xpb = 1024'h2a99de97d623b7bed7e6a83492f20b93687d7f79d75ad313fea4a2021b1f22827ffd0d4a705d2332886b71df17b0daa942b6e1688e46f7b2a429d2518034b22bb1bef806b70610731d3805d9d835a3b41680c9f963c48f75739b2dc621cc34e37528aacd176cd0c7b850e33993fde649daa37a6cadfa997f1b0914b02b66e9bb;
    5'b11100 : xpb = 1024'h60870e580e0cce30d03330c2187e0e2c42205f377d65305e10ec214afbd53a9caba0a4bcd65907a1088b596e230c2a1ae795ff0f6e6b9d67635112cf410cb56b5f882d4434313fa849bd105475ce134e00d2e28528cdab9b326bc304cbfcd8cb58067d9eab7cfc3b6bcf1d157a9a4f7545f3919750f44903e50e0103e3ca4024;
    5'b11101 : xpb = 1024'h96743e1845f5e4a2c87fb94f9e0a10c51bc33ef5236f8da82333a093dc8b52b6d7443c2f3c54ec0f88ab40fd2e67798c8c751cb64e90431c2278534d01e4b8ab0d516281b15c6edd76421acf136682e7eb24fb10edd6c7c0f13c5843762d7cb33ae450703f8d27af1f4d56f16136b8a0b143a8c1f3edf888af12ed579c2d968d;
    5'b11110 : xpb = 1024'h1bb42882bbf0c64bf5c6ca06133bcc0c83f01b81f4024a7ab79e66870a3ebdc8ff9f5628d82a51ef696ce9455664b833cd3a12770c0218853100546c87ea473946cb63107ef6a0cd902d22a718232e50e1721a042659b6d5fa805b8766337e08eeba911822d45a954c0ba9ee5002fba2cdb9e10a469c4add32a85ea6cbae868b;
    5'b11111 : xpb = 1024'h51a15842f3d9dcbdee13529398c7cea55d92fb3f9a0ca7c4c9e5e5cfeaf4d5e32b42ed9b3e26365de98cd0d461c007a57219301dec26be39f02794ea48c24a78f494984dfc21d002bcb22d21b5bb9deacbc4328feb62d2fbb950f0c6106421f0d19863e9b6e48608ff89e3ca369f64ce3909f834e995fa61fcad4afa8411dcf4;
    endcase
end

endmodule

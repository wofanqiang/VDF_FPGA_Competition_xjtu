module xpb_5_650
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8d7578144f97e61b3414ce8e4338ee0c81f014c8fb738986a6dffb8f37b7642204d58420fb58477246e37472c1dbb79e6b8fd08fce0e4fcc340b76abb425f1c2ae1ab92d35dc3e44745b1c6a510d1b9c5160ea1a58a47c8b04d9b873a5ff09564bc52278bf0f72b1a14b8c6176c56a27d0c1540702b446cf39667d7a2d8342e4;
    5'b00010 : xpb = 1024'h6a3daad2dd41976d9d242545761794c7926a2661216f7295cfe33dc8bc6c1b3c06628ac92c8a1055ee68a99ea0595e72730579397969cf4cb777adf92d796ed3e7e63dabbc277f43d61c3632093e7307aebcda9c24c2cc055426deec91d3701a6882b2c7cd55ecd5bbd731e3f5baae2652a8c92bb51d306e2c5d7fefd2241f5d;
    5'b00011 : xpb = 1024'h4705dd916aeb48c006337bfca8f63b82a2e437f9476b5ba4f8e680024120d25607ef91715dbbd93995eddeca7ed705467a7b21e324c54ecd3ae3e546a6ccebe521b1c22a4272c04337dd4ff9c16fca730c18cb1df0e11b7fa37405657da7d6de85404316db9c66f9d662d76674aff224d4903e5067861a0d1f54826576c4fbd6;
    5'b00100 : xpb = 1024'h23ce104ff894fa126f42d2b3dbd4e23db35e49916d6744b421e9c23bc5d58970097c98198eeda21d3d7313f65d54ac1a81f0ca8cd020ce4dbe501c94202068f65b7d46a8c8be0142999e69c179a121de6974bb9fbcff6af9f2c12bde697c3da2a1fdd365e9e2e11df0ee7ce8f3a536235677b37519ef03ac124b84db1b65d84f;
    5'b00101 : xpb = 1024'h96430e863eab64d852296b0eb388f8c3d85b2993632dc34aed04754a8a408a0b099ec1c01f6b00e4f849223bd252ee896673367b7c4dce41bc53e19973e6079548cb274f094241fb5f838931d27949c6d0ac21891dba74420e52575550a466bebb63b4f8295b420b7a226b729a7a21d85f2899cc57ed4b05428750c006b4c8;
    5'b00110 : xpb = 1024'h8e0bbb22d5d691800c66f7f951ec770545c86ff28ed6b749f1cd00048241a4ac0fdf22e2bb77b2732bdbbd94fdae0a8cf4f643c6498a9d9a75c7ca8d4d99d7ca4363845484e580866fba9ff382df94e61831963be1c236ff46e80acafb4fadbd0a80862db738cdf3acc5aecce95fe449a9207ca0cf0c341a3ea904caed89f7ac;
    5'b00111 : xpb = 1024'h6ad3ede1638042d275764eb084cb1dc05642818ab4d2a0591ad0423e06f65bc6116c298aeca97b56d360f2c0dc2bb160fc6bec6ff4e61d1af93401dac6ed54db7d2f08d30b30c185d17bb9bb3b10ec51758d86bdade0867996353143e7241481273e167cc57f4817c751544f685528482b07f1c581751db931a00740922ad425;
    5'b01000 : xpb = 1024'h479c209ff129f424de85a567b7a9c47b66bc9322dace896843d384778bab12e012f930331ddb443a7ae627ecbaa9583503e19519a0419c9b7ca039284040d1ecb6fa8d51917c0285333cd382f34243bcd2e9773f79fed5f3e58257bcd2f87b4543fba6cbd3c5c23be1dcf9d1e74a6c46acef66ea33de0758249709b636cbb09e;
    5'b01001 : xpb = 1024'h2464535e7ed3a5774794fc1eea886b367736a4bb00ca72776cd6c6b1105fc9fa148636db4f0d0d1e226b5d189926ff090b573dc34b9d1c1c000c7075b9944efdf0c611d017c7438494fded4aab739b28304567c1461d256e34cf7e35becce20960b9371ae20c3c5ffc689f54663fb0452ed6dc0ee646f0f7178e0c2bdb6c8d17;
    5'b01010 : xpb = 1024'h12c861d0c7d56c9b0a452d61d6711f187b0b65326c65b8695da08ea9514811416133d83803ed601c9f0924477a4a5dd12cce66cf6f89b9c8378a7c332e7cc0f2a91964e9e128483f6bf071263a4f2938da15843123b74e8841ca4aeaaa148cd7d76c769f052b68416f444d6e534f443b0be513398afda960a850ea1800d6990;
    5'b01011 : xpb = 1024'h8ea1fe315c153ce4e4b92164609ffffe09a0cb1c2239e50d3cba0479cccbe5361ae8c1a47b971d7410d406b739805d7b7e5cb6fcc506eb68b7841e6ee70dbdd1d8ac4f7bd3eec2c86b1a237cb4b20e2fdf02425d6adff17388f65d2250a05223c93be9e2af622935b83fd1385bfa5e6b817fa53a9b64216543eb8c1bad90ac74;
    5'b01100 : xpb = 1024'h6b6a30efe9beee374dc8781b937ea6b91a1adcb44835ce1c65bd46b351809c501c75c84cacc8e657b8593be317fe044f85d25fa670626ae93af055bc60613ae31277d3fa5a3a03c7ccdb3d446ce3659b3c5e32df36fe40edd843839b3c74b8e7e5f97a31bda8a359d2cb76badaefa26a03671a5f4dcd0b0436e28e91523188ed;
    5'b01101 : xpb = 1024'h483263ae77689f89b6d7ced2c65d4d742a94ee4c6e31b72b8ec088ecd635536a1e02cef4ddfaaf3b5fde710ef67bab238d4808501bbdea69be5c8d09d9b4b7f44c435878e08544c72e9c570c2514bd0699ba2361031c90682790aa1428491fac02b70a80cbef1d7ded571c3d59e4e668854e8f840035f4a329d99106f6d26566;
    5'b01110 : xpb = 1024'h24fa966d051250dc1fe72589f93bf42f3b0effe4942da03ab7c3cb265aea0a841f8fd59d0f2c781f0763a63ad4f951f794bdb0f9c71969ea41c8c45753083505860edcf766d085c6905d70d3dd461471f71613e2cf3adfe276ddd08d141d86701f749acfda3597a207e2c1bfd8da2a67073604a8b29ede421cd0937c9b7341df;
    5'b01111 : xpb = 1024'h1c2c92b92bc022e88f67c412c1a9aea4b89117cba298949e0c70d5fdf9ec19e211cdc45405e4102aee8db66b376f8cb9c3359a37274e96ac534fba4cc5bb216bfda6175ed1bc6c5f21e8a9b95776bdd547204649b592f5cc62af705fff1ed343c322b1ee87c11c6226e674257cf6e65891d79cd6507c7e10fc795f240141e58;
    5'b10000 : xpb = 1024'h8f38413fe253e849bd0b4acf6f5388f6cd792645b59d12d087a708ef175625c025f260663bb68874f5cc4fd97552b06a07c32a3340833936f94072508081a3d96df51aa322f8050a6679a705e6848779a5d2ee7ef3fdabe7cb04af79a5f0f68a87f74d97a78b8477c3b9f3a3ce94d88d59decdd467bc0eb0492e136c6d97613c;
    5'b10001 : xpb = 1024'h6c0073fe6ffd999c261aa186a2322fb1ddf337dddb98fbdfb0aa4b289c0adcda277f670e6ce851589d51850553d0573e0f38d2dcebdeb8b77caca99df9d520eaa7c09f21a9434609c83ac0cd9eb5dee5032edf00c01bfb621a51d5f291c55d4ea4b4dde6b5d1fe9bde4599264d8a1c8bdbc642f91a24f84f3c2515e212383db5;
    5'b10010 : xpb = 1024'h48c8a6bcfda74aee8f29f83dd510d66cee6d49760194e4eed9ad8d6220bf93f4290c6db69e1a1a3c44d6ba31324dfe1216ae7b86973a38380018e0eb73289dfbe18c23a02f8e870929fbda9556e73650608acf828c3a4adc699efc6b7d99c412c1726e35c41878bff8d13ea8cc7f608a5dadb81dcc8de1ee2f1c1857b6d91a2e;
    5'b10011 : xpb = 1024'h2590d97b8b50fc40f8394ef507ef7d27fee75b0e2790cdfe02b0cf9ba5744b0e2a99745ecf4be31fec5bef5d10cba4e61e2424304295b7b883851838ec7c1b0d1b57a81eb5d9c8088bbcf45d0f188dbbbde6c00458589a56b8ec22e4696e2ad6de2ffe84d25ef2e4135ce42b4b74a488df952d427ef6cb8d22131acd5b79f6a7;
    5'b10100 : xpb = 1024'h2590c3a18faad936148a5ac3ace23e30f616ca64d8cb70d2bb411d52a2902282c267b07007dac0393e12488ef494bba2599ccd9edf1373906f14f8665cf981e55232c9d3c250907ed7e0e24c749e5271b42b0862476e9d10839495d5542919afaed8ed3e0a56d082de889adca69e887617ca267315fb52c150a1d43001ad320;
    5'b10101 : xpb = 1024'h8fce844e689293ae955d743a7e0711ef9151816f49004093d2940d6461e0664a30fbff27fbd5f375dac498fbb125035891299d69bbff87053afcc63219f589e1033de5ca7201474c61d92a8f185700c36ca39aa07d1b665c0d1301d0fb419af146b2b14c9fb4dfb9cf34160f412f52af323df66e3413fbfb4e709abd2d9e1604;
    5'b10110 : xpb = 1024'h6c96b70cf63c4500fe6ccaf1b0e5b8aaa1cb93076efc29a2fb974f9de6951d64328905d02d07bc598249ce278fa2aa2c989f4613675b0685be68fd7f934906f23d096a48f84c884bc39a4456d088582ec9ff8b224939b5d65c602849e71601b56370419badfb59dde9bfbb91c02496adb4256b92e67ce59a41679d32d23ef27d;
    5'b10111 : xpb = 1024'h495ee9cb83e5f653677c21a8e3c45f65b245a49f94f812b2249a91d76b49d47e34160c785e39853d29cf03536e205100a014eebd12b6860641d534cd0c9c840376d4eec77e97c94b255b5e1e88b9af9a275b7ba415580550abad4ec2d2ea6879802dd1eabc41d402044b61143f19daac360ce0b798e5cf39345e9fa876dfcef6;
    5'b11000 : xpb = 1024'h26271c8a118fa7a5d08b786016a30620c2bfb637baf3fbc14d9dd410effe8b9835a313208f6b4e20d154387f4c9df7d4a78a9766be120586c5416c1a85f00114b0a0734604e30a4a871c77e640eb070584b76c25e17654cafafa753bbebecf3d9ceb6239ca884e261ed70696be0f1eaab7f455dc4b4eb8d82755a21e1b80ab6f;
    5'b11001 : xpb = 1024'h2ef4f489f3958f8399acf174981acdbd339c7cfe0efe4d076a1164a74b342b2373019c8c09d170478d96dab2b1b9ea8af004010696d850748ada367ff437e25ea6bf7c48b2e4b49e8dd91adf91c5e70e2135ca7ad94a4454a479bb4aa933601b9a8f288d8cec84a3962ac193d0462a939dbcb00fdb7a2771a4ca493c02187e8;
    5'b11010 : xpb = 1024'h9064c75ceed13f136daf9da58cba9ae85529dc98dc636e571d8111d9ac6aa6d43c059de9bbf55e76bfbce21decf756471a9010a0377bd4d37cb91a13b3696fe89886b0f1c10a898e5d38ae184a297a0d337446c2063920d04f21542850923f58056e150197de3afbdaae387ab3c9ccd10a9d1f08006be94653b3220deda4cacc;
    5'b11011 : xpb = 1024'h6d2cfa1b7c7af065d6bef45cbf9941a365a3ee31025f576646845413311f5dee3d92a491ed27275a67421749cb74fd1b2205b949e2d75454002551612cbcecf9d25235704755ca8dbef9c7e0025ad17890d03743d257704a9e6e7aa13c66a61c222ba550a624b51ff539ddfd32bf10cf8c84942cb2d4d2e546aa24839245a745;
    5'b11100 : xpb = 1024'h49f52cda0a24a1b83fce4b13f277e85e761dffc9285b40756f87964cb5d415083f1fab3a1e58f03e0ec74c75a9f2a3ef297b61f38e32d3d4839188aea6106a0b0c1db9eecda10b8d20bae1a7ba8c28e3ee2c27c59e75bfc4edbba11a283b0ce03ee9359fb46b2f440fc5837fb1b454ce0e6c0951653dbc8439a126f936e683be;
    5'b11101 : xpb = 1024'h26bd5f9897ce530aa8dda1cb25568f19869811614e572984988ad8863a88cc2240acb1e24f8ab921b64c81a188704ac330f10a9d398e535506fdbffc1f63e71c45e93e6d53ec4c8c827bfb6f72bd804f4b8818476a940f3f3d08c793140f73a45ba6c5eec2b1a9682a51290230a998cc90537e7617a6a6232c98296edb876037;
    5'b11110 : xpb = 1024'h38592572578045d11ecf882583535d4971222f974531293c18e1abfbf3d833c4239b88a80bc82055dd1b6cd66edf1973866b346e4e9d2d58a69f74998b7642d7fb4c2ebda378d8be43d15372aeed7baa8e408c936b25eb98c55ee0bffe3da687864563dd0f8238c44dcce84af9edccb123af39aca0f8fc21f8f2be480283cb0;
    5'b11111 : xpb = 1024'h90fb0a6b750fea784601c7109b6e23e1190237c26fc69c1a686e164ef6f4e75e470f3cab7c14c977a4b52b4028c9a935a3f683d6b2f822a1be756df54cdd55f02dcf7c191013cbd0589831a17bfbf356fa44f2e38f56db44912fa67fa5e2e3bec42978b69007963de6285ae6266446f2e2fc47a1ccc3d69158f5a95eadab7f94;
    endcase
end

endmodule

module ms_new
(
    input clk,
    input rst,
    input start,
    input [1023:0] a,

    output [1023:0] ms,
    output valid
);


localparam IDLE             = 8'b00000001;
localparam TRANS_DATA       = 8'b00000010;
localparam ACCUMLATE_1      = 8'b00000100;
localparam ACCUMLATE_2      = 8'b00001000;
localparam ACCUMLATE_3      = 8'b00010000;
localparam ACCUMLATE_4      = 8'b00100000;
localparam REDUCTION        = 8'b01000000;
localparam FINISH           = 8'b10000000;

localparam LOOPS = 31'd1073741824;

reg [7:0] state_current;
reg [7:0] state_next;

reg [1023:0] reg_a;
//reg [1023:0] reg_b;

reg reg_start;
reg reg_clear_i;




reg reg_valid;

reg [32:0] counter;



wire [1023:0] u0_al;
reg [1:0] reg_u0_sel;

assign u0_al = reg_a;
// partial_product Outputs
wire  [127:0]  u0_col_out_0;
wire  [127:0]  u0_col_out_1;
wire  [127:0]  u0_col_out_2;
wire  [127:0]  u0_col_out_3;
wire  [127:0]  u0_col_out_4;
wire  [127:0]  u0_col_out_5;
wire  [127:0]  u0_col_out_6;
wire  [127:0]  u0_col_out_7;
wire  [127:0]  u0_col_out_8;
wire  [127:0]  u0_col_out_9;
wire  [127:0]  u0_col_out_10;
wire  [127:0]  u0_col_out_11;
wire  [127:0]  u0_col_out_12;
wire  [127:0]  u0_col_out_13;
wire  [127:0]  u0_col_out_14;
wire  [127:0]  u0_col_out_15;
wire  [127:0]  u0_col_out_16;
wire  [127:0]  u0_col_out_17;
wire  [127:0]  u0_col_out_18;
wire  [127:0]  u0_col_out_19;
wire  [127:0]  u0_col_out_20;
wire  [127:0]  u0_col_out_21;
wire  [127:0]  u0_col_out_22;
wire  [127:0]  u0_col_out_23;
wire  [127:0]  u0_col_out_24;
wire  [127:0]  u0_col_out_25;
wire  [127:0]  u0_col_out_26;
wire  [127:0]  u0_col_out_27;
wire  [127:0]  u0_col_out_28;
wire  [127:0]  u0_col_out_29;
wire  [127:0]  u0_col_out_30;
wire  [127:0]  u0_col_out_31;
wire  [127:0]  u0_col_out_32;
wire  [127:0]  u0_col_out_33;
wire  [127:0]  u0_col_out_34;
wire  [127:0]  u0_col_out_35;
wire  [127:0]  u0_col_out_36;
wire  [127:0]  u0_col_out_37;
wire  [127:0]  u0_col_out_38;
wire  [127:0]  u0_col_out_39;
wire  [127:0]  u0_col_out_40;
wire  [127:0]  u0_col_out_41;
wire  [127:0]  u0_col_out_42;
wire  [127:0]  u0_col_out_43;
wire  [127:0]  u0_col_out_44;
wire  [127:0]  u0_col_out_45;
wire  [127:0]  u0_col_out_46;
wire  [127:0]  u0_col_out_47;
wire  [127:0]  u0_col_out_48;
wire  [127:0]  u0_col_out_49;
wire  [127:0]  u0_col_out_50;
wire  [127:0]  u0_col_out_51;
wire  [127:0]  u0_col_out_52;
wire  [127:0]  u0_col_out_53;
wire  [127:0]  u0_col_out_54;
wire  [127:0]  u0_col_out_55;
wire  [127:0]  u0_col_out_56;
wire  [127:0]  u0_col_out_57;
wire  [127:0]  u0_col_out_58;
wire  [127:0]  u0_col_out_59;
wire  [127:0]  u0_col_out_60;
wire  [127:0]  u0_col_out_61;
wire  [127:0]  u0_col_out_62;
wire  [127:0]  u0_col_out_63;
wire  [127:0]  u0_col_out_64;
wire  [127:0]  u0_col_out_65;
wire  [127:0]  u0_col_out_66;
wire  [127:0]  u0_col_out_67;
wire  [127:0]  u0_col_out_68;
wire  [127:0]  u0_col_out_69;
wire  [127:0]  u0_col_out_70;
wire  [127:0]  u0_col_out_71;
wire  [127:0]  u0_col_out_72;
wire  [127:0]  u0_col_out_73;
wire  [127:0]  u0_col_out_74;
wire  [127:0]  u0_col_out_75;
wire  [127:0]  u0_col_out_76;
wire  [127:0]  u0_col_out_77;
wire  [127:0]  u0_col_out_78;
wire  [127:0]  u0_col_out_79;
wire  [127:0]  u0_col_out_80;
wire  [127:0]  u0_col_out_81;
wire  [127:0]  u0_col_out_82;
wire  [127:0]  u0_col_out_83;
wire  [127:0]  u0_col_out_84;
wire  [127:0]  u0_col_out_85;
wire  [127:0]  u0_col_out_86;
wire  [127:0]  u0_col_out_87;
wire  [127:0]  u0_col_out_88;
wire  [127:0]  u0_col_out_89;
wire  [127:0]  u0_col_out_90;
wire  [127:0]  u0_col_out_91;
wire  [127:0]  u0_col_out_92;
wire  [127:0]  u0_col_out_93;
wire  [127:0]  u0_col_out_94;
wire  [127:0]  u0_col_out_95;
wire  [127:0]  u0_col_out_96;
wire  [127:0]  u0_col_out_97;
wire  [127:0]  u0_col_out_98;
wire  [127:0]  u0_col_out_99;
wire  [127:0]  u0_col_out_100;
wire  [127:0]  u0_col_out_101;
wire  [127:0]  u0_col_out_102;
wire  [127:0]  u0_col_out_103;
wire  [127:0]  u0_col_out_104;
wire  [127:0]  u0_col_out_105;
wire  [127:0]  u0_col_out_106;
wire  [127:0]  u0_col_out_107;
wire  [127:0]  u0_col_out_108;
wire  [127:0]  u0_col_out_109;
wire  [127:0]  u0_col_out_110;
wire  [127:0]  u0_col_out_111;
wire  [127:0]  u0_col_out_112;
wire  [127:0]  u0_col_out_113;
wire  [127:0]  u0_col_out_114;
wire  [127:0]  u0_col_out_115;
wire  [127:0]  u0_col_out_116;
wire  [127:0]  u0_col_out_117;
wire  [127:0]  u0_col_out_118;
wire  [127:0]  u0_col_out_119;
wire  [127:0]  u0_col_out_120;
wire  [127:0]  u0_col_out_121;
wire  [127:0]  u0_col_out_122;
wire  [127:0]  u0_col_out_123;
wire  [127:0]  u0_col_out_124;
wire  [127:0]  u0_col_out_125;
wire  [127:0]  u0_col_out_126;
wire  [127:0]  u0_col_out_127;
wire  [127:0]  u0_col_out_128;
wire  [127:0]  u0_col_out_129;
wire  [127:0]  u0_col_out_130;
wire  [127:0]  u0_col_out_131;
wire  [127:0]  u0_col_out_132;
wire  [127:0]  u0_col_out_133;
wire  [127:0]  u0_col_out_134;
wire  [127:0]  u0_col_out_135;
wire  [127:0]  u0_col_out_136;
wire  [127:0]  u0_col_out_137;
wire  [127:0]  u0_col_out_138;
wire  [127:0]  u0_col_out_139;
wire  [127:0]  u0_col_out_140;
wire  [127:0]  u0_col_out_141;
wire  [127:0]  u0_col_out_142;
wire  [127:0]  u0_col_out_143;
wire  [127:0]  u0_col_out_144;
wire  [127:0]  u0_col_out_145;
wire  [127:0]  u0_col_out_146;
wire  [127:0]  u0_col_out_147;
wire  [127:0]  u0_col_out_148;
wire  [127:0]  u0_col_out_149;
wire  [127:0]  u0_col_out_150;
wire  [127:0]  u0_col_out_151;
wire  [127:0]  u0_col_out_152;
wire  [127:0]  u0_col_out_153;
wire  [127:0]  u0_col_out_154;
wire  [127:0]  u0_col_out_155;
wire  [127:0]  u0_col_out_156;
wire  [127:0]  u0_col_out_157;
wire  [127:0]  u0_col_out_158;
wire  [127:0]  u0_col_out_159;
wire  [127:0]  u0_col_out_160;
wire  [127:0]  u0_col_out_161;
wire  [127:0]  u0_col_out_162;
wire  [127:0]  u0_col_out_163;
wire  [127:0]  u0_col_out_164;
wire  [127:0]  u0_col_out_165;
wire  [127:0]  u0_col_out_166;
wire  [127:0]  u0_col_out_167;
wire  [127:0]  u0_col_out_168;
wire  [127:0]  u0_col_out_169;
wire  [127:0]  u0_col_out_170;
wire  [127:0]  u0_col_out_171;
wire  [127:0]  u0_col_out_172;
wire  [127:0]  u0_col_out_173;
wire  [127:0]  u0_col_out_174;
wire  [127:0]  u0_col_out_175;
wire  [127:0]  u0_col_out_176;
wire  [127:0]  u0_col_out_177;
wire  [127:0]  u0_col_out_178;
wire  [127:0]  u0_col_out_179;
wire  [127:0]  u0_col_out_180;
wire  [127:0]  u0_col_out_181;
wire  [127:0]  u0_col_out_182;
wire  [127:0]  u0_col_out_183;
wire  [127:0]  u0_col_out_184;
wire  [127:0]  u0_col_out_185;
wire  [127:0]  u0_col_out_186;
wire  [127:0]  u0_col_out_187;
wire  [127:0]  u0_col_out_188;
wire  [127:0]  u0_col_out_189;
wire  [127:0]  u0_col_out_190;
wire  [127:0]  u0_col_out_191;
wire  [127:0]  u0_col_out_192;
wire  [127:0]  u0_col_out_193;
wire  [127:0]  u0_col_out_194;
wire  [127:0]  u0_col_out_195;
wire  [127:0]  u0_col_out_196;
wire  [127:0]  u0_col_out_197;
wire  [127:0]  u0_col_out_198;
wire  [127:0]  u0_col_out_199;
wire  [127:0]  u0_col_out_200;
wire  [127:0]  u0_col_out_201;
wire  [127:0]  u0_col_out_202;
wire  [127:0]  u0_col_out_203;
wire  [127:0]  u0_col_out_204;
wire  [127:0]  u0_col_out_205;
wire  [127:0]  u0_col_out_206;
wire  [127:0]  u0_col_out_207;
wire  [127:0]  u0_col_out_208;
wire  [127:0]  u0_col_out_209;
wire  [127:0]  u0_col_out_210;
wire  [127:0]  u0_col_out_211;
wire  [127:0]  u0_col_out_212;
wire  [127:0]  u0_col_out_213;
wire  [127:0]  u0_col_out_214;
wire  [127:0]  u0_col_out_215;
wire  [127:0]  u0_col_out_216;
wire  [127:0]  u0_col_out_217;
wire  [127:0]  u0_col_out_218;
wire  [127:0]  u0_col_out_219;
wire  [127:0]  u0_col_out_220;
wire  [127:0]  u0_col_out_221;
wire  [127:0]  u0_col_out_222;
wire  [127:0]  u0_col_out_223;
wire  [127:0]  u0_col_out_224;
wire  [127:0]  u0_col_out_225;
wire  [127:0]  u0_col_out_226;
wire  [127:0]  u0_col_out_227;
wire  [127:0]  u0_col_out_228;
wire  [127:0]  u0_col_out_229;
wire  [127:0]  u0_col_out_230;
wire  [127:0]  u0_col_out_231;
wire  [127:0]  u0_col_out_232;
wire  [127:0]  u0_col_out_233;
wire  [127:0]  u0_col_out_234;
wire  [127:0]  u0_col_out_235;
wire  [127:0]  u0_col_out_236;
wire  [127:0]  u0_col_out_237;
wire  [127:0]  u0_col_out_238;
wire  [127:0]  u0_col_out_239;
wire  [127:0]  u0_col_out_240;
wire  [127:0]  u0_col_out_241;
wire  [127:0]  u0_col_out_242;
wire  [127:0]  u0_col_out_243;
wire  [127:0]  u0_col_out_244;
wire  [127:0]  u0_col_out_245;
wire  [127:0]  u0_col_out_246;
wire  [127:0]  u0_col_out_247;
wire  [127:0]  u0_col_out_248;
wire  [127:0]  u0_col_out_249;
wire  [127:0]  u0_col_out_250;
wire  [127:0]  u0_col_out_251;
wire  [127:0]  u0_col_out_252;
wire  [127:0]  u0_col_out_253;
wire  [127:0]  u0_col_out_254;
wire  [127:0]  u0_col_out_255;
wire  [127:0]  u0_col_out_256;
wire  [127:0]  u0_col_out_257;
wire  [127:0]  u0_col_out_258;
wire  [127:0]  u0_col_out_259;
wire  [127:0]  u0_col_out_260;
wire  [127:0]  u0_col_out_261;
wire  [127:0]  u0_col_out_262;
wire  [127:0]  u0_col_out_263;
wire  [127:0]  u0_col_out_264;
wire  [127:0]  u0_col_out_265;
wire  [127:0]  u0_col_out_266;
wire  [127:0]  u0_col_out_267;
wire  [127:0]  u0_col_out_268;
wire  [127:0]  u0_col_out_269;
wire  [127:0]  u0_col_out_270;
wire  [127:0]  u0_col_out_271;
wire  [127:0]  u0_col_out_272;
wire  [127:0]  u0_col_out_273;
wire  [127:0]  u0_col_out_274;
wire  [127:0]  u0_col_out_275;
wire  [127:0]  u0_col_out_276;
wire  [127:0]  u0_col_out_277;
wire  [127:0]  u0_col_out_278;
wire  [127:0]  u0_col_out_279;
wire  [127:0]  u0_col_out_280;
wire  [127:0]  u0_col_out_281;
wire  [127:0]  u0_col_out_282;
wire  [127:0]  u0_col_out_283;
wire  [127:0]  u0_col_out_284;
wire  [127:0]  u0_col_out_285;
wire  [127:0]  u0_col_out_286;
wire  [127:0]  u0_col_out_287;
wire  [127:0]  u0_col_out_288;
wire  [127:0]  u0_col_out_289;
wire  [127:0]  u0_col_out_290;
wire  [127:0]  u0_col_out_291;
wire  [127:0]  u0_col_out_292;
wire  [127:0]  u0_col_out_293;
wire  [127:0]  u0_col_out_294;
wire  [127:0]  u0_col_out_295;
wire  [127:0]  u0_col_out_296;
wire  [127:0]  u0_col_out_297;
wire  [127:0]  u0_col_out_298;
wire  [127:0]  u0_col_out_299;
wire  [127:0]  u0_col_out_300;
wire  [127:0]  u0_col_out_301;
wire  [127:0]  u0_col_out_302;
wire  [127:0]  u0_col_out_303;
wire  [127:0]  u0_col_out_304;
wire  [127:0]  u0_col_out_305;
wire  [127:0]  u0_col_out_306;
wire  [127:0]  u0_col_out_307;
wire  [127:0]  u0_col_out_308;
wire  [127:0]  u0_col_out_309;
wire  [127:0]  u0_col_out_310;
wire  [127:0]  u0_col_out_311;
wire  [127:0]  u0_col_out_312;
wire  [127:0]  u0_col_out_313;
wire  [127:0]  u0_col_out_314;
wire  [127:0]  u0_col_out_315;
wire  [127:0]  u0_col_out_316;
wire  [127:0]  u0_col_out_317;
wire  [127:0]  u0_col_out_318;
wire  [127:0]  u0_col_out_319;
wire  [127:0]  u0_col_out_320;
wire  [127:0]  u0_col_out_321;
wire  [127:0]  u0_col_out_322;
wire  [127:0]  u0_col_out_323;
wire  [127:0]  u0_col_out_324;
wire  [127:0]  u0_col_out_325;
wire  [127:0]  u0_col_out_326;
wire  [127:0]  u0_col_out_327;
wire  [127:0]  u0_col_out_328;
wire  [127:0]  u0_col_out_329;
wire  [127:0]  u0_col_out_330;
wire  [127:0]  u0_col_out_331;
wire  [127:0]  u0_col_out_332;
wire  [127:0]  u0_col_out_333;
wire  [127:0]  u0_col_out_334;
wire  [127:0]  u0_col_out_335;
wire  [127:0]  u0_col_out_336;
wire  [127:0]  u0_col_out_337;
wire  [127:0]  u0_col_out_338;
wire  [127:0]  u0_col_out_339;
wire  [127:0]  u0_col_out_340;
wire  [127:0]  u0_col_out_341;
wire  [127:0]  u0_col_out_342;
wire  [127:0]  u0_col_out_343;
wire  [127:0]  u0_col_out_344;
wire  [127:0]  u0_col_out_345;
wire  [127:0]  u0_col_out_346;
wire  [127:0]  u0_col_out_347;
wire  [127:0]  u0_col_out_348;
wire  [127:0]  u0_col_out_349;
wire  [127:0]  u0_col_out_350;
wire  [127:0]  u0_col_out_351;
wire  [127:0]  u0_col_out_352;
wire  [127:0]  u0_col_out_353;
wire  [127:0]  u0_col_out_354;
wire  [127:0]  u0_col_out_355;
wire  [127:0]  u0_col_out_356;
wire  [127:0]  u0_col_out_357;
wire  [127:0]  u0_col_out_358;
wire  [127:0]  u0_col_out_359;
wire  [127:0]  u0_col_out_360;
wire  [127:0]  u0_col_out_361;
wire  [127:0]  u0_col_out_362;
wire  [127:0]  u0_col_out_363;
wire  [127:0]  u0_col_out_364;
wire  [127:0]  u0_col_out_365;
wire  [127:0]  u0_col_out_366;
wire  [127:0]  u0_col_out_367;
wire  [127:0]  u0_col_out_368;
wire  [127:0]  u0_col_out_369;
wire  [127:0]  u0_col_out_370;
wire  [127:0]  u0_col_out_371;
wire  [127:0]  u0_col_out_372;
wire  [127:0]  u0_col_out_373;
wire  [127:0]  u0_col_out_374;
wire  [127:0]  u0_col_out_375;
wire  [127:0]  u0_col_out_376;
wire  [127:0]  u0_col_out_377;
wire  [127:0]  u0_col_out_378;
wire  [127:0]  u0_col_out_379;
wire  [127:0]  u0_col_out_380;
wire  [127:0]  u0_col_out_381;
wire  [127:0]  u0_col_out_382;
wire  [127:0]  u0_col_out_383;
wire  [127:0]  u0_col_out_384;
wire  [127:0]  u0_col_out_385;
wire  [127:0]  u0_col_out_386;
wire  [127:0]  u0_col_out_387;
wire  [127:0]  u0_col_out_388;
wire  [127:0]  u0_col_out_389;
wire  [127:0]  u0_col_out_390;
wire  [127:0]  u0_col_out_391;
wire  [127:0]  u0_col_out_392;
wire  [127:0]  u0_col_out_393;
wire  [127:0]  u0_col_out_394;
wire  [127:0]  u0_col_out_395;
wire  [127:0]  u0_col_out_396;
wire  [127:0]  u0_col_out_397;
wire  [127:0]  u0_col_out_398;
wire  [127:0]  u0_col_out_399;
wire  [127:0]  u0_col_out_400;
wire  [127:0]  u0_col_out_401;
wire  [127:0]  u0_col_out_402;
wire  [127:0]  u0_col_out_403;
wire  [127:0]  u0_col_out_404;
wire  [127:0]  u0_col_out_405;
wire  [127:0]  u0_col_out_406;
wire  [127:0]  u0_col_out_407;
wire  [127:0]  u0_col_out_408;
wire  [127:0]  u0_col_out_409;
wire  [127:0]  u0_col_out_410;
wire  [127:0]  u0_col_out_411;
wire  [127:0]  u0_col_out_412;
wire  [127:0]  u0_col_out_413;
wire  [127:0]  u0_col_out_414;
wire  [127:0]  u0_col_out_415;
wire  [127:0]  u0_col_out_416;
wire  [127:0]  u0_col_out_417;
wire  [127:0]  u0_col_out_418;
wire  [127:0]  u0_col_out_419;
wire  [127:0]  u0_col_out_420;
wire  [127:0]  u0_col_out_421;
wire  [127:0]  u0_col_out_422;
wire  [127:0]  u0_col_out_423;
wire  [127:0]  u0_col_out_424;
wire  [127:0]  u0_col_out_425;
wire  [127:0]  u0_col_out_426;
wire  [127:0]  u0_col_out_427;
wire  [127:0]  u0_col_out_428;
wire  [127:0]  u0_col_out_429;
wire  [127:0]  u0_col_out_430;
wire  [127:0]  u0_col_out_431;
wire  [127:0]  u0_col_out_432;
wire  [127:0]  u0_col_out_433;
wire  [127:0]  u0_col_out_434;
wire  [127:0]  u0_col_out_435;
wire  [127:0]  u0_col_out_436;
wire  [127:0]  u0_col_out_437;
wire  [127:0]  u0_col_out_438;
wire  [127:0]  u0_col_out_439;
wire  [127:0]  u0_col_out_440;
wire  [127:0]  u0_col_out_441;
wire  [127:0]  u0_col_out_442;
wire  [127:0]  u0_col_out_443;
wire  [127:0]  u0_col_out_444;
wire  [127:0]  u0_col_out_445;
wire  [127:0]  u0_col_out_446;
wire  [127:0]  u0_col_out_447;
wire  [127:0]  u0_col_out_448;
wire  [127:0]  u0_col_out_449;
wire  [127:0]  u0_col_out_450;
wire  [127:0]  u0_col_out_451;
wire  [127:0]  u0_col_out_452;
wire  [127:0]  u0_col_out_453;
wire  [127:0]  u0_col_out_454;
wire  [127:0]  u0_col_out_455;
wire  [127:0]  u0_col_out_456;
wire  [127:0]  u0_col_out_457;
wire  [127:0]  u0_col_out_458;
wire  [127:0]  u0_col_out_459;
wire  [127:0]  u0_col_out_460;
wire  [127:0]  u0_col_out_461;
wire  [127:0]  u0_col_out_462;
wire  [127:0]  u0_col_out_463;
wire  [127:0]  u0_col_out_464;
wire  [127:0]  u0_col_out_465;
wire  [127:0]  u0_col_out_466;
wire  [127:0]  u0_col_out_467;
wire  [127:0]  u0_col_out_468;
wire  [127:0]  u0_col_out_469;
wire  [127:0]  u0_col_out_470;
wire  [127:0]  u0_col_out_471;
wire  [127:0]  u0_col_out_472;
wire  [127:0]  u0_col_out_473;
wire  [127:0]  u0_col_out_474;
wire  [127:0]  u0_col_out_475;
wire  [127:0]  u0_col_out_476;
wire  [127:0]  u0_col_out_477;
wire  [127:0]  u0_col_out_478;
wire  [127:0]  u0_col_out_479;
wire  [127:0]  u0_col_out_480;
wire  [127:0]  u0_col_out_481;
wire  [127:0]  u0_col_out_482;
wire  [127:0]  u0_col_out_483;
wire  [127:0]  u0_col_out_484;
wire  [127:0]  u0_col_out_485;
wire  [127:0]  u0_col_out_486;
wire  [127:0]  u0_col_out_487;
wire  [127:0]  u0_col_out_488;
wire  [127:0]  u0_col_out_489;
wire  [127:0]  u0_col_out_490;
wire  [127:0]  u0_col_out_491;
wire  [127:0]  u0_col_out_492;
wire  [127:0]  u0_col_out_493;
wire  [127:0]  u0_col_out_494;
wire  [127:0]  u0_col_out_495;
wire  [127:0]  u0_col_out_496;
wire  [127:0]  u0_col_out_497;
wire  [127:0]  u0_col_out_498;
wire  [127:0]  u0_col_out_499;
wire  [127:0]  u0_col_out_500;
wire  [127:0]  u0_col_out_501;
wire  [127:0]  u0_col_out_502;
wire  [127:0]  u0_col_out_503;
wire  [127:0]  u0_col_out_504;
wire  [127:0]  u0_col_out_505;
wire  [127:0]  u0_col_out_506;
wire  [127:0]  u0_col_out_507;
wire  [127:0]  u0_col_out_508;
wire  [127:0]  u0_col_out_509;
wire  [127:0]  u0_col_out_510;
wire  [127:0]  u0_col_out_511;
wire  [127:0]  u0_col_out_512;
wire  [127:0]  u0_col_out_513;
wire  [127:0]  u0_col_out_514;
wire  [127:0]  u0_col_out_515;
wire  [127:0]  u0_col_out_516;
wire  [127:0]  u0_col_out_517;
wire  [127:0]  u0_col_out_518;
wire  [127:0]  u0_col_out_519;
wire  [127:0]  u0_col_out_520;
wire  [127:0]  u0_col_out_521;
wire  [127:0]  u0_col_out_522;
wire  [127:0]  u0_col_out_523;
wire  [127:0]  u0_col_out_524;
wire  [127:0]  u0_col_out_525;
wire  [127:0]  u0_col_out_526;
wire  [127:0]  u0_col_out_527;
wire  [127:0]  u0_col_out_528;
wire  [127:0]  u0_col_out_529;
wire  [127:0]  u0_col_out_530;
wire  [127:0]  u0_col_out_531;
wire  [127:0]  u0_col_out_532;
wire  [127:0]  u0_col_out_533;
wire  [127:0]  u0_col_out_534;
wire  [127:0]  u0_col_out_535;
wire  [127:0]  u0_col_out_536;
wire  [127:0]  u0_col_out_537;
wire  [127:0]  u0_col_out_538;
wire  [127:0]  u0_col_out_539;
wire  [127:0]  u0_col_out_540;
wire  [127:0]  u0_col_out_541;
wire  [127:0]  u0_col_out_542;
wire  [127:0]  u0_col_out_543;
wire  [127:0]  u0_col_out_544;
wire  [127:0]  u0_col_out_545;
wire  [127:0]  u0_col_out_546;
wire  [127:0]  u0_col_out_547;
wire  [127:0]  u0_col_out_548;
wire  [127:0]  u0_col_out_549;
wire  [127:0]  u0_col_out_550;
wire  [127:0]  u0_col_out_551;
wire  [127:0]  u0_col_out_552;
wire  [127:0]  u0_col_out_553;
wire  [127:0]  u0_col_out_554;
wire  [127:0]  u0_col_out_555;
wire  [127:0]  u0_col_out_556;
wire  [127:0]  u0_col_out_557;
wire  [127:0]  u0_col_out_558;
wire  [127:0]  u0_col_out_559;
wire  [127:0]  u0_col_out_560;
wire  [127:0]  u0_col_out_561;
wire  [127:0]  u0_col_out_562;
wire  [127:0]  u0_col_out_563;
wire  [127:0]  u0_col_out_564;
wire  [127:0]  u0_col_out_565;
wire  [127:0]  u0_col_out_566;
wire  [127:0]  u0_col_out_567;
wire  [127:0]  u0_col_out_568;
wire  [127:0]  u0_col_out_569;
wire  [127:0]  u0_col_out_570;
wire  [127:0]  u0_col_out_571;
wire  [127:0]  u0_col_out_572;
wire  [127:0]  u0_col_out_573;
wire  [127:0]  u0_col_out_574;
wire  [127:0]  u0_col_out_575;
wire  [127:0]  u0_col_out_576;
wire  [127:0]  u0_col_out_577;
wire  [127:0]  u0_col_out_578;
wire  [127:0]  u0_col_out_579;
wire  [127:0]  u0_col_out_580;
wire  [127:0]  u0_col_out_581;
wire  [127:0]  u0_col_out_582;
wire  [127:0]  u0_col_out_583;
wire  [127:0]  u0_col_out_584;
wire  [127:0]  u0_col_out_585;
wire  [127:0]  u0_col_out_586;
wire  [127:0]  u0_col_out_587;
wire  [127:0]  u0_col_out_588;
wire  [127:0]  u0_col_out_589;
wire  [127:0]  u0_col_out_590;
wire  [127:0]  u0_col_out_591;
wire  [127:0]  u0_col_out_592;
wire  [127:0]  u0_col_out_593;
wire  [127:0]  u0_col_out_594;
wire  [127:0]  u0_col_out_595;
wire  [127:0]  u0_col_out_596;
wire  [127:0]  u0_col_out_597;
wire  [127:0]  u0_col_out_598;
wire  [127:0]  u0_col_out_599;
wire  [127:0]  u0_col_out_600;
wire  [127:0]  u0_col_out_601;
wire  [127:0]  u0_col_out_602;
wire  [127:0]  u0_col_out_603;
wire  [127:0]  u0_col_out_604;
wire  [127:0]  u0_col_out_605;
wire  [127:0]  u0_col_out_606;
wire  [127:0]  u0_col_out_607;
wire  [127:0]  u0_col_out_608;
wire  [127:0]  u0_col_out_609;
wire  [127:0]  u0_col_out_610;
wire  [127:0]  u0_col_out_611;
wire  [127:0]  u0_col_out_612;
wire  [127:0]  u0_col_out_613;
wire  [127:0]  u0_col_out_614;
wire  [127:0]  u0_col_out_615;
wire  [127:0]  u0_col_out_616;
wire  [127:0]  u0_col_out_617;
wire  [127:0]  u0_col_out_618;
wire  [127:0]  u0_col_out_619;
wire  [127:0]  u0_col_out_620;
wire  [127:0]  u0_col_out_621;
wire  [127:0]  u0_col_out_622;
wire  [127:0]  u0_col_out_623;
wire  [127:0]  u0_col_out_624;
wire  [127:0]  u0_col_out_625;
wire  [127:0]  u0_col_out_626;
wire  [127:0]  u0_col_out_627;
wire  [127:0]  u0_col_out_628;
wire  [127:0]  u0_col_out_629;
wire  [127:0]  u0_col_out_630;
wire  [127:0]  u0_col_out_631;
wire  [127:0]  u0_col_out_632;
wire  [127:0]  u0_col_out_633;
wire  [127:0]  u0_col_out_634;
wire  [127:0]  u0_col_out_635;
wire  [127:0]  u0_col_out_636;
wire  [127:0]  u0_col_out_637;
wire  [127:0]  u0_col_out_638;
wire  [127:0]  u0_col_out_639;
wire  [127:0]  u0_col_out_640;
wire  [127:0]  u0_col_out_641;
wire  [127:0]  u0_col_out_642;
wire  [127:0]  u0_col_out_643;
wire  [127:0]  u0_col_out_644;
wire  [127:0]  u0_col_out_645;
wire  [127:0]  u0_col_out_646;
wire  [127:0]  u0_col_out_647;
wire  [127:0]  u0_col_out_648;
wire  [127:0]  u0_col_out_649;
wire  [127:0]  u0_col_out_650;
wire  [127:0]  u0_col_out_651;
wire  [127:0]  u0_col_out_652;
wire  [127:0]  u0_col_out_653;
wire  [127:0]  u0_col_out_654;
wire  [127:0]  u0_col_out_655;
wire  [127:0]  u0_col_out_656;
wire  [127:0]  u0_col_out_657;
wire  [127:0]  u0_col_out_658;
wire  [127:0]  u0_col_out_659;
wire  [127:0]  u0_col_out_660;
wire  [127:0]  u0_col_out_661;
wire  [127:0]  u0_col_out_662;
wire  [127:0]  u0_col_out_663;
wire  [127:0]  u0_col_out_664;
wire  [127:0]  u0_col_out_665;
wire  [127:0]  u0_col_out_666;
wire  [127:0]  u0_col_out_667;
wire  [127:0]  u0_col_out_668;
wire  [127:0]  u0_col_out_669;
wire  [127:0]  u0_col_out_670;
wire  [127:0]  u0_col_out_671;
wire  [127:0]  u0_col_out_672;
wire  [127:0]  u0_col_out_673;
wire  [127:0]  u0_col_out_674;
wire  [127:0]  u0_col_out_675;
wire  [127:0]  u0_col_out_676;
wire  [127:0]  u0_col_out_677;
wire  [127:0]  u0_col_out_678;
wire  [127:0]  u0_col_out_679;
wire  [127:0]  u0_col_out_680;
wire  [127:0]  u0_col_out_681;
wire  [127:0]  u0_col_out_682;
wire  [127:0]  u0_col_out_683;
wire  [127:0]  u0_col_out_684;
wire  [127:0]  u0_col_out_685;
wire  [127:0]  u0_col_out_686;
wire  [127:0]  u0_col_out_687;
wire  [127:0]  u0_col_out_688;
wire  [127:0]  u0_col_out_689;
wire  [127:0]  u0_col_out_690;
wire  [127:0]  u0_col_out_691;
wire  [127:0]  u0_col_out_692;
wire  [127:0]  u0_col_out_693;
wire  [127:0]  u0_col_out_694;
wire  [127:0]  u0_col_out_695;
wire  [127:0]  u0_col_out_696;
wire  [127:0]  u0_col_out_697;
wire  [127:0]  u0_col_out_698;
wire  [127:0]  u0_col_out_699;
wire  [127:0]  u0_col_out_700;
wire  [127:0]  u0_col_out_701;
wire  [127:0]  u0_col_out_702;
wire  [127:0]  u0_col_out_703;
wire  [127:0]  u0_col_out_704;
wire  [127:0]  u0_col_out_705;
wire  [127:0]  u0_col_out_706;
wire  [127:0]  u0_col_out_707;
wire  [127:0]  u0_col_out_708;
wire  [127:0]  u0_col_out_709;
wire  [127:0]  u0_col_out_710;
wire  [127:0]  u0_col_out_711;
wire  [127:0]  u0_col_out_712;
wire  [127:0]  u0_col_out_713;
wire  [127:0]  u0_col_out_714;
wire  [127:0]  u0_col_out_715;
wire  [127:0]  u0_col_out_716;
wire  [127:0]  u0_col_out_717;
wire  [127:0]  u0_col_out_718;
wire  [127:0]  u0_col_out_719;
wire  [127:0]  u0_col_out_720;
wire  [127:0]  u0_col_out_721;
wire  [127:0]  u0_col_out_722;
wire  [127:0]  u0_col_out_723;
wire  [127:0]  u0_col_out_724;
wire  [127:0]  u0_col_out_725;
wire  [127:0]  u0_col_out_726;
wire  [127:0]  u0_col_out_727;
wire  [127:0]  u0_col_out_728;
wire  [127:0]  u0_col_out_729;
wire  [127:0]  u0_col_out_730;
wire  [127:0]  u0_col_out_731;
wire  [127:0]  u0_col_out_732;
wire  [127:0]  u0_col_out_733;
wire  [127:0]  u0_col_out_734;
wire  [127:0]  u0_col_out_735;
wire  [127:0]  u0_col_out_736;
wire  [127:0]  u0_col_out_737;
wire  [127:0]  u0_col_out_738;
wire  [127:0]  u0_col_out_739;
wire  [127:0]  u0_col_out_740;
wire  [127:0]  u0_col_out_741;
wire  [127:0]  u0_col_out_742;
wire  [127:0]  u0_col_out_743;
wire  [127:0]  u0_col_out_744;
wire  [127:0]  u0_col_out_745;
wire  [127:0]  u0_col_out_746;
wire  [127:0]  u0_col_out_747;
wire  [127:0]  u0_col_out_748;
wire  [127:0]  u0_col_out_749;
wire  [127:0]  u0_col_out_750;
wire  [127:0]  u0_col_out_751;
wire  [127:0]  u0_col_out_752;
wire  [127:0]  u0_col_out_753;
wire  [127:0]  u0_col_out_754;
wire  [127:0]  u0_col_out_755;
wire  [127:0]  u0_col_out_756;
wire  [127:0]  u0_col_out_757;
wire  [127:0]  u0_col_out_758;
wire  [127:0]  u0_col_out_759;
wire  [127:0]  u0_col_out_760;
wire  [127:0]  u0_col_out_761;
wire  [127:0]  u0_col_out_762;
wire  [127:0]  u0_col_out_763;
wire  [127:0]  u0_col_out_764;
wire  [127:0]  u0_col_out_765;
wire  [127:0]  u0_col_out_766;
wire  [127:0]  u0_col_out_767;
wire  [127:0]  u0_col_out_768;
wire  [127:0]  u0_col_out_769;
wire  [127:0]  u0_col_out_770;
wire  [127:0]  u0_col_out_771;
wire  [127:0]  u0_col_out_772;
wire  [127:0]  u0_col_out_773;
wire  [127:0]  u0_col_out_774;
wire  [127:0]  u0_col_out_775;
wire  [127:0]  u0_col_out_776;
wire  [127:0]  u0_col_out_777;
wire  [127:0]  u0_col_out_778;
wire  [127:0]  u0_col_out_779;
wire  [127:0]  u0_col_out_780;
wire  [127:0]  u0_col_out_781;
wire  [127:0]  u0_col_out_782;
wire  [127:0]  u0_col_out_783;
wire  [127:0]  u0_col_out_784;
wire  [127:0]  u0_col_out_785;
wire  [127:0]  u0_col_out_786;
wire  [127:0]  u0_col_out_787;
wire  [127:0]  u0_col_out_788;
wire  [127:0]  u0_col_out_789;
wire  [127:0]  u0_col_out_790;
wire  [127:0]  u0_col_out_791;
wire  [127:0]  u0_col_out_792;
wire  [127:0]  u0_col_out_793;
wire  [127:0]  u0_col_out_794;
wire  [127:0]  u0_col_out_795;
wire  [127:0]  u0_col_out_796;
wire  [127:0]  u0_col_out_797;
wire  [127:0]  u0_col_out_798;
wire  [127:0]  u0_col_out_799;
wire  [127:0]  u0_col_out_800;
wire  [127:0]  u0_col_out_801;
wire  [127:0]  u0_col_out_802;
wire  [127:0]  u0_col_out_803;
wire  [127:0]  u0_col_out_804;
wire  [127:0]  u0_col_out_805;
wire  [127:0]  u0_col_out_806;
wire  [127:0]  u0_col_out_807;
wire  [127:0]  u0_col_out_808;
wire  [127:0]  u0_col_out_809;
wire  [127:0]  u0_col_out_810;
wire  [127:0]  u0_col_out_811;
wire  [127:0]  u0_col_out_812;
wire  [127:0]  u0_col_out_813;
wire  [127:0]  u0_col_out_814;
wire  [127:0]  u0_col_out_815;
wire  [127:0]  u0_col_out_816;
wire  [127:0]  u0_col_out_817;
wire  [127:0]  u0_col_out_818;
wire  [127:0]  u0_col_out_819;
wire  [127:0]  u0_col_out_820;
wire  [127:0]  u0_col_out_821;
wire  [127:0]  u0_col_out_822;
wire  [127:0]  u0_col_out_823;
wire  [127:0]  u0_col_out_824;
wire  [127:0]  u0_col_out_825;
wire  [127:0]  u0_col_out_826;
wire  [127:0]  u0_col_out_827;
wire  [127:0]  u0_col_out_828;
wire  [127:0]  u0_col_out_829;
wire  [127:0]  u0_col_out_830;
wire  [127:0]  u0_col_out_831;
wire  [127:0]  u0_col_out_832;
wire  [127:0]  u0_col_out_833;
wire  [127:0]  u0_col_out_834;
wire  [127:0]  u0_col_out_835;
wire  [127:0]  u0_col_out_836;
wire  [127:0]  u0_col_out_837;
wire  [127:0]  u0_col_out_838;
wire  [127:0]  u0_col_out_839;
wire  [127:0]  u0_col_out_840;
wire  [127:0]  u0_col_out_841;
wire  [127:0]  u0_col_out_842;
wire  [127:0]  u0_col_out_843;
wire  [127:0]  u0_col_out_844;
wire  [127:0]  u0_col_out_845;
wire  [127:0]  u0_col_out_846;
wire  [127:0]  u0_col_out_847;
wire  [127:0]  u0_col_out_848;
wire  [127:0]  u0_col_out_849;
wire  [127:0]  u0_col_out_850;
wire  [127:0]  u0_col_out_851;
wire  [127:0]  u0_col_out_852;
wire  [127:0]  u0_col_out_853;
wire  [127:0]  u0_col_out_854;
wire  [127:0]  u0_col_out_855;
wire  [127:0]  u0_col_out_856;
wire  [127:0]  u0_col_out_857;
wire  [127:0]  u0_col_out_858;
wire  [127:0]  u0_col_out_859;
wire  [127:0]  u0_col_out_860;
wire  [127:0]  u0_col_out_861;
wire  [127:0]  u0_col_out_862;
wire  [127:0]  u0_col_out_863;
wire  [127:0]  u0_col_out_864;
wire  [127:0]  u0_col_out_865;
wire  [127:0]  u0_col_out_866;
wire  [127:0]  u0_col_out_867;
wire  [127:0]  u0_col_out_868;
wire  [127:0]  u0_col_out_869;
wire  [127:0]  u0_col_out_870;
wire  [127:0]  u0_col_out_871;
wire  [127:0]  u0_col_out_872;
wire  [127:0]  u0_col_out_873;
wire  [127:0]  u0_col_out_874;
wire  [127:0]  u0_col_out_875;
wire  [127:0]  u0_col_out_876;
wire  [127:0]  u0_col_out_877;
wire  [127:0]  u0_col_out_878;
wire  [127:0]  u0_col_out_879;
wire  [127:0]  u0_col_out_880;
wire  [127:0]  u0_col_out_881;
wire  [127:0]  u0_col_out_882;
wire  [127:0]  u0_col_out_883;
wire  [127:0]  u0_col_out_884;
wire  [127:0]  u0_col_out_885;
wire  [127:0]  u0_col_out_886;
wire  [127:0]  u0_col_out_887;
wire  [127:0]  u0_col_out_888;
wire  [127:0]  u0_col_out_889;
wire  [127:0]  u0_col_out_890;
wire  [127:0]  u0_col_out_891;
wire  [127:0]  u0_col_out_892;
wire  [127:0]  u0_col_out_893;
wire  [127:0]  u0_col_out_894;
wire  [127:0]  u0_col_out_895;
wire  [127:0]  u0_col_out_896;
wire  [127:0]  u0_col_out_897;
wire  [127:0]  u0_col_out_898;
wire  [127:0]  u0_col_out_899;
wire  [127:0]  u0_col_out_900;
wire  [127:0]  u0_col_out_901;
wire  [127:0]  u0_col_out_902;
wire  [127:0]  u0_col_out_903;
wire  [127:0]  u0_col_out_904;
wire  [127:0]  u0_col_out_905;
wire  [127:0]  u0_col_out_906;
wire  [127:0]  u0_col_out_907;
wire  [127:0]  u0_col_out_908;
wire  [127:0]  u0_col_out_909;
wire  [127:0]  u0_col_out_910;
wire  [127:0]  u0_col_out_911;
wire  [127:0]  u0_col_out_912;
wire  [127:0]  u0_col_out_913;
wire  [127:0]  u0_col_out_914;
wire  [127:0]  u0_col_out_915;
wire  [127:0]  u0_col_out_916;
wire  [127:0]  u0_col_out_917;
wire  [127:0]  u0_col_out_918;
wire  [127:0]  u0_col_out_919;
wire  [127:0]  u0_col_out_920;
wire  [127:0]  u0_col_out_921;
wire  [127:0]  u0_col_out_922;
wire  [127:0]  u0_col_out_923;
wire  [127:0]  u0_col_out_924;
wire  [127:0]  u0_col_out_925;
wire  [127:0]  u0_col_out_926;
wire  [127:0]  u0_col_out_927;
wire  [127:0]  u0_col_out_928;
wire  [127:0]  u0_col_out_929;
wire  [127:0]  u0_col_out_930;
wire  [127:0]  u0_col_out_931;
wire  [127:0]  u0_col_out_932;
wire  [127:0]  u0_col_out_933;
wire  [127:0]  u0_col_out_934;
wire  [127:0]  u0_col_out_935;
wire  [127:0]  u0_col_out_936;
wire  [127:0]  u0_col_out_937;
wire  [127:0]  u0_col_out_938;
wire  [127:0]  u0_col_out_939;
wire  [127:0]  u0_col_out_940;
wire  [127:0]  u0_col_out_941;
wire  [127:0]  u0_col_out_942;
wire  [127:0]  u0_col_out_943;
wire  [127:0]  u0_col_out_944;
wire  [127:0]  u0_col_out_945;
wire  [127:0]  u0_col_out_946;
wire  [127:0]  u0_col_out_947;
wire  [127:0]  u0_col_out_948;
wire  [127:0]  u0_col_out_949;
wire  [127:0]  u0_col_out_950;
wire  [127:0]  u0_col_out_951;
wire  [127:0]  u0_col_out_952;
wire  [127:0]  u0_col_out_953;
wire  [127:0]  u0_col_out_954;
wire  [127:0]  u0_col_out_955;
wire  [127:0]  u0_col_out_956;
wire  [127:0]  u0_col_out_957;
wire  [127:0]  u0_col_out_958;
wire  [127:0]  u0_col_out_959;
wire  [127:0]  u0_col_out_960;
wire  [127:0]  u0_col_out_961;
wire  [127:0]  u0_col_out_962;
wire  [127:0]  u0_col_out_963;
wire  [127:0]  u0_col_out_964;
wire  [127:0]  u0_col_out_965;
wire  [127:0]  u0_col_out_966;
wire  [127:0]  u0_col_out_967;
wire  [127:0]  u0_col_out_968;
wire  [127:0]  u0_col_out_969;
wire  [127:0]  u0_col_out_970;
wire  [127:0]  u0_col_out_971;
wire  [127:0]  u0_col_out_972;
wire  [127:0]  u0_col_out_973;
wire  [127:0]  u0_col_out_974;
wire  [127:0]  u0_col_out_975;
wire  [127:0]  u0_col_out_976;
wire  [127:0]  u0_col_out_977;
wire  [127:0]  u0_col_out_978;
wire  [127:0]  u0_col_out_979;
wire  [127:0]  u0_col_out_980;
wire  [127:0]  u0_col_out_981;
wire  [127:0]  u0_col_out_982;
wire  [127:0]  u0_col_out_983;
wire  [127:0]  u0_col_out_984;
wire  [127:0]  u0_col_out_985;
wire  [127:0]  u0_col_out_986;
wire  [127:0]  u0_col_out_987;
wire  [127:0]  u0_col_out_988;
wire  [127:0]  u0_col_out_989;
wire  [127:0]  u0_col_out_990;
wire  [127:0]  u0_col_out_991;
wire  [127:0]  u0_col_out_992;
wire  [127:0]  u0_col_out_993;
wire  [127:0]  u0_col_out_994;
wire  [127:0]  u0_col_out_995;
wire  [127:0]  u0_col_out_996;
wire  [127:0]  u0_col_out_997;
wire  [127:0]  u0_col_out_998;
wire  [127:0]  u0_col_out_999;
wire  [127:0]  u0_col_out_1000;
wire  [127:0]  u0_col_out_1001;
wire  [127:0]  u0_col_out_1002;
wire  [127:0]  u0_col_out_1003;
wire  [127:0]  u0_col_out_1004;
wire  [127:0]  u0_col_out_1005;
wire  [127:0]  u0_col_out_1006;
wire  [127:0]  u0_col_out_1007;
wire  [127:0]  u0_col_out_1008;
wire  [127:0]  u0_col_out_1009;
wire  [127:0]  u0_col_out_1010;
wire  [127:0]  u0_col_out_1011;
wire  [127:0]  u0_col_out_1012;
wire  [127:0]  u0_col_out_1013;
wire  [127:0]  u0_col_out_1014;
wire  [127:0]  u0_col_out_1015;
wire  [127:0]  u0_col_out_1016;
wire  [127:0]  u0_col_out_1017;
wire  [127:0]  u0_col_out_1018;
wire  [127:0]  u0_col_out_1019;
wire  [127:0]  u0_col_out_1020;
wire  [127:0]  u0_col_out_1021;
wire  [127:0]  u0_col_out_1022;
wire  [127:0]  u0_col_out_1023;
wire  [127:0]  u0_col_out_1024;
wire  [127:0]  u0_col_out_1025;
wire  [127:0]  u0_col_out_1026;
wire  [127:0]  u0_col_out_1027;
wire  [127:0]  u0_col_out_1028;
wire  [127:0]  u0_col_out_1029;
wire  [127:0]  u0_col_out_1030;
wire  [127:0]  u0_col_out_1031;
wire  [127:0]  u0_col_out_1032;
wire  [127:0]  u0_col_out_1033;
wire  [127:0]  u0_col_out_1034;
wire  [127:0]  u0_col_out_1035;
wire  [127:0]  u0_col_out_1036;
wire  [127:0]  u0_col_out_1037;
wire  [127:0]  u0_col_out_1038;
wire  [127:0]  u0_col_out_1039;
wire  [127:0]  u0_col_out_1040;
wire  [127:0]  u0_col_out_1041;
wire  [127:0]  u0_col_out_1042;
wire  [127:0]  u0_col_out_1043;
wire  [127:0]  u0_col_out_1044;
wire  [127:0]  u0_col_out_1045;
wire  [127:0]  u0_col_out_1046;
wire  [127:0]  u0_col_out_1047;
wire  [127:0]  u0_col_out_1048;
wire  [127:0]  u0_col_out_1049;
wire  [127:0]  u0_col_out_1050;
wire  [127:0]  u0_col_out_1051;
wire  [127:0]  u0_col_out_1052;
wire  [127:0]  u0_col_out_1053;
wire  [127:0]  u0_col_out_1054;
wire  [127:0]  u0_col_out_1055;
wire  [127:0]  u0_col_out_1056;
wire  [127:0]  u0_col_out_1057;
wire  [127:0]  u0_col_out_1058;
wire  [127:0]  u0_col_out_1059;
wire  [127:0]  u0_col_out_1060;
wire  [127:0]  u0_col_out_1061;
wire  [127:0]  u0_col_out_1062;
wire  [127:0]  u0_col_out_1063;
wire  [127:0]  u0_col_out_1064;
wire  [127:0]  u0_col_out_1065;
wire  [127:0]  u0_col_out_1066;
wire  [127:0]  u0_col_out_1067;
wire  [127:0]  u0_col_out_1068;
wire  [127:0]  u0_col_out_1069;
wire  [127:0]  u0_col_out_1070;
wire  [127:0]  u0_col_out_1071;
wire  [127:0]  u0_col_out_1072;
wire  [127:0]  u0_col_out_1073;
wire  [127:0]  u0_col_out_1074;
wire  [127:0]  u0_col_out_1075;
wire  [127:0]  u0_col_out_1076;
wire  [127:0]  u0_col_out_1077;
wire  [127:0]  u0_col_out_1078;
wire  [127:0]  u0_col_out_1079;
wire  [127:0]  u0_col_out_1080;
wire  [127:0]  u0_col_out_1081;
wire  [127:0]  u0_col_out_1082;
wire  [127:0]  u0_col_out_1083;
wire  [127:0]  u0_col_out_1084;
wire  [127:0]  u0_col_out_1085;
wire  [127:0]  u0_col_out_1086;
wire  [127:0]  u0_col_out_1087;
wire  [127:0]  u0_col_out_1088;
wire  [127:0]  u0_col_out_1089;
wire  [127:0]  u0_col_out_1090;
wire  [127:0]  u0_col_out_1091;
wire  [127:0]  u0_col_out_1092;
wire  [127:0]  u0_col_out_1093;
wire  [127:0]  u0_col_out_1094;
wire  [127:0]  u0_col_out_1095;
wire  [127:0]  u0_col_out_1096;
wire  [127:0]  u0_col_out_1097;
wire  [127:0]  u0_col_out_1098;
wire  [127:0]  u0_col_out_1099;
wire  [127:0]  u0_col_out_1100;
wire  [127:0]  u0_col_out_1101;
wire  [127:0]  u0_col_out_1102;
wire  [127:0]  u0_col_out_1103;
wire  [127:0]  u0_col_out_1104;
wire  [127:0]  u0_col_out_1105;
wire  [127:0]  u0_col_out_1106;
wire  [127:0]  u0_col_out_1107;
wire  [127:0]  u0_col_out_1108;
wire  [127:0]  u0_col_out_1109;
wire  [127:0]  u0_col_out_1110;
wire  [127:0]  u0_col_out_1111;
wire  [127:0]  u0_col_out_1112;
wire  [127:0]  u0_col_out_1113;
wire  [127:0]  u0_col_out_1114;
wire  [127:0]  u0_col_out_1115;
wire  [127:0]  u0_col_out_1116;
wire  [127:0]  u0_col_out_1117;
wire  [127:0]  u0_col_out_1118;
wire  [127:0]  u0_col_out_1119;
wire  [127:0]  u0_col_out_1120;
wire  [127:0]  u0_col_out_1121;
wire  [127:0]  u0_col_out_1122;
wire  [127:0]  u0_col_out_1123;
wire  [127:0]  u0_col_out_1124;
wire  [127:0]  u0_col_out_1125;
wire  [127:0]  u0_col_out_1126;
wire  [127:0]  u0_col_out_1127;
wire  [127:0]  u0_col_out_1128;
wire  [127:0]  u0_col_out_1129;
wire  [127:0]  u0_col_out_1130;
wire  [127:0]  u0_col_out_1131;
wire  [127:0]  u0_col_out_1132;
wire  [127:0]  u0_col_out_1133;
wire  [127:0]  u0_col_out_1134;
wire  [127:0]  u0_col_out_1135;
wire  [127:0]  u0_col_out_1136;
wire  [127:0]  u0_col_out_1137;
wire  [127:0]  u0_col_out_1138;
wire  [127:0]  u0_col_out_1139;
wire  [127:0]  u0_col_out_1140;
wire  [127:0]  u0_col_out_1141;
wire  [127:0]  u0_col_out_1142;
wire  [127:0]  u0_col_out_1143;
wire  [127:0]  u0_col_out_1144;
wire  [127:0]  u0_col_out_1145;
wire  [127:0]  u0_col_out_1146;
wire  [127:0]  u0_col_out_1147;
wire  [127:0]  u0_col_out_1148;
wire  [127:0]  u0_col_out_1149;
wire  [127:0]  u0_col_out_1150;
wire  [127:0]  u0_col_out_1151;
wire  [127:0]  u0_col_out_1152;
wire  [127:0]  u0_col_out_1153;
wire  [127:0]  u0_col_out_1154;
wire  [127:0]  u0_col_out_1155;
wire  [127:0]  u0_col_out_1156;
wire  [127:0]  u0_col_out_1157;
wire  [127:0]  u0_col_out_1158;
wire  [127:0]  u0_col_out_1159;
wire  [127:0]  u0_col_out_1160;
wire  [127:0]  u0_col_out_1161;
wire  [127:0]  u0_col_out_1162;
wire  [127:0]  u0_col_out_1163;
wire  [127:0]  u0_col_out_1164;
wire  [127:0]  u0_col_out_1165;
wire  [127:0]  u0_col_out_1166;
wire  [127:0]  u0_col_out_1167;
wire  [127:0]  u0_col_out_1168;
wire  [127:0]  u0_col_out_1169;
wire  [127:0]  u0_col_out_1170;
wire  [127:0]  u0_col_out_1171;
wire  [127:0]  u0_col_out_1172;
wire  [127:0]  u0_col_out_1173;
wire  [127:0]  u0_col_out_1174;
wire  [127:0]  u0_col_out_1175;
wire  [127:0]  u0_col_out_1176;
wire  [127:0]  u0_col_out_1177;
wire  [127:0]  u0_col_out_1178;
wire  [127:0]  u0_col_out_1179;
wire  [127:0]  u0_col_out_1180;
wire  [127:0]  u0_col_out_1181;
wire  [127:0]  u0_col_out_1182;
wire  [127:0]  u0_col_out_1183;
wire  [127:0]  u0_col_out_1184;
wire  [127:0]  u0_col_out_1185;
wire  [127:0]  u0_col_out_1186;
wire  [127:0]  u0_col_out_1187;
wire  [127:0]  u0_col_out_1188;
wire  [127:0]  u0_col_out_1189;
wire  [127:0]  u0_col_out_1190;
wire  [127:0]  u0_col_out_1191;
wire  [127:0]  u0_col_out_1192;
wire  [127:0]  u0_col_out_1193;
wire  [127:0]  u0_col_out_1194;
wire  [127:0]  u0_col_out_1195;
wire  [127:0]  u0_col_out_1196;
wire  [127:0]  u0_col_out_1197;
wire  [127:0]  u0_col_out_1198;
wire  [127:0]  u0_col_out_1199;
wire  [127:0]  u0_col_out_1200;
wire  [127:0]  u0_col_out_1201;
wire  [127:0]  u0_col_out_1202;
wire  [127:0]  u0_col_out_1203;
wire  [127:0]  u0_col_out_1204;
wire  [127:0]  u0_col_out_1205;
wire  [127:0]  u0_col_out_1206;
wire  [127:0]  u0_col_out_1207;
wire  [127:0]  u0_col_out_1208;
wire  [127:0]  u0_col_out_1209;
wire  [127:0]  u0_col_out_1210;
wire  [127:0]  u0_col_out_1211;
wire  [127:0]  u0_col_out_1212;
wire  [127:0]  u0_col_out_1213;
wire  [127:0]  u0_col_out_1214;
wire  [127:0]  u0_col_out_1215;
wire  [127:0]  u0_col_out_1216;
wire  [127:0]  u0_col_out_1217;
wire  [127:0]  u0_col_out_1218;
wire  [127:0]  u0_col_out_1219;
wire  [127:0]  u0_col_out_1220;
wire  [127:0]  u0_col_out_1221;
wire  [127:0]  u0_col_out_1222;
wire  [127:0]  u0_col_out_1223;
wire  [127:0]  u0_col_out_1224;
wire  [127:0]  u0_col_out_1225;
wire  [127:0]  u0_col_out_1226;
wire  [127:0]  u0_col_out_1227;
wire  [127:0]  u0_col_out_1228;
wire  [127:0]  u0_col_out_1229;
wire  [127:0]  u0_col_out_1230;
wire  [127:0]  u0_col_out_1231;
wire  [127:0]  u0_col_out_1232;
wire  [127:0]  u0_col_out_1233;
wire  [127:0]  u0_col_out_1234;
wire  [127:0]  u0_col_out_1235;
wire  [127:0]  u0_col_out_1236;
wire  [127:0]  u0_col_out_1237;
wire  [127:0]  u0_col_out_1238;
wire  [127:0]  u0_col_out_1239;
wire  [127:0]  u0_col_out_1240;
wire  [127:0]  u0_col_out_1241;
wire  [127:0]  u0_col_out_1242;
wire  [127:0]  u0_col_out_1243;
wire  [127:0]  u0_col_out_1244;
wire  [127:0]  u0_col_out_1245;
wire  [127:0]  u0_col_out_1246;
wire  [127:0]  u0_col_out_1247;
wire  [127:0]  u0_col_out_1248;
wire  [127:0]  u0_col_out_1249;
wire  [127:0]  u0_col_out_1250;
wire  [127:0]  u0_col_out_1251;
wire  [127:0]  u0_col_out_1252;
wire  [127:0]  u0_col_out_1253;
wire  [127:0]  u0_col_out_1254;
wire  [127:0]  u0_col_out_1255;
wire  [127:0]  u0_col_out_1256;
wire  [127:0]  u0_col_out_1257;
wire  [127:0]  u0_col_out_1258;
wire  [127:0]  u0_col_out_1259;
wire  [127:0]  u0_col_out_1260;
wire  [127:0]  u0_col_out_1261;
wire  [127:0]  u0_col_out_1262;
wire  [127:0]  u0_col_out_1263;
wire  [127:0]  u0_col_out_1264;
wire  [127:0]  u0_col_out_1265;
wire  [127:0]  u0_col_out_1266;
wire  [127:0]  u0_col_out_1267;
wire  [127:0]  u0_col_out_1268;
wire  [127:0]  u0_col_out_1269;
wire  [127:0]  u0_col_out_1270;
wire  [127:0]  u0_col_out_1271;
wire  [127:0]  u0_col_out_1272;
wire  [127:0]  u0_col_out_1273;
wire  [127:0]  u0_col_out_1274;
wire  [127:0]  u0_col_out_1275;
wire  [127:0]  u0_col_out_1276;
wire  [127:0]  u0_col_out_1277;
wire  [127:0]  u0_col_out_1278;
wire  [127:0]  u0_col_out_1279;




msq_product_period4  u0_msq_product_period4 (
    .al                      ( u0_al         ),
    .sel                     ( reg_u0_sel        ),

    .col_0                   ( u0_col_out_0      ),
    .col_1                   ( u0_col_out_1      ),
    .col_2                   ( u0_col_out_2      ),
    .col_3                   ( u0_col_out_3      ),
    .col_4                   ( u0_col_out_4      ),
    .col_5                   ( u0_col_out_5      ),
    .col_6                   ( u0_col_out_6      ),
    .col_7                   ( u0_col_out_7      ),
    .col_8                   ( u0_col_out_8      ),
    .col_9                   ( u0_col_out_9      ),
    .col_10                  ( u0_col_out_10     ),
    .col_11                  ( u0_col_out_11     ),
    .col_12                  ( u0_col_out_12     ),
    .col_13                  ( u0_col_out_13     ),
    .col_14                  ( u0_col_out_14     ),
    .col_15                  ( u0_col_out_15     ),
    .col_16                  ( u0_col_out_16     ),
    .col_17                  ( u0_col_out_17     ),
    .col_18                  ( u0_col_out_18     ),
    .col_19                  ( u0_col_out_19     ),
    .col_20                  ( u0_col_out_20     ),
    .col_21                  ( u0_col_out_21     ),
    .col_22                  ( u0_col_out_22     ),
    .col_23                  ( u0_col_out_23     ),
    .col_24                  ( u0_col_out_24     ),
    .col_25                  ( u0_col_out_25     ),
    .col_26                  ( u0_col_out_26     ),
    .col_27                  ( u0_col_out_27     ),
    .col_28                  ( u0_col_out_28     ),
    .col_29                  ( u0_col_out_29     ),
    .col_30                  ( u0_col_out_30     ),
    .col_31                  ( u0_col_out_31     ),
    .col_32                  ( u0_col_out_32     ),
    .col_33                  ( u0_col_out_33     ),
    .col_34                  ( u0_col_out_34     ),
    .col_35                  ( u0_col_out_35     ),
    .col_36                  ( u0_col_out_36     ),
    .col_37                  ( u0_col_out_37     ),
    .col_38                  ( u0_col_out_38     ),
    .col_39                  ( u0_col_out_39     ),
    .col_40                  ( u0_col_out_40     ),
    .col_41                  ( u0_col_out_41     ),
    .col_42                  ( u0_col_out_42     ),
    .col_43                  ( u0_col_out_43     ),
    .col_44                  ( u0_col_out_44     ),
    .col_45                  ( u0_col_out_45     ),
    .col_46                  ( u0_col_out_46     ),
    .col_47                  ( u0_col_out_47     ),
    .col_48                  ( u0_col_out_48     ),
    .col_49                  ( u0_col_out_49     ),
    .col_50                  ( u0_col_out_50     ),
    .col_51                  ( u0_col_out_51     ),
    .col_52                  ( u0_col_out_52     ),
    .col_53                  ( u0_col_out_53     ),
    .col_54                  ( u0_col_out_54     ),
    .col_55                  ( u0_col_out_55     ),
    .col_56                  ( u0_col_out_56     ),
    .col_57                  ( u0_col_out_57     ),
    .col_58                  ( u0_col_out_58     ),
    .col_59                  ( u0_col_out_59     ),
    .col_60                  ( u0_col_out_60     ),
    .col_61                  ( u0_col_out_61     ),
    .col_62                  ( u0_col_out_62     ),
    .col_63                  ( u0_col_out_63     ),
    .col_64                  ( u0_col_out_64     ),
    .col_65                  ( u0_col_out_65     ),
    .col_66                  ( u0_col_out_66     ),
    .col_67                  ( u0_col_out_67     ),
    .col_68                  ( u0_col_out_68     ),
    .col_69                  ( u0_col_out_69     ),
    .col_70                  ( u0_col_out_70     ),
    .col_71                  ( u0_col_out_71     ),
    .col_72                  ( u0_col_out_72     ),
    .col_73                  ( u0_col_out_73     ),
    .col_74                  ( u0_col_out_74     ),
    .col_75                  ( u0_col_out_75     ),
    .col_76                  ( u0_col_out_76     ),
    .col_77                  ( u0_col_out_77     ),
    .col_78                  ( u0_col_out_78     ),
    .col_79                  ( u0_col_out_79     ),
    .col_80                  ( u0_col_out_80     ),
    .col_81                  ( u0_col_out_81     ),
    .col_82                  ( u0_col_out_82     ),
    .col_83                  ( u0_col_out_83     ),
    .col_84                  ( u0_col_out_84     ),
    .col_85                  ( u0_col_out_85     ),
    .col_86                  ( u0_col_out_86     ),
    .col_87                  ( u0_col_out_87     ),
    .col_88                  ( u0_col_out_88     ),
    .col_89                  ( u0_col_out_89     ),
    .col_90                  ( u0_col_out_90     ),
    .col_91                  ( u0_col_out_91     ),
    .col_92                  ( u0_col_out_92     ),
    .col_93                  ( u0_col_out_93     ),
    .col_94                  ( u0_col_out_94     ),
    .col_95                  ( u0_col_out_95     ),
    .col_96                  ( u0_col_out_96     ),
    .col_97                  ( u0_col_out_97     ),
    .col_98                  ( u0_col_out_98     ),
    .col_99                  ( u0_col_out_99     ),
    .col_100                 ( u0_col_out_100    ),
    .col_101                 ( u0_col_out_101    ),
    .col_102                 ( u0_col_out_102    ),
    .col_103                 ( u0_col_out_103    ),
    .col_104                 ( u0_col_out_104    ),
    .col_105                 ( u0_col_out_105    ),
    .col_106                 ( u0_col_out_106    ),
    .col_107                 ( u0_col_out_107    ),
    .col_108                 ( u0_col_out_108    ),
    .col_109                 ( u0_col_out_109    ),
    .col_110                 ( u0_col_out_110    ),
    .col_111                 ( u0_col_out_111    ),
    .col_112                 ( u0_col_out_112    ),
    .col_113                 ( u0_col_out_113    ),
    .col_114                 ( u0_col_out_114    ),
    .col_115                 ( u0_col_out_115    ),
    .col_116                 ( u0_col_out_116    ),
    .col_117                 ( u0_col_out_117    ),
    .col_118                 ( u0_col_out_118    ),
    .col_119                 ( u0_col_out_119    ),
    .col_120                 ( u0_col_out_120    ),
    .col_121                 ( u0_col_out_121    ),
    .col_122                 ( u0_col_out_122    ),
    .col_123                 ( u0_col_out_123    ),
    .col_124                 ( u0_col_out_124    ),
    .col_125                 ( u0_col_out_125    ),
    .col_126                 ( u0_col_out_126    ),
    .col_127                 ( u0_col_out_127    ),
    .col_128                 ( u0_col_out_128    ),
    .col_129                 ( u0_col_out_129    ),
    .col_130                 ( u0_col_out_130    ),
    .col_131                 ( u0_col_out_131    ),
    .col_132                 ( u0_col_out_132    ),
    .col_133                 ( u0_col_out_133    ),
    .col_134                 ( u0_col_out_134    ),
    .col_135                 ( u0_col_out_135    ),
    .col_136                 ( u0_col_out_136    ),
    .col_137                 ( u0_col_out_137    ),
    .col_138                 ( u0_col_out_138    ),
    .col_139                 ( u0_col_out_139    ),
    .col_140                 ( u0_col_out_140    ),
    .col_141                 ( u0_col_out_141    ),
    .col_142                 ( u0_col_out_142    ),
    .col_143                 ( u0_col_out_143    ),
    .col_144                 ( u0_col_out_144    ),
    .col_145                 ( u0_col_out_145    ),
    .col_146                 ( u0_col_out_146    ),
    .col_147                 ( u0_col_out_147    ),
    .col_148                 ( u0_col_out_148    ),
    .col_149                 ( u0_col_out_149    ),
    .col_150                 ( u0_col_out_150    ),
    .col_151                 ( u0_col_out_151    ),
    .col_152                 ( u0_col_out_152    ),
    .col_153                 ( u0_col_out_153    ),
    .col_154                 ( u0_col_out_154    ),
    .col_155                 ( u0_col_out_155    ),
    .col_156                 ( u0_col_out_156    ),
    .col_157                 ( u0_col_out_157    ),
    .col_158                 ( u0_col_out_158    ),
    .col_159                 ( u0_col_out_159    ),
    .col_160                 ( u0_col_out_160    ),
    .col_161                 ( u0_col_out_161    ),
    .col_162                 ( u0_col_out_162    ),
    .col_163                 ( u0_col_out_163    ),
    .col_164                 ( u0_col_out_164    ),
    .col_165                 ( u0_col_out_165    ),
    .col_166                 ( u0_col_out_166    ),
    .col_167                 ( u0_col_out_167    ),
    .col_168                 ( u0_col_out_168    ),
    .col_169                 ( u0_col_out_169    ),
    .col_170                 ( u0_col_out_170    ),
    .col_171                 ( u0_col_out_171    ),
    .col_172                 ( u0_col_out_172    ),
    .col_173                 ( u0_col_out_173    ),
    .col_174                 ( u0_col_out_174    ),
    .col_175                 ( u0_col_out_175    ),
    .col_176                 ( u0_col_out_176    ),
    .col_177                 ( u0_col_out_177    ),
    .col_178                 ( u0_col_out_178    ),
    .col_179                 ( u0_col_out_179    ),
    .col_180                 ( u0_col_out_180    ),
    .col_181                 ( u0_col_out_181    ),
    .col_182                 ( u0_col_out_182    ),
    .col_183                 ( u0_col_out_183    ),
    .col_184                 ( u0_col_out_184    ),
    .col_185                 ( u0_col_out_185    ),
    .col_186                 ( u0_col_out_186    ),
    .col_187                 ( u0_col_out_187    ),
    .col_188                 ( u0_col_out_188    ),
    .col_189                 ( u0_col_out_189    ),
    .col_190                 ( u0_col_out_190    ),
    .col_191                 ( u0_col_out_191    ),
    .col_192                 ( u0_col_out_192    ),
    .col_193                 ( u0_col_out_193    ),
    .col_194                 ( u0_col_out_194    ),
    .col_195                 ( u0_col_out_195    ),
    .col_196                 ( u0_col_out_196    ),
    .col_197                 ( u0_col_out_197    ),
    .col_198                 ( u0_col_out_198    ),
    .col_199                 ( u0_col_out_199    ),
    .col_200                 ( u0_col_out_200    ),
    .col_201                 ( u0_col_out_201    ),
    .col_202                 ( u0_col_out_202    ),
    .col_203                 ( u0_col_out_203    ),
    .col_204                 ( u0_col_out_204    ),
    .col_205                 ( u0_col_out_205    ),
    .col_206                 ( u0_col_out_206    ),
    .col_207                 ( u0_col_out_207    ),
    .col_208                 ( u0_col_out_208    ),
    .col_209                 ( u0_col_out_209    ),
    .col_210                 ( u0_col_out_210    ),
    .col_211                 ( u0_col_out_211    ),
    .col_212                 ( u0_col_out_212    ),
    .col_213                 ( u0_col_out_213    ),
    .col_214                 ( u0_col_out_214    ),
    .col_215                 ( u0_col_out_215    ),
    .col_216                 ( u0_col_out_216    ),
    .col_217                 ( u0_col_out_217    ),
    .col_218                 ( u0_col_out_218    ),
    .col_219                 ( u0_col_out_219    ),
    .col_220                 ( u0_col_out_220    ),
    .col_221                 ( u0_col_out_221    ),
    .col_222                 ( u0_col_out_222    ),
    .col_223                 ( u0_col_out_223    ),
    .col_224                 ( u0_col_out_224    ),
    .col_225                 ( u0_col_out_225    ),
    .col_226                 ( u0_col_out_226    ),
    .col_227                 ( u0_col_out_227    ),
    .col_228                 ( u0_col_out_228    ),
    .col_229                 ( u0_col_out_229    ),
    .col_230                 ( u0_col_out_230    ),
    .col_231                 ( u0_col_out_231    ),
    .col_232                 ( u0_col_out_232    ),
    .col_233                 ( u0_col_out_233    ),
    .col_234                 ( u0_col_out_234    ),
    .col_235                 ( u0_col_out_235    ),
    .col_236                 ( u0_col_out_236    ),
    .col_237                 ( u0_col_out_237    ),
    .col_238                 ( u0_col_out_238    ),
    .col_239                 ( u0_col_out_239    ),
    .col_240                 ( u0_col_out_240    ),
    .col_241                 ( u0_col_out_241    ),
    .col_242                 ( u0_col_out_242    ),
    .col_243                 ( u0_col_out_243    ),
    .col_244                 ( u0_col_out_244    ),
    .col_245                 ( u0_col_out_245    ),
    .col_246                 ( u0_col_out_246    ),
    .col_247                 ( u0_col_out_247    ),
    .col_248                 ( u0_col_out_248    ),
    .col_249                 ( u0_col_out_249    ),
    .col_250                 ( u0_col_out_250    ),
    .col_251                 ( u0_col_out_251    ),
    .col_252                 ( u0_col_out_252    ),
    .col_253                 ( u0_col_out_253    ),
    .col_254                 ( u0_col_out_254    ),
    .col_255                 ( u0_col_out_255    ),
    .col_256                 ( u0_col_out_256    ),
    .col_257                 ( u0_col_out_257    ),
    .col_258                 ( u0_col_out_258    ),
    .col_259                 ( u0_col_out_259    ),
    .col_260                 ( u0_col_out_260    ),
    .col_261                 ( u0_col_out_261    ),
    .col_262                 ( u0_col_out_262    ),
    .col_263                 ( u0_col_out_263    ),
    .col_264                 ( u0_col_out_264    ),
    .col_265                 ( u0_col_out_265    ),
    .col_266                 ( u0_col_out_266    ),
    .col_267                 ( u0_col_out_267    ),
    .col_268                 ( u0_col_out_268    ),
    .col_269                 ( u0_col_out_269    ),
    .col_270                 ( u0_col_out_270    ),
    .col_271                 ( u0_col_out_271    ),
    .col_272                 ( u0_col_out_272    ),
    .col_273                 ( u0_col_out_273    ),
    .col_274                 ( u0_col_out_274    ),
    .col_275                 ( u0_col_out_275    ),
    .col_276                 ( u0_col_out_276    ),
    .col_277                 ( u0_col_out_277    ),
    .col_278                 ( u0_col_out_278    ),
    .col_279                 ( u0_col_out_279    ),
    .col_280                 ( u0_col_out_280    ),
    .col_281                 ( u0_col_out_281    ),
    .col_282                 ( u0_col_out_282    ),
    .col_283                 ( u0_col_out_283    ),
    .col_284                 ( u0_col_out_284    ),
    .col_285                 ( u0_col_out_285    ),
    .col_286                 ( u0_col_out_286    ),
    .col_287                 ( u0_col_out_287    ),
    .col_288                 ( u0_col_out_288    ),
    .col_289                 ( u0_col_out_289    ),
    .col_290                 ( u0_col_out_290    ),
    .col_291                 ( u0_col_out_291    ),
    .col_292                 ( u0_col_out_292    ),
    .col_293                 ( u0_col_out_293    ),
    .col_294                 ( u0_col_out_294    ),
    .col_295                 ( u0_col_out_295    ),
    .col_296                 ( u0_col_out_296    ),
    .col_297                 ( u0_col_out_297    ),
    .col_298                 ( u0_col_out_298    ),
    .col_299                 ( u0_col_out_299    ),
    .col_300                 ( u0_col_out_300    ),
    .col_301                 ( u0_col_out_301    ),
    .col_302                 ( u0_col_out_302    ),
    .col_303                 ( u0_col_out_303    ),
    .col_304                 ( u0_col_out_304    ),
    .col_305                 ( u0_col_out_305    ),
    .col_306                 ( u0_col_out_306    ),
    .col_307                 ( u0_col_out_307    ),
    .col_308                 ( u0_col_out_308    ),
    .col_309                 ( u0_col_out_309    ),
    .col_310                 ( u0_col_out_310    ),
    .col_311                 ( u0_col_out_311    ),
    .col_312                 ( u0_col_out_312    ),
    .col_313                 ( u0_col_out_313    ),
    .col_314                 ( u0_col_out_314    ),
    .col_315                 ( u0_col_out_315    ),
    .col_316                 ( u0_col_out_316    ),
    .col_317                 ( u0_col_out_317    ),
    .col_318                 ( u0_col_out_318    ),
    .col_319                 ( u0_col_out_319    ),
    .col_320                 ( u0_col_out_320    ),
    .col_321                 ( u0_col_out_321    ),
    .col_322                 ( u0_col_out_322    ),
    .col_323                 ( u0_col_out_323    ),
    .col_324                 ( u0_col_out_324    ),
    .col_325                 ( u0_col_out_325    ),
    .col_326                 ( u0_col_out_326    ),
    .col_327                 ( u0_col_out_327    ),
    .col_328                 ( u0_col_out_328    ),
    .col_329                 ( u0_col_out_329    ),
    .col_330                 ( u0_col_out_330    ),
    .col_331                 ( u0_col_out_331    ),
    .col_332                 ( u0_col_out_332    ),
    .col_333                 ( u0_col_out_333    ),
    .col_334                 ( u0_col_out_334    ),
    .col_335                 ( u0_col_out_335    ),
    .col_336                 ( u0_col_out_336    ),
    .col_337                 ( u0_col_out_337    ),
    .col_338                 ( u0_col_out_338    ),
    .col_339                 ( u0_col_out_339    ),
    .col_340                 ( u0_col_out_340    ),
    .col_341                 ( u0_col_out_341    ),
    .col_342                 ( u0_col_out_342    ),
    .col_343                 ( u0_col_out_343    ),
    .col_344                 ( u0_col_out_344    ),
    .col_345                 ( u0_col_out_345    ),
    .col_346                 ( u0_col_out_346    ),
    .col_347                 ( u0_col_out_347    ),
    .col_348                 ( u0_col_out_348    ),
    .col_349                 ( u0_col_out_349    ),
    .col_350                 ( u0_col_out_350    ),
    .col_351                 ( u0_col_out_351    ),
    .col_352                 ( u0_col_out_352    ),
    .col_353                 ( u0_col_out_353    ),
    .col_354                 ( u0_col_out_354    ),
    .col_355                 ( u0_col_out_355    ),
    .col_356                 ( u0_col_out_356    ),
    .col_357                 ( u0_col_out_357    ),
    .col_358                 ( u0_col_out_358    ),
    .col_359                 ( u0_col_out_359    ),
    .col_360                 ( u0_col_out_360    ),
    .col_361                 ( u0_col_out_361    ),
    .col_362                 ( u0_col_out_362    ),
    .col_363                 ( u0_col_out_363    ),
    .col_364                 ( u0_col_out_364    ),
    .col_365                 ( u0_col_out_365    ),
    .col_366                 ( u0_col_out_366    ),
    .col_367                 ( u0_col_out_367    ),
    .col_368                 ( u0_col_out_368    ),
    .col_369                 ( u0_col_out_369    ),
    .col_370                 ( u0_col_out_370    ),
    .col_371                 ( u0_col_out_371    ),
    .col_372                 ( u0_col_out_372    ),
    .col_373                 ( u0_col_out_373    ),
    .col_374                 ( u0_col_out_374    ),
    .col_375                 ( u0_col_out_375    ),
    .col_376                 ( u0_col_out_376    ),
    .col_377                 ( u0_col_out_377    ),
    .col_378                 ( u0_col_out_378    ),
    .col_379                 ( u0_col_out_379    ),
    .col_380                 ( u0_col_out_380    ),
    .col_381                 ( u0_col_out_381    ),
    .col_382                 ( u0_col_out_382    ),
    .col_383                 ( u0_col_out_383    ),
    .col_384                 ( u0_col_out_384    ),
    .col_385                 ( u0_col_out_385    ),
    .col_386                 ( u0_col_out_386    ),
    .col_387                 ( u0_col_out_387    ),
    .col_388                 ( u0_col_out_388    ),
    .col_389                 ( u0_col_out_389    ),
    .col_390                 ( u0_col_out_390    ),
    .col_391                 ( u0_col_out_391    ),
    .col_392                 ( u0_col_out_392    ),
    .col_393                 ( u0_col_out_393    ),
    .col_394                 ( u0_col_out_394    ),
    .col_395                 ( u0_col_out_395    ),
    .col_396                 ( u0_col_out_396    ),
    .col_397                 ( u0_col_out_397    ),
    .col_398                 ( u0_col_out_398    ),
    .col_399                 ( u0_col_out_399    ),
    .col_400                 ( u0_col_out_400    ),
    .col_401                 ( u0_col_out_401    ),
    .col_402                 ( u0_col_out_402    ),
    .col_403                 ( u0_col_out_403    ),
    .col_404                 ( u0_col_out_404    ),
    .col_405                 ( u0_col_out_405    ),
    .col_406                 ( u0_col_out_406    ),
    .col_407                 ( u0_col_out_407    ),
    .col_408                 ( u0_col_out_408    ),
    .col_409                 ( u0_col_out_409    ),
    .col_410                 ( u0_col_out_410    ),
    .col_411                 ( u0_col_out_411    ),
    .col_412                 ( u0_col_out_412    ),
    .col_413                 ( u0_col_out_413    ),
    .col_414                 ( u0_col_out_414    ),
    .col_415                 ( u0_col_out_415    ),
    .col_416                 ( u0_col_out_416    ),
    .col_417                 ( u0_col_out_417    ),
    .col_418                 ( u0_col_out_418    ),
    .col_419                 ( u0_col_out_419    ),
    .col_420                 ( u0_col_out_420    ),
    .col_421                 ( u0_col_out_421    ),
    .col_422                 ( u0_col_out_422    ),
    .col_423                 ( u0_col_out_423    ),
    .col_424                 ( u0_col_out_424    ),
    .col_425                 ( u0_col_out_425    ),
    .col_426                 ( u0_col_out_426    ),
    .col_427                 ( u0_col_out_427    ),
    .col_428                 ( u0_col_out_428    ),
    .col_429                 ( u0_col_out_429    ),
    .col_430                 ( u0_col_out_430    ),
    .col_431                 ( u0_col_out_431    ),
    .col_432                 ( u0_col_out_432    ),
    .col_433                 ( u0_col_out_433    ),
    .col_434                 ( u0_col_out_434    ),
    .col_435                 ( u0_col_out_435    ),
    .col_436                 ( u0_col_out_436    ),
    .col_437                 ( u0_col_out_437    ),
    .col_438                 ( u0_col_out_438    ),
    .col_439                 ( u0_col_out_439    ),
    .col_440                 ( u0_col_out_440    ),
    .col_441                 ( u0_col_out_441    ),
    .col_442                 ( u0_col_out_442    ),
    .col_443                 ( u0_col_out_443    ),
    .col_444                 ( u0_col_out_444    ),
    .col_445                 ( u0_col_out_445    ),
    .col_446                 ( u0_col_out_446    ),
    .col_447                 ( u0_col_out_447    ),
    .col_448                 ( u0_col_out_448    ),
    .col_449                 ( u0_col_out_449    ),
    .col_450                 ( u0_col_out_450    ),
    .col_451                 ( u0_col_out_451    ),
    .col_452                 ( u0_col_out_452    ),
    .col_453                 ( u0_col_out_453    ),
    .col_454                 ( u0_col_out_454    ),
    .col_455                 ( u0_col_out_455    ),
    .col_456                 ( u0_col_out_456    ),
    .col_457                 ( u0_col_out_457    ),
    .col_458                 ( u0_col_out_458    ),
    .col_459                 ( u0_col_out_459    ),
    .col_460                 ( u0_col_out_460    ),
    .col_461                 ( u0_col_out_461    ),
    .col_462                 ( u0_col_out_462    ),
    .col_463                 ( u0_col_out_463    ),
    .col_464                 ( u0_col_out_464    ),
    .col_465                 ( u0_col_out_465    ),
    .col_466                 ( u0_col_out_466    ),
    .col_467                 ( u0_col_out_467    ),
    .col_468                 ( u0_col_out_468    ),
    .col_469                 ( u0_col_out_469    ),
    .col_470                 ( u0_col_out_470    ),
    .col_471                 ( u0_col_out_471    ),
    .col_472                 ( u0_col_out_472    ),
    .col_473                 ( u0_col_out_473    ),
    .col_474                 ( u0_col_out_474    ),
    .col_475                 ( u0_col_out_475    ),
    .col_476                 ( u0_col_out_476    ),
    .col_477                 ( u0_col_out_477    ),
    .col_478                 ( u0_col_out_478    ),
    .col_479                 ( u0_col_out_479    ),
    .col_480                 ( u0_col_out_480    ),
    .col_481                 ( u0_col_out_481    ),
    .col_482                 ( u0_col_out_482    ),
    .col_483                 ( u0_col_out_483    ),
    .col_484                 ( u0_col_out_484    ),
    .col_485                 ( u0_col_out_485    ),
    .col_486                 ( u0_col_out_486    ),
    .col_487                 ( u0_col_out_487    ),
    .col_488                 ( u0_col_out_488    ),
    .col_489                 ( u0_col_out_489    ),
    .col_490                 ( u0_col_out_490    ),
    .col_491                 ( u0_col_out_491    ),
    .col_492                 ( u0_col_out_492    ),
    .col_493                 ( u0_col_out_493    ),
    .col_494                 ( u0_col_out_494    ),
    .col_495                 ( u0_col_out_495    ),
    .col_496                 ( u0_col_out_496    ),
    .col_497                 ( u0_col_out_497    ),
    .col_498                 ( u0_col_out_498    ),
    .col_499                 ( u0_col_out_499    ),
    .col_500                 ( u0_col_out_500    ),
    .col_501                 ( u0_col_out_501    ),
    .col_502                 ( u0_col_out_502    ),
    .col_503                 ( u0_col_out_503    ),
    .col_504                 ( u0_col_out_504    ),
    .col_505                 ( u0_col_out_505    ),
    .col_506                 ( u0_col_out_506    ),
    .col_507                 ( u0_col_out_507    ),
    .col_508                 ( u0_col_out_508    ),
    .col_509                 ( u0_col_out_509    ),
    .col_510                 ( u0_col_out_510    ),
    .col_511                 ( u0_col_out_511    ),
    .col_512                 ( u0_col_out_512    ),
    .col_513                 ( u0_col_out_513    ),
    .col_514                 ( u0_col_out_514    ),
    .col_515                 ( u0_col_out_515    ),
    .col_516                 ( u0_col_out_516    ),
    .col_517                 ( u0_col_out_517    ),
    .col_518                 ( u0_col_out_518    ),
    .col_519                 ( u0_col_out_519    ),
    .col_520                 ( u0_col_out_520    ),
    .col_521                 ( u0_col_out_521    ),
    .col_522                 ( u0_col_out_522    ),
    .col_523                 ( u0_col_out_523    ),
    .col_524                 ( u0_col_out_524    ),
    .col_525                 ( u0_col_out_525    ),
    .col_526                 ( u0_col_out_526    ),
    .col_527                 ( u0_col_out_527    ),
    .col_528                 ( u0_col_out_528    ),
    .col_529                 ( u0_col_out_529    ),
    .col_530                 ( u0_col_out_530    ),
    .col_531                 ( u0_col_out_531    ),
    .col_532                 ( u0_col_out_532    ),
    .col_533                 ( u0_col_out_533    ),
    .col_534                 ( u0_col_out_534    ),
    .col_535                 ( u0_col_out_535    ),
    .col_536                 ( u0_col_out_536    ),
    .col_537                 ( u0_col_out_537    ),
    .col_538                 ( u0_col_out_538    ),
    .col_539                 ( u0_col_out_539    ),
    .col_540                 ( u0_col_out_540    ),
    .col_541                 ( u0_col_out_541    ),
    .col_542                 ( u0_col_out_542    ),
    .col_543                 ( u0_col_out_543    ),
    .col_544                 ( u0_col_out_544    ),
    .col_545                 ( u0_col_out_545    ),
    .col_546                 ( u0_col_out_546    ),
    .col_547                 ( u0_col_out_547    ),
    .col_548                 ( u0_col_out_548    ),
    .col_549                 ( u0_col_out_549    ),
    .col_550                 ( u0_col_out_550    ),
    .col_551                 ( u0_col_out_551    ),
    .col_552                 ( u0_col_out_552    ),
    .col_553                 ( u0_col_out_553    ),
    .col_554                 ( u0_col_out_554    ),
    .col_555                 ( u0_col_out_555    ),
    .col_556                 ( u0_col_out_556    ),
    .col_557                 ( u0_col_out_557    ),
    .col_558                 ( u0_col_out_558    ),
    .col_559                 ( u0_col_out_559    ),
    .col_560                 ( u0_col_out_560    ),
    .col_561                 ( u0_col_out_561    ),
    .col_562                 ( u0_col_out_562    ),
    .col_563                 ( u0_col_out_563    ),
    .col_564                 ( u0_col_out_564    ),
    .col_565                 ( u0_col_out_565    ),
    .col_566                 ( u0_col_out_566    ),
    .col_567                 ( u0_col_out_567    ),
    .col_568                 ( u0_col_out_568    ),
    .col_569                 ( u0_col_out_569    ),
    .col_570                 ( u0_col_out_570    ),
    .col_571                 ( u0_col_out_571    ),
    .col_572                 ( u0_col_out_572    ),
    .col_573                 ( u0_col_out_573    ),
    .col_574                 ( u0_col_out_574    ),
    .col_575                 ( u0_col_out_575    ),
    .col_576                 ( u0_col_out_576    ),
    .col_577                 ( u0_col_out_577    ),
    .col_578                 ( u0_col_out_578    ),
    .col_579                 ( u0_col_out_579    ),
    .col_580                 ( u0_col_out_580    ),
    .col_581                 ( u0_col_out_581    ),
    .col_582                 ( u0_col_out_582    ),
    .col_583                 ( u0_col_out_583    ),
    .col_584                 ( u0_col_out_584    ),
    .col_585                 ( u0_col_out_585    ),
    .col_586                 ( u0_col_out_586    ),
    .col_587                 ( u0_col_out_587    ),
    .col_588                 ( u0_col_out_588    ),
    .col_589                 ( u0_col_out_589    ),
    .col_590                 ( u0_col_out_590    ),
    .col_591                 ( u0_col_out_591    ),
    .col_592                 ( u0_col_out_592    ),
    .col_593                 ( u0_col_out_593    ),
    .col_594                 ( u0_col_out_594    ),
    .col_595                 ( u0_col_out_595    ),
    .col_596                 ( u0_col_out_596    ),
    .col_597                 ( u0_col_out_597    ),
    .col_598                 ( u0_col_out_598    ),
    .col_599                 ( u0_col_out_599    ),
    .col_600                 ( u0_col_out_600    ),
    .col_601                 ( u0_col_out_601    ),
    .col_602                 ( u0_col_out_602    ),
    .col_603                 ( u0_col_out_603    ),
    .col_604                 ( u0_col_out_604    ),
    .col_605                 ( u0_col_out_605    ),
    .col_606                 ( u0_col_out_606    ),
    .col_607                 ( u0_col_out_607    ),
    .col_608                 ( u0_col_out_608    ),
    .col_609                 ( u0_col_out_609    ),
    .col_610                 ( u0_col_out_610    ),
    .col_611                 ( u0_col_out_611    ),
    .col_612                 ( u0_col_out_612    ),
    .col_613                 ( u0_col_out_613    ),
    .col_614                 ( u0_col_out_614    ),
    .col_615                 ( u0_col_out_615    ),
    .col_616                 ( u0_col_out_616    ),
    .col_617                 ( u0_col_out_617    ),
    .col_618                 ( u0_col_out_618    ),
    .col_619                 ( u0_col_out_619    ),
    .col_620                 ( u0_col_out_620    ),
    .col_621                 ( u0_col_out_621    ),
    .col_622                 ( u0_col_out_622    ),
    .col_623                 ( u0_col_out_623    ),
    .col_624                 ( u0_col_out_624    ),
    .col_625                 ( u0_col_out_625    ),
    .col_626                 ( u0_col_out_626    ),
    .col_627                 ( u0_col_out_627    ),
    .col_628                 ( u0_col_out_628    ),
    .col_629                 ( u0_col_out_629    ),
    .col_630                 ( u0_col_out_630    ),
    .col_631                 ( u0_col_out_631    ),
    .col_632                 ( u0_col_out_632    ),
    .col_633                 ( u0_col_out_633    ),
    .col_634                 ( u0_col_out_634    ),
    .col_635                 ( u0_col_out_635    ),
    .col_636                 ( u0_col_out_636    ),
    .col_637                 ( u0_col_out_637    ),
    .col_638                 ( u0_col_out_638    ),
    .col_639                 ( u0_col_out_639    ),
    .col_640                 ( u0_col_out_640    ),
    .col_641                 ( u0_col_out_641    ),
    .col_642                 ( u0_col_out_642    ),
    .col_643                 ( u0_col_out_643    ),
    .col_644                 ( u0_col_out_644    ),
    .col_645                 ( u0_col_out_645    ),
    .col_646                 ( u0_col_out_646    ),
    .col_647                 ( u0_col_out_647    ),
    .col_648                 ( u0_col_out_648    ),
    .col_649                 ( u0_col_out_649    ),
    .col_650                 ( u0_col_out_650    ),
    .col_651                 ( u0_col_out_651    ),
    .col_652                 ( u0_col_out_652    ),
    .col_653                 ( u0_col_out_653    ),
    .col_654                 ( u0_col_out_654    ),
    .col_655                 ( u0_col_out_655    ),
    .col_656                 ( u0_col_out_656    ),
    .col_657                 ( u0_col_out_657    ),
    .col_658                 ( u0_col_out_658    ),
    .col_659                 ( u0_col_out_659    ),
    .col_660                 ( u0_col_out_660    ),
    .col_661                 ( u0_col_out_661    ),
    .col_662                 ( u0_col_out_662    ),
    .col_663                 ( u0_col_out_663    ),
    .col_664                 ( u0_col_out_664    ),
    .col_665                 ( u0_col_out_665    ),
    .col_666                 ( u0_col_out_666    ),
    .col_667                 ( u0_col_out_667    ),
    .col_668                 ( u0_col_out_668    ),
    .col_669                 ( u0_col_out_669    ),
    .col_670                 ( u0_col_out_670    ),
    .col_671                 ( u0_col_out_671    ),
    .col_672                 ( u0_col_out_672    ),
    .col_673                 ( u0_col_out_673    ),
    .col_674                 ( u0_col_out_674    ),
    .col_675                 ( u0_col_out_675    ),
    .col_676                 ( u0_col_out_676    ),
    .col_677                 ( u0_col_out_677    ),
    .col_678                 ( u0_col_out_678    ),
    .col_679                 ( u0_col_out_679    ),
    .col_680                 ( u0_col_out_680    ),
    .col_681                 ( u0_col_out_681    ),
    .col_682                 ( u0_col_out_682    ),
    .col_683                 ( u0_col_out_683    ),
    .col_684                 ( u0_col_out_684    ),
    .col_685                 ( u0_col_out_685    ),
    .col_686                 ( u0_col_out_686    ),
    .col_687                 ( u0_col_out_687    ),
    .col_688                 ( u0_col_out_688    ),
    .col_689                 ( u0_col_out_689    ),
    .col_690                 ( u0_col_out_690    ),
    .col_691                 ( u0_col_out_691    ),
    .col_692                 ( u0_col_out_692    ),
    .col_693                 ( u0_col_out_693    ),
    .col_694                 ( u0_col_out_694    ),
    .col_695                 ( u0_col_out_695    ),
    .col_696                 ( u0_col_out_696    ),
    .col_697                 ( u0_col_out_697    ),
    .col_698                 ( u0_col_out_698    ),
    .col_699                 ( u0_col_out_699    ),
    .col_700                 ( u0_col_out_700    ),
    .col_701                 ( u0_col_out_701    ),
    .col_702                 ( u0_col_out_702    ),
    .col_703                 ( u0_col_out_703    ),
    .col_704                 ( u0_col_out_704    ),
    .col_705                 ( u0_col_out_705    ),
    .col_706                 ( u0_col_out_706    ),
    .col_707                 ( u0_col_out_707    ),
    .col_708                 ( u0_col_out_708    ),
    .col_709                 ( u0_col_out_709    ),
    .col_710                 ( u0_col_out_710    ),
    .col_711                 ( u0_col_out_711    ),
    .col_712                 ( u0_col_out_712    ),
    .col_713                 ( u0_col_out_713    ),
    .col_714                 ( u0_col_out_714    ),
    .col_715                 ( u0_col_out_715    ),
    .col_716                 ( u0_col_out_716    ),
    .col_717                 ( u0_col_out_717    ),
    .col_718                 ( u0_col_out_718    ),
    .col_719                 ( u0_col_out_719    ),
    .col_720                 ( u0_col_out_720    ),
    .col_721                 ( u0_col_out_721    ),
    .col_722                 ( u0_col_out_722    ),
    .col_723                 ( u0_col_out_723    ),
    .col_724                 ( u0_col_out_724    ),
    .col_725                 ( u0_col_out_725    ),
    .col_726                 ( u0_col_out_726    ),
    .col_727                 ( u0_col_out_727    ),
    .col_728                 ( u0_col_out_728    ),
    .col_729                 ( u0_col_out_729    ),
    .col_730                 ( u0_col_out_730    ),
    .col_731                 ( u0_col_out_731    ),
    .col_732                 ( u0_col_out_732    ),
    .col_733                 ( u0_col_out_733    ),
    .col_734                 ( u0_col_out_734    ),
    .col_735                 ( u0_col_out_735    ),
    .col_736                 ( u0_col_out_736    ),
    .col_737                 ( u0_col_out_737    ),
    .col_738                 ( u0_col_out_738    ),
    .col_739                 ( u0_col_out_739    ),
    .col_740                 ( u0_col_out_740    ),
    .col_741                 ( u0_col_out_741    ),
    .col_742                 ( u0_col_out_742    ),
    .col_743                 ( u0_col_out_743    ),
    .col_744                 ( u0_col_out_744    ),
    .col_745                 ( u0_col_out_745    ),
    .col_746                 ( u0_col_out_746    ),
    .col_747                 ( u0_col_out_747    ),
    .col_748                 ( u0_col_out_748    ),
    .col_749                 ( u0_col_out_749    ),
    .col_750                 ( u0_col_out_750    ),
    .col_751                 ( u0_col_out_751    ),
    .col_752                 ( u0_col_out_752    ),
    .col_753                 ( u0_col_out_753    ),
    .col_754                 ( u0_col_out_754    ),
    .col_755                 ( u0_col_out_755    ),
    .col_756                 ( u0_col_out_756    ),
    .col_757                 ( u0_col_out_757    ),
    .col_758                 ( u0_col_out_758    ),
    .col_759                 ( u0_col_out_759    ),
    .col_760                 ( u0_col_out_760    ),
    .col_761                 ( u0_col_out_761    ),
    .col_762                 ( u0_col_out_762    ),
    .col_763                 ( u0_col_out_763    ),
    .col_764                 ( u0_col_out_764    ),
    .col_765                 ( u0_col_out_765    ),
    .col_766                 ( u0_col_out_766    ),
    .col_767                 ( u0_col_out_767    ),
    .col_768                 ( u0_col_out_768    ),
    .col_769                 ( u0_col_out_769    ),
    .col_770                 ( u0_col_out_770    ),
    .col_771                 ( u0_col_out_771    ),
    .col_772                 ( u0_col_out_772    ),
    .col_773                 ( u0_col_out_773    ),
    .col_774                 ( u0_col_out_774    ),
    .col_775                 ( u0_col_out_775    ),
    .col_776                 ( u0_col_out_776    ),
    .col_777                 ( u0_col_out_777    ),
    .col_778                 ( u0_col_out_778    ),
    .col_779                 ( u0_col_out_779    ),
    .col_780                 ( u0_col_out_780    ),
    .col_781                 ( u0_col_out_781    ),
    .col_782                 ( u0_col_out_782    ),
    .col_783                 ( u0_col_out_783    ),
    .col_784                 ( u0_col_out_784    ),
    .col_785                 ( u0_col_out_785    ),
    .col_786                 ( u0_col_out_786    ),
    .col_787                 ( u0_col_out_787    ),
    .col_788                 ( u0_col_out_788    ),
    .col_789                 ( u0_col_out_789    ),
    .col_790                 ( u0_col_out_790    ),
    .col_791                 ( u0_col_out_791    ),
    .col_792                 ( u0_col_out_792    ),
    .col_793                 ( u0_col_out_793    ),
    .col_794                 ( u0_col_out_794    ),
    .col_795                 ( u0_col_out_795    ),
    .col_796                 ( u0_col_out_796    ),
    .col_797                 ( u0_col_out_797    ),
    .col_798                 ( u0_col_out_798    ),
    .col_799                 ( u0_col_out_799    ),
    .col_800                 ( u0_col_out_800    ),
    .col_801                 ( u0_col_out_801    ),
    .col_802                 ( u0_col_out_802    ),
    .col_803                 ( u0_col_out_803    ),
    .col_804                 ( u0_col_out_804    ),
    .col_805                 ( u0_col_out_805    ),
    .col_806                 ( u0_col_out_806    ),
    .col_807                 ( u0_col_out_807    ),
    .col_808                 ( u0_col_out_808    ),
    .col_809                 ( u0_col_out_809    ),
    .col_810                 ( u0_col_out_810    ),
    .col_811                 ( u0_col_out_811    ),
    .col_812                 ( u0_col_out_812    ),
    .col_813                 ( u0_col_out_813    ),
    .col_814                 ( u0_col_out_814    ),
    .col_815                 ( u0_col_out_815    ),
    .col_816                 ( u0_col_out_816    ),
    .col_817                 ( u0_col_out_817    ),
    .col_818                 ( u0_col_out_818    ),
    .col_819                 ( u0_col_out_819    ),
    .col_820                 ( u0_col_out_820    ),
    .col_821                 ( u0_col_out_821    ),
    .col_822                 ( u0_col_out_822    ),
    .col_823                 ( u0_col_out_823    ),
    .col_824                 ( u0_col_out_824    ),
    .col_825                 ( u0_col_out_825    ),
    .col_826                 ( u0_col_out_826    ),
    .col_827                 ( u0_col_out_827    ),
    .col_828                 ( u0_col_out_828    ),
    .col_829                 ( u0_col_out_829    ),
    .col_830                 ( u0_col_out_830    ),
    .col_831                 ( u0_col_out_831    ),
    .col_832                 ( u0_col_out_832    ),
    .col_833                 ( u0_col_out_833    ),
    .col_834                 ( u0_col_out_834    ),
    .col_835                 ( u0_col_out_835    ),
    .col_836                 ( u0_col_out_836    ),
    .col_837                 ( u0_col_out_837    ),
    .col_838                 ( u0_col_out_838    ),
    .col_839                 ( u0_col_out_839    ),
    .col_840                 ( u0_col_out_840    ),
    .col_841                 ( u0_col_out_841    ),
    .col_842                 ( u0_col_out_842    ),
    .col_843                 ( u0_col_out_843    ),
    .col_844                 ( u0_col_out_844    ),
    .col_845                 ( u0_col_out_845    ),
    .col_846                 ( u0_col_out_846    ),
    .col_847                 ( u0_col_out_847    ),
    .col_848                 ( u0_col_out_848    ),
    .col_849                 ( u0_col_out_849    ),
    .col_850                 ( u0_col_out_850    ),
    .col_851                 ( u0_col_out_851    ),
    .col_852                 ( u0_col_out_852    ),
    .col_853                 ( u0_col_out_853    ),
    .col_854                 ( u0_col_out_854    ),
    .col_855                 ( u0_col_out_855    ),
    .col_856                 ( u0_col_out_856    ),
    .col_857                 ( u0_col_out_857    ),
    .col_858                 ( u0_col_out_858    ),
    .col_859                 ( u0_col_out_859    ),
    .col_860                 ( u0_col_out_860    ),
    .col_861                 ( u0_col_out_861    ),
    .col_862                 ( u0_col_out_862    ),
    .col_863                 ( u0_col_out_863    ),
    .col_864                 ( u0_col_out_864    ),
    .col_865                 ( u0_col_out_865    ),
    .col_866                 ( u0_col_out_866    ),
    .col_867                 ( u0_col_out_867    ),
    .col_868                 ( u0_col_out_868    ),
    .col_869                 ( u0_col_out_869    ),
    .col_870                 ( u0_col_out_870    ),
    .col_871                 ( u0_col_out_871    ),
    .col_872                 ( u0_col_out_872    ),
    .col_873                 ( u0_col_out_873    ),
    .col_874                 ( u0_col_out_874    ),
    .col_875                 ( u0_col_out_875    ),
    .col_876                 ( u0_col_out_876    ),
    .col_877                 ( u0_col_out_877    ),
    .col_878                 ( u0_col_out_878    ),
    .col_879                 ( u0_col_out_879    ),
    .col_880                 ( u0_col_out_880    ),
    .col_881                 ( u0_col_out_881    ),
    .col_882                 ( u0_col_out_882    ),
    .col_883                 ( u0_col_out_883    ),
    .col_884                 ( u0_col_out_884    ),
    .col_885                 ( u0_col_out_885    ),
    .col_886                 ( u0_col_out_886    ),
    .col_887                 ( u0_col_out_887    ),
    .col_888                 ( u0_col_out_888    ),
    .col_889                 ( u0_col_out_889    ),
    .col_890                 ( u0_col_out_890    ),
    .col_891                 ( u0_col_out_891    ),
    .col_892                 ( u0_col_out_892    ),
    .col_893                 ( u0_col_out_893    ),
    .col_894                 ( u0_col_out_894    ),
    .col_895                 ( u0_col_out_895    ),
    .col_896                 ( u0_col_out_896    ),
    .col_897                 ( u0_col_out_897    ),
    .col_898                 ( u0_col_out_898    ),
    .col_899                 ( u0_col_out_899    ),
    .col_900                 ( u0_col_out_900    ),
    .col_901                 ( u0_col_out_901    ),
    .col_902                 ( u0_col_out_902    ),
    .col_903                 ( u0_col_out_903    ),
    .col_904                 ( u0_col_out_904    ),
    .col_905                 ( u0_col_out_905    ),
    .col_906                 ( u0_col_out_906    ),
    .col_907                 ( u0_col_out_907    ),
    .col_908                 ( u0_col_out_908    ),
    .col_909                 ( u0_col_out_909    ),
    .col_910                 ( u0_col_out_910    ),
    .col_911                 ( u0_col_out_911    ),
    .col_912                 ( u0_col_out_912    ),
    .col_913                 ( u0_col_out_913    ),
    .col_914                 ( u0_col_out_914    ),
    .col_915                 ( u0_col_out_915    ),
    .col_916                 ( u0_col_out_916    ),
    .col_917                 ( u0_col_out_917    ),
    .col_918                 ( u0_col_out_918    ),
    .col_919                 ( u0_col_out_919    ),
    .col_920                 ( u0_col_out_920    ),
    .col_921                 ( u0_col_out_921    ),
    .col_922                 ( u0_col_out_922    ),
    .col_923                 ( u0_col_out_923    ),
    .col_924                 ( u0_col_out_924    ),
    .col_925                 ( u0_col_out_925    ),
    .col_926                 ( u0_col_out_926    ),
    .col_927                 ( u0_col_out_927    ),
    .col_928                 ( u0_col_out_928    ),
    .col_929                 ( u0_col_out_929    ),
    .col_930                 ( u0_col_out_930    ),
    .col_931                 ( u0_col_out_931    ),
    .col_932                 ( u0_col_out_932    ),
    .col_933                 ( u0_col_out_933    ),
    .col_934                 ( u0_col_out_934    ),
    .col_935                 ( u0_col_out_935    ),
    .col_936                 ( u0_col_out_936    ),
    .col_937                 ( u0_col_out_937    ),
    .col_938                 ( u0_col_out_938    ),
    .col_939                 ( u0_col_out_939    ),
    .col_940                 ( u0_col_out_940    ),
    .col_941                 ( u0_col_out_941    ),
    .col_942                 ( u0_col_out_942    ),
    .col_943                 ( u0_col_out_943    ),
    .col_944                 ( u0_col_out_944    ),
    .col_945                 ( u0_col_out_945    ),
    .col_946                 ( u0_col_out_946    ),
    .col_947                 ( u0_col_out_947    ),
    .col_948                 ( u0_col_out_948    ),
    .col_949                 ( u0_col_out_949    ),
    .col_950                 ( u0_col_out_950    ),
    .col_951                 ( u0_col_out_951    ),
    .col_952                 ( u0_col_out_952    ),
    .col_953                 ( u0_col_out_953    ),
    .col_954                 ( u0_col_out_954    ),
    .col_955                 ( u0_col_out_955    ),
    .col_956                 ( u0_col_out_956    ),
    .col_957                 ( u0_col_out_957    ),
    .col_958                 ( u0_col_out_958    ),
    .col_959                 ( u0_col_out_959    ),
    .col_960                 ( u0_col_out_960    ),
    .col_961                 ( u0_col_out_961    ),
    .col_962                 ( u0_col_out_962    ),
    .col_963                 ( u0_col_out_963    ),
    .col_964                 ( u0_col_out_964    ),
    .col_965                 ( u0_col_out_965    ),
    .col_966                 ( u0_col_out_966    ),
    .col_967                 ( u0_col_out_967    ),
    .col_968                 ( u0_col_out_968    ),
    .col_969                 ( u0_col_out_969    ),
    .col_970                 ( u0_col_out_970    ),
    .col_971                 ( u0_col_out_971    ),
    .col_972                 ( u0_col_out_972    ),
    .col_973                 ( u0_col_out_973    ),
    .col_974                 ( u0_col_out_974    ),
    .col_975                 ( u0_col_out_975    ),
    .col_976                 ( u0_col_out_976    ),
    .col_977                 ( u0_col_out_977    ),
    .col_978                 ( u0_col_out_978    ),
    .col_979                 ( u0_col_out_979    ),
    .col_980                 ( u0_col_out_980    ),
    .col_981                 ( u0_col_out_981    ),
    .col_982                 ( u0_col_out_982    ),
    .col_983                 ( u0_col_out_983    ),
    .col_984                 ( u0_col_out_984    ),
    .col_985                 ( u0_col_out_985    ),
    .col_986                 ( u0_col_out_986    ),
    .col_987                 ( u0_col_out_987    ),
    .col_988                 ( u0_col_out_988    ),
    .col_989                 ( u0_col_out_989    ),
    .col_990                 ( u0_col_out_990    ),
    .col_991                 ( u0_col_out_991    ),
    .col_992                 ( u0_col_out_992    ),
    .col_993                 ( u0_col_out_993    ),
    .col_994                 ( u0_col_out_994    ),
    .col_995                 ( u0_col_out_995    ),
    .col_996                 ( u0_col_out_996    ),
    .col_997                 ( u0_col_out_997    ),
    .col_998                 ( u0_col_out_998    ),
    .col_999                 ( u0_col_out_999    ),
    .col_1000                ( u0_col_out_1000   ),
    .col_1001                ( u0_col_out_1001   ),
    .col_1002                ( u0_col_out_1002   ),
    .col_1003                ( u0_col_out_1003   ),
    .col_1004                ( u0_col_out_1004   ),
    .col_1005                ( u0_col_out_1005   ),
    .col_1006                ( u0_col_out_1006   ),
    .col_1007                ( u0_col_out_1007   ),
    .col_1008                ( u0_col_out_1008   ),
    .col_1009                ( u0_col_out_1009   ),
    .col_1010                ( u0_col_out_1010   ),
    .col_1011                ( u0_col_out_1011   ),
    .col_1012                ( u0_col_out_1012   ),
    .col_1013                ( u0_col_out_1013   ),
    .col_1014                ( u0_col_out_1014   ),
    .col_1015                ( u0_col_out_1015   ),
    .col_1016                ( u0_col_out_1016   ),
    .col_1017                ( u0_col_out_1017   ),
    .col_1018                ( u0_col_out_1018   ),
    .col_1019                ( u0_col_out_1019   ),
    .col_1020                ( u0_col_out_1020   ),
    .col_1021                ( u0_col_out_1021   ),
    .col_1022                ( u0_col_out_1022   ),
    .col_1023                ( u0_col_out_1023   ),
    .col_1024                ( u0_col_out_1024   ),
    .col_1025                ( u0_col_out_1025   ),
    .col_1026                ( u0_col_out_1026   ),
    .col_1027                ( u0_col_out_1027   ),
    .col_1028                ( u0_col_out_1028   ),
    .col_1029                ( u0_col_out_1029   ),
    .col_1030                ( u0_col_out_1030   ),
    .col_1031                ( u0_col_out_1031   ),
    .col_1032                ( u0_col_out_1032   ),
    .col_1033                ( u0_col_out_1033   ),
    .col_1034                ( u0_col_out_1034   ),
    .col_1035                ( u0_col_out_1035   ),
    .col_1036                ( u0_col_out_1036   ),
    .col_1037                ( u0_col_out_1037   ),
    .col_1038                ( u0_col_out_1038   ),
    .col_1039                ( u0_col_out_1039   ),
    .col_1040                ( u0_col_out_1040   ),
    .col_1041                ( u0_col_out_1041   ),
    .col_1042                ( u0_col_out_1042   ),
    .col_1043                ( u0_col_out_1043   ),
    .col_1044                ( u0_col_out_1044   ),
    .col_1045                ( u0_col_out_1045   ),
    .col_1046                ( u0_col_out_1046   ),
    .col_1047                ( u0_col_out_1047   ),
    .col_1048                ( u0_col_out_1048   ),
    .col_1049                ( u0_col_out_1049   ),
    .col_1050                ( u0_col_out_1050   ),
    .col_1051                ( u0_col_out_1051   ),
    .col_1052                ( u0_col_out_1052   ),
    .col_1053                ( u0_col_out_1053   ),
    .col_1054                ( u0_col_out_1054   ),
    .col_1055                ( u0_col_out_1055   ),
    .col_1056                ( u0_col_out_1056   ),
    .col_1057                ( u0_col_out_1057   ),
    .col_1058                ( u0_col_out_1058   ),
    .col_1059                ( u0_col_out_1059   ),
    .col_1060                ( u0_col_out_1060   ),
    .col_1061                ( u0_col_out_1061   ),
    .col_1062                ( u0_col_out_1062   ),
    .col_1063                ( u0_col_out_1063   ),
    .col_1064                ( u0_col_out_1064   ),
    .col_1065                ( u0_col_out_1065   ),
    .col_1066                ( u0_col_out_1066   ),
    .col_1067                ( u0_col_out_1067   ),
    .col_1068                ( u0_col_out_1068   ),
    .col_1069                ( u0_col_out_1069   ),
    .col_1070                ( u0_col_out_1070   ),
    .col_1071                ( u0_col_out_1071   ),
    .col_1072                ( u0_col_out_1072   ),
    .col_1073                ( u0_col_out_1073   ),
    .col_1074                ( u0_col_out_1074   ),
    .col_1075                ( u0_col_out_1075   ),
    .col_1076                ( u0_col_out_1076   ),
    .col_1077                ( u0_col_out_1077   ),
    .col_1078                ( u0_col_out_1078   ),
    .col_1079                ( u0_col_out_1079   ),
    .col_1080                ( u0_col_out_1080   ),
    .col_1081                ( u0_col_out_1081   ),
    .col_1082                ( u0_col_out_1082   ),
    .col_1083                ( u0_col_out_1083   ),
    .col_1084                ( u0_col_out_1084   ),
    .col_1085                ( u0_col_out_1085   ),
    .col_1086                ( u0_col_out_1086   ),
    .col_1087                ( u0_col_out_1087   ),
    .col_1088                ( u0_col_out_1088   ),
    .col_1089                ( u0_col_out_1089   ),
    .col_1090                ( u0_col_out_1090   ),
    .col_1091                ( u0_col_out_1091   ),
    .col_1092                ( u0_col_out_1092   ),
    .col_1093                ( u0_col_out_1093   ),
    .col_1094                ( u0_col_out_1094   ),
    .col_1095                ( u0_col_out_1095   ),
    .col_1096                ( u0_col_out_1096   ),
    .col_1097                ( u0_col_out_1097   ),
    .col_1098                ( u0_col_out_1098   ),
    .col_1099                ( u0_col_out_1099   ),
    .col_1100                ( u0_col_out_1100   ),
    .col_1101                ( u0_col_out_1101   ),
    .col_1102                ( u0_col_out_1102   ),
    .col_1103                ( u0_col_out_1103   ),
    .col_1104                ( u0_col_out_1104   ),
    .col_1105                ( u0_col_out_1105   ),
    .col_1106                ( u0_col_out_1106   ),
    .col_1107                ( u0_col_out_1107   ),
    .col_1108                ( u0_col_out_1108   ),
    .col_1109                ( u0_col_out_1109   ),
    .col_1110                ( u0_col_out_1110   ),
    .col_1111                ( u0_col_out_1111   ),
    .col_1112                ( u0_col_out_1112   ),
    .col_1113                ( u0_col_out_1113   ),
    .col_1114                ( u0_col_out_1114   ),
    .col_1115                ( u0_col_out_1115   ),
    .col_1116                ( u0_col_out_1116   ),
    .col_1117                ( u0_col_out_1117   ),
    .col_1118                ( u0_col_out_1118   ),
    .col_1119                ( u0_col_out_1119   ),
    .col_1120                ( u0_col_out_1120   ),
    .col_1121                ( u0_col_out_1121   ),
    .col_1122                ( u0_col_out_1122   ),
    .col_1123                ( u0_col_out_1123   ),
    .col_1124                ( u0_col_out_1124   ),
    .col_1125                ( u0_col_out_1125   ),
    .col_1126                ( u0_col_out_1126   ),
    .col_1127                ( u0_col_out_1127   ),
    .col_1128                ( u0_col_out_1128   ),
    .col_1129                ( u0_col_out_1129   ),
    .col_1130                ( u0_col_out_1130   ),
    .col_1131                ( u0_col_out_1131   ),
    .col_1132                ( u0_col_out_1132   ),
    .col_1133                ( u0_col_out_1133   ),
    .col_1134                ( u0_col_out_1134   ),
    .col_1135                ( u0_col_out_1135   ),
    .col_1136                ( u0_col_out_1136   ),
    .col_1137                ( u0_col_out_1137   ),
    .col_1138                ( u0_col_out_1138   ),
    .col_1139                ( u0_col_out_1139   ),
    .col_1140                ( u0_col_out_1140   ),
    .col_1141                ( u0_col_out_1141   ),
    .col_1142                ( u0_col_out_1142   ),
    .col_1143                ( u0_col_out_1143   ),
    .col_1144                ( u0_col_out_1144   ),
    .col_1145                ( u0_col_out_1145   ),
    .col_1146                ( u0_col_out_1146   ),
    .col_1147                ( u0_col_out_1147   ),
    .col_1148                ( u0_col_out_1148   ),
    .col_1149                ( u0_col_out_1149   ),
    .col_1150                ( u0_col_out_1150   ),
    .col_1151                ( u0_col_out_1151   ),
    .col_1152                ( u0_col_out_1152   ),
    .col_1153                ( u0_col_out_1153   ),
    .col_1154                ( u0_col_out_1154   ),
    .col_1155                ( u0_col_out_1155   ),
    .col_1156                ( u0_col_out_1156   ),
    .col_1157                ( u0_col_out_1157   ),
    .col_1158                ( u0_col_out_1158   ),
    .col_1159                ( u0_col_out_1159   ),
    .col_1160                ( u0_col_out_1160   ),
    .col_1161                ( u0_col_out_1161   ),
    .col_1162                ( u0_col_out_1162   ),
    .col_1163                ( u0_col_out_1163   ),
    .col_1164                ( u0_col_out_1164   ),
    .col_1165                ( u0_col_out_1165   ),
    .col_1166                ( u0_col_out_1166   ),
    .col_1167                ( u0_col_out_1167   ),
    .col_1168                ( u0_col_out_1168   ),
    .col_1169                ( u0_col_out_1169   ),
    .col_1170                ( u0_col_out_1170   ),
    .col_1171                ( u0_col_out_1171   ),
    .col_1172                ( u0_col_out_1172   ),
    .col_1173                ( u0_col_out_1173   ),
    .col_1174                ( u0_col_out_1174   ),
    .col_1175                ( u0_col_out_1175   ),
    .col_1176                ( u0_col_out_1176   ),
    .col_1177                ( u0_col_out_1177   ),
    .col_1178                ( u0_col_out_1178   ),
    .col_1179                ( u0_col_out_1179   ),
    .col_1180                ( u0_col_out_1180   ),
    .col_1181                ( u0_col_out_1181   ),
    .col_1182                ( u0_col_out_1182   ),
    .col_1183                ( u0_col_out_1183   ),
    .col_1184                ( u0_col_out_1184   ),
    .col_1185                ( u0_col_out_1185   ),
    .col_1186                ( u0_col_out_1186   ),
    .col_1187                ( u0_col_out_1187   ),
    .col_1188                ( u0_col_out_1188   ),
    .col_1189                ( u0_col_out_1189   ),
    .col_1190                ( u0_col_out_1190   ),
    .col_1191                ( u0_col_out_1191   ),
    .col_1192                ( u0_col_out_1192   ),
    .col_1193                ( u0_col_out_1193   ),
    .col_1194                ( u0_col_out_1194   ),
    .col_1195                ( u0_col_out_1195   ),
    .col_1196                ( u0_col_out_1196   ),
    .col_1197                ( u0_col_out_1197   ),
    .col_1198                ( u0_col_out_1198   ),
    .col_1199                ( u0_col_out_1199   ),
    .col_1200                ( u0_col_out_1200   ),
    .col_1201                ( u0_col_out_1201   ),
    .col_1202                ( u0_col_out_1202   ),
    .col_1203                ( u0_col_out_1203   ),
    .col_1204                ( u0_col_out_1204   ),
    .col_1205                ( u0_col_out_1205   ),
    .col_1206                ( u0_col_out_1206   ),
    .col_1207                ( u0_col_out_1207   ),
    .col_1208                ( u0_col_out_1208   ),
    .col_1209                ( u0_col_out_1209   ),
    .col_1210                ( u0_col_out_1210   ),
    .col_1211                ( u0_col_out_1211   ),
    .col_1212                ( u0_col_out_1212   ),
    .col_1213                ( u0_col_out_1213   ),
    .col_1214                ( u0_col_out_1214   ),
    .col_1215                ( u0_col_out_1215   ),
    .col_1216                ( u0_col_out_1216   ),
    .col_1217                ( u0_col_out_1217   ),
    .col_1218                ( u0_col_out_1218   ),
    .col_1219                ( u0_col_out_1219   ),
    .col_1220                ( u0_col_out_1220   ),
    .col_1221                ( u0_col_out_1221   ),
    .col_1222                ( u0_col_out_1222   ),
    .col_1223                ( u0_col_out_1223   ),
    .col_1224                ( u0_col_out_1224   ),
    .col_1225                ( u0_col_out_1225   ),
    .col_1226                ( u0_col_out_1226   ),
    .col_1227                ( u0_col_out_1227   ),
    .col_1228                ( u0_col_out_1228   ),
    .col_1229                ( u0_col_out_1229   ),
    .col_1230                ( u0_col_out_1230   ),
    .col_1231                ( u0_col_out_1231   ),
    .col_1232                ( u0_col_out_1232   ),
    .col_1233                ( u0_col_out_1233   ),
    .col_1234                ( u0_col_out_1234   ),
    .col_1235                ( u0_col_out_1235   ),
    .col_1236                ( u0_col_out_1236   ),
    .col_1237                ( u0_col_out_1237   ),
    .col_1238                ( u0_col_out_1238   ),
    .col_1239                ( u0_col_out_1239   ),
    .col_1240                ( u0_col_out_1240   ),
    .col_1241                ( u0_col_out_1241   ),
    .col_1242                ( u0_col_out_1242   ),
    .col_1243                ( u0_col_out_1243   ),
    .col_1244                ( u0_col_out_1244   ),
    .col_1245                ( u0_col_out_1245   ),
    .col_1246                ( u0_col_out_1246   ),
    .col_1247                ( u0_col_out_1247   ),
    .col_1248                ( u0_col_out_1248   ),
    .col_1249                ( u0_col_out_1249   ),
    .col_1250                ( u0_col_out_1250   ),
    .col_1251                ( u0_col_out_1251   ),
    .col_1252                ( u0_col_out_1252   ),
    .col_1253                ( u0_col_out_1253   ),
    .col_1254                ( u0_col_out_1254   ),
    .col_1255                ( u0_col_out_1255   ),
    .col_1256                ( u0_col_out_1256   ),
    .col_1257                ( u0_col_out_1257   ),
    .col_1258                ( u0_col_out_1258   ),
    .col_1259                ( u0_col_out_1259   ),
    .col_1260                ( u0_col_out_1260   ),
    .col_1261                ( u0_col_out_1261   ),
    .col_1262                ( u0_col_out_1262   ),
    .col_1263                ( u0_col_out_1263   ),
    .col_1264                ( u0_col_out_1264   ),
    .col_1265                ( u0_col_out_1265   ),
    .col_1266                ( u0_col_out_1266   ),
    .col_1267                ( u0_col_out_1267   ),
    .col_1268                ( u0_col_out_1268   ),
    .col_1269                ( u0_col_out_1269   ),
    .col_1270                ( u0_col_out_1270   ),
    .col_1271                ( u0_col_out_1271   ),
    .col_1272                ( u0_col_out_1272   ),
    .col_1273                ( u0_col_out_1273   ),
    .col_1274                ( u0_col_out_1274   ),
    .col_1275                ( u0_col_out_1275   ),
    .col_1276                ( u0_col_out_1276   ),
    .col_1277                ( u0_col_out_1277   ),
    .col_1278                ( u0_col_out_1278   ),
    .col_1279                ( u0_col_out_1279   )
);





wire [1023:0] u1_ms;

alu  u1_alu (
    .clk                     ( clk                   ),
    .rst                     ( {rst  | reg_clear_i}  ),
    .col_in_0                ( u0_col_out_0     [127:0]  ),
    .col_in_1                ( u0_col_out_1     [127:0]  ),
    .col_in_2                ( u0_col_out_2     [127:0]  ),
    .col_in_3                ( u0_col_out_3     [127:0]  ),
    .col_in_4                ( u0_col_out_4     [127:0]  ),
    .col_in_5                ( u0_col_out_5     [127:0]  ),
    .col_in_6                ( u0_col_out_6     [127:0]  ),
    .col_in_7                ( u0_col_out_7     [127:0]  ),
    .col_in_8                ( u0_col_out_8     [127:0]  ),
    .col_in_9                ( u0_col_out_9     [127:0]  ),
    .col_in_10               ( u0_col_out_10    [127:0]  ),
    .col_in_11               ( u0_col_out_11    [127:0]  ),
    .col_in_12               ( u0_col_out_12    [127:0]  ),
    .col_in_13               ( u0_col_out_13    [127:0]  ),
    .col_in_14               ( u0_col_out_14    [127:0]  ),
    .col_in_15               ( u0_col_out_15    [127:0]  ),
    .col_in_16               ( u0_col_out_16    [127:0]  ),
    .col_in_17               ( u0_col_out_17    [127:0]  ),
    .col_in_18               ( u0_col_out_18    [127:0]  ),
    .col_in_19               ( u0_col_out_19    [127:0]  ),
    .col_in_20               ( u0_col_out_20    [127:0]  ),
    .col_in_21               ( u0_col_out_21    [127:0]  ),
    .col_in_22               ( u0_col_out_22    [127:0]  ),
    .col_in_23               ( u0_col_out_23    [127:0]  ),
    .col_in_24               ( u0_col_out_24    [127:0]  ),
    .col_in_25               ( u0_col_out_25    [127:0]  ),
    .col_in_26               ( u0_col_out_26    [127:0]  ),
    .col_in_27               ( u0_col_out_27    [127:0]  ),
    .col_in_28               ( u0_col_out_28    [127:0]  ),
    .col_in_29               ( u0_col_out_29    [127:0]  ),
    .col_in_30               ( u0_col_out_30    [127:0]  ),
    .col_in_31               ( u0_col_out_31    [127:0]  ),
    .col_in_32               ( u0_col_out_32    [127:0]  ),
    .col_in_33               ( u0_col_out_33    [127:0]  ),
    .col_in_34               ( u0_col_out_34    [127:0]  ),
    .col_in_35               ( u0_col_out_35    [127:0]  ),
    .col_in_36               ( u0_col_out_36    [127:0]  ),
    .col_in_37               ( u0_col_out_37    [127:0]  ),
    .col_in_38               ( u0_col_out_38    [127:0]  ),
    .col_in_39               ( u0_col_out_39    [127:0]  ),
    .col_in_40               ( u0_col_out_40    [127:0]  ),
    .col_in_41               ( u0_col_out_41    [127:0]  ),
    .col_in_42               ( u0_col_out_42    [127:0]  ),
    .col_in_43               ( u0_col_out_43    [127:0]  ),
    .col_in_44               ( u0_col_out_44    [127:0]  ),
    .col_in_45               ( u0_col_out_45    [127:0]  ),
    .col_in_46               ( u0_col_out_46    [127:0]  ),
    .col_in_47               ( u0_col_out_47    [127:0]  ),
    .col_in_48               ( u0_col_out_48    [127:0]  ),
    .col_in_49               ( u0_col_out_49    [127:0]  ),
    .col_in_50               ( u0_col_out_50    [127:0]  ),
    .col_in_51               ( u0_col_out_51    [127:0]  ),
    .col_in_52               ( u0_col_out_52    [127:0]  ),
    .col_in_53               ( u0_col_out_53    [127:0]  ),
    .col_in_54               ( u0_col_out_54    [127:0]  ),
    .col_in_55               ( u0_col_out_55    [127:0]  ),
    .col_in_56               ( u0_col_out_56    [127:0]  ),
    .col_in_57               ( u0_col_out_57    [127:0]  ),
    .col_in_58               ( u0_col_out_58    [127:0]  ),
    .col_in_59               ( u0_col_out_59    [127:0]  ),
    .col_in_60               ( u0_col_out_60    [127:0]  ),
    .col_in_61               ( u0_col_out_61    [127:0]  ),
    .col_in_62               ( u0_col_out_62    [127:0]  ),
    .col_in_63               ( u0_col_out_63    [127:0]  ),
    .col_in_64               ( u0_col_out_64    [127:0]  ),
    .col_in_65               ( u0_col_out_65    [127:0]  ),
    .col_in_66               ( u0_col_out_66    [127:0]  ),
    .col_in_67               ( u0_col_out_67    [127:0]  ),
    .col_in_68               ( u0_col_out_68    [127:0]  ),
    .col_in_69               ( u0_col_out_69    [127:0]  ),
    .col_in_70               ( u0_col_out_70    [127:0]  ),
    .col_in_71               ( u0_col_out_71    [127:0]  ),
    .col_in_72               ( u0_col_out_72    [127:0]  ),
    .col_in_73               ( u0_col_out_73    [127:0]  ),
    .col_in_74               ( u0_col_out_74    [127:0]  ),
    .col_in_75               ( u0_col_out_75    [127:0]  ),
    .col_in_76               ( u0_col_out_76    [127:0]  ),
    .col_in_77               ( u0_col_out_77    [127:0]  ),
    .col_in_78               ( u0_col_out_78    [127:0]  ),
    .col_in_79               ( u0_col_out_79    [127:0]  ),
    .col_in_80               ( u0_col_out_80    [127:0]  ),
    .col_in_81               ( u0_col_out_81    [127:0]  ),
    .col_in_82               ( u0_col_out_82    [127:0]  ),
    .col_in_83               ( u0_col_out_83    [127:0]  ),
    .col_in_84               ( u0_col_out_84    [127:0]  ),
    .col_in_85               ( u0_col_out_85    [127:0]  ),
    .col_in_86               ( u0_col_out_86    [127:0]  ),
    .col_in_87               ( u0_col_out_87    [127:0]  ),
    .col_in_88               ( u0_col_out_88    [127:0]  ),
    .col_in_89               ( u0_col_out_89    [127:0]  ),
    .col_in_90               ( u0_col_out_90    [127:0]  ),
    .col_in_91               ( u0_col_out_91    [127:0]  ),
    .col_in_92               ( u0_col_out_92    [127:0]  ),
    .col_in_93               ( u0_col_out_93    [127:0]  ),
    .col_in_94               ( u0_col_out_94    [127:0]  ),
    .col_in_95               ( u0_col_out_95    [127:0]  ),
    .col_in_96               ( u0_col_out_96    [127:0]  ),
    .col_in_97               ( u0_col_out_97    [127:0]  ),
    .col_in_98               ( u0_col_out_98    [127:0]  ),
    .col_in_99               ( u0_col_out_99    [127:0]  ),
    .col_in_100              ( u0_col_out_100   [127:0]  ),
    .col_in_101              ( u0_col_out_101   [127:0]  ),
    .col_in_102              ( u0_col_out_102   [127:0]  ),
    .col_in_103              ( u0_col_out_103   [127:0]  ),
    .col_in_104              ( u0_col_out_104   [127:0]  ),
    .col_in_105              ( u0_col_out_105   [127:0]  ),
    .col_in_106              ( u0_col_out_106   [127:0]  ),
    .col_in_107              ( u0_col_out_107   [127:0]  ),
    .col_in_108              ( u0_col_out_108   [127:0]  ),
    .col_in_109              ( u0_col_out_109   [127:0]  ),
    .col_in_110              ( u0_col_out_110   [127:0]  ),
    .col_in_111              ( u0_col_out_111   [127:0]  ),
    .col_in_112              ( u0_col_out_112   [127:0]  ),
    .col_in_113              ( u0_col_out_113   [127:0]  ),
    .col_in_114              ( u0_col_out_114   [127:0]  ),
    .col_in_115              ( u0_col_out_115   [127:0]  ),
    .col_in_116              ( u0_col_out_116   [127:0]  ),
    .col_in_117              ( u0_col_out_117   [127:0]  ),
    .col_in_118              ( u0_col_out_118   [127:0]  ),
    .col_in_119              ( u0_col_out_119   [127:0]  ),
    .col_in_120              ( u0_col_out_120   [127:0]  ),
    .col_in_121              ( u0_col_out_121   [127:0]  ),
    .col_in_122              ( u0_col_out_122   [127:0]  ),
    .col_in_123              ( u0_col_out_123   [127:0]  ),
    .col_in_124              ( u0_col_out_124   [127:0]  ),
    .col_in_125              ( u0_col_out_125   [127:0]  ),
    .col_in_126              ( u0_col_out_126   [127:0]  ),
    .col_in_127              ( u0_col_out_127   [127:0]  ),
    .col_in_128              ( u0_col_out_128   [127:0]  ),
    .col_in_129              ( u0_col_out_129   [127:0]  ),
    .col_in_130              ( u0_col_out_130   [127:0]  ),
    .col_in_131              ( u0_col_out_131   [127:0]  ),
    .col_in_132              ( u0_col_out_132   [127:0]  ),
    .col_in_133              ( u0_col_out_133   [127:0]  ),
    .col_in_134              ( u0_col_out_134   [127:0]  ),
    .col_in_135              ( u0_col_out_135   [127:0]  ),
    .col_in_136              ( u0_col_out_136   [127:0]  ),
    .col_in_137              ( u0_col_out_137   [127:0]  ),
    .col_in_138              ( u0_col_out_138   [127:0]  ),
    .col_in_139              ( u0_col_out_139   [127:0]  ),
    .col_in_140              ( u0_col_out_140   [127:0]  ),
    .col_in_141              ( u0_col_out_141   [127:0]  ),
    .col_in_142              ( u0_col_out_142   [127:0]  ),
    .col_in_143              ( u0_col_out_143   [127:0]  ),
    .col_in_144              ( u0_col_out_144   [127:0]  ),
    .col_in_145              ( u0_col_out_145   [127:0]  ),
    .col_in_146              ( u0_col_out_146   [127:0]  ),
    .col_in_147              ( u0_col_out_147   [127:0]  ),
    .col_in_148              ( u0_col_out_148   [127:0]  ),
    .col_in_149              ( u0_col_out_149   [127:0]  ),
    .col_in_150              ( u0_col_out_150   [127:0]  ),
    .col_in_151              ( u0_col_out_151   [127:0]  ),
    .col_in_152              ( u0_col_out_152   [127:0]  ),
    .col_in_153              ( u0_col_out_153   [127:0]  ),
    .col_in_154              ( u0_col_out_154   [127:0]  ),
    .col_in_155              ( u0_col_out_155   [127:0]  ),
    .col_in_156              ( u0_col_out_156   [127:0]  ),
    .col_in_157              ( u0_col_out_157   [127:0]  ),
    .col_in_158              ( u0_col_out_158   [127:0]  ),
    .col_in_159              ( u0_col_out_159   [127:0]  ),
    .col_in_160              ( u0_col_out_160   [127:0]  ),
    .col_in_161              ( u0_col_out_161   [127:0]  ),
    .col_in_162              ( u0_col_out_162   [127:0]  ),
    .col_in_163              ( u0_col_out_163   [127:0]  ),
    .col_in_164              ( u0_col_out_164   [127:0]  ),
    .col_in_165              ( u0_col_out_165   [127:0]  ),
    .col_in_166              ( u0_col_out_166   [127:0]  ),
    .col_in_167              ( u0_col_out_167   [127:0]  ),
    .col_in_168              ( u0_col_out_168   [127:0]  ),
    .col_in_169              ( u0_col_out_169   [127:0]  ),
    .col_in_170              ( u0_col_out_170   [127:0]  ),
    .col_in_171              ( u0_col_out_171   [127:0]  ),
    .col_in_172              ( u0_col_out_172   [127:0]  ),
    .col_in_173              ( u0_col_out_173   [127:0]  ),
    .col_in_174              ( u0_col_out_174   [127:0]  ),
    .col_in_175              ( u0_col_out_175   [127:0]  ),
    .col_in_176              ( u0_col_out_176   [127:0]  ),
    .col_in_177              ( u0_col_out_177   [127:0]  ),
    .col_in_178              ( u0_col_out_178   [127:0]  ),
    .col_in_179              ( u0_col_out_179   [127:0]  ),
    .col_in_180              ( u0_col_out_180   [127:0]  ),
    .col_in_181              ( u0_col_out_181   [127:0]  ),
    .col_in_182              ( u0_col_out_182   [127:0]  ),
    .col_in_183              ( u0_col_out_183   [127:0]  ),
    .col_in_184              ( u0_col_out_184   [127:0]  ),
    .col_in_185              ( u0_col_out_185   [127:0]  ),
    .col_in_186              ( u0_col_out_186   [127:0]  ),
    .col_in_187              ( u0_col_out_187   [127:0]  ),
    .col_in_188              ( u0_col_out_188   [127:0]  ),
    .col_in_189              ( u0_col_out_189   [127:0]  ),
    .col_in_190              ( u0_col_out_190   [127:0]  ),
    .col_in_191              ( u0_col_out_191   [127:0]  ),
    .col_in_192              ( u0_col_out_192   [127:0]  ),
    .col_in_193              ( u0_col_out_193   [127:0]  ),
    .col_in_194              ( u0_col_out_194   [127:0]  ),
    .col_in_195              ( u0_col_out_195   [127:0]  ),
    .col_in_196              ( u0_col_out_196   [127:0]  ),
    .col_in_197              ( u0_col_out_197   [127:0]  ),
    .col_in_198              ( u0_col_out_198   [127:0]  ),
    .col_in_199              ( u0_col_out_199   [127:0]  ),
    .col_in_200              ( u0_col_out_200   [127:0]  ),
    .col_in_201              ( u0_col_out_201   [127:0]  ),
    .col_in_202              ( u0_col_out_202   [127:0]  ),
    .col_in_203              ( u0_col_out_203   [127:0]  ),
    .col_in_204              ( u0_col_out_204   [127:0]  ),
    .col_in_205              ( u0_col_out_205   [127:0]  ),
    .col_in_206              ( u0_col_out_206   [127:0]  ),
    .col_in_207              ( u0_col_out_207   [127:0]  ),
    .col_in_208              ( u0_col_out_208   [127:0]  ),
    .col_in_209              ( u0_col_out_209   [127:0]  ),
    .col_in_210              ( u0_col_out_210   [127:0]  ),
    .col_in_211              ( u0_col_out_211   [127:0]  ),
    .col_in_212              ( u0_col_out_212   [127:0]  ),
    .col_in_213              ( u0_col_out_213   [127:0]  ),
    .col_in_214              ( u0_col_out_214   [127:0]  ),
    .col_in_215              ( u0_col_out_215   [127:0]  ),
    .col_in_216              ( u0_col_out_216   [127:0]  ),
    .col_in_217              ( u0_col_out_217   [127:0]  ),
    .col_in_218              ( u0_col_out_218   [127:0]  ),
    .col_in_219              ( u0_col_out_219   [127:0]  ),
    .col_in_220              ( u0_col_out_220   [127:0]  ),
    .col_in_221              ( u0_col_out_221   [127:0]  ),
    .col_in_222              ( u0_col_out_222   [127:0]  ),
    .col_in_223              ( u0_col_out_223   [127:0]  ),
    .col_in_224              ( u0_col_out_224   [127:0]  ),
    .col_in_225              ( u0_col_out_225   [127:0]  ),
    .col_in_226              ( u0_col_out_226   [127:0]  ),
    .col_in_227              ( u0_col_out_227   [127:0]  ),
    .col_in_228              ( u0_col_out_228   [127:0]  ),
    .col_in_229              ( u0_col_out_229   [127:0]  ),
    .col_in_230              ( u0_col_out_230   [127:0]  ),
    .col_in_231              ( u0_col_out_231   [127:0]  ),
    .col_in_232              ( u0_col_out_232   [127:0]  ),
    .col_in_233              ( u0_col_out_233   [127:0]  ),
    .col_in_234              ( u0_col_out_234   [127:0]  ),
    .col_in_235              ( u0_col_out_235   [127:0]  ),
    .col_in_236              ( u0_col_out_236   [127:0]  ),
    .col_in_237              ( u0_col_out_237   [127:0]  ),
    .col_in_238              ( u0_col_out_238   [127:0]  ),
    .col_in_239              ( u0_col_out_239   [127:0]  ),
    .col_in_240              ( u0_col_out_240   [127:0]  ),
    .col_in_241              ( u0_col_out_241   [127:0]  ),
    .col_in_242              ( u0_col_out_242   [127:0]  ),
    .col_in_243              ( u0_col_out_243   [127:0]  ),
    .col_in_244              ( u0_col_out_244   [127:0]  ),
    .col_in_245              ( u0_col_out_245   [127:0]  ),
    .col_in_246              ( u0_col_out_246   [127:0]  ),
    .col_in_247              ( u0_col_out_247   [127:0]  ),
    .col_in_248              ( u0_col_out_248   [127:0]  ),
    .col_in_249              ( u0_col_out_249   [127:0]  ),
    .col_in_250              ( u0_col_out_250   [127:0]  ),
    .col_in_251              ( u0_col_out_251   [127:0]  ),
    .col_in_252              ( u0_col_out_252   [127:0]  ),
    .col_in_253              ( u0_col_out_253   [127:0]  ),
    .col_in_254              ( u0_col_out_254   [127:0]  ),
    .col_in_255              ( u0_col_out_255   [127:0]  ),
    .col_in_256              ( u0_col_out_256   [127:0]  ),
    .col_in_257              ( u0_col_out_257   [127:0]  ),
    .col_in_258              ( u0_col_out_258   [127:0]  ),
    .col_in_259              ( u0_col_out_259   [127:0]  ),
    .col_in_260              ( u0_col_out_260   [127:0]  ),
    .col_in_261              ( u0_col_out_261   [127:0]  ),
    .col_in_262              ( u0_col_out_262   [127:0]  ),
    .col_in_263              ( u0_col_out_263   [127:0]  ),
    .col_in_264              ( u0_col_out_264   [127:0]  ),
    .col_in_265              ( u0_col_out_265   [127:0]  ),
    .col_in_266              ( u0_col_out_266   [127:0]  ),
    .col_in_267              ( u0_col_out_267   [127:0]  ),
    .col_in_268              ( u0_col_out_268   [127:0]  ),
    .col_in_269              ( u0_col_out_269   [127:0]  ),
    .col_in_270              ( u0_col_out_270   [127:0]  ),
    .col_in_271              ( u0_col_out_271   [127:0]  ),
    .col_in_272              ( u0_col_out_272   [127:0]  ),
    .col_in_273              ( u0_col_out_273   [127:0]  ),
    .col_in_274              ( u0_col_out_274   [127:0]  ),
    .col_in_275              ( u0_col_out_275   [127:0]  ),
    .col_in_276              ( u0_col_out_276   [127:0]  ),
    .col_in_277              ( u0_col_out_277   [127:0]  ),
    .col_in_278              ( u0_col_out_278   [127:0]  ),
    .col_in_279              ( u0_col_out_279   [127:0]  ),
    .col_in_280              ( u0_col_out_280   [127:0]  ),
    .col_in_281              ( u0_col_out_281   [127:0]  ),
    .col_in_282              ( u0_col_out_282   [127:0]  ),
    .col_in_283              ( u0_col_out_283   [127:0]  ),
    .col_in_284              ( u0_col_out_284   [127:0]  ),
    .col_in_285              ( u0_col_out_285   [127:0]  ),
    .col_in_286              ( u0_col_out_286   [127:0]  ),
    .col_in_287              ( u0_col_out_287   [127:0]  ),
    .col_in_288              ( u0_col_out_288   [127:0]  ),
    .col_in_289              ( u0_col_out_289   [127:0]  ),
    .col_in_290              ( u0_col_out_290   [127:0]  ),
    .col_in_291              ( u0_col_out_291   [127:0]  ),
    .col_in_292              ( u0_col_out_292   [127:0]  ),
    .col_in_293              ( u0_col_out_293   [127:0]  ),
    .col_in_294              ( u0_col_out_294   [127:0]  ),
    .col_in_295              ( u0_col_out_295   [127:0]  ),
    .col_in_296              ( u0_col_out_296   [127:0]  ),
    .col_in_297              ( u0_col_out_297   [127:0]  ),
    .col_in_298              ( u0_col_out_298   [127:0]  ),
    .col_in_299              ( u0_col_out_299   [127:0]  ),
    .col_in_300              ( u0_col_out_300   [127:0]  ),
    .col_in_301              ( u0_col_out_301   [127:0]  ),
    .col_in_302              ( u0_col_out_302   [127:0]  ),
    .col_in_303              ( u0_col_out_303   [127:0]  ),
    .col_in_304              ( u0_col_out_304   [127:0]  ),
    .col_in_305              ( u0_col_out_305   [127:0]  ),
    .col_in_306              ( u0_col_out_306   [127:0]  ),
    .col_in_307              ( u0_col_out_307   [127:0]  ),
    .col_in_308              ( u0_col_out_308   [127:0]  ),
    .col_in_309              ( u0_col_out_309   [127:0]  ),
    .col_in_310              ( u0_col_out_310   [127:0]  ),
    .col_in_311              ( u0_col_out_311   [127:0]  ),
    .col_in_312              ( u0_col_out_312   [127:0]  ),
    .col_in_313              ( u0_col_out_313   [127:0]  ),
    .col_in_314              ( u0_col_out_314   [127:0]  ),
    .col_in_315              ( u0_col_out_315   [127:0]  ),
    .col_in_316              ( u0_col_out_316   [127:0]  ),
    .col_in_317              ( u0_col_out_317   [127:0]  ),
    .col_in_318              ( u0_col_out_318   [127:0]  ),
    .col_in_319              ( u0_col_out_319   [127:0]  ),
    .col_in_320              ( u0_col_out_320   [127:0]  ),
    .col_in_321              ( u0_col_out_321   [127:0]  ),
    .col_in_322              ( u0_col_out_322   [127:0]  ),
    .col_in_323              ( u0_col_out_323   [127:0]  ),
    .col_in_324              ( u0_col_out_324   [127:0]  ),
    .col_in_325              ( u0_col_out_325   [127:0]  ),
    .col_in_326              ( u0_col_out_326   [127:0]  ),
    .col_in_327              ( u0_col_out_327   [127:0]  ),
    .col_in_328              ( u0_col_out_328   [127:0]  ),
    .col_in_329              ( u0_col_out_329   [127:0]  ),
    .col_in_330              ( u0_col_out_330   [127:0]  ),
    .col_in_331              ( u0_col_out_331   [127:0]  ),
    .col_in_332              ( u0_col_out_332   [127:0]  ),
    .col_in_333              ( u0_col_out_333   [127:0]  ),
    .col_in_334              ( u0_col_out_334   [127:0]  ),
    .col_in_335              ( u0_col_out_335   [127:0]  ),
    .col_in_336              ( u0_col_out_336   [127:0]  ),
    .col_in_337              ( u0_col_out_337   [127:0]  ),
    .col_in_338              ( u0_col_out_338   [127:0]  ),
    .col_in_339              ( u0_col_out_339   [127:0]  ),
    .col_in_340              ( u0_col_out_340   [127:0]  ),
    .col_in_341              ( u0_col_out_341   [127:0]  ),
    .col_in_342              ( u0_col_out_342   [127:0]  ),
    .col_in_343              ( u0_col_out_343   [127:0]  ),
    .col_in_344              ( u0_col_out_344   [127:0]  ),
    .col_in_345              ( u0_col_out_345   [127:0]  ),
    .col_in_346              ( u0_col_out_346   [127:0]  ),
    .col_in_347              ( u0_col_out_347   [127:0]  ),
    .col_in_348              ( u0_col_out_348   [127:0]  ),
    .col_in_349              ( u0_col_out_349   [127:0]  ),
    .col_in_350              ( u0_col_out_350   [127:0]  ),
    .col_in_351              ( u0_col_out_351   [127:0]  ),
    .col_in_352              ( u0_col_out_352   [127:0]  ),
    .col_in_353              ( u0_col_out_353   [127:0]  ),
    .col_in_354              ( u0_col_out_354   [127:0]  ),
    .col_in_355              ( u0_col_out_355   [127:0]  ),
    .col_in_356              ( u0_col_out_356   [127:0]  ),
    .col_in_357              ( u0_col_out_357   [127:0]  ),
    .col_in_358              ( u0_col_out_358   [127:0]  ),
    .col_in_359              ( u0_col_out_359   [127:0]  ),
    .col_in_360              ( u0_col_out_360   [127:0]  ),
    .col_in_361              ( u0_col_out_361   [127:0]  ),
    .col_in_362              ( u0_col_out_362   [127:0]  ),
    .col_in_363              ( u0_col_out_363   [127:0]  ),
    .col_in_364              ( u0_col_out_364   [127:0]  ),
    .col_in_365              ( u0_col_out_365   [127:0]  ),
    .col_in_366              ( u0_col_out_366   [127:0]  ),
    .col_in_367              ( u0_col_out_367   [127:0]  ),
    .col_in_368              ( u0_col_out_368   [127:0]  ),
    .col_in_369              ( u0_col_out_369   [127:0]  ),
    .col_in_370              ( u0_col_out_370   [127:0]  ),
    .col_in_371              ( u0_col_out_371   [127:0]  ),
    .col_in_372              ( u0_col_out_372   [127:0]  ),
    .col_in_373              ( u0_col_out_373   [127:0]  ),
    .col_in_374              ( u0_col_out_374   [127:0]  ),
    .col_in_375              ( u0_col_out_375   [127:0]  ),
    .col_in_376              ( u0_col_out_376   [127:0]  ),
    .col_in_377              ( u0_col_out_377   [127:0]  ),
    .col_in_378              ( u0_col_out_378   [127:0]  ),
    .col_in_379              ( u0_col_out_379   [127:0]  ),
    .col_in_380              ( u0_col_out_380   [127:0]  ),
    .col_in_381              ( u0_col_out_381   [127:0]  ),
    .col_in_382              ( u0_col_out_382   [127:0]  ),
    .col_in_383              ( u0_col_out_383   [127:0]  ),
    .col_in_384              ( u0_col_out_384   [127:0]  ),
    .col_in_385              ( u0_col_out_385   [127:0]  ),
    .col_in_386              ( u0_col_out_386   [127:0]  ),
    .col_in_387              ( u0_col_out_387   [127:0]  ),
    .col_in_388              ( u0_col_out_388   [127:0]  ),
    .col_in_389              ( u0_col_out_389   [127:0]  ),
    .col_in_390              ( u0_col_out_390   [127:0]  ),
    .col_in_391              ( u0_col_out_391   [127:0]  ),
    .col_in_392              ( u0_col_out_392   [127:0]  ),
    .col_in_393              ( u0_col_out_393   [127:0]  ),
    .col_in_394              ( u0_col_out_394   [127:0]  ),
    .col_in_395              ( u0_col_out_395   [127:0]  ),
    .col_in_396              ( u0_col_out_396   [127:0]  ),
    .col_in_397              ( u0_col_out_397   [127:0]  ),
    .col_in_398              ( u0_col_out_398   [127:0]  ),
    .col_in_399              ( u0_col_out_399   [127:0]  ),
    .col_in_400              ( u0_col_out_400   [127:0]  ),
    .col_in_401              ( u0_col_out_401   [127:0]  ),
    .col_in_402              ( u0_col_out_402   [127:0]  ),
    .col_in_403              ( u0_col_out_403   [127:0]  ),
    .col_in_404              ( u0_col_out_404   [127:0]  ),
    .col_in_405              ( u0_col_out_405   [127:0]  ),
    .col_in_406              ( u0_col_out_406   [127:0]  ),
    .col_in_407              ( u0_col_out_407   [127:0]  ),
    .col_in_408              ( u0_col_out_408   [127:0]  ),
    .col_in_409              ( u0_col_out_409   [127:0]  ),
    .col_in_410              ( u0_col_out_410   [127:0]  ),
    .col_in_411              ( u0_col_out_411   [127:0]  ),
    .col_in_412              ( u0_col_out_412   [127:0]  ),
    .col_in_413              ( u0_col_out_413   [127:0]  ),
    .col_in_414              ( u0_col_out_414   [127:0]  ),
    .col_in_415              ( u0_col_out_415   [127:0]  ),
    .col_in_416              ( u0_col_out_416   [127:0]  ),
    .col_in_417              ( u0_col_out_417   [127:0]  ),
    .col_in_418              ( u0_col_out_418   [127:0]  ),
    .col_in_419              ( u0_col_out_419   [127:0]  ),
    .col_in_420              ( u0_col_out_420   [127:0]  ),
    .col_in_421              ( u0_col_out_421   [127:0]  ),
    .col_in_422              ( u0_col_out_422   [127:0]  ),
    .col_in_423              ( u0_col_out_423   [127:0]  ),
    .col_in_424              ( u0_col_out_424   [127:0]  ),
    .col_in_425              ( u0_col_out_425   [127:0]  ),
    .col_in_426              ( u0_col_out_426   [127:0]  ),
    .col_in_427              ( u0_col_out_427   [127:0]  ),
    .col_in_428              ( u0_col_out_428   [127:0]  ),
    .col_in_429              ( u0_col_out_429   [127:0]  ),
    .col_in_430              ( u0_col_out_430   [127:0]  ),
    .col_in_431              ( u0_col_out_431   [127:0]  ),
    .col_in_432              ( u0_col_out_432   [127:0]  ),
    .col_in_433              ( u0_col_out_433   [127:0]  ),
    .col_in_434              ( u0_col_out_434   [127:0]  ),
    .col_in_435              ( u0_col_out_435   [127:0]  ),
    .col_in_436              ( u0_col_out_436   [127:0]  ),
    .col_in_437              ( u0_col_out_437   [127:0]  ),
    .col_in_438              ( u0_col_out_438   [127:0]  ),
    .col_in_439              ( u0_col_out_439   [127:0]  ),
    .col_in_440              ( u0_col_out_440   [127:0]  ),
    .col_in_441              ( u0_col_out_441   [127:0]  ),
    .col_in_442              ( u0_col_out_442   [127:0]  ),
    .col_in_443              ( u0_col_out_443   [127:0]  ),
    .col_in_444              ( u0_col_out_444   [127:0]  ),
    .col_in_445              ( u0_col_out_445   [127:0]  ),
    .col_in_446              ( u0_col_out_446   [127:0]  ),
    .col_in_447              ( u0_col_out_447   [127:0]  ),
    .col_in_448              ( u0_col_out_448   [127:0]  ),
    .col_in_449              ( u0_col_out_449   [127:0]  ),
    .col_in_450              ( u0_col_out_450   [127:0]  ),
    .col_in_451              ( u0_col_out_451   [127:0]  ),
    .col_in_452              ( u0_col_out_452   [127:0]  ),
    .col_in_453              ( u0_col_out_453   [127:0]  ),
    .col_in_454              ( u0_col_out_454   [127:0]  ),
    .col_in_455              ( u0_col_out_455   [127:0]  ),
    .col_in_456              ( u0_col_out_456   [127:0]  ),
    .col_in_457              ( u0_col_out_457   [127:0]  ),
    .col_in_458              ( u0_col_out_458   [127:0]  ),
    .col_in_459              ( u0_col_out_459   [127:0]  ),
    .col_in_460              ( u0_col_out_460   [127:0]  ),
    .col_in_461              ( u0_col_out_461   [127:0]  ),
    .col_in_462              ( u0_col_out_462   [127:0]  ),
    .col_in_463              ( u0_col_out_463   [127:0]  ),
    .col_in_464              ( u0_col_out_464   [127:0]  ),
    .col_in_465              ( u0_col_out_465   [127:0]  ),
    .col_in_466              ( u0_col_out_466   [127:0]  ),
    .col_in_467              ( u0_col_out_467   [127:0]  ),
    .col_in_468              ( u0_col_out_468   [127:0]  ),
    .col_in_469              ( u0_col_out_469   [127:0]  ),
    .col_in_470              ( u0_col_out_470   [127:0]  ),
    .col_in_471              ( u0_col_out_471   [127:0]  ),
    .col_in_472              ( u0_col_out_472   [127:0]  ),
    .col_in_473              ( u0_col_out_473   [127:0]  ),
    .col_in_474              ( u0_col_out_474   [127:0]  ),
    .col_in_475              ( u0_col_out_475   [127:0]  ),
    .col_in_476              ( u0_col_out_476   [127:0]  ),
    .col_in_477              ( u0_col_out_477   [127:0]  ),
    .col_in_478              ( u0_col_out_478   [127:0]  ),
    .col_in_479              ( u0_col_out_479   [127:0]  ),
    .col_in_480              ( u0_col_out_480   [127:0]  ),
    .col_in_481              ( u0_col_out_481   [127:0]  ),
    .col_in_482              ( u0_col_out_482   [127:0]  ),
    .col_in_483              ( u0_col_out_483   [127:0]  ),
    .col_in_484              ( u0_col_out_484   [127:0]  ),
    .col_in_485              ( u0_col_out_485   [127:0]  ),
    .col_in_486              ( u0_col_out_486   [127:0]  ),
    .col_in_487              ( u0_col_out_487   [127:0]  ),
    .col_in_488              ( u0_col_out_488   [127:0]  ),
    .col_in_489              ( u0_col_out_489   [127:0]  ),
    .col_in_490              ( u0_col_out_490   [127:0]  ),
    .col_in_491              ( u0_col_out_491   [127:0]  ),
    .col_in_492              ( u0_col_out_492   [127:0]  ),
    .col_in_493              ( u0_col_out_493   [127:0]  ),
    .col_in_494              ( u0_col_out_494   [127:0]  ),
    .col_in_495              ( u0_col_out_495   [127:0]  ),
    .col_in_496              ( u0_col_out_496   [127:0]  ),
    .col_in_497              ( u0_col_out_497   [127:0]  ),
    .col_in_498              ( u0_col_out_498   [127:0]  ),
    .col_in_499              ( u0_col_out_499   [127:0]  ),
    .col_in_500              ( u0_col_out_500   [127:0]  ),
    .col_in_501              ( u0_col_out_501   [127:0]  ),
    .col_in_502              ( u0_col_out_502   [127:0]  ),
    .col_in_503              ( u0_col_out_503   [127:0]  ),
    .col_in_504              ( u0_col_out_504   [127:0]  ),
    .col_in_505              ( u0_col_out_505   [127:0]  ),
    .col_in_506              ( u0_col_out_506   [127:0]  ),
    .col_in_507              ( u0_col_out_507   [127:0]  ),
    .col_in_508              ( u0_col_out_508   [127:0]  ),
    .col_in_509              ( u0_col_out_509   [127:0]  ),
    .col_in_510              ( u0_col_out_510   [127:0]  ),
    .col_in_511              ( u0_col_out_511   [127:0]  ),
    .col_in_512              ( u0_col_out_512   [127:0]  ),
    .col_in_513              ( u0_col_out_513   [127:0]  ),
    .col_in_514              ( u0_col_out_514   [127:0]  ),
    .col_in_515              ( u0_col_out_515   [127:0]  ),
    .col_in_516              ( u0_col_out_516   [127:0]  ),
    .col_in_517              ( u0_col_out_517   [127:0]  ),
    .col_in_518              ( u0_col_out_518   [127:0]  ),
    .col_in_519              ( u0_col_out_519   [127:0]  ),
    .col_in_520              ( u0_col_out_520   [127:0]  ),
    .col_in_521              ( u0_col_out_521   [127:0]  ),
    .col_in_522              ( u0_col_out_522   [127:0]  ),
    .col_in_523              ( u0_col_out_523   [127:0]  ),
    .col_in_524              ( u0_col_out_524   [127:0]  ),
    .col_in_525              ( u0_col_out_525   [127:0]  ),
    .col_in_526              ( u0_col_out_526   [127:0]  ),
    .col_in_527              ( u0_col_out_527   [127:0]  ),
    .col_in_528              ( u0_col_out_528   [127:0]  ),
    .col_in_529              ( u0_col_out_529   [127:0]  ),
    .col_in_530              ( u0_col_out_530   [127:0]  ),
    .col_in_531              ( u0_col_out_531   [127:0]  ),
    .col_in_532              ( u0_col_out_532   [127:0]  ),
    .col_in_533              ( u0_col_out_533   [127:0]  ),
    .col_in_534              ( u0_col_out_534   [127:0]  ),
    .col_in_535              ( u0_col_out_535   [127:0]  ),
    .col_in_536              ( u0_col_out_536   [127:0]  ),
    .col_in_537              ( u0_col_out_537   [127:0]  ),
    .col_in_538              ( u0_col_out_538   [127:0]  ),
    .col_in_539              ( u0_col_out_539   [127:0]  ),
    .col_in_540              ( u0_col_out_540   [127:0]  ),
    .col_in_541              ( u0_col_out_541   [127:0]  ),
    .col_in_542              ( u0_col_out_542   [127:0]  ),
    .col_in_543              ( u0_col_out_543   [127:0]  ),
    .col_in_544              ( u0_col_out_544   [127:0]  ),
    .col_in_545              ( u0_col_out_545   [127:0]  ),
    .col_in_546              ( u0_col_out_546   [127:0]  ),
    .col_in_547              ( u0_col_out_547   [127:0]  ),
    .col_in_548              ( u0_col_out_548   [127:0]  ),
    .col_in_549              ( u0_col_out_549   [127:0]  ),
    .col_in_550              ( u0_col_out_550   [127:0]  ),
    .col_in_551              ( u0_col_out_551   [127:0]  ),
    .col_in_552              ( u0_col_out_552   [127:0]  ),
    .col_in_553              ( u0_col_out_553   [127:0]  ),
    .col_in_554              ( u0_col_out_554   [127:0]  ),
    .col_in_555              ( u0_col_out_555   [127:0]  ),
    .col_in_556              ( u0_col_out_556   [127:0]  ),
    .col_in_557              ( u0_col_out_557   [127:0]  ),
    .col_in_558              ( u0_col_out_558   [127:0]  ),
    .col_in_559              ( u0_col_out_559   [127:0]  ),
    .col_in_560              ( u0_col_out_560   [127:0]  ),
    .col_in_561              ( u0_col_out_561   [127:0]  ),
    .col_in_562              ( u0_col_out_562   [127:0]  ),
    .col_in_563              ( u0_col_out_563   [127:0]  ),
    .col_in_564              ( u0_col_out_564   [127:0]  ),
    .col_in_565              ( u0_col_out_565   [127:0]  ),
    .col_in_566              ( u0_col_out_566   [127:0]  ),
    .col_in_567              ( u0_col_out_567   [127:0]  ),
    .col_in_568              ( u0_col_out_568   [127:0]  ),
    .col_in_569              ( u0_col_out_569   [127:0]  ),
    .col_in_570              ( u0_col_out_570   [127:0]  ),
    .col_in_571              ( u0_col_out_571   [127:0]  ),
    .col_in_572              ( u0_col_out_572   [127:0]  ),
    .col_in_573              ( u0_col_out_573   [127:0]  ),
    .col_in_574              ( u0_col_out_574   [127:0]  ),
    .col_in_575              ( u0_col_out_575   [127:0]  ),
    .col_in_576              ( u0_col_out_576   [127:0]  ),
    .col_in_577              ( u0_col_out_577   [127:0]  ),
    .col_in_578              ( u0_col_out_578   [127:0]  ),
    .col_in_579              ( u0_col_out_579   [127:0]  ),
    .col_in_580              ( u0_col_out_580   [127:0]  ),
    .col_in_581              ( u0_col_out_581   [127:0]  ),
    .col_in_582              ( u0_col_out_582   [127:0]  ),
    .col_in_583              ( u0_col_out_583   [127:0]  ),
    .col_in_584              ( u0_col_out_584   [127:0]  ),
    .col_in_585              ( u0_col_out_585   [127:0]  ),
    .col_in_586              ( u0_col_out_586   [127:0]  ),
    .col_in_587              ( u0_col_out_587   [127:0]  ),
    .col_in_588              ( u0_col_out_588   [127:0]  ),
    .col_in_589              ( u0_col_out_589   [127:0]  ),
    .col_in_590              ( u0_col_out_590   [127:0]  ),
    .col_in_591              ( u0_col_out_591   [127:0]  ),
    .col_in_592              ( u0_col_out_592   [127:0]  ),
    .col_in_593              ( u0_col_out_593   [127:0]  ),
    .col_in_594              ( u0_col_out_594   [127:0]  ),
    .col_in_595              ( u0_col_out_595   [127:0]  ),
    .col_in_596              ( u0_col_out_596   [127:0]  ),
    .col_in_597              ( u0_col_out_597   [127:0]  ),
    .col_in_598              ( u0_col_out_598   [127:0]  ),
    .col_in_599              ( u0_col_out_599   [127:0]  ),
    .col_in_600              ( u0_col_out_600   [127:0]  ),
    .col_in_601              ( u0_col_out_601   [127:0]  ),
    .col_in_602              ( u0_col_out_602   [127:0]  ),
    .col_in_603              ( u0_col_out_603   [127:0]  ),
    .col_in_604              ( u0_col_out_604   [127:0]  ),
    .col_in_605              ( u0_col_out_605   [127:0]  ),
    .col_in_606              ( u0_col_out_606   [127:0]  ),
    .col_in_607              ( u0_col_out_607   [127:0]  ),
    .col_in_608              ( u0_col_out_608   [127:0]  ),
    .col_in_609              ( u0_col_out_609   [127:0]  ),
    .col_in_610              ( u0_col_out_610   [127:0]  ),
    .col_in_611              ( u0_col_out_611   [127:0]  ),
    .col_in_612              ( u0_col_out_612   [127:0]  ),
    .col_in_613              ( u0_col_out_613   [127:0]  ),
    .col_in_614              ( u0_col_out_614   [127:0]  ),
    .col_in_615              ( u0_col_out_615   [127:0]  ),
    .col_in_616              ( u0_col_out_616   [127:0]  ),
    .col_in_617              ( u0_col_out_617   [127:0]  ),
    .col_in_618              ( u0_col_out_618   [127:0]  ),
    .col_in_619              ( u0_col_out_619   [127:0]  ),
    .col_in_620              ( u0_col_out_620   [127:0]  ),
    .col_in_621              ( u0_col_out_621   [127:0]  ),
    .col_in_622              ( u0_col_out_622   [127:0]  ),
    .col_in_623              ( u0_col_out_623   [127:0]  ),
    .col_in_624              ( u0_col_out_624   [127:0]  ),
    .col_in_625              ( u0_col_out_625   [127:0]  ),
    .col_in_626              ( u0_col_out_626   [127:0]  ),
    .col_in_627              ( u0_col_out_627   [127:0]  ),
    .col_in_628              ( u0_col_out_628   [127:0]  ),
    .col_in_629              ( u0_col_out_629   [127:0]  ),
    .col_in_630              ( u0_col_out_630   [127:0]  ),
    .col_in_631              ( u0_col_out_631   [127:0]  ),
    .col_in_632              ( u0_col_out_632   [127:0]  ),
    .col_in_633              ( u0_col_out_633   [127:0]  ),
    .col_in_634              ( u0_col_out_634   [127:0]  ),
    .col_in_635              ( u0_col_out_635   [127:0]  ),
    .col_in_636              ( u0_col_out_636   [127:0]  ),
    .col_in_637              ( u0_col_out_637   [127:0]  ),
    .col_in_638              ( u0_col_out_638   [127:0]  ),
    .col_in_639              ( u0_col_out_639   [127:0]  ),
    .col_in_640              ( u0_col_out_640   [127:0]  ),
    .col_in_641              ( u0_col_out_641   [127:0]  ),
    .col_in_642              ( u0_col_out_642   [127:0]  ),
    .col_in_643              ( u0_col_out_643   [127:0]  ),
    .col_in_644              ( u0_col_out_644   [127:0]  ),
    .col_in_645              ( u0_col_out_645   [127:0]  ),
    .col_in_646              ( u0_col_out_646   [127:0]  ),
    .col_in_647              ( u0_col_out_647   [127:0]  ),
    .col_in_648              ( u0_col_out_648   [127:0]  ),
    .col_in_649              ( u0_col_out_649   [127:0]  ),
    .col_in_650              ( u0_col_out_650   [127:0]  ),
    .col_in_651              ( u0_col_out_651   [127:0]  ),
    .col_in_652              ( u0_col_out_652   [127:0]  ),
    .col_in_653              ( u0_col_out_653   [127:0]  ),
    .col_in_654              ( u0_col_out_654   [127:0]  ),
    .col_in_655              ( u0_col_out_655   [127:0]  ),
    .col_in_656              ( u0_col_out_656   [127:0]  ),
    .col_in_657              ( u0_col_out_657   [127:0]  ),
    .col_in_658              ( u0_col_out_658   [127:0]  ),
    .col_in_659              ( u0_col_out_659   [127:0]  ),
    .col_in_660              ( u0_col_out_660   [127:0]  ),
    .col_in_661              ( u0_col_out_661   [127:0]  ),
    .col_in_662              ( u0_col_out_662   [127:0]  ),
    .col_in_663              ( u0_col_out_663   [127:0]  ),
    .col_in_664              ( u0_col_out_664   [127:0]  ),
    .col_in_665              ( u0_col_out_665   [127:0]  ),
    .col_in_666              ( u0_col_out_666   [127:0]  ),
    .col_in_667              ( u0_col_out_667   [127:0]  ),
    .col_in_668              ( u0_col_out_668   [127:0]  ),
    .col_in_669              ( u0_col_out_669   [127:0]  ),
    .col_in_670              ( u0_col_out_670   [127:0]  ),
    .col_in_671              ( u0_col_out_671   [127:0]  ),
    .col_in_672              ( u0_col_out_672   [127:0]  ),
    .col_in_673              ( u0_col_out_673   [127:0]  ),
    .col_in_674              ( u0_col_out_674   [127:0]  ),
    .col_in_675              ( u0_col_out_675   [127:0]  ),
    .col_in_676              ( u0_col_out_676   [127:0]  ),
    .col_in_677              ( u0_col_out_677   [127:0]  ),
    .col_in_678              ( u0_col_out_678   [127:0]  ),
    .col_in_679              ( u0_col_out_679   [127:0]  ),
    .col_in_680              ( u0_col_out_680   [127:0]  ),
    .col_in_681              ( u0_col_out_681   [127:0]  ),
    .col_in_682              ( u0_col_out_682   [127:0]  ),
    .col_in_683              ( u0_col_out_683   [127:0]  ),
    .col_in_684              ( u0_col_out_684   [127:0]  ),
    .col_in_685              ( u0_col_out_685   [127:0]  ),
    .col_in_686              ( u0_col_out_686   [127:0]  ),
    .col_in_687              ( u0_col_out_687   [127:0]  ),
    .col_in_688              ( u0_col_out_688   [127:0]  ),
    .col_in_689              ( u0_col_out_689   [127:0]  ),
    .col_in_690              ( u0_col_out_690   [127:0]  ),
    .col_in_691              ( u0_col_out_691   [127:0]  ),
    .col_in_692              ( u0_col_out_692   [127:0]  ),
    .col_in_693              ( u0_col_out_693   [127:0]  ),
    .col_in_694              ( u0_col_out_694   [127:0]  ),
    .col_in_695              ( u0_col_out_695   [127:0]  ),
    .col_in_696              ( u0_col_out_696   [127:0]  ),
    .col_in_697              ( u0_col_out_697   [127:0]  ),
    .col_in_698              ( u0_col_out_698   [127:0]  ),
    .col_in_699              ( u0_col_out_699   [127:0]  ),
    .col_in_700              ( u0_col_out_700   [127:0]  ),
    .col_in_701              ( u0_col_out_701   [127:0]  ),
    .col_in_702              ( u0_col_out_702   [127:0]  ),
    .col_in_703              ( u0_col_out_703   [127:0]  ),
    .col_in_704              ( u0_col_out_704   [127:0]  ),
    .col_in_705              ( u0_col_out_705   [127:0]  ),
    .col_in_706              ( u0_col_out_706   [127:0]  ),
    .col_in_707              ( u0_col_out_707   [127:0]  ),
    .col_in_708              ( u0_col_out_708   [127:0]  ),
    .col_in_709              ( u0_col_out_709   [127:0]  ),
    .col_in_710              ( u0_col_out_710   [127:0]  ),
    .col_in_711              ( u0_col_out_711   [127:0]  ),
    .col_in_712              ( u0_col_out_712   [127:0]  ),
    .col_in_713              ( u0_col_out_713   [127:0]  ),
    .col_in_714              ( u0_col_out_714   [127:0]  ),
    .col_in_715              ( u0_col_out_715   [127:0]  ),
    .col_in_716              ( u0_col_out_716   [127:0]  ),
    .col_in_717              ( u0_col_out_717   [127:0]  ),
    .col_in_718              ( u0_col_out_718   [127:0]  ),
    .col_in_719              ( u0_col_out_719   [127:0]  ),
    .col_in_720              ( u0_col_out_720   [127:0]  ),
    .col_in_721              ( u0_col_out_721   [127:0]  ),
    .col_in_722              ( u0_col_out_722   [127:0]  ),
    .col_in_723              ( u0_col_out_723   [127:0]  ),
    .col_in_724              ( u0_col_out_724   [127:0]  ),
    .col_in_725              ( u0_col_out_725   [127:0]  ),
    .col_in_726              ( u0_col_out_726   [127:0]  ),
    .col_in_727              ( u0_col_out_727   [127:0]  ),
    .col_in_728              ( u0_col_out_728   [127:0]  ),
    .col_in_729              ( u0_col_out_729   [127:0]  ),
    .col_in_730              ( u0_col_out_730   [127:0]  ),
    .col_in_731              ( u0_col_out_731   [127:0]  ),
    .col_in_732              ( u0_col_out_732   [127:0]  ),
    .col_in_733              ( u0_col_out_733   [127:0]  ),
    .col_in_734              ( u0_col_out_734   [127:0]  ),
    .col_in_735              ( u0_col_out_735   [127:0]  ),
    .col_in_736              ( u0_col_out_736   [127:0]  ),
    .col_in_737              ( u0_col_out_737   [127:0]  ),
    .col_in_738              ( u0_col_out_738   [127:0]  ),
    .col_in_739              ( u0_col_out_739   [127:0]  ),
    .col_in_740              ( u0_col_out_740   [127:0]  ),
    .col_in_741              ( u0_col_out_741   [127:0]  ),
    .col_in_742              ( u0_col_out_742   [127:0]  ),
    .col_in_743              ( u0_col_out_743   [127:0]  ),
    .col_in_744              ( u0_col_out_744   [127:0]  ),
    .col_in_745              ( u0_col_out_745   [127:0]  ),
    .col_in_746              ( u0_col_out_746   [127:0]  ),
    .col_in_747              ( u0_col_out_747   [127:0]  ),
    .col_in_748              ( u0_col_out_748   [127:0]  ),
    .col_in_749              ( u0_col_out_749   [127:0]  ),
    .col_in_750              ( u0_col_out_750   [127:0]  ),
    .col_in_751              ( u0_col_out_751   [127:0]  ),
    .col_in_752              ( u0_col_out_752   [127:0]  ),
    .col_in_753              ( u0_col_out_753   [127:0]  ),
    .col_in_754              ( u0_col_out_754   [127:0]  ),
    .col_in_755              ( u0_col_out_755   [127:0]  ),
    .col_in_756              ( u0_col_out_756   [127:0]  ),
    .col_in_757              ( u0_col_out_757   [127:0]  ),
    .col_in_758              ( u0_col_out_758   [127:0]  ),
    .col_in_759              ( u0_col_out_759   [127:0]  ),
    .col_in_760              ( u0_col_out_760   [127:0]  ),
    .col_in_761              ( u0_col_out_761   [127:0]  ),
    .col_in_762              ( u0_col_out_762   [127:0]  ),
    .col_in_763              ( u0_col_out_763   [127:0]  ),
    .col_in_764              ( u0_col_out_764   [127:0]  ),
    .col_in_765              ( u0_col_out_765   [127:0]  ),
    .col_in_766              ( u0_col_out_766   [127:0]  ),
    .col_in_767              ( u0_col_out_767   [127:0]  ),
    .col_in_768              ( u0_col_out_768   [127:0]  ),
    .col_in_769              ( u0_col_out_769   [127:0]  ),
    .col_in_770              ( u0_col_out_770   [127:0]  ),
    .col_in_771              ( u0_col_out_771   [127:0]  ),
    .col_in_772              ( u0_col_out_772   [127:0]  ),
    .col_in_773              ( u0_col_out_773   [127:0]  ),
    .col_in_774              ( u0_col_out_774   [127:0]  ),
    .col_in_775              ( u0_col_out_775   [127:0]  ),
    .col_in_776              ( u0_col_out_776   [127:0]  ),
    .col_in_777              ( u0_col_out_777   [127:0]  ),
    .col_in_778              ( u0_col_out_778   [127:0]  ),
    .col_in_779              ( u0_col_out_779   [127:0]  ),
    .col_in_780              ( u0_col_out_780   [127:0]  ),
    .col_in_781              ( u0_col_out_781   [127:0]  ),
    .col_in_782              ( u0_col_out_782   [127:0]  ),
    .col_in_783              ( u0_col_out_783   [127:0]  ),
    .col_in_784              ( u0_col_out_784   [127:0]  ),
    .col_in_785              ( u0_col_out_785   [127:0]  ),
    .col_in_786              ( u0_col_out_786   [127:0]  ),
    .col_in_787              ( u0_col_out_787   [127:0]  ),
    .col_in_788              ( u0_col_out_788   [127:0]  ),
    .col_in_789              ( u0_col_out_789   [127:0]  ),
    .col_in_790              ( u0_col_out_790   [127:0]  ),
    .col_in_791              ( u0_col_out_791   [127:0]  ),
    .col_in_792              ( u0_col_out_792   [127:0]  ),
    .col_in_793              ( u0_col_out_793   [127:0]  ),
    .col_in_794              ( u0_col_out_794   [127:0]  ),
    .col_in_795              ( u0_col_out_795   [127:0]  ),
    .col_in_796              ( u0_col_out_796   [127:0]  ),
    .col_in_797              ( u0_col_out_797   [127:0]  ),
    .col_in_798              ( u0_col_out_798   [127:0]  ),
    .col_in_799              ( u0_col_out_799   [127:0]  ),
    .col_in_800              ( u0_col_out_800   [127:0]  ),
    .col_in_801              ( u0_col_out_801   [127:0]  ),
    .col_in_802              ( u0_col_out_802   [127:0]  ),
    .col_in_803              ( u0_col_out_803   [127:0]  ),
    .col_in_804              ( u0_col_out_804   [127:0]  ),
    .col_in_805              ( u0_col_out_805   [127:0]  ),
    .col_in_806              ( u0_col_out_806   [127:0]  ),
    .col_in_807              ( u0_col_out_807   [127:0]  ),
    .col_in_808              ( u0_col_out_808   [127:0]  ),
    .col_in_809              ( u0_col_out_809   [127:0]  ),
    .col_in_810              ( u0_col_out_810   [127:0]  ),
    .col_in_811              ( u0_col_out_811   [127:0]  ),
    .col_in_812              ( u0_col_out_812   [127:0]  ),
    .col_in_813              ( u0_col_out_813   [127:0]  ),
    .col_in_814              ( u0_col_out_814   [127:0]  ),
    .col_in_815              ( u0_col_out_815   [127:0]  ),
    .col_in_816              ( u0_col_out_816   [127:0]  ),
    .col_in_817              ( u0_col_out_817   [127:0]  ),
    .col_in_818              ( u0_col_out_818   [127:0]  ),
    .col_in_819              ( u0_col_out_819   [127:0]  ),
    .col_in_820              ( u0_col_out_820   [127:0]  ),
    .col_in_821              ( u0_col_out_821   [127:0]  ),
    .col_in_822              ( u0_col_out_822   [127:0]  ),
    .col_in_823              ( u0_col_out_823   [127:0]  ),
    .col_in_824              ( u0_col_out_824   [127:0]  ),
    .col_in_825              ( u0_col_out_825   [127:0]  ),
    .col_in_826              ( u0_col_out_826   [127:0]  ),
    .col_in_827              ( u0_col_out_827   [127:0]  ),
    .col_in_828              ( u0_col_out_828   [127:0]  ),
    .col_in_829              ( u0_col_out_829   [127:0]  ),
    .col_in_830              ( u0_col_out_830   [127:0]  ),
    .col_in_831              ( u0_col_out_831   [127:0]  ),
    .col_in_832              ( u0_col_out_832   [127:0]  ),
    .col_in_833              ( u0_col_out_833   [127:0]  ),
    .col_in_834              ( u0_col_out_834   [127:0]  ),
    .col_in_835              ( u0_col_out_835   [127:0]  ),
    .col_in_836              ( u0_col_out_836   [127:0]  ),
    .col_in_837              ( u0_col_out_837   [127:0]  ),
    .col_in_838              ( u0_col_out_838   [127:0]  ),
    .col_in_839              ( u0_col_out_839   [127:0]  ),
    .col_in_840              ( u0_col_out_840   [127:0]  ),
    .col_in_841              ( u0_col_out_841   [127:0]  ),
    .col_in_842              ( u0_col_out_842   [127:0]  ),
    .col_in_843              ( u0_col_out_843   [127:0]  ),
    .col_in_844              ( u0_col_out_844   [127:0]  ),
    .col_in_845              ( u0_col_out_845   [127:0]  ),
    .col_in_846              ( u0_col_out_846   [127:0]  ),
    .col_in_847              ( u0_col_out_847   [127:0]  ),
    .col_in_848              ( u0_col_out_848   [127:0]  ),
    .col_in_849              ( u0_col_out_849   [127:0]  ),
    .col_in_850              ( u0_col_out_850   [127:0]  ),
    .col_in_851              ( u0_col_out_851   [127:0]  ),
    .col_in_852              ( u0_col_out_852   [127:0]  ),
    .col_in_853              ( u0_col_out_853   [127:0]  ),
    .col_in_854              ( u0_col_out_854   [127:0]  ),
    .col_in_855              ( u0_col_out_855   [127:0]  ),
    .col_in_856              ( u0_col_out_856   [127:0]  ),
    .col_in_857              ( u0_col_out_857   [127:0]  ),
    .col_in_858              ( u0_col_out_858   [127:0]  ),
    .col_in_859              ( u0_col_out_859   [127:0]  ),
    .col_in_860              ( u0_col_out_860   [127:0]  ),
    .col_in_861              ( u0_col_out_861   [127:0]  ),
    .col_in_862              ( u0_col_out_862   [127:0]  ),
    .col_in_863              ( u0_col_out_863   [127:0]  ),
    .col_in_864              ( u0_col_out_864   [127:0]  ),
    .col_in_865              ( u0_col_out_865   [127:0]  ),
    .col_in_866              ( u0_col_out_866   [127:0]  ),
    .col_in_867              ( u0_col_out_867   [127:0]  ),
    .col_in_868              ( u0_col_out_868   [127:0]  ),
    .col_in_869              ( u0_col_out_869   [127:0]  ),
    .col_in_870              ( u0_col_out_870   [127:0]  ),
    .col_in_871              ( u0_col_out_871   [127:0]  ),
    .col_in_872              ( u0_col_out_872   [127:0]  ),
    .col_in_873              ( u0_col_out_873   [127:0]  ),
    .col_in_874              ( u0_col_out_874   [127:0]  ),
    .col_in_875              ( u0_col_out_875   [127:0]  ),
    .col_in_876              ( u0_col_out_876   [127:0]  ),
    .col_in_877              ( u0_col_out_877   [127:0]  ),
    .col_in_878              ( u0_col_out_878   [127:0]  ),
    .col_in_879              ( u0_col_out_879   [127:0]  ),
    .col_in_880              ( u0_col_out_880   [127:0]  ),
    .col_in_881              ( u0_col_out_881   [127:0]  ),
    .col_in_882              ( u0_col_out_882   [127:0]  ),
    .col_in_883              ( u0_col_out_883   [127:0]  ),
    .col_in_884              ( u0_col_out_884   [127:0]  ),
    .col_in_885              ( u0_col_out_885   [127:0]  ),
    .col_in_886              ( u0_col_out_886   [127:0]  ),
    .col_in_887              ( u0_col_out_887   [127:0]  ),
    .col_in_888              ( u0_col_out_888   [127:0]  ),
    .col_in_889              ( u0_col_out_889   [127:0]  ),
    .col_in_890              ( u0_col_out_890   [127:0]  ),
    .col_in_891              ( u0_col_out_891   [127:0]  ),
    .col_in_892              ( u0_col_out_892   [127:0]  ),
    .col_in_893              ( u0_col_out_893   [127:0]  ),
    .col_in_894              ( u0_col_out_894   [127:0]  ),
    .col_in_895              ( u0_col_out_895   [127:0]  ),
    .col_in_896              ( u0_col_out_896   [127:0]  ),
    .col_in_897              ( u0_col_out_897   [127:0]  ),
    .col_in_898              ( u0_col_out_898   [127:0]  ),
    .col_in_899              ( u0_col_out_899   [127:0]  ),
    .col_in_900              ( u0_col_out_900   [127:0]  ),
    .col_in_901              ( u0_col_out_901   [127:0]  ),
    .col_in_902              ( u0_col_out_902   [127:0]  ),
    .col_in_903              ( u0_col_out_903   [127:0]  ),
    .col_in_904              ( u0_col_out_904   [127:0]  ),
    .col_in_905              ( u0_col_out_905   [127:0]  ),
    .col_in_906              ( u0_col_out_906   [127:0]  ),
    .col_in_907              ( u0_col_out_907   [127:0]  ),
    .col_in_908              ( u0_col_out_908   [127:0]  ),
    .col_in_909              ( u0_col_out_909   [127:0]  ),
    .col_in_910              ( u0_col_out_910   [127:0]  ),
    .col_in_911              ( u0_col_out_911   [127:0]  ),
    .col_in_912              ( u0_col_out_912   [127:0]  ),
    .col_in_913              ( u0_col_out_913   [127:0]  ),
    .col_in_914              ( u0_col_out_914   [127:0]  ),
    .col_in_915              ( u0_col_out_915   [127:0]  ),
    .col_in_916              ( u0_col_out_916   [127:0]  ),
    .col_in_917              ( u0_col_out_917   [127:0]  ),
    .col_in_918              ( u0_col_out_918   [127:0]  ),
    .col_in_919              ( u0_col_out_919   [127:0]  ),
    .col_in_920              ( u0_col_out_920   [127:0]  ),
    .col_in_921              ( u0_col_out_921   [127:0]  ),
    .col_in_922              ( u0_col_out_922   [127:0]  ),
    .col_in_923              ( u0_col_out_923   [127:0]  ),
    .col_in_924              ( u0_col_out_924   [127:0]  ),
    .col_in_925              ( u0_col_out_925   [127:0]  ),
    .col_in_926              ( u0_col_out_926   [127:0]  ),
    .col_in_927              ( u0_col_out_927   [127:0]  ),
    .col_in_928              ( u0_col_out_928   [127:0]  ),
    .col_in_929              ( u0_col_out_929   [127:0]  ),
    .col_in_930              ( u0_col_out_930   [127:0]  ),
    .col_in_931              ( u0_col_out_931   [127:0]  ),
    .col_in_932              ( u0_col_out_932   [127:0]  ),
    .col_in_933              ( u0_col_out_933   [127:0]  ),
    .col_in_934              ( u0_col_out_934   [127:0]  ),
    .col_in_935              ( u0_col_out_935   [127:0]  ),
    .col_in_936              ( u0_col_out_936   [127:0]  ),
    .col_in_937              ( u0_col_out_937   [127:0]  ),
    .col_in_938              ( u0_col_out_938   [127:0]  ),
    .col_in_939              ( u0_col_out_939   [127:0]  ),
    .col_in_940              ( u0_col_out_940   [127:0]  ),
    .col_in_941              ( u0_col_out_941   [127:0]  ),
    .col_in_942              ( u0_col_out_942   [127:0]  ),
    .col_in_943              ( u0_col_out_943   [127:0]  ),
    .col_in_944              ( u0_col_out_944   [127:0]  ),
    .col_in_945              ( u0_col_out_945   [127:0]  ),
    .col_in_946              ( u0_col_out_946   [127:0]  ),
    .col_in_947              ( u0_col_out_947   [127:0]  ),
    .col_in_948              ( u0_col_out_948   [127:0]  ),
    .col_in_949              ( u0_col_out_949   [127:0]  ),
    .col_in_950              ( u0_col_out_950   [127:0]  ),
    .col_in_951              ( u0_col_out_951   [127:0]  ),
    .col_in_952              ( u0_col_out_952   [127:0]  ),
    .col_in_953              ( u0_col_out_953   [127:0]  ),
    .col_in_954              ( u0_col_out_954   [127:0]  ),
    .col_in_955              ( u0_col_out_955   [127:0]  ),
    .col_in_956              ( u0_col_out_956   [127:0]  ),
    .col_in_957              ( u0_col_out_957   [127:0]  ),
    .col_in_958              ( u0_col_out_958   [127:0]  ),
    .col_in_959              ( u0_col_out_959   [127:0]  ),
    .col_in_960              ( u0_col_out_960   [127:0]  ),
    .col_in_961              ( u0_col_out_961   [127:0]  ),
    .col_in_962              ( u0_col_out_962   [127:0]  ),
    .col_in_963              ( u0_col_out_963   [127:0]  ),
    .col_in_964              ( u0_col_out_964   [127:0]  ),
    .col_in_965              ( u0_col_out_965   [127:0]  ),
    .col_in_966              ( u0_col_out_966   [127:0]  ),
    .col_in_967              ( u0_col_out_967   [127:0]  ),
    .col_in_968              ( u0_col_out_968   [127:0]  ),
    .col_in_969              ( u0_col_out_969   [127:0]  ),
    .col_in_970              ( u0_col_out_970   [127:0]  ),
    .col_in_971              ( u0_col_out_971   [127:0]  ),
    .col_in_972              ( u0_col_out_972   [127:0]  ),
    .col_in_973              ( u0_col_out_973   [127:0]  ),
    .col_in_974              ( u0_col_out_974   [127:0]  ),
    .col_in_975              ( u0_col_out_975   [127:0]  ),
    .col_in_976              ( u0_col_out_976   [127:0]  ),
    .col_in_977              ( u0_col_out_977   [127:0]  ),
    .col_in_978              ( u0_col_out_978   [127:0]  ),
    .col_in_979              ( u0_col_out_979   [127:0]  ),
    .col_in_980              ( u0_col_out_980   [127:0]  ),
    .col_in_981              ( u0_col_out_981   [127:0]  ),
    .col_in_982              ( u0_col_out_982   [127:0]  ),
    .col_in_983              ( u0_col_out_983   [127:0]  ),
    .col_in_984              ( u0_col_out_984   [127:0]  ),
    .col_in_985              ( u0_col_out_985   [127:0]  ),
    .col_in_986              ( u0_col_out_986   [127:0]  ),
    .col_in_987              ( u0_col_out_987   [127:0]  ),
    .col_in_988              ( u0_col_out_988   [127:0]  ),
    .col_in_989              ( u0_col_out_989   [127:0]  ),
    .col_in_990              ( u0_col_out_990   [127:0]  ),
    .col_in_991              ( u0_col_out_991   [127:0]  ),
    .col_in_992              ( u0_col_out_992   [127:0]  ),
    .col_in_993              ( u0_col_out_993   [127:0]  ),
    .col_in_994              ( u0_col_out_994   [127:0]  ),
    .col_in_995              ( u0_col_out_995   [127:0]  ),
    .col_in_996              ( u0_col_out_996   [127:0]  ),
    .col_in_997              ( u0_col_out_997   [127:0]  ),
    .col_in_998              ( u0_col_out_998   [127:0]  ),
    .col_in_999              ( u0_col_out_999   [127:0]  ),
    .col_in_1000             ( u0_col_out_1000  [127:0]  ),
    .col_in_1001             ( u0_col_out_1001  [127:0]  ),
    .col_in_1002             ( u0_col_out_1002  [127:0]  ),
    .col_in_1003             ( u0_col_out_1003  [127:0]  ),
    .col_in_1004             ( u0_col_out_1004  [127:0]  ),
    .col_in_1005             ( u0_col_out_1005  [127:0]  ),
    .col_in_1006             ( u0_col_out_1006  [127:0]  ),
    .col_in_1007             ( u0_col_out_1007  [127:0]  ),
    .col_in_1008             ( u0_col_out_1008  [127:0]  ),
    .col_in_1009             ( u0_col_out_1009  [127:0]  ),
    .col_in_1010             ( u0_col_out_1010  [127:0]  ),
    .col_in_1011             ( u0_col_out_1011  [127:0]  ),
    .col_in_1012             ( u0_col_out_1012  [127:0]  ),
    .col_in_1013             ( u0_col_out_1013  [127:0]  ),
    .col_in_1014             ( u0_col_out_1014  [127:0]  ),
    .col_in_1015             ( u0_col_out_1015  [127:0]  ),
    .col_in_1016             ( u0_col_out_1016  [127:0]  ),
    .col_in_1017             ( u0_col_out_1017  [127:0]  ),
    .col_in_1018             ( u0_col_out_1018  [127:0]  ),
    .col_in_1019             ( u0_col_out_1019  [127:0]  ),
    .col_in_1020             ( u0_col_out_1020  [127:0]  ),
    .col_in_1021             ( u0_col_out_1021  [127:0]  ),
    .col_in_1022             ( u0_col_out_1022  [127:0]  ),
    .col_in_1023             ( u0_col_out_1023  [127:0]  ),
    .col_in_1024             ( u0_col_out_1024  [127:0]  ),
    .col_in_1025             ( u0_col_out_1025  [127:0]  ),
    .col_in_1026             ( u0_col_out_1026  [127:0]  ),
    .col_in_1027             ( u0_col_out_1027  [127:0]  ),
    .col_in_1028             ( u0_col_out_1028  [127:0]  ),
    .col_in_1029             ( u0_col_out_1029  [127:0]  ),
    .col_in_1030             ( u0_col_out_1030  [127:0]  ),
    .col_in_1031             ( u0_col_out_1031  [127:0]  ),
    .col_in_1032             ( u0_col_out_1032  [127:0]  ),
    .col_in_1033             ( u0_col_out_1033  [127:0]  ),
    .col_in_1034             ( u0_col_out_1034  [127:0]  ),
    .col_in_1035             ( u0_col_out_1035  [127:0]  ),
    .col_in_1036             ( u0_col_out_1036  [127:0]  ),
    .col_in_1037             ( u0_col_out_1037  [127:0]  ),
    .col_in_1038             ( u0_col_out_1038  [127:0]  ),
    .col_in_1039             ( u0_col_out_1039  [127:0]  ),
    .col_in_1040             ( u0_col_out_1040  [127:0]  ),
    .col_in_1041             ( u0_col_out_1041  [127:0]  ),
    .col_in_1042             ( u0_col_out_1042  [127:0]  ),
    .col_in_1043             ( u0_col_out_1043  [127:0]  ),
    .col_in_1044             ( u0_col_out_1044  [127:0]  ),
    .col_in_1045             ( u0_col_out_1045  [127:0]  ),
    .col_in_1046             ( u0_col_out_1046  [127:0]  ),
    .col_in_1047             ( u0_col_out_1047  [127:0]  ),
    .col_in_1048             ( u0_col_out_1048  [127:0]  ),
    .col_in_1049             ( u0_col_out_1049  [127:0]  ),
    .col_in_1050             ( u0_col_out_1050  [127:0]  ),
    .col_in_1051             ( u0_col_out_1051  [127:0]  ),
    .col_in_1052             ( u0_col_out_1052  [127:0]  ),
    .col_in_1053             ( u0_col_out_1053  [127:0]  ),
    .col_in_1054             ( u0_col_out_1054  [127:0]  ),
    .col_in_1055             ( u0_col_out_1055  [127:0]  ),
    .col_in_1056             ( u0_col_out_1056  [127:0]  ),
    .col_in_1057             ( u0_col_out_1057  [127:0]  ),
    .col_in_1058             ( u0_col_out_1058  [127:0]  ),
    .col_in_1059             ( u0_col_out_1059  [127:0]  ),
    .col_in_1060             ( u0_col_out_1060  [127:0]  ),
    .col_in_1061             ( u0_col_out_1061  [127:0]  ),
    .col_in_1062             ( u0_col_out_1062  [127:0]  ),
    .col_in_1063             ( u0_col_out_1063  [127:0]  ),
    .col_in_1064             ( u0_col_out_1064  [127:0]  ),
    .col_in_1065             ( u0_col_out_1065  [127:0]  ),
    .col_in_1066             ( u0_col_out_1066  [127:0]  ),
    .col_in_1067             ( u0_col_out_1067  [127:0]  ),
    .col_in_1068             ( u0_col_out_1068  [127:0]  ),
    .col_in_1069             ( u0_col_out_1069  [127:0]  ),
    .col_in_1070             ( u0_col_out_1070  [127:0]  ),
    .col_in_1071             ( u0_col_out_1071  [127:0]  ),
    .col_in_1072             ( u0_col_out_1072  [127:0]  ),
    .col_in_1073             ( u0_col_out_1073  [127:0]  ),
    .col_in_1074             ( u0_col_out_1074  [127:0]  ),
    .col_in_1075             ( u0_col_out_1075  [127:0]  ),
    .col_in_1076             ( u0_col_out_1076  [127:0]  ),
    .col_in_1077             ( u0_col_out_1077  [127:0]  ),
    .col_in_1078             ( u0_col_out_1078  [127:0]  ),
    .col_in_1079             ( u0_col_out_1079  [127:0]  ),
    .col_in_1080             ( u0_col_out_1080  [127:0]  ),
    .col_in_1081             ( u0_col_out_1081  [127:0]  ),
    .col_in_1082             ( u0_col_out_1082  [127:0]  ),
    .col_in_1083             ( u0_col_out_1083  [127:0]  ),
    .col_in_1084             ( u0_col_out_1084  [127:0]  ),
    .col_in_1085             ( u0_col_out_1085  [127:0]  ),
    .col_in_1086             ( u0_col_out_1086  [127:0]  ),
    .col_in_1087             ( u0_col_out_1087  [127:0]  ),
    .col_in_1088             ( u0_col_out_1088  [127:0]  ),
    .col_in_1089             ( u0_col_out_1089  [127:0]  ),
    .col_in_1090             ( u0_col_out_1090  [127:0]  ),
    .col_in_1091             ( u0_col_out_1091  [127:0]  ),
    .col_in_1092             ( u0_col_out_1092  [127:0]  ),
    .col_in_1093             ( u0_col_out_1093  [127:0]  ),
    .col_in_1094             ( u0_col_out_1094  [127:0]  ),
    .col_in_1095             ( u0_col_out_1095  [127:0]  ),
    .col_in_1096             ( u0_col_out_1096  [127:0]  ),
    .col_in_1097             ( u0_col_out_1097  [127:0]  ),
    .col_in_1098             ( u0_col_out_1098  [127:0]  ),
    .col_in_1099             ( u0_col_out_1099  [127:0]  ),
    .col_in_1100             ( u0_col_out_1100  [127:0]  ),
    .col_in_1101             ( u0_col_out_1101  [127:0]  ),
    .col_in_1102             ( u0_col_out_1102  [127:0]  ),
    .col_in_1103             ( u0_col_out_1103  [127:0]  ),
    .col_in_1104             ( u0_col_out_1104  [127:0]  ),
    .col_in_1105             ( u0_col_out_1105  [127:0]  ),
    .col_in_1106             ( u0_col_out_1106  [127:0]  ),
    .col_in_1107             ( u0_col_out_1107  [127:0]  ),
    .col_in_1108             ( u0_col_out_1108  [127:0]  ),
    .col_in_1109             ( u0_col_out_1109  [127:0]  ),
    .col_in_1110             ( u0_col_out_1110  [127:0]  ),
    .col_in_1111             ( u0_col_out_1111  [127:0]  ),
    .col_in_1112             ( u0_col_out_1112  [127:0]  ),
    .col_in_1113             ( u0_col_out_1113  [127:0]  ),
    .col_in_1114             ( u0_col_out_1114  [127:0]  ),
    .col_in_1115             ( u0_col_out_1115  [127:0]  ),
    .col_in_1116             ( u0_col_out_1116  [127:0]  ),
    .col_in_1117             ( u0_col_out_1117  [127:0]  ),
    .col_in_1118             ( u0_col_out_1118  [127:0]  ),
    .col_in_1119             ( u0_col_out_1119  [127:0]  ),
    .col_in_1120             ( u0_col_out_1120  [127:0]  ),
    .col_in_1121             ( u0_col_out_1121  [127:0]  ),
    .col_in_1122             ( u0_col_out_1122  [127:0]  ),
    .col_in_1123             ( u0_col_out_1123  [127:0]  ),
    .col_in_1124             ( u0_col_out_1124  [127:0]  ),
    .col_in_1125             ( u0_col_out_1125  [127:0]  ),
    .col_in_1126             ( u0_col_out_1126  [127:0]  ),
    .col_in_1127             ( u0_col_out_1127  [127:0]  ),
    .col_in_1128             ( u0_col_out_1128  [127:0]  ),
    .col_in_1129             ( u0_col_out_1129  [127:0]  ),
    .col_in_1130             ( u0_col_out_1130  [127:0]  ),
    .col_in_1131             ( u0_col_out_1131  [127:0]  ),
    .col_in_1132             ( u0_col_out_1132  [127:0]  ),
    .col_in_1133             ( u0_col_out_1133  [127:0]  ),
    .col_in_1134             ( u0_col_out_1134  [127:0]  ),
    .col_in_1135             ( u0_col_out_1135  [127:0]  ),
    .col_in_1136             ( u0_col_out_1136  [127:0]  ),
    .col_in_1137             ( u0_col_out_1137  [127:0]  ),
    .col_in_1138             ( u0_col_out_1138  [127:0]  ),
    .col_in_1139             ( u0_col_out_1139  [127:0]  ),
    .col_in_1140             ( u0_col_out_1140  [127:0]  ),
    .col_in_1141             ( u0_col_out_1141  [127:0]  ),
    .col_in_1142             ( u0_col_out_1142  [127:0]  ),
    .col_in_1143             ( u0_col_out_1143  [127:0]  ),
    .col_in_1144             ( u0_col_out_1144  [127:0]  ),
    .col_in_1145             ( u0_col_out_1145  [127:0]  ),
    .col_in_1146             ( u0_col_out_1146  [127:0]  ),
    .col_in_1147             ( u0_col_out_1147  [127:0]  ),
    .col_in_1148             ( u0_col_out_1148  [127:0]  ),
    .col_in_1149             ( u0_col_out_1149  [127:0]  ),
    .col_in_1150             ( u0_col_out_1150  [127:0]  ),
    .col_in_1151             ( u0_col_out_1151  [127:0]  ),
    .col_in_1152             ( u0_col_out_1152  [127:0]  ),
    .col_in_1153             ( u0_col_out_1153  [127:0]  ),
    .col_in_1154             ( u0_col_out_1154  [127:0]  ),
    .col_in_1155             ( u0_col_out_1155  [127:0]  ),
    .col_in_1156             ( u0_col_out_1156  [127:0]  ),
    .col_in_1157             ( u0_col_out_1157  [127:0]  ),
    .col_in_1158             ( u0_col_out_1158  [127:0]  ),
    .col_in_1159             ( u0_col_out_1159  [127:0]  ),
    .col_in_1160             ( u0_col_out_1160  [127:0]  ),
    .col_in_1161             ( u0_col_out_1161  [127:0]  ),
    .col_in_1162             ( u0_col_out_1162  [127:0]  ),
    .col_in_1163             ( u0_col_out_1163  [127:0]  ),
    .col_in_1164             ( u0_col_out_1164  [127:0]  ),
    .col_in_1165             ( u0_col_out_1165  [127:0]  ),
    .col_in_1166             ( u0_col_out_1166  [127:0]  ),
    .col_in_1167             ( u0_col_out_1167  [127:0]  ),
    .col_in_1168             ( u0_col_out_1168  [127:0]  ),
    .col_in_1169             ( u0_col_out_1169  [127:0]  ),
    .col_in_1170             ( u0_col_out_1170  [127:0]  ),
    .col_in_1171             ( u0_col_out_1171  [127:0]  ),
    .col_in_1172             ( u0_col_out_1172  [127:0]  ),
    .col_in_1173             ( u0_col_out_1173  [127:0]  ),
    .col_in_1174             ( u0_col_out_1174  [127:0]  ),
    .col_in_1175             ( u0_col_out_1175  [127:0]  ),
    .col_in_1176             ( u0_col_out_1176  [127:0]  ),
    .col_in_1177             ( u0_col_out_1177  [127:0]  ),
    .col_in_1178             ( u0_col_out_1178  [127:0]  ),
    .col_in_1179             ( u0_col_out_1179  [127:0]  ),
    .col_in_1180             ( u0_col_out_1180  [127:0]  ),
    .col_in_1181             ( u0_col_out_1181  [127:0]  ),
    .col_in_1182             ( u0_col_out_1182  [127:0]  ),
    .col_in_1183             ( u0_col_out_1183  [127:0]  ),
    .col_in_1184             ( u0_col_out_1184  [127:0]  ),
    .col_in_1185             ( u0_col_out_1185  [127:0]  ),
    .col_in_1186             ( u0_col_out_1186  [127:0]  ),
    .col_in_1187             ( u0_col_out_1187  [127:0]  ),
    .col_in_1188             ( u0_col_out_1188  [127:0]  ),
    .col_in_1189             ( u0_col_out_1189  [127:0]  ),
    .col_in_1190             ( u0_col_out_1190  [127:0]  ),
    .col_in_1191             ( u0_col_out_1191  [127:0]  ),
    .col_in_1192             ( u0_col_out_1192  [127:0]  ),
    .col_in_1193             ( u0_col_out_1193  [127:0]  ),
    .col_in_1194             ( u0_col_out_1194  [127:0]  ),
    .col_in_1195             ( u0_col_out_1195  [127:0]  ),
    .col_in_1196             ( u0_col_out_1196  [127:0]  ),
    .col_in_1197             ( u0_col_out_1197  [127:0]  ),
    .col_in_1198             ( u0_col_out_1198  [127:0]  ),
    .col_in_1199             ( u0_col_out_1199  [127:0]  ),
    .col_in_1200             ( u0_col_out_1200  [127:0]  ),
    .col_in_1201             ( u0_col_out_1201  [127:0]  ),
    .col_in_1202             ( u0_col_out_1202  [127:0]  ),
    .col_in_1203             ( u0_col_out_1203  [127:0]  ),
    .col_in_1204             ( u0_col_out_1204  [127:0]  ),
    .col_in_1205             ( u0_col_out_1205  [127:0]  ),
    .col_in_1206             ( u0_col_out_1206  [127:0]  ),
    .col_in_1207             ( u0_col_out_1207  [127:0]  ),
    .col_in_1208             ( u0_col_out_1208  [127:0]  ),
    .col_in_1209             ( u0_col_out_1209  [127:0]  ),
    .col_in_1210             ( u0_col_out_1210  [127:0]  ),
    .col_in_1211             ( u0_col_out_1211  [127:0]  ),
    .col_in_1212             ( u0_col_out_1212  [127:0]  ),
    .col_in_1213             ( u0_col_out_1213  [127:0]  ),
    .col_in_1214             ( u0_col_out_1214  [127:0]  ),
    .col_in_1215             ( u0_col_out_1215  [127:0]  ),
    .col_in_1216             ( u0_col_out_1216  [127:0]  ),
    .col_in_1217             ( u0_col_out_1217  [127:0]  ),
    .col_in_1218             ( u0_col_out_1218  [127:0]  ),
    .col_in_1219             ( u0_col_out_1219  [127:0]  ),
    .col_in_1220             ( u0_col_out_1220  [127:0]  ),
    .col_in_1221             ( u0_col_out_1221  [127:0]  ),
    .col_in_1222             ( u0_col_out_1222  [127:0]  ),
    .col_in_1223             ( u0_col_out_1223  [127:0]  ),
    .col_in_1224             ( u0_col_out_1224  [127:0]  ),
    .col_in_1225             ( u0_col_out_1225  [127:0]  ),
    .col_in_1226             ( u0_col_out_1226  [127:0]  ),
    .col_in_1227             ( u0_col_out_1227  [127:0]  ),
    .col_in_1228             ( u0_col_out_1228  [127:0]  ),
    .col_in_1229             ( u0_col_out_1229  [127:0]  ),
    .col_in_1230             ( u0_col_out_1230  [127:0]  ),
    .col_in_1231             ( u0_col_out_1231  [127:0]  ),
    .col_in_1232             ( u0_col_out_1232  [127:0]  ),
    .col_in_1233             ( u0_col_out_1233  [127:0]  ),
    .col_in_1234             ( u0_col_out_1234  [127:0]  ),
    .col_in_1235             ( u0_col_out_1235  [127:0]  ),
    .col_in_1236             ( u0_col_out_1236  [127:0]  ),
    .col_in_1237             ( u0_col_out_1237  [127:0]  ),
    .col_in_1238             ( u0_col_out_1238  [127:0]  ),
    .col_in_1239             ( u0_col_out_1239  [127:0]  ),
    .col_in_1240             ( u0_col_out_1240  [127:0]  ),
    .col_in_1241             ( u0_col_out_1241  [127:0]  ),
    .col_in_1242             ( u0_col_out_1242  [127:0]  ),
    .col_in_1243             ( u0_col_out_1243  [127:0]  ),
    .col_in_1244             ( u0_col_out_1244  [127:0]  ),
    .col_in_1245             ( u0_col_out_1245  [127:0]  ),
    .col_in_1246             ( u0_col_out_1246  [127:0]  ),
    .col_in_1247             ( u0_col_out_1247  [127:0]  ),
    .col_in_1248             ( u0_col_out_1248  [127:0]  ),
    .col_in_1249             ( u0_col_out_1249  [127:0]  ),
    .col_in_1250             ( u0_col_out_1250  [127:0]  ),
    .col_in_1251             ( u0_col_out_1251  [127:0]  ),
    .col_in_1252             ( u0_col_out_1252  [127:0]  ),
    .col_in_1253             ( u0_col_out_1253  [127:0]  ),
    .col_in_1254             ( u0_col_out_1254  [127:0]  ),
    .col_in_1255             ( u0_col_out_1255  [127:0]  ),
    .col_in_1256             ( u0_col_out_1256  [127:0]  ),
    .col_in_1257             ( u0_col_out_1257  [127:0]  ),
    .col_in_1258             ( u0_col_out_1258  [127:0]  ),
    .col_in_1259             ( u0_col_out_1259  [127:0]  ),
    .col_in_1260             ( u0_col_out_1260  [127:0]  ),
    .col_in_1261             ( u0_col_out_1261  [127:0]  ),
    .col_in_1262             ( u0_col_out_1262  [127:0]  ),
    .col_in_1263             ( u0_col_out_1263  [127:0]  ),
    .col_in_1264             ( u0_col_out_1264  [127:0]  ),
    .col_in_1265             ( u0_col_out_1265  [127:0]  ),
    .col_in_1266             ( u0_col_out_1266  [127:0]  ),
    .col_in_1267             ( u0_col_out_1267  [127:0]  ),
    .col_in_1268             ( u0_col_out_1268  [127:0]  ),
    .col_in_1269             ( u0_col_out_1269  [127:0]  ),
    .col_in_1270             ( u0_col_out_1270  [127:0]  ),
    .col_in_1271             ( u0_col_out_1271  [127:0]  ),
    .col_in_1272             ( u0_col_out_1272  [127:0]  ),
    .col_in_1273             ( u0_col_out_1273  [127:0]  ),
    .col_in_1274             ( u0_col_out_1274  [127:0]  ),
    .col_in_1275             ( u0_col_out_1275  [127:0]  ),
    .col_in_1276             ( u0_col_out_1276  [127:0]  ),
    .col_in_1277             ( u0_col_out_1277  [127:0]  ),
    .col_in_1278             ( u0_col_out_1278  [127:0]  ),
    .col_in_1279             ( u0_col_out_1279  [127:0]  ),

    .ms                      ( u1_ms           [1023:0] )
);











always@(posedge clk) begin
    if(rst) begin 
        state_current <= IDLE;
    end
    else begin
        state_current <= state_next;
    end
end

always@(posedge clk) begin
    if(rst) begin 
        counter <= 31'b0;
    end
    else begin
        if(valid) counter <= counter + 1'b1;
        else counter <= counter;

    end
end


always@(*)begin
    case(state_current)
    IDLE: 
        begin
            if(reg_start)
                state_next <= TRANS_DATA;
            else
                state_next <= IDLE;
        end

    TRANS_DATA: 
        begin
            state_next <= ACCUMLATE_1;
        end

    ACCUMLATE_1:
        begin 
            state_next <= ACCUMLATE_2;
        end

    ACCUMLATE_2: 
        begin
            state_next <= ACCUMLATE_3;
        end
    ACCUMLATE_3: 
        begin
            state_next <= ACCUMLATE_4;
        end
    ACCUMLATE_4: 
        begin
            state_next <= REDUCTION;
        end

    REDUCTION: 
        begin
            state_next <= FINISH;
        end

    FINISH: 
        begin
            if(counter < LOOPS)
                state_next <= ACCUMLATE_1;
            else
                state_next <= IDLE;
        end

    default: 
        begin
            state_next <= IDLE;
        end
    endcase
end


always@(posedge clk)begin
    case(state_next)
    IDLE: 
        begin
            reg_a           <= 1024'b0;
            //reg_b           <= 1024'b0;
            reg_u0_sel      <= 2'b00;
            reg_start       <= start;
            reg_clear_i     <= 1'b1;
            reg_valid       <= 1'b0;
        end

    TRANS_DATA: 
        begin
            reg_a           <= a;
            //reg_b           <= a;
            reg_u0_sel      <= 2'b00;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b0;
        end

    ACCUMLATE_1:
        begin 
            reg_a           <= {reg_a[895:0], reg_a[1023:896]};
            //reg_b           <= reg_b << 256;
            reg_u0_sel      <= 2'b01;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b0;
        end

    ACCUMLATE_2: 
        begin
            reg_a           <= {reg_a[895:0], reg_a[1023:896]};
            //reg_b           <= reg_b << 256;
            reg_u0_sel      <= 2'b10;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b0;
        end
    ACCUMLATE_3: 
        begin
            reg_a           <= {reg_a[895:0], reg_a[1023:896]};
            //reg_b           <= reg_b << 256;
            reg_u0_sel      <= 2'b11;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b0;            
        end
    ACCUMLATE_4: 
        begin
            reg_a           <= 1024'h0;
            //reg_b           <= reg_b << 256;
            reg_u0_sel      <= 2'b00;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b0;
        end

    REDUCTION: 
        begin
            reg_a           <= 1204'h0;
            //reg_b           <= reg_b << 256;
            reg_u0_sel      <= 2'b00;
            reg_start       <= start;
            reg_clear_i     <= 1'b1;
            reg_valid       <= 1'b0;
        end

    FINISH: 
        begin
            reg_a           <= u1_ms;
            //reg_b           <= u1_ms;
            reg_u0_sel      <= 2'b00;
            reg_start       <= start;
            reg_clear_i     <= 1'b0;
            reg_valid       <= 1'b1;
        end

    default: 
        begin
            reg_a           <= 1024'b0;
            //reg_b           <= 1024'b0;
            reg_start       <= start;
            reg_clear_i     <= 1'b1;
            reg_valid       <= 1'b0;
        end
    endcase
end



assign ms = reg_a;
assign valid = reg_valid;

endmodule
module xpb_5_410
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4a339bb343616408b061ca7a3f9e943e06b14b41118e5b610fed6874a0e1ee4fa1681080af2b3e40b84d13ff062e782c7a789f3509a8ca4fd50a3d8cc5b51ea35d198a937c2f947b5b98d025bd12da5907fdd74eaca7e2ccfadb6475e988c7d6d690202a1b90dfd9288290ddeaf9c6331c1fa892e0eaef0893385b223980a9bf;
    5'b00010 : xpb = 1024'h9467376686c2c81160c394f47f3d287c0d629682231cb6c21fdad0e941c3dc9f42d021015e567c81709a27fe0c5cf058f4f13e6a1351949faa147b198b6a3d46ba331526f85f28f6b731a04b7a25b4b20ffbae9d594fc599f5b6c8ebd3118fadad2040543721bfb2510521bbd5f38c66383f5125c1d5de112670b6447301537e;
    5'b00011 : xpb = 1024'h2ded8dc40835f751461fe797ae817568a29dde925f3371abb1eb80082fa31de6e0efb409435b3c338988fcb62f2d57bb0b4fb5b8fa478ea3ce7f7948164ce738a2fd6b0bc4fdc02d00306dce9e5ccada23f48c5379717b563b059b67026fb4f254a8ce54a1e9a6fdf2c7cbbac91d2c7005851ad652756fe973399662239f96d2;
    5'b00100 : xpb = 1024'h782129774b975b59f681b211ee2009a6a94f29d370c1cd0cc1d8e87cd0850c368257c489f2867a7441d610b5355bcfe785c854ee03f058f3a389b6d4dc0205dc0016f59f412d54a85bc93df45b6fa5332bf263a226195e2335e0ffdcebf87cc92b38ee7ebd7a86d71b4a5c98b416f2a321a4c36933605ef20671f1845d204091;
    5'b00101 : xpb = 1024'h11a77fd4cd0a8a99dbde04b51d6456933e8a71e3acd887f653e9979bbe644d7e20775791d78b3a265ac4e56d582c37499c26cc3ceae652f7c7f4b50366e4afcde8e14b840dcbebdea4c80b777fa6bb5b3feb4158463b13df7b2fd2581b56a20dd2c17c7f28426e22bd0d0697a74092aceeea8d19c3fff0ca533ad1a20dbe83e5;
    5'b00110 : xpb = 1024'h5bdb1b88106beea28c3fcf2f5d02ead1453bbd24be66e35763d700105f463bcdc1df681286b678671311f96c5e5aaf76169f6b71f48f1d479cfef2902c99ce7145fad61789fb805a0060db9d3cb995b447e918a6f2e2f6ac760b36ce04df69e4a9519ca943d34dfbe58f9775923a58e00b0a35aca4eadfd2e6732cc4473f2da4;
    5'b00111 : xpb = 1024'ha60eb73b53cd52ab3ca199a99ca17f0f4bed0865cff53eb873c4688500282a1d6347789335e1b6a7cb5f0d6b648927a291180aa6fe37e7977209301cf24eed14a31460ab062b14d55bf9abc2f9cc700d4fe6eff59f8ad97970e69b43ee6831bb7fe1bcd35f642dd50e1228537d341f132729de3f85d5cedb79ab87e680bfd763;
    5'b01000 : xpb = 1024'h3f950d98d54081eb21fdec4ccbe5cbfbe12850760c0bf9a205d517a3ee076b6501670b9b1ae67659e44de22387598f04a77681f5e52de19b96742e4b7d3197068bdeb68fd2c9ac0ba4f879461e03863563dfcdabbfac8f35b6356dbf1dc65700276a4ad3ca2c1520afd4d252705dbf1cf46fa7f0167560b3c6746804315e1ab7;
    5'b01001 : xpb = 1024'h89c8a94c18a1e5f3d25fb6c70b846039e7d99bb71d9a550315c280188ee959b4a2cf1c1bca11b49a9c9af6228d88073121ef212aeed6abeb6b7e6bd842e6b5a9e8f841234ef940870091496bdb16608e6bdda4fa6c547202b110d235074f1ed6fdfa6afde5bcf4f9d85763305b578550108f5082f7604fbc59acc3266adec476;
    5'b01010 : xpb = 1024'h234effa99a151533b7bc096a3ac8ad267d14e3c759b10feca7d32f377cc89afc40eeaf23af16744cb589cadab0586e93384d9879d5cca5ef8fe96a06cdc95f9bd1c297081b97d7bd499016eeff4d76b67fd682b08c7627bef65fa4b036ad441ba582f8fe5084dc457a1a0d2f4e812559ddd51a3387ffe194a675a3441b7d07ca;
    5'b01011 : xpb = 1024'h6d829b5cdd76793c681dd3e47a67416483c62f086b3f6b4db7c097ac1daa894be256bfa45e41b28d6dd6ded9b686e6bfb2c637aedf75703f64f3a793937e7e3f2edc219b97c76c38a528e714bc60510f87d459ff391e0a8bf13b092620360bf27c1319286c15bc1ea29c9e0d397aeb8cf9f4c2c668ead09d39adfe6654fdb189;
    5'b01100 : xpb = 1024'h708f1ba5ee9a87c4d7a2687a9ab8e5119017718a756263749d146cb0b89ca93807652ac4346723f86c5b391d9574e21c924aefdc66b6a43895ea5c21e61283117a677806466036eee27b497e09767379bcd37b5593fc0483689dba14f943137239ba728d6dda36a445f480c2ca48b96c73a8c76f98a62758676de84059bf4dd;
    5'b01101 : xpb = 1024'h513c8d6da24b0c84fddbf101e94a228f1fb2c259b8e4819859beaf3fac6bb8e321de632cf271b0803f12c790df85c64e439d4e32d01434935e68e34ee41646d474c00213e09597ea49c084bd9daa4190a3cb0f0405e7a31531654017391cf90dfa2bc752f26e83436ce1d8ea179e51c9e35a3509da75517e19af39a63f1c9e9c;
    5'b01110 : xpb = 1024'h9b702920e5ac708dae3dbb7c28e8b6cd26640d9aca72dcf969ac17b44d4da732c34673ada19ceec0f75fdb8fe5b43e7abe15ed67d9bcfee3337320dba9cb6577d1d98ca75cc52c65a55954e35abd1be9abc8e652b28f85e22c40a48d22a5c0e4d0bbe77d0dff631c956469c8029817fcff79dd9cbb604086ace794c8789d485b;
    5'b01111 : xpb = 1024'h34f67f7e671f9fcd939a0e1f582d03b9bb9f55ab068997e2fbbcc6d33b2ce87a616606b586a1ae73104eb0480884a5dcd47464b6c0b2f8e757de1f0a34ae0f69baa3e28c2963c39bee5822667ef43211bfc1c408d2b13b9e718f77085203e6297844757d78c74a68372713c6f5c1b806ccbfa74d4bffd25ef9b074e6293b8baf;
    5'b10000 : xpb = 1024'h7f2a1b31aa8103d643fbd89997cb97f7c250a0ec1817f3440baa2f47dc0ed6ca02ce173635ccecb3c89bc4470eb31e094eed03ebca5bc3372ce85c96fa632e0d17bd6d1fa593581749f0f28c3c070c6ac7bf9b577f591e6b6c6adb7e3b8cae004ed495a794582a415fa9a4a4e0bb7e39e8df4fe02ceac1678ce8d00862bc356e;
    5'b10001 : xpb = 1024'h18b0718f2bf4331629582b3cc70fe4e4578be8fc542eae2d9dbade66c9ee1811a0edaa3e1ad1ac65e18a98ff3183856b654b7b3ab151bd3b51535ac58545d7ff0087c3047231ef4d92efc00f603e2292dbb8790d9f7ad427b1b9adf96aead344f65d23a7ff20118d016c4ea3d3e51e43b6251990bd8a533fd9b1b026135a78c2;
    5'b10010 : xpb = 1024'h62e40d426f55971ed9b9f5b706ae79225e3d343d65bd098eada846db6ad006614255babec9fceaa699d7acfe37b1fd97dfc41a6fbafa878b265d98524afaf6a25da14d97ee6183c8ee8890351d50fcebe3b6505c4c22b6f4ac95126f54739b1bcced43d21ab0f16629eedf81bedee476d244c2239e7542486cea0b484cdb2281;
    5'b10011 : xpb = 1024'had17a8f5b2b6fb278a1bc031464d0d6064ee7f7e774b64efbd95af500bb1f4b0e3bdcb3f792828e75224c0fd3de075c45a3cb9a4c4a351dafb67d5df10b01545babad82b6a9118444a21605ada63d744ebb427aaf8ca99c1a77076e53dfc62f2a37d63fc3641d13f5271705fa9d8aaa9ee646ab67f6031510022666a865bcc40;
    5'b10100 : xpb = 1024'h469dff53342a2a676f7812d475915a4cfa29c78eb3621fd94fa65e6ef99135f881dd5e475e2ce8996b1395b560b0dd26709b30f3ab994bdf1fd2d40d9b92bf37a3852e10372faf7a93202dddfe9aed6cffad056118ec4f7decbf49606d5a88374b05f1fca109b88af4341a5e9d024ab3bbaa34670fffc3294ceb468836fa0f94;
    5'b10101 : xpb = 1024'h90d19b06778b8e701fd9dd4eb52fee8b00db12cfc4f07b3a5f93c6e39a73244823456ec80d5826da2360a9b466df5552eb13d028b542162ef4dd119a6147dddb009eb8a3b35f43f5eeb8fe03bbadc7c607aadcafc594324ae79aadd656e3500e21961226bc9a98641cb6ab3c87fc10e6d7c9dcf9f0eab231e023a1aa707ab953;
    5'b10110 : xpb = 1024'h2a57f163f8febdb005362ff1e4743b7796165ae001073623f1a476028852658fc16501cff25ce68c3c4f7e6c89afbcb5017247779c38103319480fc8ec2a87cce9690e887ffddb2c37b7cb86dfe4ddee1ba3ba65e5b5e8072ce9805186417552c91ea02727627fafbe79553b7b25b0f0a50fa6aa818a440a2cec81c82118fca7;
    5'b10111 : xpb = 1024'h748b8d173c6021b8b597fa6c2412cfb59cc7a621129591850191de77293453df62cd1250a18824ccf49c926b8fde34e17beae6aca5e0da82ee524d55b1dfa6704682991bfc2d6fa793509bac9cf7b84723a191b4925dcad427c4e4c76fca3d299faec05142f35f88e6fbe619661f7723c12f4f3d62753312c024dcea5a99a666;
    5'b11000 : xpb = 1024'he11e374bdd350f89af44d0f53571ca23202ee314eac4c6e93a28d961713952700eca558868ce47f0d8b6723b2ae9c4392495dfb8cd6d48712bd4b843cc250622f4cef00c8cc06dddc4f692fc12ece6f379a6f6ab27f80906d13b7429f28626e47374e51adbb46d488be90185949172d8e7518edf314c4eb0cedbd080b37e9ba;
    5'b11001 : xpb = 1024'h58457f280134b5014b56178992f5b0e038b43972603aa7cfa38ff60ab7f58376a254b5d935b822bfc5d87b22b8dd14700cc1fd30967f9ed6e7c7891102776f058c66799444fb9b5937e839557e41a8c83f9846b95f27635d67ef1bb888b12a451dc76e7bc94c26adb14120f64442dd60aa94c180d3ffb3f3a026182a44b89379;
    5'b11010 : xpb = 1024'ha2791adb44961909fbb7e203d294451e3f6584b371c90330b37d5e7f58d771c643bcc659e4e361007e258f21bf0b8c9c873a9c65a0286926bcd1c69dc82c8da8e9800427c12b2fd49381097b3b54832147961e080bcf462a62ca802e7239f21bf4578ea5e4dd0686d9c3b1d42f3ca393c6b46a13b4eaa2fc335e734c7e393d38;
    5'b11011 : xpb = 1024'h3bff7138c6094849e11434a701d8920ad4a0ccc3addfbe1a458e0d9e46b6b30de1dc5961c9e820b2971463d9e1dbf3fe9d9913b4871e632ae13cc4cc530f379ad24a5a0c8dc9c70adc7fd6fe5f8b99495b8efbbe2bf0fbe6a81952a9a19817609be01ca64fa4edd27b865bd32266439d93fa33c4458a34d48027536a2ed7808c;
    5'b11100 : xpb = 1024'h86330cec096aac529175ff2141772648db521804bf6e197b557b7612e798a15d834469e279135ef34f6177d8e80a6c2b1811b2e990c72d7ab647025918c4563e2f63e4a009f95b863818a7241c9e73a2638cd30cd898deb3a2f4b71f8b20df3772703cd06b35cdaba408ecb10d6009d0b019dc57267523dd135fae8c68582a4b;
    5'b11101 : xpb = 1024'h1fb963498adddb9276d251c470bb7335708d6014fb84d464e78c2531d577e2a52163fcea5e181ea568504c910adad38d2e702a3877bd277edab20087a3a70030182e3a84d697f2bc811774a740d589ca7785b0c2f8ba946fe843899aba7f047c19f8cad0d5fdb4f745cb96b00089a9da7d5fa607b714b5b560288eaa18f66d9f;
    5'b11110 : xpb = 1024'h69ecfefcce3f3f9b27341c3eb05a0773773eab560d132fc5f7798da67659d0f4c2cc0d6b0d435ce6209d609011094bb9a8e8c96d8165f1ceafbc3e14695c1ed37547c51852c78737dcb044ccfde864237f838811a562773ce31eee10a407cc52f088eafaf18e94d06e4e278deb83700d997f4e9a97ffa4bdf360e9cc5277175e;
    5'b11111 : xpb = 1024'h373555a4fb26edb0c906ee1df9e54600c79f3664929eaaf898a3cc56439123c60eba072f2481c98398c354833d9b31bbf4740bc685bebd2d4273c42f43ec8c55e121afd1f661e6e25af1250221f7a4b937c65c7c5842cf9286dc08bd365f197981178fb5c567c1c1010d18cdead101766c5184b289f36964029c9ea03155ab2;
    endcase
end

endmodule

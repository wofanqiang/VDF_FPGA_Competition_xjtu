module xpb_5_800
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h489139defb7ea23aaf96056241b51944cf0cae579d82d196324e1afdf4925174c5970c5d41f47ceb98484595525c10bb46a71b087f2fc05364d1a3e26ebf495af2406d6e65b98a794507c5a66066fcb43da571f9fcf269e34aecdfdd9488ac9e1ce0792cda9bd8d56b70727446cf854d2fea0064ee5db2469ad326aa480876ae;
    5'b00010 : xpb = 1024'h912273bdf6fd44755f2c0ac4836a32899e195caf3b05a32c649c35fbe924a2e98b2e18ba83e8f9d730908b2aa4b821768d4e3610fe5f80a6c9a347c4dd7e92b5e480dadccb7314f28a0f8b4cc0cdf9687b4ae3f3f9e4d3c695d9bfbb2911593c39c0f259b537b1aad6e0e4e88d9f0a9a5fd400c9dcbb648d35a64d549010ed5c;
    5'b00011 : xpb = 1024'h29066847308db1e743bc984fb4c5047cfbb007d60310d44b190d97a42ab447564d7ca79efbb6f834297a917913b621676fdb29335adc70ae7dd5ac49116b675f6272139c819ba226bc7d4e50885931ebc4eb5c556a5110992b3a0d9e036f63482799d95cdf0a91f2bb91707ddc9e69be40e4224c7acdb9a38a09f8fa4f36fd9f;
    5'b00100 : xpb = 1024'h7197a2262c0c5421f3529db1f67a1dc1cabcb62da093a5e14b5bb2a21f4698cb1313b3fc3dab751fc1c2d70e66123222b682443bda0c3101e2a7502b802ab0ba54b2810ae7552ca0018513f6e8c02ea00290ce4f67437a7c7626ed7b97f80fe6447a5289b9a66ac82701e2f2236def0b70ce22b1692b6bea24dd1fa4973f744d;
    5'b00101 : xpb = 1024'h97b96af659cc193d7e32b3d27d4efb528536154689ed6ffffcd144a60d63d37d56242e0b579737cbaacdd5cd5103213990f375e3689210996d9b4afb4178563d2a3b9ca9d7db9d433f2d6fab04b67234c3146b0d7afb74f0b873b5e725619f23253398ce3794b100bb26e87726d4e2f51de4434073dc1007940cb4a56658490;
    5'b00110 : xpb = 1024'h520cd08e611b63ce8779309f698a08f9f7600fac0621a896321b2f4855688eac9af94f3df76df06852f522f2276c42cedfb65266b5b8e15cfbab589222d6cebec4e427390337444d78fa9ca110b263d789d6b8aad4a2213256741b3c06dec6904f33b2b9be1523e57722e0fbb93cd37c81c84498f59b73471413f1f49e6dfb3e;
    5'b00111 : xpb = 1024'h9a9e0a6d5c9a0609370f3601ab3f223ec66cbe03a3a47a2c64694a4649fae02160905b9b39626d53eb3d688779c8538a265d6d6f34e8a1b0607cfc7491961819b72494a768f0cec6be0262477119608bc77c2aa4d1948b15a160fb199b67732e6c142be698b0fcbae2935370000c58c9b1b244fde3f9258daee7189ee67671ec;
    5'b01000 : xpb = 1024'h3281fef6962a737b1b9fc38cdc99f4322403692a6bafab4b18daabee8b8a848e22deea7fb1306bb0e4276ed5e8c6537b08ea6091916591b814af60f8c582ecc33515cd671f195bfaf070254b38a4990f111ca3064200c7e836c148fc75c57d3a59ed12e9c283dd02c743df054f0bb7ed92c26680820b7aa4034ac444a59c822f;
    5'b01001 : xpb = 1024'h7b1338d591a915b5cb35c8ef1e4f0d76f310178209327ce14b28c6ec801cd602e875f6dcf324e89c7c6fb46b3b2264364f917b9a1095520b798104db3442361e27563ad584d2e6743577eaf1990b95c34ec215003ef331cb81ae28da0a4e29d876cd8c169d1fb5d832b4517995db3d3ac2ac66e570692cea9e1deaeeeda4f8dd;
    5'b01010 : xpb = 1024'h12f72d5ecb398327afc6567a4fa9df6a50a6c2a8d13dadffff9a2894c1ac7a6faac485c16af2e6f97559bab9aa206427321e6ebc6d1242132db3695f682f0ac7a54773953afb73a867e5adf56096ce4698628d61af5f6e9e170e76bce4ac33e464a67319c6f296201764dd0ee4da9c5ea3bc88680e7b8200f2819694accb0920;
    5'b01011 : xpb = 1024'h5b88673dc6b825625f5c5bdc915ef8af1fb371006ec07f9631e84392b63ecbe4705b921eace763e50da2004efc7c74e278c589c4ec42026692850d41d6ee54229787e103a0b4fe21aced739bc0fdcafad607ff5bac51d88161fb569a7934e0828186ec46a18e6ef582d54f832baa21abd3a688ccfcd934478d54bd3ef4d37fce;
    5'b01100 : xpb = 1024'ha419a11cc236c79d0ef2613ed31411f3eec01f580c43512c64365e90aad11d5935f29e7beedbe0d0a5ea45e44ed8859dbf6ca4cd6b71c2b9f756b12445ad9d7d89c84e72066e889af1f539422164c7af13ad7155a9444264ace836780dbd8d209e6765737c2a47caee45c1f77279a6f903908931eb36e68e2827e3e93cdbf67c;
    5'b01101 : xpb = 1024'h3bfd95a5fbc7350ef382eeca046ee3e74c56ca7ed44e824b18a7c038ec60c1c5f8412d6066a9df2d9ed44c32bdd6858ea1f997efc7eeb2c1ab8915a8799a722707b98731bc9715cf2462fc45e8f000325d4de9b719b07f374248845ae81b972c8c404c76a5fd2812d2f64d8cc179061ce4a0aab489493ba47c8b8f8efc0206bf;
    5'b01110 : xpb = 1024'h848ecf84f745d749a318f42c4623fd2c1b6378d671d153e14af5db36e0f3133abdd839bda89e5c19371c91c810329649e8a0b2f8471e7315105ab98ae859bb81f9f9f4a02250a048696ac1ec4956fce69af35bb116a2e91a8d3564387ca443caa920c5a3809900e83e66c00108488b6a148aab1977a6edeb175eb639440a7d6d;
    5'b01111 : xpb = 1024'h1c72c40e30d644bb87a981b7777ecf1f78fa23fd39dc84ffff673cdf2282b7a78026c8a2206c5a76300698167f30963acb2da61aa39b631cc48d1e0f1c46902b77eb2d5fd8792d7c9bd884f010e23569e493d412870f25ed2295b21b57024dd696f9aca6aa6be13023174b965747ea8df59acc9c15b943016bc261df03308db0;
    5'b10000 : xpb = 1024'h6503fded2c54e6f6373f8719b933e8644806d254d75f569631b557dd1715091c45bdd4ff6260d761c84eddabd18ca6f611d4c12322cb2370295ec1f18b05d9866a2b9ace3e32b7f5e0e04a967149321e2239460c84018fd06d8291f8eb8afa74b3da25d38507ba058e87be0a9e176fdb2584cd010416f548069588894b39045e;
    5'b10001 : xpb = 1024'had9537cc27d38930e6d58c7bfae901a9171380ac74e2282c640372db0ba75a910b54e15ca455544d6097234123e8b7b1587bdc2ba1fae3c38e3065d3f9c522e15c6c083ca3ec426f25e8103cd1b02ed25fdeb80680f3f9b3b86f71d68013a712d0ba9f005fa392daf9f8307ee4e6f528556ecd65f274a78ea168af3393417b0c;
    5'b10010 : xpb = 1024'h45792c556163f6a2cb661a072c43d39c74aa2bd33ced594b1874d4834d36fefdcda370411c2352aa5981298f92e6b7a23b08cf4dfe77d3cb4262ca582db1f78ada5d40fc5a14cfa35855d340993b6755a97f3067f16036864dcfbfb95a71b11ebe93860389767322dea8bc1433e6544c367eeee89086fca4f5cc5ad952678b4f;
    5'b10011 : xpb = 1024'h8e0a66345ce298dd7afc1f696df8ece143b6da2ada702ae14ac2ef8141c95072933a7c9e5e17cf95f1c96f24e542c85d81afea567da7941ea7346e3a9c7140e5cc9dae6abfce5a1c9d5d98e6f9a26409e724a261ee52a06998bc9f96eefa5dbcdb73ff3064124bf84a192e887ab5d9996668ef4d7ee4aeeb909f81839a7001fd;
    5'b10100 : xpb = 1024'h25ee5abd9673064f5f8cacf49f53bed4a14d8551a27b5bffff3451298358f4df55890b82d5e5cdf2eab375735440c84e643cdd78da2484265b66d2bed05e158f4a8ee72a75f6e750cfcb5beac12d9c8d30c51ac35ebedd3c2e1ced79c95867c8c94ce6338de52c402ec9ba1dc9b538bd477910d01cf70401e5032d2959961240;
    5'b10101 : xpb = 1024'h6e7f949c91f1a88a0f22b256e108d819705a33a93ffe2d9631826c2777eb46541b2017e017da4ade82fbbb08a69cd909aae3f88159544479c03876a13f1d5eea3ccf5498dbb071ca14d32191219499416e6a8cbd5bb1471f7909cd575de11466e62d5f60688105159a3a2c921084be0a776311350b54b6487fd653d3a19e88ee;
    5'b10110 : xpb = 1024'h6638925cb8215fbf3b33fe21263aa0ccdf0ded008095eb4e5f3cdcfb97aeac0dd6ea6c48fa8493b7be5c157159ad8fa8d70eba3b5d13481746adb25730a3393bac08d5891d8fefe4740e494e91fd1c4b80b051ecc1d83f20e6a1b3a383f1e72d40646639253e55d7eeab8275f841d2e587332b7a9670b5ed439ff7960c49931;
    5'b10111 : xpb = 1024'h4ef4c304c700b836a34945445418c3519cfd8d27a58c304b1841e8cdae0d3c35a305b321d19cc627142e06ec67f6e9b5d41806ac3500f4d4d93c7f07e1c97ceead00fac6f79289778c48aa3b4986ce78f5b07718c90fedd55956fb17ccc7cb10f0e6bf906cefbe32ea5b2a9ba653a27b885d331c97c4bda56f0d2623a8cd0fdf;
    5'b11000 : xpb = 1024'h9785fce3c27f5a7152df4aa695cddc966c0a3b7f430f01e14a9003cba29f8daa689cbf7f13914312ac764c81ba52fa711abf21b4b430b5283e0e22ea5088c6499f4168355d4c13f0d1506fe1a9edcb2d3355e912c60257b8a443daf5615077af0dc738bd478b970855cb9d0fed2327c8b847338186226fec09e04ccdf0d5868d;
    5'b11001 : xpb = 1024'h2f69f16cfc0fc7e3376fd831c728ae89c9a0e6a60b1a32ffff016573e42f32172aeb4e638b5f416fa56052d02950fa61fd4c14d710ada52ff240876e84759af31d32a0f51374a12503be32e5717903b07cf66174366e948b39a428d83bae81bafba01fc0715e77503a7c28a53c2286ec995755042434c5025e43f873affb96d0;
    5'b11010 : xpb = 1024'h77fb2b4bf78e6a1de705dd9408ddc7ce98ad94fda89d0496314f8071d8c1838bf0825ac0cd53be5b3da898657bad0b1d43f32fdf8fdd658357122b50f334e44e0f730e63792e2b9e48c5f88bd1e00064ba9bd36e3360fe6e849108b5d0372e59188098ed4bfa5025a5ec9b1982f20c39c941556912927748f9171f1df8040d7e;
    5'b11011 : xpb = 1024'hfdf1fd5311ed78fcb966b1f3a3899c1f644402470a835b4e5c0e21a1a5127f8b2d0e9a54521bcb836929eb3eaab0b0e26802301ec5a558b0b448fd52721b8f78d6447232f56b8d27b33bb8f996b38e8043c4bcfa3cd3b4119f15698aa95386506597ff075cd306d8a9d26aed1f16b5daa5176ebb0a4cc5f4d7acac3b72a1dc1;
    5'b11100 : xpb = 1024'h587059b42c9d79ca7b2c70817bedb306c550ee7c0e2b074b180efd180ee3796d7867f602871639a3cedae4493d071bc96d273e0a6b8a15de701633b795e102527fa4b4919510434bc03b8135f9d2359c41e1bdc9a0bfa52464de36763f1de5032339f91d50690942f60d992318c0f0aada3b77509f027ea5e84df16dff32946f;
    5'b11101 : xpb = 1024'ha1019393281c1c052ac275e3bda2cc4b945d9cd3abadd8e14a5d18160375cae23dff025fc90ab68f672329de8f632c84b3ce5912eab9d631d4e7d79a04a04bad71e521fffac9cdc5054346dc5a3932507f872fc39db20f07afcb1653d3a691a1401a724a2b04e218617e0b975f9075f80a2577b58d6030ec83211818473b0b1d;
    5'b11110 : xpb = 1024'h38e5881c61ac89770f53036eeefd9e3ef1f447fa73b909fffece79be45056f4f004d914440d8b4ec600d302cfe612c75965b4c354736c639891a3c1e388d2056efd65abfb0f25af937b109e021c46ad3c927a8250e1e4bda452b6436ae049bad2df3594d54d7c260462e972cae8fd51beb3599382b728602d784c3be06611b60;
    5'b11111 : xpb = 1024'h8176c1fb5d2b2bb1bee908d130b2b783c100f652113bdb96311c94bc3997c0c3c5e49da182cd31d7f85575c250bd3d30dd02673dc666868cedebe000a74c69b1e216c82e16abe5727cb8cf86822b678806cd1a1f0b10b5bd90184414428d484b4ad3d27a2f739b35b19f09a0f55f5a691b1f999d19d038497257ea684e69920e;
    endcase
end

endmodule

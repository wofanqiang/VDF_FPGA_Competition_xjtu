module xpb_5_360
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h25623133aa605d5237dc7303e9fb7a7141feafebfa1bba2cfff615575786868f25c1944a0bf14237f3be2857bfeb534d1a1acc381becff5b70957c22b01f9ee2381f9f6d80c275a604e8898b4b1a4821b6cc3e1d634af5d643d0408ca0f421d3d9b5ed4f4043af0dcbe6b99a2605a79a87a173d250ec0fba0fc196d8ba1a4028;
    5'b00010 : xpb = 1024'h4ac4626754c0baa46fb8e607d3f6f4e283fd5fd7f4377459ffec2aaeaf0d0d1e4b83289417e2846fe77c50af7fd6a69a3435987037d9feb6e12af845603f3dc4703f3edb0184eb4c09d11316963490436d987c3ac695ebac87a0811941e843a7b36bda9e80875e1b97cd73344c0b4f350f42e7a4a1d81f741f832db174348050;
    5'b00011 : xpb = 1024'h7026939aff2117f6a795590bbdf26f53c5fc0fc3ee532e86ffe24006069393ad7144bcde23d3c6a7db3a79073fc1f9e74e5064a853c6fe1251c07468105edca6a85ede48824760f20eb99ca1e14ed8652464ba5829e0e182cb70c1a5e2dc657b8d21c7edc0cb0d2963b42cce7210f6cf96e45b76f2c42f2e2f44c48a2e4ec078;
    5'b00100 : xpb = 1024'h9588c4cea9817548df71cc0fa7ede9c507fabfafe86ee8b3ffd8555d5e1a1a3c970651282fc508dfcef8a15effad4d34686b30e06fb3fd6dc255f08ac07e7b88e07e7db60309d69813a2262d2c692086db30f8758d2bd7590f41023283d0874f66d7b53d010ebc372f9ae66898169e6a1e85cf4943b03ee83f065b62e86900a0;
    5'b00101 : xpb = 1024'ha3db0ac91f39dd24c48c73c818f1ce4d8836c6b0d13026981f1b15f029df3c3b97f67f9718fcc8923588a6fdc3a8fb71e6bd53268ee2c7d824c2d4f35cba5b9a44ee874d43b4ef905f0ad15dea7a4779df83cfa63f0a01e9d84b0c46a9a069111861062908972b774c1b923c64c1fdb574d64394450f1720858773719a0da5d;
    5'b00110 : xpb = 1024'h2f9fe1e03c53fb2484253a406b8a97561a821c57072ebc9681e7c6b65a247a52df40fc437d810ec11716b2c79c25e3043886a16a84db2bd8f2e1a971e5eb449bdc6e87e254fdc49f0ad936a129c1ec9954c47b17c73b95f4e154f1510b8e2864eb3bfdb1d0cd21c540a872bdec51c775deeed80b953d012c181a0e0fd3bb1a85;
    5'b00111 : xpb = 1024'h55021313e6b45876bc01ad44558611c75c80cc43014a76c381dddc0db1ab00e20502908d897250f90ad4db1f5c11365152a16da2a0c82b3463772594960ae37e148e274fd5c03a450fc1c02c74dc34bb0b90b9352a868bcb252531ddac824a38c4f1eb011110d0d30c8f2c5812576f1066904bdde62910e627dba4e88dd55aad;
    5'b01000 : xpb = 1024'h7a6444479114b5c8f3de20483f818c389e7f7c2efb6630f081d3f165093187712ac424d795639330fe9303771bfc899e6cbc39dabcb52a8fd40ca1b7462a82604cadc6bd5682afeb14aa49b7bff67cdcc25cf7528dd181a168f5726a4d766c0c9ea7d85051547fe0d875e5f2385d16aaee31bfb0371520a0379d3bc147ef9ad5;
    5'b01001 : xpb = 1024'h9fc6757b3b75131b2bba934c297d06a9e07e2c1af581eb1d81ca06bc60b80e005085b921a154d568f2512bcedbe7dceb86d70612d8a229eb44a21dd9f64a214284cd662ad74525911992d3430b10c4fe7929356ff11c7777acc5b2f6ee6a8de0785dc59f91982eeea45c9f8c5e62be4575d333828801305a475ed29a0209dafd;
    5'b01010 : xpb = 1024'h147b615923e73ba498918e79031e39c9b106d8d61a2604d303e362be053be78772fecff2e31f991246b114dfb8751f6e3cd7aa64d1dc58fb04985a9e6b974b73489dd0e9a8769df20be15a2bbd4f48ef3bf079f4c7e1403d3b096188d5340d22230c20c52112e56ee98372478c983fb6ae9ac87288a1e2e410b0ee6e3341b4ba;
    5'b01011 : xpb = 1024'h39dd928cce4798f6d06e017ced19b43af30588c21441bf0003d978155cc26e1698c0643cef10db4a3a6f3d37786072bb56f2769cedc95856752dd6c11bb6ea5580bd70572939139810c9e3b708699110f2bcb8122b2c36137ed9a21576282ef5fcc20e146156947cb56a2be1b29de751363c3c44d98df29e20728546ed5bf4e2;
    5'b01100 : xpb = 1024'h5f3fc3c078a7f649084a7480d7152eac350438ae0e5d792d03cf8d6cb448f4a5be81f886fb021d822e2d658f384bc608710d42d509b657b1e5c352e3cbd68937b8dd0fc4a9fb893e15b26d425383d932a988f62f8e772be9c2a9e2a2171c50c9d677fb63a19a438a8150e57bd8a38eebbdddb0172a7a025830341c1fa776350a;
    5'b01101 : xpb = 1024'h84a1f4f42308539b4026e784c110a91d7702e89a0879335a03c5a2c40bcf7b34e4438cd106f35fba21eb8de6f83719558b280f0d25a3570d5658cf067bf62819f0fcaf322abdfee41a9af6cd9e9e21546055344cf1c221c0067a232eb810729db02de8b2e1ddf2984d379f15fea93686457f23e97b6612123ff5b2f861907532;
    5'b01110 : xpb = 1024'haa042627cd68b0ed78035a88ab0c238eb90198860294ed8703bbb81b635601c40a05211b12e4a1f215a9b63eb8226ca2a542db4541905668c6ee4b292c15c6fc291c4e9fab80748a1f838058e9b869761721726a550d17964a4a63bb5904947189e3d6022221a1a6191e58b024aede20cd2097bbcc5221cc4fb749d11baab55a;
    5'b01111 : xpb = 1024'h1eb91205b5dad976e4da55b584ad56ae898a45412739073c85d5141d07d9db4b2c7e37ec54af659b6a099f4f94afaf255b437f973aca857886e487eda162f12cececb95e7cb1eceb11d207419bf6ed66d9e8b6ef2bd1e05bd88e124d3fce13b334923127b19c58265e452b6b52e45f9205e82cabccf2d456190965a54ce28f17;
    5'b10000 : xpb = 1024'h441b4339603b36c91cb6c8b96ea8d11fcb88f52d2154c16985cb29745f6061da523fcc3660a0a7d35dc7c7a7549b0272755e4bcf56b784d3f77a04105182900f250c58cbfd74629116ba90cce711358890b4f50c8f1cd6321c5e52d9e0c235870e481e76f1e007342a2be50578ea072c8d89a07e1ddee41028cafc7e06fccf3f;
    5'b10001 : xpb = 1024'h697d746d0a9b941b54933bbd58a44b910d87a5191b707b9685c13ecbb6e6e869780160806c91ea0b5185efff148655bf8f79180772a4842f680f803301a22ef15d2bf8397e36d8371ba31a58322b7daa47813329f267cc08602e936681b6575ae7fe0bc63223b641f6129e9f9eefaec7152b14506ecaf3ca388c9356c1170f67;
    5'b10010 : xpb = 1024'h8edfa5a0b4fbf16d8c6faec1429fc6024f865505158c35c385b754230e6d6ef89dc2f4ca78832c4345441856d471a90ca993e43f8e91838ad8a4fc55b1c1cdd3954b97a6fef94ddd208ba3e37d45c5cbfe4d714755b2c1dea3fed3f322aa792ec1b3f9157267654fc1f95839c4f556619ccc8822bfb70384484e2a2f7b314f8f;
    5'b10011 : xpb = 1024'h394917e9d6e19f6f946a9ee1c40f922200f01c03a304f7907d0b024b2f1487fc03c0b9bba4defec99a40167b0feeb8f5f94889187cbb29a989b391a270ef804591c0265d02ac63e12da2acc2f8449bcc114b5cc2c778aa4324282850973f8706c62543b01e21bd007202af4f32ad7d2d5941d12c057b60e11a04603ac69294c;
    5'b10100 : xpb = 1024'h28f6c2b247ce774931231cf2063c7393620db1ac344c09a607c6c57c0a77cf0ee5fd9fe5c63f32248d6229bf70ea3edc79af54c9a3b8b1f60930b53cd72e96e6913ba1d350ed3be417c2b4577a9e91de77e0f3e98fc2807a7612c311aa681a444618418a4225caddd306e48f19307f6d5d3590e51143c5c82161dcdc66836974;
    5'b10101 : xpb = 1024'h4e58f3e5f22ed49b68ff8ff5f037ee04a40c61982e67c3d307bcdad361fe559e0bbf342fd230745c8120521730d5922993ca2101bfa5b15179c6315f874e35c8c95b4140d1afb18a1cab3de2c5b8da002ead3206f30d7650b9e3039e4b5c3c181fce2ed9826979eb9eed9e293f362707e4d704b7622fd582312373b5209da99c;
    5'b10110 : xpb = 1024'h73bb25199c8f31eda0dc02f9da336875e60b118428837e0007b2f02ab984dc2d3180c879de21b69474de7a6ef0c0e576ade4ed39db92b0acea5bad82376dd4ab017ae0ae527227302193c76e10d32221e579702456586c26fdb3442aec505debf9841c28c2ad28f96ad457c3653bcea26c787889b31be53c40e50a8ddab7e9c4;
    5'b10111 : xpb = 1024'h991d564d46ef8f3fd8b875fdc42ee2e72809c170229f382d07a90582110b62bc57425cc3ea12f8cc689ca2c6b0ac38c3c7ffb971f77fb0085af129a4e78d738d399a801bd3349cd6267c50f95bed6a439c45ae41b9a361fd418384b78d447fbfd33a097802f0d80736bb115d8b41763cf419ec5c0407f4f650a6a16694d229ec;
    5'b11000 : xpb = 1024'hdd2422b2f61b7c9458f712a9dd01606f8926e2b474351e289c26183b58f3c4379bb73952bddbc75bcfc8bd78d397b467e005dc3f0b9df181ae766695cda9dbdfd6aeadaa466153718cad7e20e2bee345f0cf2c690682ac2cfc73349740dff017de8649d926b8e877be1e418b976f7ae2ce1814c04a8a78019f8bd3ac60a03a9;
    5'b11001 : xpb = 1024'h3334735ed9c2151b7d6be42e87cb90783a911e17415f0c0f89b876db0d15c2d29f7d07df37cefeadb0bab42f4d24ce93981b29fc0ca6de738b7ce28c0cfa3ca0358a8a4825288add1db3616d5946365615d930e3f3b32099139773d6150220d5579e51ecd2af3d9547c89db2df7c9f48b482f51e5594b73a29ba5413802443d1;
    5'b11010 : xpb = 1024'h5896a4928422726db548573271c70ae97c8fce033b7ac63c89ae8c32649c4961c53e9c2943c040e5a478dc870d1021e0b235f6342893ddcefc125eaebd19db826daa29b5a5eb0083229beaf8a4607e77cca56f0156fe166f5767b462b5f642a931543f3c12f2eca313af574d058246e33c2468f0a680c6f4397beaec3a3e83f9;
    5'b11011 : xpb = 1024'h7df8d5c62e82cfbfed24ca365bc2855abe8e7def3596806989a4a189bc22cff0eb0030734fb1831d983704deccfb752dcc50c26c4480dd2a6ca7dad16d397a64a5c9c92326ad762927847483ef7ac6998371ad1eba490c459b37f4ef56ea647d0b0a2c8b53369bb0df9610e72b87ee7dc3c5dcc2f76cd6ae493d81c4f458c421;
    5'b11100 : xpb = 1024'ha35b06f9d8e32d1225013d3a45bdffcc008d2ddb2fb23a96899ab6e113a9568010c1c4bd5ba2c5558bf52d368ce6c87ae66b8ea4606ddc85dd3d56f41d591946dde96890a76febcf2c6cfe0f3a950ebb3a3deb3c1d94021bdf08357bf7de8650e4c019da937a4abeab7cca81518d96184b6750954858e66858ff189dae730449;
    5'b11101 : xpb = 1024'h180ff2d7c155559b91d838671f5f32ebd115da965456544c0bb412e2b82d3007333adb8e9d6d88fee055164769740afd9c6c32f659a80b959d3393b892a64377a1b9d34f78a164301ebb84f7ecd392abfd052fc0f458cae16d4be40ddea805928f6e750022f5013ef0a39d3c7fc31789842ee58548f998f222513471dfaade06;
    5'b11110 : xpb = 1024'h3d72240b6bb5b2edc9b4ab6b095aad5d13148a824e720e790baa283a0fb3b69658fc6fd8a95ecb36d4133e9f295f5e4ab686ff2e75950af10dc90fdb42c5e259d9d972bcf963d9d623a40e8337eddacdb3d16dde57a3c0b7b11c249a7f9c27666924624f6338b04cbc8a56d6a5c8bf240bd0595799e5a8ac3212cb4a99c51e2e;
    5'b11111 : xpb = 1024'h62d4553f1616104001911e6ef35627ce55133a6e488dc8a60ba03d91673a3d257ebe0422b5500d6ec7d166f6e94ab197d0a1cb6691820a4c7e5e8bfdf2e5813c11f9122a7a264f7c288c980e830822ef6a9dabfbbaeeb68df4ec65272090493a42da4f9ea37c5f5a88711070cbce66be9371cd29ead1b86641d4622353df5e56;
    endcase
end

endmodule

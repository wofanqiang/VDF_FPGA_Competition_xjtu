module xpb_2048
(
    input [1023:0] data_in0, 
    input [1023:0] data_in1, 

    output [1023:0] data_out_0,
    output [1023:0] data_out_1,
    output [1023:0] data_out_2,
    output [1023:0] data_out_3,
    output [1023:0] data_out_4,
    output [1023:0] data_out_5,
    output [1023:0] data_out_6,
    output [1023:0] data_out_7,
    output [1023:0] data_out_8,
    output [1023:0] data_out_9,
    output [1023:0] data_out_10,
    output [1023:0] data_out_11,
    output [1023:0] data_out_12,
    output [1023:0] data_out_13,
    output [1023:0] data_out_14,
    output [1023:0] data_out_15,
    output [1023:0] data_out_16,
    output [1023:0] data_out_17,
    output [1023:0] data_out_18,
    output [1023:0] data_out_19,
    output [1023:0] data_out_20,
    output [1023:0] data_out_21,
    output [1023:0] data_out_22,
    output [1023:0] data_out_23,
    output [1023:0] data_out_24,
    output [1023:0] data_out_25,
    output [1023:0] data_out_26,
    output [1023:0] data_out_27,
    output [1023:0] data_out_28,
    output [1023:0] data_out_29,
    output [1023:0] data_out_30,
    output [1023:0] data_out_31,
    output [1023:0] data_out_32,
    output [1023:0] data_out_33,
    output [1023:0] data_out_34,
    output [1023:0] data_out_35,
    output [1023:0] data_out_36,
    output [1023:0] data_out_37,
    output [1023:0] data_out_38,
    output [1023:0] data_out_39,
    output [1023:0] data_out_40,
    output [1023:0] data_out_41,
    output [1023:0] data_out_42,
    output [1023:0] data_out_43,
    output [1023:0] data_out_44,
    output [1023:0] data_out_45,
    output [1023:0] data_out_46,
    output [1023:0] data_out_47,
    output [1023:0] data_out_48,
    output [1023:0] data_out_49,
    output [1023:0] data_out_50,
    output [1023:0] data_out_51,
    output [1023:0] data_out_52,
    output [1023:0] data_out_53,
    output [1023:0] data_out_54,
    output [1023:0] data_out_55,
    output [1023:0] data_out_56,
    output [1023:0] data_out_57,
    output [1023:0] data_out_58,
    output [1023:0] data_out_59,
    output [1023:0] data_out_60,
    output [1023:0] data_out_61,
    output [1023:0] data_out_62,
    output [1023:0] data_out_63,
    output [1023:0] data_out_64,
    output [1023:0] data_out_65,
    output [1023:0] data_out_66,
    output [1023:0] data_out_67,
    output [1023:0] data_out_68,
    output [1023:0] data_out_69,
    output [1023:0] data_out_70,
    output [1023:0] data_out_71,
    output [1023:0] data_out_72,
    output [1023:0] data_out_73,
    output [1023:0] data_out_74,
    output [1023:0] data_out_75,
    output [1023:0] data_out_76,
    output [1023:0] data_out_77,
    output [1023:0] data_out_78,
    output [1023:0] data_out_79,
    output [1023:0] data_out_80,
    output [1023:0] data_out_81,
    output [1023:0] data_out_82,
    output [1023:0] data_out_83,
    output [1023:0] data_out_84,
    output [1023:0] data_out_85,
    output [1023:0] data_out_86,
    output [1023:0] data_out_87,
    output [1023:0] data_out_88,
    output [1023:0] data_out_89,
    output [1023:0] data_out_90,
    output [1023:0] data_out_91,
    output [1023:0] data_out_92,
    output [1023:0] data_out_93,
    output [1023:0] data_out_94,
    output [1023:0] data_out_95,
    output [1023:0] data_out_96,
    output [1023:0] data_out_97,
    output [1023:0] data_out_98,
    output [1023:0] data_out_99,
    output [1023:0] data_out_100,
    output [1023:0] data_out_101,
    output [1023:0] data_out_102,
    output [1023:0] data_out_103,
    output [1023:0] data_out_104,
    output [1023:0] data_out_105,
    output [1023:0] data_out_106,
    output [1023:0] data_out_107,
    output [1023:0] data_out_108,
    output [1023:0] data_out_109,
    output [1023:0] data_out_110,
    output [1023:0] data_out_111,
    output [1023:0] data_out_112,
    output [1023:0] data_out_113,
    output [1023:0] data_out_114,
    output [1023:0] data_out_115,
    output [1023:0] data_out_116,
    output [1023:0] data_out_117,
    output [1023:0] data_out_118,
    output [1023:0] data_out_119,
    output [1023:0] data_out_120,
    output [1023:0] data_out_121,
    output [1023:0] data_out_122,
    output [1023:0] data_out_123,
    output [1023:0] data_out_124,
    output [1023:0] data_out_125,
    output [1023:0] data_out_126,
    output [1023:0] data_out_127,
    output [1023:0] data_out_128,
    output [1023:0] data_out_129,
    output [1023:0] data_out_130,
    output [1023:0] data_out_131,
    output [1023:0] data_out_132,
    output [1023:0] data_out_133,
    output [1023:0] data_out_134,
    output [1023:0] data_out_135,
    output [1023:0] data_out_136,
    output [1023:0] data_out_137,
    output [1023:0] data_out_138,
    output [1023:0] data_out_139,
    output [1023:0] data_out_140,
    output [1023:0] data_out_141,
    output [1023:0] data_out_142,
    output [1023:0] data_out_143,
    output [1023:0] data_out_144,
    output [1023:0] data_out_145,
    output [1023:0] data_out_146,
    output [1023:0] data_out_147,
    output [1023:0] data_out_148,
    output [1023:0] data_out_149,
    output [1023:0] data_out_150,
    output [1023:0] data_out_151,
    output [1023:0] data_out_152,
    output [1023:0] data_out_153,
    output [1023:0] data_out_154,
    output [1023:0] data_out_155,
    output [1023:0] data_out_156,
    output [1023:0] data_out_157,
    output [1023:0] data_out_158,
    output [1023:0] data_out_159,
    output [1023:0] data_out_160,
    output [1023:0] data_out_161,
    output [1023:0] data_out_162,
    output [1023:0] data_out_163,
    output [1023:0] data_out_164,
    output [1023:0] data_out_165,
    output [1023:0] data_out_166,
    output [1023:0] data_out_167,
    output [1023:0] data_out_168,
    output [1023:0] data_out_169,
    output [1023:0] data_out_170,
    output [1023:0] data_out_171,
    output [1023:0] data_out_172,
    output [1023:0] data_out_173,
    output [1023:0] data_out_174,
    output [1023:0] data_out_175,
    output [1023:0] data_out_176,
    output [1023:0] data_out_177,
    output [1023:0] data_out_178,
    output [1023:0] data_out_179,
    output [1023:0] data_out_180,
    output [1023:0] data_out_181,
    output [1023:0] data_out_182,
    output [1023:0] data_out_183,
    output [1023:0] data_out_184,
    output [1023:0] data_out_185,
    output [1023:0] data_out_186,
    output [1023:0] data_out_187,
    output [1023:0] data_out_188,
    output [1023:0] data_out_189,
    output [1023:0] data_out_190,
    output [1023:0] data_out_191,
    output [1023:0] data_out_192,
    output [1023:0] data_out_193,
    output [1023:0] data_out_194,
    output [1023:0] data_out_195,
    output [1023:0] data_out_196,
    output [1023:0] data_out_197,
    output [1023:0] data_out_198,
    output [1023:0] data_out_199,
    output [1023:0] data_out_200,
    output [1023:0] data_out_201,
    output [1023:0] data_out_202,
    output [1023:0] data_out_203,
    output [1023:0] data_out_204,
    output [1023:0] data_out_205,
    output [1023:0] data_out_206,
    output [1023:0] data_out_207,
    output [1023:0] data_out_208,
    output [1023:0] data_out_209,
    output [1023:0] data_out_210,
    output [1023:0] data_out_211,
    output [1023:0] data_out_212,
    output [1023:0] data_out_213,
    output [1023:0] data_out_214,
    output [1023:0] data_out_215,
    output [1023:0] data_out_216,
    output [1023:0] data_out_217,
    output [1023:0] data_out_218,
    output [1023:0] data_out_219,
    output [1023:0] data_out_220,
    output [1023:0] data_out_221,
    output [1023:0] data_out_222,
    output [1023:0] data_out_223,
    output [1023:0] data_out_224,
    output [1023:0] data_out_225,
    output [1023:0] data_out_226,
    output [1023:0] data_out_227,
    output [1023:0] data_out_228,
    output [1023:0] data_out_229,
    output [1023:0] data_out_230,
    output [1023:0] data_out_231,
    output [1023:0] data_out_232,
    output [1023:0] data_out_233,
    output [1023:0] data_out_234,
    output [1023:0] data_out_235,
    output [1023:0] data_out_236,
    output [1023:0] data_out_237,
    output [1023:0] data_out_238,
    output [1023:0] data_out_239,
    output [1023:0] data_out_240,
    output [1023:0] data_out_241,
    output [1023:0] data_out_242,
    output [1023:0] data_out_243,
    output [1023:0] data_out_244,
    output [1023:0] data_out_245,
    output [1023:0] data_out_246,
    output [1023:0] data_out_247,
    output [1023:0] data_out_248,
    output [1023:0] data_out_249,
    output [1023:0] data_out_250,
    output [1023:0] data_out_251,
    output [1023:0] data_out_252,
    output [1023:0] data_out_253,
    output [1023:0] data_out_254,
    output [1023:0] data_out_255,
    output [1023:0] data_out_256,
    output [1023:0] data_out_257,
    output [1023:0] data_out_258,
    output [1023:0] data_out_259,
    output [1023:0] data_out_260,
    output [1023:0] data_out_261,
    output [1023:0] data_out_262,
    output [1023:0] data_out_263,
    output [1023:0] data_out_264,
    output [1023:0] data_out_265,
    output [1023:0] data_out_266,
    output [1023:0] data_out_267,
    output [1023:0] data_out_268,
    output [1023:0] data_out_269,
    output [1023:0] data_out_270,
    output [1023:0] data_out_271,
    output [1023:0] data_out_272,
    output [1023:0] data_out_273,
    output [1023:0] data_out_274,
    output [1023:0] data_out_275,
    output [1023:0] data_out_276,
    output [1023:0] data_out_277,
    output [1023:0] data_out_278,
    output [1023:0] data_out_279,
    output [1023:0] data_out_280,
    output [1023:0] data_out_281,
    output [1023:0] data_out_282,
    output [1023:0] data_out_283,
    output [1023:0] data_out_284,
    output [1023:0] data_out_285,
    output [1023:0] data_out_286,
    output [1023:0] data_out_287,
    output [1023:0] data_out_288,
    output [1023:0] data_out_289,
    output [1023:0] data_out_290,
    output [1023:0] data_out_291,
    output [1023:0] data_out_292,
    output [1023:0] data_out_293,
    output [1023:0] data_out_294,
    output [1023:0] data_out_295,
    output [1023:0] data_out_296,
    output [1023:0] data_out_297,
    output [1023:0] data_out_298,
    output [1023:0] data_out_299,
    output [1023:0] data_out_300,
    output [1023:0] data_out_301,
    output [1023:0] data_out_302,
    output [1023:0] data_out_303,
    output [1023:0] data_out_304,
    output [1023:0] data_out_305,
    output [1023:0] data_out_306,
    output [1023:0] data_out_307,
    output [1023:0] data_out_308,
    output [1023:0] data_out_309,
    output [1023:0] data_out_310,
    output [1023:0] data_out_311,
    output [1023:0] data_out_312,
    output [1023:0] data_out_313,
    output [1023:0] data_out_314,
    output [1023:0] data_out_315,
    output [1023:0] data_out_316,
    output [1023:0] data_out_317,
    output [1023:0] data_out_318,
    output [1023:0] data_out_319,
    output [1023:0] data_out_320,
    output [1023:0] data_out_321,
    output [1023:0] data_out_322,
    output [1023:0] data_out_323,
    output [1023:0] data_out_324,
    output [1023:0] data_out_325,
    output [1023:0] data_out_326,
    output [1023:0] data_out_327,
    output [1023:0] data_out_328,
    output [1023:0] data_out_329,
    output [1023:0] data_out_330,
    output [1023:0] data_out_331,
    output [1023:0] data_out_332,
    output [1023:0] data_out_333,
    output [1023:0] data_out_334,
    output [1023:0] data_out_335,
    output [1023:0] data_out_336,
    output [1023:0] data_out_337,
    output [1023:0] data_out_338,
    output [1023:0] data_out_339,
    output [1023:0] data_out_340,
    output [1023:0] data_out_341,
    output [1023:0] data_out_342,
    output [1023:0] data_out_343,
    output [1023:0] data_out_344,
    output [1023:0] data_out_345,
    output [1023:0] data_out_346,
    output [1023:0] data_out_347,
    output [1023:0] data_out_348,
    output [1023:0] data_out_349,
    output [1023:0] data_out_350,
    output [1023:0] data_out_351,
    output [1023:0] data_out_352,
    output [1023:0] data_out_353,
    output [1023:0] data_out_354,
    output [1023:0] data_out_355,
    output [1023:0] data_out_356,
    output [1023:0] data_out_357,
    output [1023:0] data_out_358,
    output [1023:0] data_out_359,
    output [1023:0] data_out_360,
    output [1023:0] data_out_361,
    output [1023:0] data_out_362,
    output [1023:0] data_out_363,
    output [1023:0] data_out_364,
    output [1023:0] data_out_365,
    output [1023:0] data_out_366,
    output [1023:0] data_out_367,
    output [1023:0] data_out_368,
    output [1023:0] data_out_369,
    output [1023:0] data_out_370,
    output [1023:0] data_out_371,
    output [1023:0] data_out_372,
    output [1023:0] data_out_373,
    output [1023:0] data_out_374,
    output [1023:0] data_out_375,
    output [1023:0] data_out_376,
    output [1023:0] data_out_377,
    output [1023:0] data_out_378,
    output [1023:0] data_out_379,
    output [1023:0] data_out_380,
    output [1023:0] data_out_381,
    output [1023:0] data_out_382,
    output [1023:0] data_out_383,
    output [1023:0] data_out_384,
    output [1023:0] data_out_385,
    output [1023:0] data_out_386,
    output [1023:0] data_out_387,
    output [1023:0] data_out_388,
    output [1023:0] data_out_389,
    output [1023:0] data_out_390,
    output [1023:0] data_out_391,
    output [1023:0] data_out_392,
    output [1023:0] data_out_393,
    output [1023:0] data_out_394,
    output [1023:0] data_out_395,
    output [1023:0] data_out_396,
    output [1023:0] data_out_397,
    output [1023:0] data_out_398,
    output [1023:0] data_out_399,
    output [1023:0] data_out_400,
    output [1023:0] data_out_401,
    output [1023:0] data_out_402,
    output [1023:0] data_out_403,
    output [1023:0] data_out_404,
    output [1023:0] data_out_405,
    output [1023:0] data_out_406,
    output [1023:0] data_out_407,
    output [1023:0] data_out_408,
    output [1023:0] data_out_409


);




xpb_1024 u0_xpb_1024(
.data_in(data_in0),


.data_out_0(data_out_0),
.data_out_1(data_out_1),
.data_out_2(data_out_2),
.data_out_3(data_out_3),
.data_out_4(data_out_4),
.data_out_5(data_out_5),
.data_out_6(data_out_6),
.data_out_7(data_out_7),
.data_out_8(data_out_8),
.data_out_9(data_out_9),
.data_out_10(data_out_10),
.data_out_11(data_out_11),
.data_out_12(data_out_12),
.data_out_13(data_out_13),
.data_out_14(data_out_14),
.data_out_15(data_out_15),
.data_out_16(data_out_16),
.data_out_17(data_out_17),
.data_out_18(data_out_18),
.data_out_19(data_out_19),
.data_out_20(data_out_20),
.data_out_21(data_out_21),
.data_out_22(data_out_22),
.data_out_23(data_out_23),
.data_out_24(data_out_24),
.data_out_25(data_out_25),
.data_out_26(data_out_26),
.data_out_27(data_out_27),
.data_out_28(data_out_28),
.data_out_29(data_out_29),
.data_out_30(data_out_30),
.data_out_31(data_out_31),
.data_out_32(data_out_32),
.data_out_33(data_out_33),
.data_out_34(data_out_34),
.data_out_35(data_out_35),
.data_out_36(data_out_36),
.data_out_37(data_out_37),
.data_out_38(data_out_38),
.data_out_39(data_out_39),
.data_out_40(data_out_40),
.data_out_41(data_out_41),
.data_out_42(data_out_42),
.data_out_43(data_out_43),
.data_out_44(data_out_44),
.data_out_45(data_out_45),
.data_out_46(data_out_46),
.data_out_47(data_out_47),
.data_out_48(data_out_48),
.data_out_49(data_out_49),
.data_out_50(data_out_50),
.data_out_51(data_out_51),
.data_out_52(data_out_52),
.data_out_53(data_out_53),
.data_out_54(data_out_54),
.data_out_55(data_out_55),
.data_out_56(data_out_56),
.data_out_57(data_out_57),
.data_out_58(data_out_58),
.data_out_59(data_out_59),
.data_out_60(data_out_60),
.data_out_61(data_out_61),
.data_out_62(data_out_62),
.data_out_63(data_out_63),
.data_out_64(data_out_64),
.data_out_65(data_out_65),
.data_out_66(data_out_66),
.data_out_67(data_out_67),
.data_out_68(data_out_68),
.data_out_69(data_out_69),
.data_out_70(data_out_70),
.data_out_71(data_out_71),
.data_out_72(data_out_72),
.data_out_73(data_out_73),
.data_out_74(data_out_74),
.data_out_75(data_out_75),
.data_out_76(data_out_76),
.data_out_77(data_out_77),
.data_out_78(data_out_78),
.data_out_79(data_out_79),
.data_out_80(data_out_80),
.data_out_81(data_out_81),
.data_out_82(data_out_82),
.data_out_83(data_out_83),
.data_out_84(data_out_84),
.data_out_85(data_out_85),
.data_out_86(data_out_86),
.data_out_87(data_out_87),
.data_out_88(data_out_88),
.data_out_89(data_out_89),
.data_out_90(data_out_90),
.data_out_91(data_out_91),
.data_out_92(data_out_92),
.data_out_93(data_out_93),
.data_out_94(data_out_94),
.data_out_95(data_out_95),
.data_out_96(data_out_96),
.data_out_97(data_out_97),
.data_out_98(data_out_98),
.data_out_99(data_out_99),
.data_out_100(data_out_100),
.data_out_101(data_out_101),
.data_out_102(data_out_102),
.data_out_103(data_out_103),
.data_out_104(data_out_104),
.data_out_105(data_out_105),
.data_out_106(data_out_106),
.data_out_107(data_out_107),
.data_out_108(data_out_108),
.data_out_109(data_out_109),
.data_out_110(data_out_110),
.data_out_111(data_out_111),
.data_out_112(data_out_112),
.data_out_113(data_out_113),
.data_out_114(data_out_114),
.data_out_115(data_out_115),
.data_out_116(data_out_116),
.data_out_117(data_out_117),
.data_out_118(data_out_118),
.data_out_119(data_out_119),
.data_out_120(data_out_120),
.data_out_121(data_out_121),
.data_out_122(data_out_122),
.data_out_123(data_out_123),
.data_out_124(data_out_124),
.data_out_125(data_out_125),
.data_out_126(data_out_126),
.data_out_127(data_out_127),
.data_out_128(data_out_128),
.data_out_129(data_out_129),
.data_out_130(data_out_130),
.data_out_131(data_out_131),
.data_out_132(data_out_132),
.data_out_133(data_out_133),
.data_out_134(data_out_134),
.data_out_135(data_out_135),
.data_out_136(data_out_136),
.data_out_137(data_out_137),
.data_out_138(data_out_138),
.data_out_139(data_out_139),
.data_out_140(data_out_140),
.data_out_141(data_out_141),
.data_out_142(data_out_142),
.data_out_143(data_out_143),
.data_out_144(data_out_144),
.data_out_145(data_out_145),
.data_out_146(data_out_146),
.data_out_147(data_out_147),
.data_out_148(data_out_148),
.data_out_149(data_out_149),
.data_out_150(data_out_150),
.data_out_151(data_out_151),
.data_out_152(data_out_152),
.data_out_153(data_out_153),
.data_out_154(data_out_154),
.data_out_155(data_out_155),
.data_out_156(data_out_156),
.data_out_157(data_out_157),
.data_out_158(data_out_158),
.data_out_159(data_out_159),
.data_out_160(data_out_160),
.data_out_161(data_out_161),
.data_out_162(data_out_162),
.data_out_163(data_out_163),
.data_out_164(data_out_164),
.data_out_165(data_out_165),
.data_out_166(data_out_166),
.data_out_167(data_out_167),
.data_out_168(data_out_168),
.data_out_169(data_out_169),
.data_out_170(data_out_170),
.data_out_171(data_out_171),
.data_out_172(data_out_172),
.data_out_173(data_out_173),
.data_out_174(data_out_174),
.data_out_175(data_out_175),
.data_out_176(data_out_176),
.data_out_177(data_out_177),
.data_out_178(data_out_178),
.data_out_179(data_out_179),
.data_out_180(data_out_180),
.data_out_181(data_out_181),
.data_out_182(data_out_182),
.data_out_183(data_out_183),
.data_out_184(data_out_184),
.data_out_185(data_out_185),
.data_out_186(data_out_186),
.data_out_187(data_out_187),
.data_out_188(data_out_188),
.data_out_189(data_out_189),
.data_out_190(data_out_190),
.data_out_191(data_out_191),
.data_out_192(data_out_192),
.data_out_193(data_out_193),
.data_out_194(data_out_194),
.data_out_195(data_out_195),
.data_out_196(data_out_196),
.data_out_197(data_out_197),
.data_out_198(data_out_198),
.data_out_199(data_out_199),
.data_out_200(data_out_200),
.data_out_201(data_out_201),
.data_out_202(data_out_202),
.data_out_203(data_out_203),
.data_out_204(data_out_204)

);

xpb_1024 u1_xpb_1024(
.data_in(data_in1),


.data_out_0(data_out_205),
.data_out_1(data_out_206),
.data_out_2(data_out_207),
.data_out_3(data_out_208),
.data_out_4(data_out_209),
.data_out_5(data_out_210),
.data_out_6(data_out_211),
.data_out_7(data_out_212),
.data_out_8(data_out_213),
.data_out_9(data_out_214),
.data_out_10(data_out_215),
.data_out_11(data_out_216),
.data_out_12(data_out_217),
.data_out_13(data_out_218),
.data_out_14(data_out_219),
.data_out_15(data_out_220),
.data_out_16(data_out_221),
.data_out_17(data_out_222),
.data_out_18(data_out_223),
.data_out_19(data_out_224),
.data_out_20(data_out_225),
.data_out_21(data_out_226),
.data_out_22(data_out_227),
.data_out_23(data_out_228),
.data_out_24(data_out_229),
.data_out_25(data_out_230),
.data_out_26(data_out_231),
.data_out_27(data_out_232),
.data_out_28(data_out_233),
.data_out_29(data_out_234),
.data_out_30(data_out_235),
.data_out_31(data_out_236),
.data_out_32(data_out_237),
.data_out_33(data_out_238),
.data_out_34(data_out_239),
.data_out_35(data_out_240),
.data_out_36(data_out_241),
.data_out_37(data_out_242),
.data_out_38(data_out_243),
.data_out_39(data_out_244),
.data_out_40(data_out_245),
.data_out_41(data_out_246),
.data_out_42(data_out_247),
.data_out_43(data_out_248),
.data_out_44(data_out_249),
.data_out_45(data_out_250),
.data_out_46(data_out_251),
.data_out_47(data_out_252),
.data_out_48(data_out_253),
.data_out_49(data_out_254),
.data_out_50(data_out_255),
.data_out_51(data_out_256),
.data_out_52(data_out_257),
.data_out_53(data_out_258),
.data_out_54(data_out_259),
.data_out_55(data_out_260),
.data_out_56(data_out_261),
.data_out_57(data_out_262),
.data_out_58(data_out_263),
.data_out_59(data_out_264),
.data_out_60(data_out_265),
.data_out_61(data_out_266),
.data_out_62(data_out_267),
.data_out_63(data_out_268),
.data_out_64(data_out_269),
.data_out_65(data_out_270),
.data_out_66(data_out_271),
.data_out_67(data_out_272),
.data_out_68(data_out_273),
.data_out_69(data_out_274),
.data_out_70(data_out_275),
.data_out_71(data_out_276),
.data_out_72(data_out_277),
.data_out_73(data_out_278),
.data_out_74(data_out_279),
.data_out_75(data_out_280),
.data_out_76(data_out_281),
.data_out_77(data_out_282),
.data_out_78(data_out_283),
.data_out_79(data_out_284),
.data_out_80(data_out_285),
.data_out_81(data_out_286),
.data_out_82(data_out_287),
.data_out_83(data_out_288),
.data_out_84(data_out_289),
.data_out_85(data_out_290),
.data_out_86(data_out_291),
.data_out_87(data_out_292),
.data_out_88(data_out_293),
.data_out_89(data_out_294),
.data_out_90(data_out_295),
.data_out_91(data_out_296),
.data_out_92(data_out_297),
.data_out_93(data_out_298),
.data_out_94(data_out_299),
.data_out_95(data_out_300),
.data_out_96(data_out_301),
.data_out_97(data_out_302),
.data_out_98(data_out_303),
.data_out_99(data_out_304),
.data_out_100(data_out_305),
.data_out_101(data_out_306),
.data_out_102(data_out_307),
.data_out_103(data_out_308),
.data_out_104(data_out_309),
.data_out_105(data_out_310),
.data_out_106(data_out_311),
.data_out_107(data_out_312),
.data_out_108(data_out_313),
.data_out_109(data_out_314),
.data_out_110(data_out_315),
.data_out_111(data_out_316),
.data_out_112(data_out_317),
.data_out_113(data_out_318),
.data_out_114(data_out_319),
.data_out_115(data_out_320),
.data_out_116(data_out_321),
.data_out_117(data_out_322),
.data_out_118(data_out_323),
.data_out_119(data_out_324),
.data_out_120(data_out_325),
.data_out_121(data_out_326),
.data_out_122(data_out_327),
.data_out_123(data_out_328),
.data_out_124(data_out_329),
.data_out_125(data_out_330),
.data_out_126(data_out_331),
.data_out_127(data_out_332),
.data_out_128(data_out_333),
.data_out_129(data_out_334),
.data_out_130(data_out_335),
.data_out_131(data_out_336),
.data_out_132(data_out_337),
.data_out_133(data_out_338),
.data_out_134(data_out_339),
.data_out_135(data_out_340),
.data_out_136(data_out_341),
.data_out_137(data_out_342),
.data_out_138(data_out_343),
.data_out_139(data_out_344),
.data_out_140(data_out_345),
.data_out_141(data_out_346),
.data_out_142(data_out_347),
.data_out_143(data_out_348),
.data_out_144(data_out_349),
.data_out_145(data_out_350),
.data_out_146(data_out_351),
.data_out_147(data_out_352),
.data_out_148(data_out_353),
.data_out_149(data_out_354),
.data_out_150(data_out_355),
.data_out_151(data_out_356),
.data_out_152(data_out_357),
.data_out_153(data_out_358),
.data_out_154(data_out_359),
.data_out_155(data_out_360),
.data_out_156(data_out_361),
.data_out_157(data_out_362),
.data_out_158(data_out_363),
.data_out_159(data_out_364),
.data_out_160(data_out_365),
.data_out_161(data_out_366),
.data_out_162(data_out_367),
.data_out_163(data_out_368),
.data_out_164(data_out_369),
.data_out_165(data_out_370),
.data_out_166(data_out_371),
.data_out_167(data_out_372),
.data_out_168(data_out_373),
.data_out_169(data_out_374),
.data_out_170(data_out_375),
.data_out_171(data_out_376),
.data_out_172(data_out_377),
.data_out_173(data_out_378),
.data_out_174(data_out_379),
.data_out_175(data_out_380),
.data_out_176(data_out_381),
.data_out_177(data_out_382),
.data_out_178(data_out_383),
.data_out_179(data_out_384),
.data_out_180(data_out_385),
.data_out_181(data_out_386),
.data_out_182(data_out_387),
.data_out_183(data_out_388),
.data_out_184(data_out_389),
.data_out_185(data_out_390),
.data_out_186(data_out_391),
.data_out_187(data_out_392),
.data_out_188(data_out_393),
.data_out_189(data_out_394),
.data_out_190(data_out_395),
.data_out_191(data_out_396),
.data_out_192(data_out_397),
.data_out_193(data_out_398),
.data_out_194(data_out_399),
.data_out_195(data_out_400),
.data_out_196(data_out_401),
.data_out_197(data_out_402),
.data_out_198(data_out_403),
.data_out_199(data_out_404),
.data_out_200(data_out_405),
.data_out_201(data_out_406),
.data_out_202(data_out_407),
.data_out_203(data_out_408),
.data_out_204(data_out_409)

);


endmodule
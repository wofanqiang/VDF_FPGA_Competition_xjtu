module xpb_264
(
    input [263:0] data_in,

    output [1023:0] data_out_0,
    output [1023:0] data_out_1,
    output [1023:0] data_out_2,
    output [1023:0] data_out_3,
    output [1023:0] data_out_4,
    output [1023:0] data_out_5,
    output [1023:0] data_out_6,
    output [1023:0] data_out_7,
    output [1023:0] data_out_8,
    output [1023:0] data_out_9,
    output [1023:0] data_out_10,
    output [1023:0] data_out_11,
    output [1023:0] data_out_12,
    output [1023:0] data_out_13,
    output [1023:0] data_out_14,
    output [1023:0] data_out_15,
    output [1023:0] data_out_16,
    output [1023:0] data_out_17,
    output [1023:0] data_out_18,
    output [1023:0] data_out_19,
    output [1023:0] data_out_20,
    output [1023:0] data_out_21,
    output [1023:0] data_out_22,
    output [1023:0] data_out_23,
    output [1023:0] data_out_24,
    output [1023:0] data_out_25,
    output [1023:0] data_out_26,
    output [1023:0] data_out_27,
    output [1023:0] data_out_28,
    output [1023:0] data_out_29,
    output [1023:0] data_out_30,
    output [1023:0] data_out_31,
    output [1023:0] data_out_32,
    output [1023:0] data_out_33,
    output [1023:0] data_out_34,
    output [1023:0] data_out_35,
    output [1023:0] data_out_36,
    output [1023:0] data_out_37,
    output [1023:0] data_out_38,
    output [1023:0] data_out_39,
    output [1023:0] data_out_40,
    output [1023:0] data_out_41,
    output [1023:0] data_out_42,
    output [1023:0] data_out_43,
    output [1023:0] data_out_44,
    output [1023:0] data_out_45,
    output [1023:0] data_out_46,
    output [1023:0] data_out_47,
    output [1023:0] data_out_48,
    output [1023:0] data_out_49,
    output [1023:0] data_out_50,
    output [1023:0] data_out_51,
    output [1023:0] data_out_52
);





xpb_5_0 u_xpb_5_0(.data_in(data_in[ 4 : 0] ), .data_out(data_out_0));
xpb_5_5 u_xpb_5_5(.data_in(data_in[ 9 : 5] ), .data_out(data_out_1));
xpb_5_10 u_xpb_5_10(.data_in(data_in[ 14 : 10] ), .data_out(data_out_2));
xpb_5_15 u_xpb_5_15(.data_in(data_in[ 19 : 15] ), .data_out(data_out_3));
xpb_5_20 u_xpb_5_20(.data_in(data_in[ 24 : 20] ), .data_out(data_out_4));
xpb_5_25 u_xpb_5_25(.data_in(data_in[ 29 : 25] ), .data_out(data_out_5));
xpb_5_30 u_xpb_5_30(.data_in(data_in[ 34 : 30] ), .data_out(data_out_6));
xpb_5_35 u_xpb_5_35(.data_in(data_in[ 39 : 35] ), .data_out(data_out_7));
xpb_5_40 u_xpb_5_40(.data_in(data_in[ 44 : 40] ), .data_out(data_out_8));
xpb_5_45 u_xpb_5_45(.data_in(data_in[ 49 : 45] ), .data_out(data_out_9));
xpb_5_50 u_xpb_5_50(.data_in(data_in[ 54 : 50] ), .data_out(data_out_10));
xpb_5_55 u_xpb_5_55(.data_in(data_in[ 59 : 55] ), .data_out(data_out_11));
xpb_5_60 u_xpb_5_60(.data_in(data_in[ 64 : 60] ), .data_out(data_out_12));
xpb_5_65 u_xpb_5_65(.data_in(data_in[ 69 : 65] ), .data_out(data_out_13));
xpb_5_70 u_xpb_5_70(.data_in(data_in[ 74 : 70] ), .data_out(data_out_14));
xpb_5_75 u_xpb_5_75(.data_in(data_in[ 79 : 75] ), .data_out(data_out_15));
xpb_5_80 u_xpb_5_80(.data_in(data_in[ 84 : 80] ), .data_out(data_out_16));
xpb_5_85 u_xpb_5_85(.data_in(data_in[ 89 : 85] ), .data_out(data_out_17));
xpb_5_90 u_xpb_5_90(.data_in(data_in[ 94 : 90] ), .data_out(data_out_18));
xpb_5_95 u_xpb_5_95(.data_in(data_in[ 99 : 95] ), .data_out(data_out_19));
xpb_5_100 u_xpb_5_100(.data_in(data_in[ 104 : 100] ), .data_out(data_out_20));
xpb_5_105 u_xpb_5_105(.data_in(data_in[ 109 : 105] ), .data_out(data_out_21));
xpb_5_110 u_xpb_5_110(.data_in(data_in[ 114 : 110] ), .data_out(data_out_22));
xpb_5_115 u_xpb_5_115(.data_in(data_in[ 119 : 115] ), .data_out(data_out_23));
xpb_5_120 u_xpb_5_120(.data_in(data_in[ 124 : 120] ), .data_out(data_out_24));
xpb_5_125 u_xpb_5_125(.data_in(data_in[ 129 : 125] ), .data_out(data_out_25));
xpb_5_130 u_xpb_5_130(.data_in(data_in[ 134 : 130] ), .data_out(data_out_26));
xpb_5_135 u_xpb_5_135(.data_in(data_in[ 139 : 135] ), .data_out(data_out_27));
xpb_5_140 u_xpb_5_140(.data_in(data_in[ 144 : 140] ), .data_out(data_out_28));
xpb_5_145 u_xpb_5_145(.data_in(data_in[ 149 : 145] ), .data_out(data_out_29));
xpb_5_150 u_xpb_5_150(.data_in(data_in[ 154 : 150] ), .data_out(data_out_30));
xpb_5_155 u_xpb_5_155(.data_in(data_in[ 159 : 155] ), .data_out(data_out_31));
xpb_5_160 u_xpb_5_160(.data_in(data_in[ 164 : 160] ), .data_out(data_out_32));
xpb_5_165 u_xpb_5_165(.data_in(data_in[ 169 : 165] ), .data_out(data_out_33));
xpb_5_170 u_xpb_5_170(.data_in(data_in[ 174 : 170] ), .data_out(data_out_34));
xpb_5_175 u_xpb_5_175(.data_in(data_in[ 179 : 175] ), .data_out(data_out_35));
xpb_5_180 u_xpb_5_180(.data_in(data_in[ 184 : 180] ), .data_out(data_out_36));
xpb_5_185 u_xpb_5_185(.data_in(data_in[ 189 : 185] ), .data_out(data_out_37));
xpb_5_190 u_xpb_5_190(.data_in(data_in[ 194 : 190] ), .data_out(data_out_38));
xpb_5_195 u_xpb_5_195(.data_in(data_in[ 199 : 195] ), .data_out(data_out_39));
xpb_5_200 u_xpb_5_200(.data_in(data_in[ 204 : 200] ), .data_out(data_out_40));
xpb_5_205 u_xpb_5_205(.data_in(data_in[ 209 : 205] ), .data_out(data_out_41));
xpb_5_210 u_xpb_5_210(.data_in(data_in[ 214 : 210] ), .data_out(data_out_42));
xpb_5_215 u_xpb_5_215(.data_in(data_in[ 219 : 215] ), .data_out(data_out_43));
xpb_5_220 u_xpb_5_220(.data_in(data_in[ 224 : 220] ), .data_out(data_out_44));
xpb_5_225 u_xpb_5_225(.data_in(data_in[ 229 : 225] ), .data_out(data_out_45));
xpb_5_230 u_xpb_5_230(.data_in(data_in[ 234 : 230] ), .data_out(data_out_46));
xpb_5_235 u_xpb_5_235(.data_in(data_in[ 239 : 235] ), .data_out(data_out_47));
xpb_5_240 u_xpb_5_240(.data_in(data_in[ 244 : 240] ), .data_out(data_out_48));
xpb_5_245 u_xpb_5_245(.data_in(data_in[ 249 : 245] ), .data_out(data_out_49));
xpb_5_250 u_xpb_5_250(.data_in(data_in[ 254 : 250] ), .data_out(data_out_50));
xpb_5_255 u_xpb_5_255(.data_in(data_in[ 259 : 255] ), .data_out(data_out_51));
xpb_4_260 u_xpb_4_260(.data_in(data_in[263 : 260]), .data_out(data_out_52));


endmodule



module xpb_5_230
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9557bf8b5b7368950d03e30c6b0dc228b09955e22d07bf9927a2227194c394793de59529a1ed3d38daf9022cd386eccfefdef290a8e4c9c6172250029b12aecba71835e996506170f1f200798b21f5969e6ee643fafd161aad690bad40846be07538f52d8ba8be3d6f1287d0553ae4d0654932642b86491fe7dae08f619a0619;
    5'b00010 : xpb = 1024'h7a0239c0f4f89c614f024e41c5c13cffefbca8938497debad1678b8d76847bea7882acda79b3fbe31693c512c3afc8d57ba3bd3b2f16c3407da560a6fb52e8e5d9e137247d0fc59cd149fe507d6826fc48d8d2ef6973ff24a545855fc6de352ebb6a5831668883ed576528c1b2a5a3777bb885e606c1350f8946461a3a51a5c7;
    5'b00011 : xpb = 1024'h5eacb3f68e7dd02d9100b9772074b7d72edffb44dc27fddc7b2cf4a95845635bb31fc48b517aba8d522e87f8b3d8a4db076887e5b548bcbae428714b5b9323000caa385f63cf29c8b0a1fc276fae5861f342bf9ad7eae82e9d21ff124d37fe7d019bbb354168499d3fb7c9b31010621e9227d967e1fc20ff2ab1aba513094575;
    5'b00100 : xpb = 1024'h43572e2c280303f9d2ff24ac7b2832ae6e034df633b81cfe24f25dc53a064accedbcdc3c294179378dc94adea40180e0932d52903b7ab6354aab81efbbd35d1a3f73399a4a8e8df48ff9f9fe61f489c79dacac464661d13894fe78c4d391c7cb47cd1e391c480f4d280a6aa46d7b20c5a8972ce9bd370ceecc1d112febc0e523;
    5'b00101 : xpb = 1024'h2801a861c18837c614fd8fe1d5dbad85ad26a0a78b483c1fceb7c6e11bc7323e2859f3ed010837e1c9640dc4942a5ce61ef21d3ac1acafafb12e92941c139734723c3ad5314df2206f51f7d5543abb2d481698f1b4d8ba428cdaf27759eb91198dfe813cf727d4fd105d0b95cae5df6cbf06806b9871f8de6d8876bac47884d1;
    5'b00110 : xpb = 1024'hcac22975b0d6b9256fbfb17308f285cec49f358e2d85b41787d2ffcfd8819af62f70b9dd8cef68c04fed0aa845338ebaab6e7e547dea92a17b1a3387c53d14ea5053c10180d564c4ea9f5ac4680ec92f280859d234fa34c84b76c29e0455a67d42fe440d2079aacf8afac8728509e13d575d3ed73ace4ce0ef3dc459d30247f;
    5'b00111 : xpb = 1024'ha203e222b680d42763ffde239b9cea859ce3493b0fe01adaa01f526e924bae28a0dca0c77abc33c4dff7d2d757da25bb9a95da75f0c372f02ed3f33b1766801a4c1d71f9ae5db7bd409bf625d1a2e22990ef6be11e4cb967322077d720c9c6484968d96e5db058ea67c234577d8b82e43abf06519f332dedf6cebcd4feca2a98;
    5'b01000 : xpb = 1024'h86ae5c58500607f3a5fe4958f650655cdc069bec677039fc49e4bb8a740c9599db79b8785282f26f1b9295bd480301c1265aa52076f56c6a955703df77a6ba347ee67334951d1be91ff3f3fcc3e9138f3b59588c8cc3a27129fcf189a7238f968f9a3c7238901e9a5014d548daf6418b512e59d37a6e19dd983a225fd781ca46;
    5'b01001 : xpb = 1024'h6b58d68de98b3bbfe7fcb48e5103e0341b29ee9dbf00591df3aa24a655cd7d0b1616d0292a49b119572d58a3382bddc6b21f6fcafd2765e4fbda1483d7e6f44eb1af746f7bdc8014ff4bf1d3b62f44f4e5c34537fb3a8b7b21d96b3c2d7d58e4d5cb9f76136fe44a3867763a38610032679dad5555a905cd39a587eab03969f4;
    5'b01010 : xpb = 1024'h500350c383106f8c29fb1fc3abb75b0b5a4d414f1690783f9d6f8dc2378e647c50b3e7da02106fc392c81b892854b9cc3de43a7583595f5f625d252838272e68e47875aa629be440dea3efaaa875765a902d31e369b1748519b5e4eeb3d722331bfd0279ee4fa9fa20ba172b95cbbed97e0d00d730e3f1bcdb10ed7588f109a2;
    5'b01011 : xpb = 1024'h34adcaf91c95a3586bf98af9066ad5e2997094006e2097614734f6de194f4bed8b50ff8ad9d72e6dce62de6f187d95d1c9a90520098b58d9c8e035cc98676883174176e5495b486cbdfbed819abba7c03a971e8ed8285d8f11925ea13a30eb81622e657dc92f6faa090cb81cf3367d80947c54590c1eddac7c7c530061a8a950;
    5'b01100 : xpb = 1024'h1958452eb61ad724adf7f62e611e50b9d893e6b1c5b0b682f0fa5ff9fb10335ec5ee173bb19ded1809fda15508a671d7556dcfca8fbd52542f634670f8a7a29d4a0a7820301aac989d53eb588d01d925e5010b3a469f4699096ed853c08ab4cfa85fc881a40f3559f15f590e50a13c27aaeba7dae759c99c1de7b88b3a6048fe;
    5'b01101 : xpb = 1024'haeb004ba118e3fb9bafbd93acc2c12e2892d3c93f2b8761c189c826b8fd3c7d803d3ac65538b2a50e4f6a381dc2d5ea7454cc25b38a21c1a4685967393ba5168f122ae09c66b0e098f45ebd21823cebc836ff17e419c5cb3b6d7e401010f20b01d98bdaf2fb7f3976071e0dea5dc20f81034da3f12e012bc05c2991a9bfa4f17;
    5'b01110 : xpb = 1024'h935a7eefab137385fcfa447026df8db9c8508f454a48953dc261eb877194af493e70c4162b51e8fb20916667cc563aacd1118d05bed41594ad08a717f3fa8b8323ebaf44ad2a72356e9de9a90a6a00222dd9de29b01345bdaeb45db38768e9fe63ca20b30a97b94748c481d00346df9f26a42dc0ee1afeaba72dfea574b1eec5;
    5'b01111 : xpb = 1024'h7804f9254498a7523ef8afa5819308910773e1f6a1d8b45f6c2754a3535596ba790ddbc70318a7a55c2c294dbc7f16b25cd657b045060f0f138bb7bc543ac59d56b4b07f93e9d6614df5e77ffcb03187d843cad51e8a2ec7a690d7660dc2b34ca9fb83b6e5777ef7311722c160b19e463d138142c955ea9b489964304d698e73;
    5'b10000 : xpb = 1024'h5caf735ade1ddb1e80f71adadc468368469734a7f968d38115ecbdbf35167e2bb3aaf377dadf664f97c6ec33aca7f2b7e89b225acb3808897a0ec860b47affb7897db1ba7aa93a8d2d4de556eef662ed82adb7808d0117d19e6d5118941c7c9af02ce6bac05744a71969c3b2be1c5ced5382d4c4a490d68aea04c9bb26212e21;
    5'b10001 : xpb = 1024'h4159ed9077a30eeac2f5861036f9fe3f85ba875950f8f2a2bfb226db16d7659cee480b28b2a624f9d361af199cd0cebd745fed05516a0203e091d90514bb39d1bc46b2f561689eb90ca5e32de13c94532d17a42bfb7800db9649cacb1a7645e9365e49be9b370a5701bc64a41b871b9469f228467fcbc27a8b702f45fed8cdcf;
    5'b10010 : xpb = 1024'h260467c6112842b704f3f14591ad7916c4ddda0aa88911c469778ff6f8984d0e28e522d98a6ce3a40efc71ff8cf9aac30024b7afd79bfb7e4714e9a974fb73ebef0fb430482802e4ebfde104d382c5b8d78190d769eee9e58e26447da0d00f377c8facc27616d006ea0f059578f1da3b80617bc85b06ae6a2cdb94d0d7906d7d;
    5'b10011 : xpb = 1024'haaee1fbaaad768346f25c7aec60f3ee04012cbc001930e6133cf912da59347f63823a8a6233a24e4a9734e57d2286c88be9825a5dcdf4f8ad97fa4dd53bae0621d8b56b2ee76710cb55dedbc5c8f71e81eb7d82d865d2ef8602be302729d885c2c10fc650f695b6d261a686d65c98e296d0cf4a36419a59ce46fa5bb0480d2b;
    5'b10100 : xpb = 1024'ha006a1870620df1853f63f87576eb616b49a829e2d20f07f3adf1b846f1cc8f8a167cfb40420df872590371250a973987bc874eb06b2bebec4ba4a50704e5cd1c8f0eb54c537c881bd47df5550eaecb5205a63c6d362e90a336bc9dd67ae446637fa04f3dc9f53f441742e572b977db2fc1a01ae61c7e379b621daeb11e21344;
    5'b10101 : xpb = 1024'h84b11bbc9fa612e495f4aabcb22230edf3bdd54f84b10fa0e4a484a050ddb069dc04e764dbe79e31612af9f840d24f9e078d3f958ce4b8392b3d5af4d08e96ebfbb9ec8fabf72cad9c9fdd2c43311e1acac4507241d9d2142b48438fee080db47e2b67f7b77f19a429c6cf4889023c5a128955303d02cf69578d4075ea99b2f2;
    5'b10110 : xpb = 1024'h695b95f2392b46b0d7f315f20cd5abc532e12800dc412ec28e69edbc329e97db16a1ff15b3ae5cdb9cc5bcde30fb2ba393520a401316b1b391c06b9930ced1062e82edca92b690d97bf7db0335774f80752e3d1db050bb1e2324bd427461d702c45ccafb925edf5412197039e66cfb0128f8a8b2183dbb58f8f8a600c35152a0;
    5'b10111 : xpb = 1024'h4e061027d2b07a7d19f181276789269c72047ab233d14de4382f56d8145f7f4c513f16c68b751b85d8607fc4212407a91f16d4ea9948ab2df8437c3d910f0b20614bef057975f5055b4fd8da27bd80e61f9829c91ec7a4281b0136f4fabba0510a8e2dff6d3ea503fa6c112b43d7b9a83f67fc33f378a7489a640b8b9c08f24e;
    5'b11000 : xpb = 1024'h32b08a5d6c35ae495befec5cc23ca173b127cd638b616d05e1f4bff3f62066bd8bdc2e77633bda3013fb42aa114ce3aeaadb9f951f7aa4a85ec68ce1f14f453a9414f040603559313aa7d6b11a03b24bca0216748d3e8d3212ddb0a78115699f50bf9103481e6ab3e2beb21ca142784f55d74fb5ceb393383bcf711674c091fc;
    5'b11001 : xpb = 1024'h175b049305bae2159dee57921cf01c4af04b2014e2f18c278bba290fd7e14e2ec67946283b0298da4f9605900175bfb436a06a3fa5ac9e22c5499d86518f7f54c6ddf17b46f4bd5d19ffd4880c49e3b1746c031ffbb5763c0aba2a5a076f32ed96f0f40722fe3063cb11530dfead36f66c46a337a9ee7f27dd3ad6a14d7831aa;
    5'b11010 : xpb = 1024'hacb2c41e612e4aaaaaf23a9e87fdde73a0e475f70ff94bc0b35c4b816ca4e2a8045edb51dcefd6132a8f07bcd4fcac84267f5cd04e9167e8dc6bed88eca22e206df62764dd451ece0bf1d501976bd94812dae963f6b28c56b823360747f39ece0c29e934aea6eea13a23dade53e81bc6d18fd59bd574c847c515b730af1237c3;
    5'b11011 : xpb = 1024'h915d3e53fab37e76ecf0a5d3e2b1594ae007c8a867896ae25d21b49d4e65ca193efbf302b4b694bd6629caa2c5258889b244277ad4c3616342eefe2d4ce2683aa0bf289fc40482f9eb49d2d889b20aadbd44d60f65297560afffafb9ce4d681c525b4c388986b45122767bcfb152da6de7ff291db0afb43766811cbb87c9d771;
    5'b11100 : xpb = 1024'h7607b8899438b2432eef11093d64d4221f2b1b59bf198a0406e71db93026b18a79990ab38c7d5367a1c48d88b54e648f3e08f2255af55adda9720ed1ad22a254d38829daaac3e725caa1d0af7bf83c1367aec2bad3a05e6aa7dc296c54a7316a988caf3c64667a010ac91cc10ebd9914fe6e7c9f8beaa02707ec82466081771f;
    5'b11101 : xpb = 1024'h5ab232bf2dbde60f70ed7c3e98184ef95e4e6e0b16a9a925b0ac86d511e798fbb436226464441211dd5f506ea5774094c9cdbccfe12754580ff51f760d62dc6f06512b1591834b51a9f9ce866e3e6d791218af66421747749fb8a31edb00fab8debe12403f463fb0f31bbdb26c2857bc14ddd02167258c16a957e7d1393916cd;
    5'b11110 : xpb = 1024'h3f5cacf4c74319dbb2ebe773f2cbc9d09d71c0bc6e39c8475a71eff0f3a8806ceed33a153c0ad0bc18fa135495a01c9a5592877a67594dd27678301a6da31689391a2c507842af7d8951cc5d60849edebc829c11b08e307e97951cd1615ac40724ef75441a260560db6e5ea3c99316632b4d23a3426078064ac34d5c11f0b67b;
    5'b11111 : xpb = 1024'h2407272a60c84da7f4ea52a94d7f44a7dc95136dc5c9e7690437590cd56967de297051c613d18f665494d63a85c8f89fe1575224ed8b474cdcfb40becde350a36be32d8b5f0213a968a9ca3452cad04466ec88bd1f0519888f719683e7b48d556b20d847f505cb10c3c0ff9526fdd50a41bc77251d9b63f5ec2eb2e6eaa85629;
    endcase
end

endmodule

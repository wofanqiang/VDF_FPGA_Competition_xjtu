`timescale 1ns/1ns
/*******************************************************************************
    Institute:   Xi'an Jiaotong University
    Department:  Microelectronic
    Author :     Li Xiaocong

    Unless you get the permission of the Author, you can't modify,
    distribute or use for commercial purposes.
*******************************************************************************/
module msq_half_product_gene
(
	input wire [1023:0] a,
	input wire sel,
	output wire [511:0] col_0,
	output wire [511:0] col_1,
	output wire [511:0] col_2,
	output wire [511:0] col_3,
	output wire [511:0] col_4,
	output wire [511:0] col_5,
	output wire [511:0] col_6,
	output wire [511:0] col_7,
	output wire [511:0] col_8,
	output wire [511:0] col_9,
	output wire [511:0] col_10,
	output wire [511:0] col_11,
	output wire [511:0] col_12,
	output wire [511:0] col_13,
	output wire [511:0] col_14,
	output wire [511:0] col_15,
	output wire [511:0] col_16,
	output wire [511:0] col_17,
	output wire [511:0] col_18,
	output wire [511:0] col_19,
	output wire [511:0] col_20,
	output wire [511:0] col_21,
	output wire [511:0] col_22,
	output wire [511:0] col_23,
	output wire [511:0] col_24,
	output wire [511:0] col_25,
	output wire [511:0] col_26,
	output wire [511:0] col_27,
	output wire [511:0] col_28,
	output wire [511:0] col_29,
	output wire [511:0] col_30,
	output wire [511:0] col_31,
	output wire [511:0] col_32,
	output wire [511:0] col_33,
	output wire [511:0] col_34,
	output wire [511:0] col_35,
	output wire [511:0] col_36,
	output wire [511:0] col_37,
	output wire [511:0] col_38,
	output wire [511:0] col_39,
	output wire [511:0] col_40,
	output wire [511:0] col_41,
	output wire [511:0] col_42,
	output wire [511:0] col_43,
	output wire [511:0] col_44,
	output wire [511:0] col_45,
	output wire [511:0] col_46,
	output wire [511:0] col_47,
	output wire [511:0] col_48,
	output wire [511:0] col_49,
	output wire [511:0] col_50,
	output wire [511:0] col_51,
	output wire [511:0] col_52,
	output wire [511:0] col_53,
	output wire [511:0] col_54,
	output wire [511:0] col_55,
	output wire [511:0] col_56,
	output wire [511:0] col_57,
	output wire [511:0] col_58,
	output wire [511:0] col_59,
	output wire [511:0] col_60,
	output wire [511:0] col_61,
	output wire [511:0] col_62,
	output wire [511:0] col_63,
	output wire [511:0] col_64,
	output wire [511:0] col_65,
	output wire [511:0] col_66,
	output wire [511:0] col_67,
	output wire [511:0] col_68,
	output wire [511:0] col_69,
	output wire [511:0] col_70,
	output wire [511:0] col_71,
	output wire [511:0] col_72,
	output wire [511:0] col_73,
	output wire [511:0] col_74,
	output wire [511:0] col_75,
	output wire [511:0] col_76,
	output wire [511:0] col_77,
	output wire [511:0] col_78,
	output wire [511:0] col_79,
	output wire [511:0] col_80,
	output wire [511:0] col_81,
	output wire [511:0] col_82,
	output wire [511:0] col_83,
	output wire [511:0] col_84,
	output wire [511:0] col_85,
	output wire [511:0] col_86,
	output wire [511:0] col_87,
	output wire [511:0] col_88,
	output wire [511:0] col_89,
	output wire [511:0] col_90,
	output wire [511:0] col_91,
	output wire [511:0] col_92,
	output wire [511:0] col_93,
	output wire [511:0] col_94,
	output wire [511:0] col_95,
	output wire [511:0] col_96,
	output wire [511:0] col_97,
	output wire [511:0] col_98,
	output wire [511:0] col_99,
	output wire [511:0] col_100,
	output wire [511:0] col_101,
	output wire [511:0] col_102,
	output wire [511:0] col_103,
	output wire [511:0] col_104,
	output wire [511:0] col_105,
	output wire [511:0] col_106,
	output wire [511:0] col_107,
	output wire [511:0] col_108,
	output wire [511:0] col_109,
	output wire [511:0] col_110,
	output wire [511:0] col_111,
	output wire [511:0] col_112,
	output wire [511:0] col_113,
	output wire [511:0] col_114,
	output wire [511:0] col_115,
	output wire [511:0] col_116,
	output wire [511:0] col_117,
	output wire [511:0] col_118,
	output wire [511:0] col_119,
	output wire [511:0] col_120,
	output wire [511:0] col_121,
	output wire [511:0] col_122,
	output wire [511:0] col_123,
	output wire [511:0] col_124,
	output wire [511:0] col_125,
	output wire [511:0] col_126,
	output wire [511:0] col_127,
	output wire [511:0] col_128,
	output wire [511:0] col_129,
	output wire [511:0] col_130,
	output wire [511:0] col_131,
	output wire [511:0] col_132,
	output wire [511:0] col_133,
	output wire [511:0] col_134,
	output wire [511:0] col_135,
	output wire [511:0] col_136,
	output wire [511:0] col_137,
	output wire [511:0] col_138,
	output wire [511:0] col_139,
	output wire [511:0] col_140,
	output wire [511:0] col_141,
	output wire [511:0] col_142,
	output wire [511:0] col_143,
	output wire [511:0] col_144,
	output wire [511:0] col_145,
	output wire [511:0] col_146,
	output wire [511:0] col_147,
	output wire [511:0] col_148,
	output wire [511:0] col_149,
	output wire [511:0] col_150,
	output wire [511:0] col_151,
	output wire [511:0] col_152,
	output wire [511:0] col_153,
	output wire [511:0] col_154,
	output wire [511:0] col_155,
	output wire [511:0] col_156,
	output wire [511:0] col_157,
	output wire [511:0] col_158,
	output wire [511:0] col_159,
	output wire [511:0] col_160,
	output wire [511:0] col_161,
	output wire [511:0] col_162,
	output wire [511:0] col_163,
	output wire [511:0] col_164,
	output wire [511:0] col_165,
	output wire [511:0] col_166,
	output wire [511:0] col_167,
	output wire [511:0] col_168,
	output wire [511:0] col_169,
	output wire [511:0] col_170,
	output wire [511:0] col_171,
	output wire [511:0] col_172,
	output wire [511:0] col_173,
	output wire [511:0] col_174,
	output wire [511:0] col_175,
	output wire [511:0] col_176,
	output wire [511:0] col_177,
	output wire [511:0] col_178,
	output wire [511:0] col_179,
	output wire [511:0] col_180,
	output wire [511:0] col_181,
	output wire [511:0] col_182,
	output wire [511:0] col_183,
	output wire [511:0] col_184,
	output wire [511:0] col_185,
	output wire [511:0] col_186,
	output wire [511:0] col_187,
	output wire [511:0] col_188,
	output wire [511:0] col_189,
	output wire [511:0] col_190,
	output wire [511:0] col_191,
	output wire [511:0] col_192,
	output wire [511:0] col_193,
	output wire [511:0] col_194,
	output wire [511:0] col_195,
	output wire [511:0] col_196,
	output wire [511:0] col_197,
	output wire [511:0] col_198,
	output wire [511:0] col_199,
	output wire [511:0] col_200,
	output wire [511:0] col_201,
	output wire [511:0] col_202,
	output wire [511:0] col_203,
	output wire [511:0] col_204,
	output wire [511:0] col_205,
	output wire [511:0] col_206,
	output wire [511:0] col_207,
	output wire [511:0] col_208,
	output wire [511:0] col_209,
	output wire [511:0] col_210,
	output wire [511:0] col_211,
	output wire [511:0] col_212,
	output wire [511:0] col_213,
	output wire [511:0] col_214,
	output wire [511:0] col_215,
	output wire [511:0] col_216,
	output wire [511:0] col_217,
	output wire [511:0] col_218,
	output wire [511:0] col_219,
	output wire [511:0] col_220,
	output wire [511:0] col_221,
	output wire [511:0] col_222,
	output wire [511:0] col_223,
	output wire [511:0] col_224,
	output wire [511:0] col_225,
	output wire [511:0] col_226,
	output wire [511:0] col_227,
	output wire [511:0] col_228,
	output wire [511:0] col_229,
	output wire [511:0] col_230,
	output wire [511:0] col_231,
	output wire [511:0] col_232,
	output wire [511:0] col_233,
	output wire [511:0] col_234,
	output wire [511:0] col_235,
	output wire [511:0] col_236,
	output wire [511:0] col_237,
	output wire [511:0] col_238,
	output wire [511:0] col_239,
	output wire [511:0] col_240,
	output wire [511:0] col_241,
	output wire [511:0] col_242,
	output wire [511:0] col_243,
	output wire [511:0] col_244,
	output wire [511:0] col_245,
	output wire [511:0] col_246,
	output wire [511:0] col_247,
	output wire [511:0] col_248,
	output wire [511:0] col_249,
	output wire [511:0] col_250,
	output wire [511:0] col_251,
	output wire [511:0] col_252,
	output wire [511:0] col_253,
	output wire [511:0] col_254,
	output wire [511:0] col_255,
	output wire [511:0] col_256,
	output wire [511:0] col_257,
	output wire [511:0] col_258,
	output wire [511:0] col_259,
	output wire [511:0] col_260,
	output wire [511:0] col_261,
	output wire [511:0] col_262,
	output wire [511:0] col_263,
	output wire [511:0] col_264,
	output wire [511:0] col_265,
	output wire [511:0] col_266,
	output wire [511:0] col_267,
	output wire [511:0] col_268,
	output wire [511:0] col_269,
	output wire [511:0] col_270,
	output wire [511:0] col_271,
	output wire [511:0] col_272,
	output wire [511:0] col_273,
	output wire [511:0] col_274,
	output wire [511:0] col_275,
	output wire [511:0] col_276,
	output wire [511:0] col_277,
	output wire [511:0] col_278,
	output wire [511:0] col_279,
	output wire [511:0] col_280,
	output wire [511:0] col_281,
	output wire [511:0] col_282,
	output wire [511:0] col_283,
	output wire [511:0] col_284,
	output wire [511:0] col_285,
	output wire [511:0] col_286,
	output wire [511:0] col_287,
	output wire [511:0] col_288,
	output wire [511:0] col_289,
	output wire [511:0] col_290,
	output wire [511:0] col_291,
	output wire [511:0] col_292,
	output wire [511:0] col_293,
	output wire [511:0] col_294,
	output wire [511:0] col_295,
	output wire [511:0] col_296,
	output wire [511:0] col_297,
	output wire [511:0] col_298,
	output wire [511:0] col_299,
	output wire [511:0] col_300,
	output wire [511:0] col_301,
	output wire [511:0] col_302,
	output wire [511:0] col_303,
	output wire [511:0] col_304,
	output wire [511:0] col_305,
	output wire [511:0] col_306,
	output wire [511:0] col_307,
	output wire [511:0] col_308,
	output wire [511:0] col_309,
	output wire [511:0] col_310,
	output wire [511:0] col_311,
	output wire [511:0] col_312,
	output wire [511:0] col_313,
	output wire [511:0] col_314,
	output wire [511:0] col_315,
	output wire [511:0] col_316,
	output wire [511:0] col_317,
	output wire [511:0] col_318,
	output wire [511:0] col_319,
	output wire [511:0] col_320,
	output wire [511:0] col_321,
	output wire [511:0] col_322,
	output wire [511:0] col_323,
	output wire [511:0] col_324,
	output wire [511:0] col_325,
	output wire [511:0] col_326,
	output wire [511:0] col_327,
	output wire [511:0] col_328,
	output wire [511:0] col_329,
	output wire [511:0] col_330,
	output wire [511:0] col_331,
	output wire [511:0] col_332,
	output wire [511:0] col_333,
	output wire [511:0] col_334,
	output wire [511:0] col_335,
	output wire [511:0] col_336,
	output wire [511:0] col_337,
	output wire [511:0] col_338,
	output wire [511:0] col_339,
	output wire [511:0] col_340,
	output wire [511:0] col_341,
	output wire [511:0] col_342,
	output wire [511:0] col_343,
	output wire [511:0] col_344,
	output wire [511:0] col_345,
	output wire [511:0] col_346,
	output wire [511:0] col_347,
	output wire [511:0] col_348,
	output wire [511:0] col_349,
	output wire [511:0] col_350,
	output wire [511:0] col_351,
	output wire [511:0] col_352,
	output wire [511:0] col_353,
	output wire [511:0] col_354,
	output wire [511:0] col_355,
	output wire [511:0] col_356,
	output wire [511:0] col_357,
	output wire [511:0] col_358,
	output wire [511:0] col_359,
	output wire [511:0] col_360,
	output wire [511:0] col_361,
	output wire [511:0] col_362,
	output wire [511:0] col_363,
	output wire [511:0] col_364,
	output wire [511:0] col_365,
	output wire [511:0] col_366,
	output wire [511:0] col_367,
	output wire [511:0] col_368,
	output wire [511:0] col_369,
	output wire [511:0] col_370,
	output wire [511:0] col_371,
	output wire [511:0] col_372,
	output wire [511:0] col_373,
	output wire [511:0] col_374,
	output wire [511:0] col_375,
	output wire [511:0] col_376,
	output wire [511:0] col_377,
	output wire [511:0] col_378,
	output wire [511:0] col_379,
	output wire [511:0] col_380,
	output wire [511:0] col_381,
	output wire [511:0] col_382,
	output wire [511:0] col_383,
	output wire [511:0] col_384,
	output wire [511:0] col_385,
	output wire [511:0] col_386,
	output wire [511:0] col_387,
	output wire [511:0] col_388,
	output wire [511:0] col_389,
	output wire [511:0] col_390,
	output wire [511:0] col_391,
	output wire [511:0] col_392,
	output wire [511:0] col_393,
	output wire [511:0] col_394,
	output wire [511:0] col_395,
	output wire [511:0] col_396,
	output wire [511:0] col_397,
	output wire [511:0] col_398,
	output wire [511:0] col_399,
	output wire [511:0] col_400,
	output wire [511:0] col_401,
	output wire [511:0] col_402,
	output wire [511:0] col_403,
	output wire [511:0] col_404,
	output wire [511:0] col_405,
	output wire [511:0] col_406,
	output wire [511:0] col_407,
	output wire [511:0] col_408,
	output wire [511:0] col_409,
	output wire [511:0] col_410,
	output wire [511:0] col_411,
	output wire [511:0] col_412,
	output wire [511:0] col_413,
	output wire [511:0] col_414,
	output wire [511:0] col_415,
	output wire [511:0] col_416,
	output wire [511:0] col_417,
	output wire [511:0] col_418,
	output wire [511:0] col_419,
	output wire [511:0] col_420,
	output wire [511:0] col_421,
	output wire [511:0] col_422,
	output wire [511:0] col_423,
	output wire [511:0] col_424,
	output wire [511:0] col_425,
	output wire [511:0] col_426,
	output wire [511:0] col_427,
	output wire [511:0] col_428,
	output wire [511:0] col_429,
	output wire [511:0] col_430,
	output wire [511:0] col_431,
	output wire [511:0] col_432,
	output wire [511:0] col_433,
	output wire [511:0] col_434,
	output wire [511:0] col_435,
	output wire [511:0] col_436,
	output wire [511:0] col_437,
	output wire [511:0] col_438,
	output wire [511:0] col_439,
	output wire [511:0] col_440,
	output wire [511:0] col_441,
	output wire [511:0] col_442,
	output wire [511:0] col_443,
	output wire [511:0] col_444,
	output wire [511:0] col_445,
	output wire [511:0] col_446,
	output wire [511:0] col_447,
	output wire [511:0] col_448,
	output wire [511:0] col_449,
	output wire [511:0] col_450,
	output wire [511:0] col_451,
	output wire [511:0] col_452,
	output wire [511:0] col_453,
	output wire [511:0] col_454,
	output wire [511:0] col_455,
	output wire [511:0] col_456,
	output wire [511:0] col_457,
	output wire [511:0] col_458,
	output wire [511:0] col_459,
	output wire [511:0] col_460,
	output wire [511:0] col_461,
	output wire [511:0] col_462,
	output wire [511:0] col_463,
	output wire [511:0] col_464,
	output wire [511:0] col_465,
	output wire [511:0] col_466,
	output wire [511:0] col_467,
	output wire [511:0] col_468,
	output wire [511:0] col_469,
	output wire [511:0] col_470,
	output wire [511:0] col_471,
	output wire [511:0] col_472,
	output wire [511:0] col_473,
	output wire [511:0] col_474,
	output wire [511:0] col_475,
	output wire [511:0] col_476,
	output wire [511:0] col_477,
	output wire [511:0] col_478,
	output wire [511:0] col_479,
	output wire [511:0] col_480,
	output wire [511:0] col_481,
	output wire [511:0] col_482,
	output wire [511:0] col_483,
	output wire [511:0] col_484,
	output wire [511:0] col_485,
	output wire [511:0] col_486,
	output wire [511:0] col_487,
	output wire [511:0] col_488,
	output wire [511:0] col_489,
	output wire [511:0] col_490,
	output wire [511:0] col_491,
	output wire [511:0] col_492,
	output wire [511:0] col_493,
	output wire [511:0] col_494,
	output wire [511:0] col_495,
	output wire [511:0] col_496,
	output wire [511:0] col_497,
	output wire [511:0] col_498,
	output wire [511:0] col_499,
	output wire [511:0] col_500,
	output wire [511:0] col_501,
	output wire [511:0] col_502,
	output wire [511:0] col_503,
	output wire [511:0] col_504,
	output wire [511:0] col_505,
	output wire [511:0] col_506,
	output wire [511:0] col_507,
	output wire [511:0] col_508,
	output wire [511:0] col_509,
	output wire [511:0] col_510,
	output wire [511:0] col_511,
	output wire [511:0] col_512,
	output wire [511:0] col_513,
	output wire [511:0] col_514,
	output wire [511:0] col_515,
	output wire [511:0] col_516,
	output wire [511:0] col_517,
	output wire [511:0] col_518,
	output wire [511:0] col_519,
	output wire [511:0] col_520,
	output wire [511:0] col_521,
	output wire [511:0] col_522,
	output wire [511:0] col_523,
	output wire [511:0] col_524,
	output wire [511:0] col_525,
	output wire [511:0] col_526,
	output wire [511:0] col_527,
	output wire [511:0] col_528,
	output wire [511:0] col_529,
	output wire [511:0] col_530,
	output wire [511:0] col_531,
	output wire [511:0] col_532,
	output wire [511:0] col_533,
	output wire [511:0] col_534,
	output wire [511:0] col_535,
	output wire [511:0] col_536,
	output wire [511:0] col_537,
	output wire [511:0] col_538,
	output wire [511:0] col_539,
	output wire [511:0] col_540,
	output wire [511:0] col_541,
	output wire [511:0] col_542,
	output wire [511:0] col_543,
	output wire [511:0] col_544,
	output wire [511:0] col_545,
	output wire [511:0] col_546,
	output wire [511:0] col_547,
	output wire [511:0] col_548,
	output wire [511:0] col_549,
	output wire [511:0] col_550,
	output wire [511:0] col_551,
	output wire [511:0] col_552,
	output wire [511:0] col_553,
	output wire [511:0] col_554,
	output wire [511:0] col_555,
	output wire [511:0] col_556,
	output wire [511:0] col_557,
	output wire [511:0] col_558,
	output wire [511:0] col_559,
	output wire [511:0] col_560,
	output wire [511:0] col_561,
	output wire [511:0] col_562,
	output wire [511:0] col_563,
	output wire [511:0] col_564,
	output wire [511:0] col_565,
	output wire [511:0] col_566,
	output wire [511:0] col_567,
	output wire [511:0] col_568,
	output wire [511:0] col_569,
	output wire [511:0] col_570,
	output wire [511:0] col_571,
	output wire [511:0] col_572,
	output wire [511:0] col_573,
	output wire [511:0] col_574,
	output wire [511:0] col_575,
	output wire [511:0] col_576,
	output wire [511:0] col_577,
	output wire [511:0] col_578,
	output wire [511:0] col_579,
	output wire [511:0] col_580,
	output wire [511:0] col_581,
	output wire [511:0] col_582,
	output wire [511:0] col_583,
	output wire [511:0] col_584,
	output wire [511:0] col_585,
	output wire [511:0] col_586,
	output wire [511:0] col_587,
	output wire [511:0] col_588,
	output wire [511:0] col_589,
	output wire [511:0] col_590,
	output wire [511:0] col_591,
	output wire [511:0] col_592,
	output wire [511:0] col_593,
	output wire [511:0] col_594,
	output wire [511:0] col_595,
	output wire [511:0] col_596,
	output wire [511:0] col_597,
	output wire [511:0] col_598,
	output wire [511:0] col_599,
	output wire [511:0] col_600,
	output wire [511:0] col_601,
	output wire [511:0] col_602,
	output wire [511:0] col_603,
	output wire [511:0] col_604,
	output wire [511:0] col_605,
	output wire [511:0] col_606,
	output wire [511:0] col_607,
	output wire [511:0] col_608,
	output wire [511:0] col_609,
	output wire [511:0] col_610,
	output wire [511:0] col_611,
	output wire [511:0] col_612,
	output wire [511:0] col_613,
	output wire [511:0] col_614,
	output wire [511:0] col_615,
	output wire [511:0] col_616,
	output wire [511:0] col_617,
	output wire [511:0] col_618,
	output wire [511:0] col_619,
	output wire [511:0] col_620,
	output wire [511:0] col_621,
	output wire [511:0] col_622,
	output wire [511:0] col_623,
	output wire [511:0] col_624,
	output wire [511:0] col_625,
	output wire [511:0] col_626,
	output wire [511:0] col_627,
	output wire [511:0] col_628,
	output wire [511:0] col_629,
	output wire [511:0] col_630,
	output wire [511:0] col_631,
	output wire [511:0] col_632,
	output wire [511:0] col_633,
	output wire [511:0] col_634,
	output wire [511:0] col_635,
	output wire [511:0] col_636,
	output wire [511:0] col_637,
	output wire [511:0] col_638,
	output wire [511:0] col_639,
	output wire [511:0] col_640,
	output wire [511:0] col_641,
	output wire [511:0] col_642,
	output wire [511:0] col_643,
	output wire [511:0] col_644,
	output wire [511:0] col_645,
	output wire [511:0] col_646,
	output wire [511:0] col_647,
	output wire [511:0] col_648,
	output wire [511:0] col_649,
	output wire [511:0] col_650,
	output wire [511:0] col_651,
	output wire [511:0] col_652,
	output wire [511:0] col_653,
	output wire [511:0] col_654,
	output wire [511:0] col_655,
	output wire [511:0] col_656,
	output wire [511:0] col_657,
	output wire [511:0] col_658,
	output wire [511:0] col_659,
	output wire [511:0] col_660,
	output wire [511:0] col_661,
	output wire [511:0] col_662,
	output wire [511:0] col_663,
	output wire [511:0] col_664,
	output wire [511:0] col_665,
	output wire [511:0] col_666,
	output wire [511:0] col_667,
	output wire [511:0] col_668,
	output wire [511:0] col_669,
	output wire [511:0] col_670,
	output wire [511:0] col_671,
	output wire [511:0] col_672,
	output wire [511:0] col_673,
	output wire [511:0] col_674,
	output wire [511:0] col_675,
	output wire [511:0] col_676,
	output wire [511:0] col_677,
	output wire [511:0] col_678,
	output wire [511:0] col_679,
	output wire [511:0] col_680,
	output wire [511:0] col_681,
	output wire [511:0] col_682,
	output wire [511:0] col_683,
	output wire [511:0] col_684,
	output wire [511:0] col_685,
	output wire [511:0] col_686,
	output wire [511:0] col_687,
	output wire [511:0] col_688,
	output wire [511:0] col_689,
	output wire [511:0] col_690,
	output wire [511:0] col_691,
	output wire [511:0] col_692,
	output wire [511:0] col_693,
	output wire [511:0] col_694,
	output wire [511:0] col_695,
	output wire [511:0] col_696,
	output wire [511:0] col_697,
	output wire [511:0] col_698,
	output wire [511:0] col_699,
	output wire [511:0] col_700,
	output wire [511:0] col_701,
	output wire [511:0] col_702,
	output wire [511:0] col_703,
	output wire [511:0] col_704,
	output wire [511:0] col_705,
	output wire [511:0] col_706,
	output wire [511:0] col_707,
	output wire [511:0] col_708,
	output wire [511:0] col_709,
	output wire [511:0] col_710,
	output wire [511:0] col_711,
	output wire [511:0] col_712,
	output wire [511:0] col_713,
	output wire [511:0] col_714,
	output wire [511:0] col_715,
	output wire [511:0] col_716,
	output wire [511:0] col_717,
	output wire [511:0] col_718,
	output wire [511:0] col_719,
	output wire [511:0] col_720,
	output wire [511:0] col_721,
	output wire [511:0] col_722,
	output wire [511:0] col_723,
	output wire [511:0] col_724,
	output wire [511:0] col_725,
	output wire [511:0] col_726,
	output wire [511:0] col_727,
	output wire [511:0] col_728,
	output wire [511:0] col_729,
	output wire [511:0] col_730,
	output wire [511:0] col_731,
	output wire [511:0] col_732,
	output wire [511:0] col_733,
	output wire [511:0] col_734,
	output wire [511:0] col_735,
	output wire [511:0] col_736,
	output wire [511:0] col_737,
	output wire [511:0] col_738,
	output wire [511:0] col_739,
	output wire [511:0] col_740,
	output wire [511:0] col_741,
	output wire [511:0] col_742,
	output wire [511:0] col_743,
	output wire [511:0] col_744,
	output wire [511:0] col_745,
	output wire [511:0] col_746,
	output wire [511:0] col_747,
	output wire [511:0] col_748,
	output wire [511:0] col_749,
	output wire [511:0] col_750,
	output wire [511:0] col_751,
	output wire [511:0] col_752,
	output wire [511:0] col_753,
	output wire [511:0] col_754,
	output wire [511:0] col_755,
	output wire [511:0] col_756,
	output wire [511:0] col_757,
	output wire [511:0] col_758,
	output wire [511:0] col_759,
	output wire [511:0] col_760,
	output wire [511:0] col_761,
	output wire [511:0] col_762,
	output wire [511:0] col_763,
	output wire [511:0] col_764,
	output wire [511:0] col_765,
	output wire [511:0] col_766,
	output wire [511:0] col_767,
	output wire [511:0] col_768,
	output wire [511:0] col_769,
	output wire [511:0] col_770,
	output wire [511:0] col_771,
	output wire [511:0] col_772,
	output wire [511:0] col_773,
	output wire [511:0] col_774,
	output wire [511:0] col_775,
	output wire [511:0] col_776,
	output wire [511:0] col_777,
	output wire [511:0] col_778,
	output wire [511:0] col_779,
	output wire [511:0] col_780,
	output wire [511:0] col_781,
	output wire [511:0] col_782,
	output wire [511:0] col_783,
	output wire [511:0] col_784,
	output wire [511:0] col_785,
	output wire [511:0] col_786,
	output wire [511:0] col_787,
	output wire [511:0] col_788,
	output wire [511:0] col_789,
	output wire [511:0] col_790,
	output wire [511:0] col_791,
	output wire [511:0] col_792,
	output wire [511:0] col_793,
	output wire [511:0] col_794,
	output wire [511:0] col_795,
	output wire [511:0] col_796,
	output wire [511:0] col_797,
	output wire [511:0] col_798,
	output wire [511:0] col_799,
	output wire [511:0] col_800,
	output wire [511:0] col_801,
	output wire [511:0] col_802,
	output wire [511:0] col_803,
	output wire [511:0] col_804,
	output wire [511:0] col_805,
	output wire [511:0] col_806,
	output wire [511:0] col_807,
	output wire [511:0] col_808,
	output wire [511:0] col_809,
	output wire [511:0] col_810,
	output wire [511:0] col_811,
	output wire [511:0] col_812,
	output wire [511:0] col_813,
	output wire [511:0] col_814,
	output wire [511:0] col_815,
	output wire [511:0] col_816,
	output wire [511:0] col_817,
	output wire [511:0] col_818,
	output wire [511:0] col_819,
	output wire [511:0] col_820,
	output wire [511:0] col_821,
	output wire [511:0] col_822,
	output wire [511:0] col_823,
	output wire [511:0] col_824,
	output wire [511:0] col_825,
	output wire [511:0] col_826,
	output wire [511:0] col_827,
	output wire [511:0] col_828,
	output wire [511:0] col_829,
	output wire [511:0] col_830,
	output wire [511:0] col_831,
	output wire [511:0] col_832,
	output wire [511:0] col_833,
	output wire [511:0] col_834,
	output wire [511:0] col_835,
	output wire [511:0] col_836,
	output wire [511:0] col_837,
	output wire [511:0] col_838,
	output wire [511:0] col_839,
	output wire [511:0] col_840,
	output wire [511:0] col_841,
	output wire [511:0] col_842,
	output wire [511:0] col_843,
	output wire [511:0] col_844,
	output wire [511:0] col_845,
	output wire [511:0] col_846,
	output wire [511:0] col_847,
	output wire [511:0] col_848,
	output wire [511:0] col_849,
	output wire [511:0] col_850,
	output wire [511:0] col_851,
	output wire [511:0] col_852,
	output wire [511:0] col_853,
	output wire [511:0] col_854,
	output wire [511:0] col_855,
	output wire [511:0] col_856,
	output wire [511:0] col_857,
	output wire [511:0] col_858,
	output wire [511:0] col_859,
	output wire [511:0] col_860,
	output wire [511:0] col_861,
	output wire [511:0] col_862,
	output wire [511:0] col_863,
	output wire [511:0] col_864,
	output wire [511:0] col_865,
	output wire [511:0] col_866,
	output wire [511:0] col_867,
	output wire [511:0] col_868,
	output wire [511:0] col_869,
	output wire [511:0] col_870,
	output wire [511:0] col_871,
	output wire [511:0] col_872,
	output wire [511:0] col_873,
	output wire [511:0] col_874,
	output wire [511:0] col_875,
	output wire [511:0] col_876,
	output wire [511:0] col_877,
	output wire [511:0] col_878,
	output wire [511:0] col_879,
	output wire [511:0] col_880,
	output wire [511:0] col_881,
	output wire [511:0] col_882,
	output wire [511:0] col_883,
	output wire [511:0] col_884,
	output wire [511:0] col_885,
	output wire [511:0] col_886,
	output wire [511:0] col_887,
	output wire [511:0] col_888,
	output wire [511:0] col_889,
	output wire [511:0] col_890,
	output wire [511:0] col_891,
	output wire [511:0] col_892,
	output wire [511:0] col_893,
	output wire [511:0] col_894,
	output wire [511:0] col_895,
	output wire [511:0] col_896,
	output wire [511:0] col_897,
	output wire [511:0] col_898,
	output wire [511:0] col_899,
	output wire [511:0] col_900,
	output wire [511:0] col_901,
	output wire [511:0] col_902,
	output wire [511:0] col_903,
	output wire [511:0] col_904,
	output wire [511:0] col_905,
	output wire [511:0] col_906,
	output wire [511:0] col_907,
	output wire [511:0] col_908,
	output wire [511:0] col_909,
	output wire [511:0] col_910,
	output wire [511:0] col_911,
	output wire [511:0] col_912,
	output wire [511:0] col_913,
	output wire [511:0] col_914,
	output wire [511:0] col_915,
	output wire [511:0] col_916,
	output wire [511:0] col_917,
	output wire [511:0] col_918,
	output wire [511:0] col_919,
	output wire [511:0] col_920,
	output wire [511:0] col_921,
	output wire [511:0] col_922,
	output wire [511:0] col_923,
	output wire [511:0] col_924,
	output wire [511:0] col_925,
	output wire [511:0] col_926,
	output wire [511:0] col_927,
	output wire [511:0] col_928,
	output wire [511:0] col_929,
	output wire [511:0] col_930,
	output wire [511:0] col_931,
	output wire [511:0] col_932,
	output wire [511:0] col_933,
	output wire [511:0] col_934,
	output wire [511:0] col_935,
	output wire [511:0] col_936,
	output wire [511:0] col_937,
	output wire [511:0] col_938,
	output wire [511:0] col_939,
	output wire [511:0] col_940,
	output wire [511:0] col_941,
	output wire [511:0] col_942,
	output wire [511:0] col_943,
	output wire [511:0] col_944,
	output wire [511:0] col_945,
	output wire [511:0] col_946,
	output wire [511:0] col_947,
	output wire [511:0] col_948,
	output wire [511:0] col_949,
	output wire [511:0] col_950,
	output wire [511:0] col_951,
	output wire [511:0] col_952,
	output wire [511:0] col_953,
	output wire [511:0] col_954,
	output wire [511:0] col_955,
	output wire [511:0] col_956,
	output wire [511:0] col_957,
	output wire [511:0] col_958,
	output wire [511:0] col_959,
	output wire [511:0] col_960,
	output wire [511:0] col_961,
	output wire [511:0] col_962,
	output wire [511:0] col_963,
	output wire [511:0] col_964,
	output wire [511:0] col_965,
	output wire [511:0] col_966,
	output wire [511:0] col_967,
	output wire [511:0] col_968,
	output wire [511:0] col_969,
	output wire [511:0] col_970,
	output wire [511:0] col_971,
	output wire [511:0] col_972,
	output wire [511:0] col_973,
	output wire [511:0] col_974,
	output wire [511:0] col_975,
	output wire [511:0] col_976,
	output wire [511:0] col_977,
	output wire [511:0] col_978,
	output wire [511:0] col_979,
	output wire [511:0] col_980,
	output wire [511:0] col_981,
	output wire [511:0] col_982,
	output wire [511:0] col_983,
	output wire [511:0] col_984,
	output wire [511:0] col_985,
	output wire [511:0] col_986,
	output wire [511:0] col_987,
	output wire [511:0] col_988,
	output wire [511:0] col_989,
	output wire [511:0] col_990,
	output wire [511:0] col_991,
	output wire [511:0] col_992,
	output wire [511:0] col_993,
	output wire [511:0] col_994,
	output wire [511:0] col_995,
	output wire [511:0] col_996,
	output wire [511:0] col_997,
	output wire [511:0] col_998,
	output wire [511:0] col_999,
	output wire [511:0] col_1000,
	output wire [511:0] col_1001,
	output wire [511:0] col_1002,
	output wire [511:0] col_1003,
	output wire [511:0] col_1004,
	output wire [511:0] col_1005,
	output wire [511:0] col_1006,
	output wire [511:0] col_1007,
	output wire [511:0] col_1008,
	output wire [511:0] col_1009,
	output wire [511:0] col_1010,
	output wire [511:0] col_1011,
	output wire [511:0] col_1012,
	output wire [511:0] col_1013,
	output wire [511:0] col_1014,
	output wire [511:0] col_1015,
	output wire [511:0] col_1016,
	output wire [511:0] col_1017,
	output wire [511:0] col_1018,
	output wire [511:0] col_1019,
	output wire [511:0] col_1020,
	output wire [511:0] col_1021,
	output wire [511:0] col_1022,
	output wire [511:0] col_1023
);


wire [1023:0] ta;

wire [510:0] t_col_2;
wire [510:0] t_col_3;
wire [510:0] t_col_4;
wire [510:0] t_col_5;
wire [510:0] t_col_6;
wire [510:0] t_col_7;
wire [510:0] t_col_8;
wire [510:0] t_col_9;
wire [510:0] t_col_10;
wire [510:0] t_col_11;
wire [510:0] t_col_12;
wire [510:0] t_col_13;
wire [510:0] t_col_14;
wire [510:0] t_col_15;
wire [510:0] t_col_16;
wire [510:0] t_col_17;
wire [510:0] t_col_18;
wire [510:0] t_col_19;
wire [510:0] t_col_20;
wire [510:0] t_col_21;
wire [510:0] t_col_22;
wire [510:0] t_col_23;
wire [510:0] t_col_24;
wire [510:0] t_col_25;
wire [510:0] t_col_26;
wire [510:0] t_col_27;
wire [510:0] t_col_28;
wire [510:0] t_col_29;
wire [510:0] t_col_30;
wire [510:0] t_col_31;
wire [510:0] t_col_32;
wire [510:0] t_col_33;
wire [510:0] t_col_34;
wire [510:0] t_col_35;
wire [510:0] t_col_36;
wire [510:0] t_col_37;
wire [510:0] t_col_38;
wire [510:0] t_col_39;
wire [510:0] t_col_40;
wire [510:0] t_col_41;
wire [510:0] t_col_42;
wire [510:0] t_col_43;
wire [510:0] t_col_44;
wire [510:0] t_col_45;
wire [510:0] t_col_46;
wire [510:0] t_col_47;
wire [510:0] t_col_48;
wire [510:0] t_col_49;
wire [510:0] t_col_50;
wire [510:0] t_col_51;
wire [510:0] t_col_52;
wire [510:0] t_col_53;
wire [510:0] t_col_54;
wire [510:0] t_col_55;
wire [510:0] t_col_56;
wire [510:0] t_col_57;
wire [510:0] t_col_58;
wire [510:0] t_col_59;
wire [510:0] t_col_60;
wire [510:0] t_col_61;
wire [510:0] t_col_62;
wire [510:0] t_col_63;
wire [510:0] t_col_64;
wire [510:0] t_col_65;
wire [510:0] t_col_66;
wire [510:0] t_col_67;
wire [510:0] t_col_68;
wire [510:0] t_col_69;
wire [510:0] t_col_70;
wire [510:0] t_col_71;
wire [510:0] t_col_72;
wire [510:0] t_col_73;
wire [510:0] t_col_74;
wire [510:0] t_col_75;
wire [510:0] t_col_76;
wire [510:0] t_col_77;
wire [510:0] t_col_78;
wire [510:0] t_col_79;
wire [510:0] t_col_80;
wire [510:0] t_col_81;
wire [510:0] t_col_82;
wire [510:0] t_col_83;
wire [510:0] t_col_84;
wire [510:0] t_col_85;
wire [510:0] t_col_86;
wire [510:0] t_col_87;
wire [510:0] t_col_88;
wire [510:0] t_col_89;
wire [510:0] t_col_90;
wire [510:0] t_col_91;
wire [510:0] t_col_92;
wire [510:0] t_col_93;
wire [510:0] t_col_94;
wire [510:0] t_col_95;
wire [510:0] t_col_96;
wire [510:0] t_col_97;
wire [510:0] t_col_98;
wire [510:0] t_col_99;
wire [510:0] t_col_100;
wire [510:0] t_col_101;
wire [510:0] t_col_102;
wire [510:0] t_col_103;
wire [510:0] t_col_104;
wire [510:0] t_col_105;
wire [510:0] t_col_106;
wire [510:0] t_col_107;
wire [510:0] t_col_108;
wire [510:0] t_col_109;
wire [510:0] t_col_110;
wire [510:0] t_col_111;
wire [510:0] t_col_112;
wire [510:0] t_col_113;
wire [510:0] t_col_114;
wire [510:0] t_col_115;
wire [510:0] t_col_116;
wire [510:0] t_col_117;
wire [510:0] t_col_118;
wire [510:0] t_col_119;
wire [510:0] t_col_120;
wire [510:0] t_col_121;
wire [510:0] t_col_122;
wire [510:0] t_col_123;
wire [510:0] t_col_124;
wire [510:0] t_col_125;
wire [510:0] t_col_126;
wire [510:0] t_col_127;
wire [510:0] t_col_128;
wire [510:0] t_col_129;
wire [510:0] t_col_130;
wire [510:0] t_col_131;
wire [510:0] t_col_132;
wire [510:0] t_col_133;
wire [510:0] t_col_134;
wire [510:0] t_col_135;
wire [510:0] t_col_136;
wire [510:0] t_col_137;
wire [510:0] t_col_138;
wire [510:0] t_col_139;
wire [510:0] t_col_140;
wire [510:0] t_col_141;
wire [510:0] t_col_142;
wire [510:0] t_col_143;
wire [510:0] t_col_144;
wire [510:0] t_col_145;
wire [510:0] t_col_146;
wire [510:0] t_col_147;
wire [510:0] t_col_148;
wire [510:0] t_col_149;
wire [510:0] t_col_150;
wire [510:0] t_col_151;
wire [510:0] t_col_152;
wire [510:0] t_col_153;
wire [510:0] t_col_154;
wire [510:0] t_col_155;
wire [510:0] t_col_156;
wire [510:0] t_col_157;
wire [510:0] t_col_158;
wire [510:0] t_col_159;
wire [510:0] t_col_160;
wire [510:0] t_col_161;
wire [510:0] t_col_162;
wire [510:0] t_col_163;
wire [510:0] t_col_164;
wire [510:0] t_col_165;
wire [510:0] t_col_166;
wire [510:0] t_col_167;
wire [510:0] t_col_168;
wire [510:0] t_col_169;
wire [510:0] t_col_170;
wire [510:0] t_col_171;
wire [510:0] t_col_172;
wire [510:0] t_col_173;
wire [510:0] t_col_174;
wire [510:0] t_col_175;
wire [510:0] t_col_176;
wire [510:0] t_col_177;
wire [510:0] t_col_178;
wire [510:0] t_col_179;
wire [510:0] t_col_180;
wire [510:0] t_col_181;
wire [510:0] t_col_182;
wire [510:0] t_col_183;
wire [510:0] t_col_184;
wire [510:0] t_col_185;
wire [510:0] t_col_186;
wire [510:0] t_col_187;
wire [510:0] t_col_188;
wire [510:0] t_col_189;
wire [510:0] t_col_190;
wire [510:0] t_col_191;
wire [510:0] t_col_192;
wire [510:0] t_col_193;
wire [510:0] t_col_194;
wire [510:0] t_col_195;
wire [510:0] t_col_196;
wire [510:0] t_col_197;
wire [510:0] t_col_198;
wire [510:0] t_col_199;
wire [510:0] t_col_200;
wire [510:0] t_col_201;
wire [510:0] t_col_202;
wire [510:0] t_col_203;
wire [510:0] t_col_204;
wire [510:0] t_col_205;
wire [510:0] t_col_206;
wire [510:0] t_col_207;
wire [510:0] t_col_208;
wire [510:0] t_col_209;
wire [510:0] t_col_210;
wire [510:0] t_col_211;
wire [510:0] t_col_212;
wire [510:0] t_col_213;
wire [510:0] t_col_214;
wire [510:0] t_col_215;
wire [510:0] t_col_216;
wire [510:0] t_col_217;
wire [510:0] t_col_218;
wire [510:0] t_col_219;
wire [510:0] t_col_220;
wire [510:0] t_col_221;
wire [510:0] t_col_222;
wire [510:0] t_col_223;
wire [510:0] t_col_224;
wire [510:0] t_col_225;
wire [510:0] t_col_226;
wire [510:0] t_col_227;
wire [510:0] t_col_228;
wire [510:0] t_col_229;
wire [510:0] t_col_230;
wire [510:0] t_col_231;
wire [510:0] t_col_232;
wire [510:0] t_col_233;
wire [510:0] t_col_234;
wire [510:0] t_col_235;
wire [510:0] t_col_236;
wire [510:0] t_col_237;
wire [510:0] t_col_238;
wire [510:0] t_col_239;
wire [510:0] t_col_240;
wire [510:0] t_col_241;
wire [510:0] t_col_242;
wire [510:0] t_col_243;
wire [510:0] t_col_244;
wire [510:0] t_col_245;
wire [510:0] t_col_246;
wire [510:0] t_col_247;
wire [510:0] t_col_248;
wire [510:0] t_col_249;
wire [510:0] t_col_250;
wire [510:0] t_col_251;
wire [510:0] t_col_252;
wire [510:0] t_col_253;
wire [510:0] t_col_254;
wire [510:0] t_col_255;
wire [510:0] t_col_256;
wire [510:0] t_col_257;
wire [510:0] t_col_258;
wire [510:0] t_col_259;
wire [510:0] t_col_260;
wire [510:0] t_col_261;
wire [510:0] t_col_262;
wire [510:0] t_col_263;
wire [510:0] t_col_264;
wire [510:0] t_col_265;
wire [510:0] t_col_266;
wire [510:0] t_col_267;
wire [510:0] t_col_268;
wire [510:0] t_col_269;
wire [510:0] t_col_270;
wire [510:0] t_col_271;
wire [510:0] t_col_272;
wire [510:0] t_col_273;
wire [510:0] t_col_274;
wire [510:0] t_col_275;
wire [510:0] t_col_276;
wire [510:0] t_col_277;
wire [510:0] t_col_278;
wire [510:0] t_col_279;
wire [510:0] t_col_280;
wire [510:0] t_col_281;
wire [510:0] t_col_282;
wire [510:0] t_col_283;
wire [510:0] t_col_284;
wire [510:0] t_col_285;
wire [510:0] t_col_286;
wire [510:0] t_col_287;
wire [510:0] t_col_288;
wire [510:0] t_col_289;
wire [510:0] t_col_290;
wire [510:0] t_col_291;
wire [510:0] t_col_292;
wire [510:0] t_col_293;
wire [510:0] t_col_294;
wire [510:0] t_col_295;
wire [510:0] t_col_296;
wire [510:0] t_col_297;
wire [510:0] t_col_298;
wire [510:0] t_col_299;
wire [510:0] t_col_300;
wire [510:0] t_col_301;
wire [510:0] t_col_302;
wire [510:0] t_col_303;
wire [510:0] t_col_304;
wire [510:0] t_col_305;
wire [510:0] t_col_306;
wire [510:0] t_col_307;
wire [510:0] t_col_308;
wire [510:0] t_col_309;
wire [510:0] t_col_310;
wire [510:0] t_col_311;
wire [510:0] t_col_312;
wire [510:0] t_col_313;
wire [510:0] t_col_314;
wire [510:0] t_col_315;
wire [510:0] t_col_316;
wire [510:0] t_col_317;
wire [510:0] t_col_318;
wire [510:0] t_col_319;
wire [510:0] t_col_320;
wire [510:0] t_col_321;
wire [510:0] t_col_322;
wire [510:0] t_col_323;
wire [510:0] t_col_324;
wire [510:0] t_col_325;
wire [510:0] t_col_326;
wire [510:0] t_col_327;
wire [510:0] t_col_328;
wire [510:0] t_col_329;
wire [510:0] t_col_330;
wire [510:0] t_col_331;
wire [510:0] t_col_332;
wire [510:0] t_col_333;
wire [510:0] t_col_334;
wire [510:0] t_col_335;
wire [510:0] t_col_336;
wire [510:0] t_col_337;
wire [510:0] t_col_338;
wire [510:0] t_col_339;
wire [510:0] t_col_340;
wire [510:0] t_col_341;
wire [510:0] t_col_342;
wire [510:0] t_col_343;
wire [510:0] t_col_344;
wire [510:0] t_col_345;
wire [510:0] t_col_346;
wire [510:0] t_col_347;
wire [510:0] t_col_348;
wire [510:0] t_col_349;
wire [510:0] t_col_350;
wire [510:0] t_col_351;
wire [510:0] t_col_352;
wire [510:0] t_col_353;
wire [510:0] t_col_354;
wire [510:0] t_col_355;
wire [510:0] t_col_356;
wire [510:0] t_col_357;
wire [510:0] t_col_358;
wire [510:0] t_col_359;
wire [510:0] t_col_360;
wire [510:0] t_col_361;
wire [510:0] t_col_362;
wire [510:0] t_col_363;
wire [510:0] t_col_364;
wire [510:0] t_col_365;
wire [510:0] t_col_366;
wire [510:0] t_col_367;
wire [510:0] t_col_368;
wire [510:0] t_col_369;
wire [510:0] t_col_370;
wire [510:0] t_col_371;
wire [510:0] t_col_372;
wire [510:0] t_col_373;
wire [510:0] t_col_374;
wire [510:0] t_col_375;
wire [510:0] t_col_376;
wire [510:0] t_col_377;
wire [510:0] t_col_378;
wire [510:0] t_col_379;
wire [510:0] t_col_380;
wire [510:0] t_col_381;
wire [510:0] t_col_382;
wire [510:0] t_col_383;
wire [510:0] t_col_384;
wire [510:0] t_col_385;
wire [510:0] t_col_386;
wire [510:0] t_col_387;
wire [510:0] t_col_388;
wire [510:0] t_col_389;
wire [510:0] t_col_390;
wire [510:0] t_col_391;
wire [510:0] t_col_392;
wire [510:0] t_col_393;
wire [510:0] t_col_394;
wire [510:0] t_col_395;
wire [510:0] t_col_396;
wire [510:0] t_col_397;
wire [510:0] t_col_398;
wire [510:0] t_col_399;
wire [510:0] t_col_400;
wire [510:0] t_col_401;
wire [510:0] t_col_402;
wire [510:0] t_col_403;
wire [510:0] t_col_404;
wire [510:0] t_col_405;
wire [510:0] t_col_406;
wire [510:0] t_col_407;
wire [510:0] t_col_408;
wire [510:0] t_col_409;
wire [510:0] t_col_410;
wire [510:0] t_col_411;
wire [510:0] t_col_412;
wire [510:0] t_col_413;
wire [510:0] t_col_414;
wire [510:0] t_col_415;
wire [510:0] t_col_416;
wire [510:0] t_col_417;
wire [510:0] t_col_418;
wire [510:0] t_col_419;
wire [510:0] t_col_420;
wire [510:0] t_col_421;
wire [510:0] t_col_422;
wire [510:0] t_col_423;
wire [510:0] t_col_424;
wire [510:0] t_col_425;
wire [510:0] t_col_426;
wire [510:0] t_col_427;
wire [510:0] t_col_428;
wire [510:0] t_col_429;
wire [510:0] t_col_430;
wire [510:0] t_col_431;
wire [510:0] t_col_432;
wire [510:0] t_col_433;
wire [510:0] t_col_434;
wire [510:0] t_col_435;
wire [510:0] t_col_436;
wire [510:0] t_col_437;
wire [510:0] t_col_438;
wire [510:0] t_col_439;
wire [510:0] t_col_440;
wire [510:0] t_col_441;
wire [510:0] t_col_442;
wire [510:0] t_col_443;
wire [510:0] t_col_444;
wire [510:0] t_col_445;
wire [510:0] t_col_446;
wire [510:0] t_col_447;
wire [510:0] t_col_448;
wire [510:0] t_col_449;
wire [510:0] t_col_450;
wire [510:0] t_col_451;
wire [510:0] t_col_452;
wire [510:0] t_col_453;
wire [510:0] t_col_454;
wire [510:0] t_col_455;
wire [510:0] t_col_456;
wire [510:0] t_col_457;
wire [510:0] t_col_458;
wire [510:0] t_col_459;
wire [510:0] t_col_460;
wire [510:0] t_col_461;
wire [510:0] t_col_462;
wire [510:0] t_col_463;
wire [510:0] t_col_464;
wire [510:0] t_col_465;
wire [510:0] t_col_466;
wire [510:0] t_col_467;
wire [510:0] t_col_468;
wire [510:0] t_col_469;
wire [510:0] t_col_470;
wire [510:0] t_col_471;
wire [510:0] t_col_472;
wire [510:0] t_col_473;
wire [510:0] t_col_474;
wire [510:0] t_col_475;
wire [510:0] t_col_476;
wire [510:0] t_col_477;
wire [510:0] t_col_478;
wire [510:0] t_col_479;
wire [510:0] t_col_480;
wire [510:0] t_col_481;
wire [510:0] t_col_482;
wire [510:0] t_col_483;
wire [510:0] t_col_484;
wire [510:0] t_col_485;
wire [510:0] t_col_486;
wire [510:0] t_col_487;
wire [510:0] t_col_488;
wire [510:0] t_col_489;
wire [510:0] t_col_490;
wire [510:0] t_col_491;
wire [510:0] t_col_492;
wire [510:0] t_col_493;
wire [510:0] t_col_494;
wire [510:0] t_col_495;
wire [510:0] t_col_496;
wire [510:0] t_col_497;
wire [510:0] t_col_498;
wire [510:0] t_col_499;
wire [510:0] t_col_500;
wire [510:0] t_col_501;
wire [510:0] t_col_502;
wire [510:0] t_col_503;
wire [510:0] t_col_504;
wire [510:0] t_col_505;
wire [510:0] t_col_506;
wire [510:0] t_col_507;
wire [510:0] t_col_508;
wire [510:0] t_col_509;
wire [510:0] t_col_510;
wire [510:0] t_col_511;
wire [510:0] t_col_512;
wire [510:0] t_col_513;
wire [510:0] t_col_514;
wire [510:0] t_col_515;
wire [510:0] t_col_516;
wire [510:0] t_col_517;
wire [510:0] t_col_518;
wire [510:0] t_col_519;
wire [510:0] t_col_520;
wire [510:0] t_col_521;
wire [510:0] t_col_522;
wire [510:0] t_col_523;
wire [510:0] t_col_524;
wire [510:0] t_col_525;
wire [510:0] t_col_526;
wire [510:0] t_col_527;
wire [510:0] t_col_528;
wire [510:0] t_col_529;
wire [510:0] t_col_530;
wire [510:0] t_col_531;
wire [510:0] t_col_532;
wire [510:0] t_col_533;
wire [510:0] t_col_534;
wire [510:0] t_col_535;
wire [510:0] t_col_536;
wire [510:0] t_col_537;
wire [510:0] t_col_538;
wire [510:0] t_col_539;
wire [510:0] t_col_540;
wire [510:0] t_col_541;
wire [510:0] t_col_542;
wire [510:0] t_col_543;
wire [510:0] t_col_544;
wire [510:0] t_col_545;
wire [510:0] t_col_546;
wire [510:0] t_col_547;
wire [510:0] t_col_548;
wire [510:0] t_col_549;
wire [510:0] t_col_550;
wire [510:0] t_col_551;
wire [510:0] t_col_552;
wire [510:0] t_col_553;
wire [510:0] t_col_554;
wire [510:0] t_col_555;
wire [510:0] t_col_556;
wire [510:0] t_col_557;
wire [510:0] t_col_558;
wire [510:0] t_col_559;
wire [510:0] t_col_560;
wire [510:0] t_col_561;
wire [510:0] t_col_562;
wire [510:0] t_col_563;
wire [510:0] t_col_564;
wire [510:0] t_col_565;
wire [510:0] t_col_566;
wire [510:0] t_col_567;
wire [510:0] t_col_568;
wire [510:0] t_col_569;
wire [510:0] t_col_570;
wire [510:0] t_col_571;
wire [510:0] t_col_572;
wire [510:0] t_col_573;
wire [510:0] t_col_574;
wire [510:0] t_col_575;
wire [510:0] t_col_576;
wire [510:0] t_col_577;
wire [510:0] t_col_578;
wire [510:0] t_col_579;
wire [510:0] t_col_580;
wire [510:0] t_col_581;
wire [510:0] t_col_582;
wire [510:0] t_col_583;
wire [510:0] t_col_584;
wire [510:0] t_col_585;
wire [510:0] t_col_586;
wire [510:0] t_col_587;
wire [510:0] t_col_588;
wire [510:0] t_col_589;
wire [510:0] t_col_590;
wire [510:0] t_col_591;
wire [510:0] t_col_592;
wire [510:0] t_col_593;
wire [510:0] t_col_594;
wire [510:0] t_col_595;
wire [510:0] t_col_596;
wire [510:0] t_col_597;
wire [510:0] t_col_598;
wire [510:0] t_col_599;
wire [510:0] t_col_600;
wire [510:0] t_col_601;
wire [510:0] t_col_602;
wire [510:0] t_col_603;
wire [510:0] t_col_604;
wire [510:0] t_col_605;
wire [510:0] t_col_606;
wire [510:0] t_col_607;
wire [510:0] t_col_608;
wire [510:0] t_col_609;
wire [510:0] t_col_610;
wire [510:0] t_col_611;
wire [510:0] t_col_612;
wire [510:0] t_col_613;
wire [510:0] t_col_614;
wire [510:0] t_col_615;
wire [510:0] t_col_616;
wire [510:0] t_col_617;
wire [510:0] t_col_618;
wire [510:0] t_col_619;
wire [510:0] t_col_620;
wire [510:0] t_col_621;
wire [510:0] t_col_622;
wire [510:0] t_col_623;
wire [510:0] t_col_624;
wire [510:0] t_col_625;
wire [510:0] t_col_626;
wire [510:0] t_col_627;
wire [510:0] t_col_628;
wire [510:0] t_col_629;
wire [510:0] t_col_630;
wire [510:0] t_col_631;
wire [510:0] t_col_632;
wire [510:0] t_col_633;
wire [510:0] t_col_634;
wire [510:0] t_col_635;
wire [510:0] t_col_636;
wire [510:0] t_col_637;
wire [510:0] t_col_638;
wire [510:0] t_col_639;
wire [510:0] t_col_640;
wire [510:0] t_col_641;
wire [510:0] t_col_642;
wire [510:0] t_col_643;
wire [510:0] t_col_644;
wire [510:0] t_col_645;
wire [510:0] t_col_646;
wire [510:0] t_col_647;
wire [510:0] t_col_648;
wire [510:0] t_col_649;
wire [510:0] t_col_650;
wire [510:0] t_col_651;
wire [510:0] t_col_652;
wire [510:0] t_col_653;
wire [510:0] t_col_654;
wire [510:0] t_col_655;
wire [510:0] t_col_656;
wire [510:0] t_col_657;
wire [510:0] t_col_658;
wire [510:0] t_col_659;
wire [510:0] t_col_660;
wire [510:0] t_col_661;
wire [510:0] t_col_662;
wire [510:0] t_col_663;
wire [510:0] t_col_664;
wire [510:0] t_col_665;
wire [510:0] t_col_666;
wire [510:0] t_col_667;
wire [510:0] t_col_668;
wire [510:0] t_col_669;
wire [510:0] t_col_670;
wire [510:0] t_col_671;
wire [510:0] t_col_672;
wire [510:0] t_col_673;
wire [510:0] t_col_674;
wire [510:0] t_col_675;
wire [510:0] t_col_676;
wire [510:0] t_col_677;
wire [510:0] t_col_678;
wire [510:0] t_col_679;
wire [510:0] t_col_680;
wire [510:0] t_col_681;
wire [510:0] t_col_682;
wire [510:0] t_col_683;
wire [510:0] t_col_684;
wire [510:0] t_col_685;
wire [510:0] t_col_686;
wire [510:0] t_col_687;
wire [510:0] t_col_688;
wire [510:0] t_col_689;
wire [510:0] t_col_690;
wire [510:0] t_col_691;
wire [510:0] t_col_692;
wire [510:0] t_col_693;
wire [510:0] t_col_694;
wire [510:0] t_col_695;
wire [510:0] t_col_696;
wire [510:0] t_col_697;
wire [510:0] t_col_698;
wire [510:0] t_col_699;
wire [510:0] t_col_700;
wire [510:0] t_col_701;
wire [510:0] t_col_702;
wire [510:0] t_col_703;
wire [510:0] t_col_704;
wire [510:0] t_col_705;
wire [510:0] t_col_706;
wire [510:0] t_col_707;
wire [510:0] t_col_708;
wire [510:0] t_col_709;
wire [510:0] t_col_710;
wire [510:0] t_col_711;
wire [510:0] t_col_712;
wire [510:0] t_col_713;
wire [510:0] t_col_714;
wire [510:0] t_col_715;
wire [510:0] t_col_716;
wire [510:0] t_col_717;
wire [510:0] t_col_718;
wire [510:0] t_col_719;
wire [510:0] t_col_720;
wire [510:0] t_col_721;
wire [510:0] t_col_722;
wire [510:0] t_col_723;
wire [510:0] t_col_724;
wire [510:0] t_col_725;
wire [510:0] t_col_726;
wire [510:0] t_col_727;
wire [510:0] t_col_728;
wire [510:0] t_col_729;
wire [510:0] t_col_730;
wire [510:0] t_col_731;
wire [510:0] t_col_732;
wire [510:0] t_col_733;
wire [510:0] t_col_734;
wire [510:0] t_col_735;
wire [510:0] t_col_736;
wire [510:0] t_col_737;
wire [510:0] t_col_738;
wire [510:0] t_col_739;
wire [510:0] t_col_740;
wire [510:0] t_col_741;
wire [510:0] t_col_742;
wire [510:0] t_col_743;
wire [510:0] t_col_744;
wire [510:0] t_col_745;
wire [510:0] t_col_746;
wire [510:0] t_col_747;
wire [510:0] t_col_748;
wire [510:0] t_col_749;
wire [510:0] t_col_750;
wire [510:0] t_col_751;
wire [510:0] t_col_752;
wire [510:0] t_col_753;
wire [510:0] t_col_754;
wire [510:0] t_col_755;
wire [510:0] t_col_756;
wire [510:0] t_col_757;
wire [510:0] t_col_758;
wire [510:0] t_col_759;
wire [510:0] t_col_760;
wire [510:0] t_col_761;
wire [510:0] t_col_762;
wire [510:0] t_col_763;
wire [510:0] t_col_764;
wire [510:0] t_col_765;
wire [510:0] t_col_766;
wire [510:0] t_col_767;
wire [510:0] t_col_768;
wire [510:0] t_col_769;
wire [510:0] t_col_770;
wire [510:0] t_col_771;
wire [510:0] t_col_772;
wire [510:0] t_col_773;
wire [510:0] t_col_774;
wire [510:0] t_col_775;
wire [510:0] t_col_776;
wire [510:0] t_col_777;
wire [510:0] t_col_778;
wire [510:0] t_col_779;
wire [510:0] t_col_780;
wire [510:0] t_col_781;
wire [510:0] t_col_782;
wire [510:0] t_col_783;
wire [510:0] t_col_784;
wire [510:0] t_col_785;
wire [510:0] t_col_786;
wire [510:0] t_col_787;
wire [510:0] t_col_788;
wire [510:0] t_col_789;
wire [510:0] t_col_790;
wire [510:0] t_col_791;
wire [510:0] t_col_792;
wire [510:0] t_col_793;
wire [510:0] t_col_794;
wire [510:0] t_col_795;
wire [510:0] t_col_796;
wire [510:0] t_col_797;
wire [510:0] t_col_798;
wire [510:0] t_col_799;
wire [510:0] t_col_800;
wire [510:0] t_col_801;
wire [510:0] t_col_802;
wire [510:0] t_col_803;
wire [510:0] t_col_804;
wire [510:0] t_col_805;
wire [510:0] t_col_806;
wire [510:0] t_col_807;
wire [510:0] t_col_808;
wire [510:0] t_col_809;
wire [510:0] t_col_810;
wire [510:0] t_col_811;
wire [510:0] t_col_812;
wire [510:0] t_col_813;
wire [510:0] t_col_814;
wire [510:0] t_col_815;
wire [510:0] t_col_816;
wire [510:0] t_col_817;
wire [510:0] t_col_818;
wire [510:0] t_col_819;
wire [510:0] t_col_820;
wire [510:0] t_col_821;
wire [510:0] t_col_822;
wire [510:0] t_col_823;
wire [510:0] t_col_824;
wire [510:0] t_col_825;
wire [510:0] t_col_826;
wire [510:0] t_col_827;
wire [510:0] t_col_828;
wire [510:0] t_col_829;
wire [510:0] t_col_830;
wire [510:0] t_col_831;
wire [510:0] t_col_832;
wire [510:0] t_col_833;
wire [510:0] t_col_834;
wire [510:0] t_col_835;
wire [510:0] t_col_836;
wire [510:0] t_col_837;
wire [510:0] t_col_838;
wire [510:0] t_col_839;
wire [510:0] t_col_840;
wire [510:0] t_col_841;
wire [510:0] t_col_842;
wire [510:0] t_col_843;
wire [510:0] t_col_844;
wire [510:0] t_col_845;
wire [510:0] t_col_846;
wire [510:0] t_col_847;
wire [510:0] t_col_848;
wire [510:0] t_col_849;
wire [510:0] t_col_850;
wire [510:0] t_col_851;
wire [510:0] t_col_852;
wire [510:0] t_col_853;
wire [510:0] t_col_854;
wire [510:0] t_col_855;
wire [510:0] t_col_856;
wire [510:0] t_col_857;
wire [510:0] t_col_858;
wire [510:0] t_col_859;
wire [510:0] t_col_860;
wire [510:0] t_col_861;
wire [510:0] t_col_862;
wire [510:0] t_col_863;
wire [510:0] t_col_864;
wire [510:0] t_col_865;
wire [510:0] t_col_866;
wire [510:0] t_col_867;
wire [510:0] t_col_868;
wire [510:0] t_col_869;
wire [510:0] t_col_870;
wire [510:0] t_col_871;
wire [510:0] t_col_872;
wire [510:0] t_col_873;
wire [510:0] t_col_874;
wire [510:0] t_col_875;
wire [510:0] t_col_876;
wire [510:0] t_col_877;
wire [510:0] t_col_878;
wire [510:0] t_col_879;
wire [510:0] t_col_880;
wire [510:0] t_col_881;
wire [510:0] t_col_882;
wire [510:0] t_col_883;
wire [510:0] t_col_884;
wire [510:0] t_col_885;
wire [510:0] t_col_886;
wire [510:0] t_col_887;
wire [510:0] t_col_888;
wire [510:0] t_col_889;
wire [510:0] t_col_890;
wire [510:0] t_col_891;
wire [510:0] t_col_892;
wire [510:0] t_col_893;
wire [510:0] t_col_894;
wire [510:0] t_col_895;
wire [510:0] t_col_896;
wire [510:0] t_col_897;
wire [510:0] t_col_898;
wire [510:0] t_col_899;
wire [510:0] t_col_900;
wire [510:0] t_col_901;
wire [510:0] t_col_902;
wire [510:0] t_col_903;
wire [510:0] t_col_904;
wire [510:0] t_col_905;
wire [510:0] t_col_906;
wire [510:0] t_col_907;
wire [510:0] t_col_908;
wire [510:0] t_col_909;
wire [510:0] t_col_910;
wire [510:0] t_col_911;
wire [510:0] t_col_912;
wire [510:0] t_col_913;
wire [510:0] t_col_914;
wire [510:0] t_col_915;
wire [510:0] t_col_916;
wire [510:0] t_col_917;
wire [510:0] t_col_918;
wire [510:0] t_col_919;
wire [510:0] t_col_920;
wire [510:0] t_col_921;
wire [510:0] t_col_922;
wire [510:0] t_col_923;
wire [510:0] t_col_924;
wire [510:0] t_col_925;
wire [510:0] t_col_926;
wire [510:0] t_col_927;
wire [510:0] t_col_928;
wire [510:0] t_col_929;
wire [510:0] t_col_930;
wire [510:0] t_col_931;
wire [510:0] t_col_932;
wire [510:0] t_col_933;
wire [510:0] t_col_934;
wire [510:0] t_col_935;
wire [510:0] t_col_936;
wire [510:0] t_col_937;
wire [510:0] t_col_938;
wire [510:0] t_col_939;
wire [510:0] t_col_940;
wire [510:0] t_col_941;
wire [510:0] t_col_942;
wire [510:0] t_col_943;
wire [510:0] t_col_944;
wire [510:0] t_col_945;
wire [510:0] t_col_946;
wire [510:0] t_col_947;
wire [510:0] t_col_948;
wire [510:0] t_col_949;
wire [510:0] t_col_950;
wire [510:0] t_col_951;
wire [510:0] t_col_952;
wire [510:0] t_col_953;
wire [510:0] t_col_954;
wire [510:0] t_col_955;
wire [510:0] t_col_956;
wire [510:0] t_col_957;
wire [510:0] t_col_958;
wire [510:0] t_col_959;
wire [510:0] t_col_960;
wire [510:0] t_col_961;
wire [510:0] t_col_962;
wire [510:0] t_col_963;
wire [510:0] t_col_964;
wire [510:0] t_col_965;
wire [510:0] t_col_966;
wire [510:0] t_col_967;
wire [510:0] t_col_968;
wire [510:0] t_col_969;
wire [510:0] t_col_970;
wire [510:0] t_col_971;
wire [510:0] t_col_972;
wire [510:0] t_col_973;
wire [510:0] t_col_974;
wire [510:0] t_col_975;
wire [510:0] t_col_976;
wire [510:0] t_col_977;
wire [510:0] t_col_978;
wire [510:0] t_col_979;
wire [510:0] t_col_980;
wire [510:0] t_col_981;
wire [510:0] t_col_982;
wire [510:0] t_col_983;
wire [510:0] t_col_984;
wire [510:0] t_col_985;
wire [510:0] t_col_986;
wire [510:0] t_col_987;
wire [510:0] t_col_988;
wire [510:0] t_col_989;
wire [510:0] t_col_990;
wire [510:0] t_col_991;
wire [510:0] t_col_992;
wire [510:0] t_col_993;
wire [510:0] t_col_994;
wire [510:0] t_col_995;
wire [510:0] t_col_996;
wire [510:0] t_col_997;
wire [510:0] t_col_998;
wire [510:0] t_col_999;
wire [510:0] t_col_1000;
wire [510:0] t_col_1001;
wire [510:0] t_col_1002;
wire [510:0] t_col_1003;
wire [510:0] t_col_1004;
wire [510:0] t_col_1005;
wire [510:0] t_col_1006;
wire [510:0] t_col_1007;
wire [510:0] t_col_1008;
wire [510:0] t_col_1009;
wire [510:0] t_col_1010;
wire [510:0] t_col_1011;
wire [510:0] t_col_1012;
wire [510:0] t_col_1013;
wire [510:0] t_col_1014;
wire [510:0] t_col_1015;
wire [510:0] t_col_1016;
wire [510:0] t_col_1017;
wire [510:0] t_col_1018;
wire [510:0] t_col_1019;
wire [510:0] t_col_1020;
wire [510:0] t_col_1021;
wire [510:0] t_col_1022;
wire [510:0] t_col_1023;

msq_common_array msq_common_array (
	.a(ta),
	.col_2(t_col_2),
	.col_3(t_col_3),
	.col_4(t_col_4),
	.col_5(t_col_5),
	.col_6(t_col_6),
	.col_7(t_col_7),
	.col_8(t_col_8),
	.col_9(t_col_9),
	.col_10(t_col_10),
	.col_11(t_col_11),
	.col_12(t_col_12),
	.col_13(t_col_13),
	.col_14(t_col_14),
	.col_15(t_col_15),
	.col_16(t_col_16),
	.col_17(t_col_17),
	.col_18(t_col_18),
	.col_19(t_col_19),
	.col_20(t_col_20),
	.col_21(t_col_21),
	.col_22(t_col_22),
	.col_23(t_col_23),
	.col_24(t_col_24),
	.col_25(t_col_25),
	.col_26(t_col_26),
	.col_27(t_col_27),
	.col_28(t_col_28),
	.col_29(t_col_29),
	.col_30(t_col_30),
	.col_31(t_col_31),
	.col_32(t_col_32),
	.col_33(t_col_33),
	.col_34(t_col_34),
	.col_35(t_col_35),
	.col_36(t_col_36),
	.col_37(t_col_37),
	.col_38(t_col_38),
	.col_39(t_col_39),
	.col_40(t_col_40),
	.col_41(t_col_41),
	.col_42(t_col_42),
	.col_43(t_col_43),
	.col_44(t_col_44),
	.col_45(t_col_45),
	.col_46(t_col_46),
	.col_47(t_col_47),
	.col_48(t_col_48),
	.col_49(t_col_49),
	.col_50(t_col_50),
	.col_51(t_col_51),
	.col_52(t_col_52),
	.col_53(t_col_53),
	.col_54(t_col_54),
	.col_55(t_col_55),
	.col_56(t_col_56),
	.col_57(t_col_57),
	.col_58(t_col_58),
	.col_59(t_col_59),
	.col_60(t_col_60),
	.col_61(t_col_61),
	.col_62(t_col_62),
	.col_63(t_col_63),
	.col_64(t_col_64),
	.col_65(t_col_65),
	.col_66(t_col_66),
	.col_67(t_col_67),
	.col_68(t_col_68),
	.col_69(t_col_69),
	.col_70(t_col_70),
	.col_71(t_col_71),
	.col_72(t_col_72),
	.col_73(t_col_73),
	.col_74(t_col_74),
	.col_75(t_col_75),
	.col_76(t_col_76),
	.col_77(t_col_77),
	.col_78(t_col_78),
	.col_79(t_col_79),
	.col_80(t_col_80),
	.col_81(t_col_81),
	.col_82(t_col_82),
	.col_83(t_col_83),
	.col_84(t_col_84),
	.col_85(t_col_85),
	.col_86(t_col_86),
	.col_87(t_col_87),
	.col_88(t_col_88),
	.col_89(t_col_89),
	.col_90(t_col_90),
	.col_91(t_col_91),
	.col_92(t_col_92),
	.col_93(t_col_93),
	.col_94(t_col_94),
	.col_95(t_col_95),
	.col_96(t_col_96),
	.col_97(t_col_97),
	.col_98(t_col_98),
	.col_99(t_col_99),
	.col_100(t_col_100),
	.col_101(t_col_101),
	.col_102(t_col_102),
	.col_103(t_col_103),
	.col_104(t_col_104),
	.col_105(t_col_105),
	.col_106(t_col_106),
	.col_107(t_col_107),
	.col_108(t_col_108),
	.col_109(t_col_109),
	.col_110(t_col_110),
	.col_111(t_col_111),
	.col_112(t_col_112),
	.col_113(t_col_113),
	.col_114(t_col_114),
	.col_115(t_col_115),
	.col_116(t_col_116),
	.col_117(t_col_117),
	.col_118(t_col_118),
	.col_119(t_col_119),
	.col_120(t_col_120),
	.col_121(t_col_121),
	.col_122(t_col_122),
	.col_123(t_col_123),
	.col_124(t_col_124),
	.col_125(t_col_125),
	.col_126(t_col_126),
	.col_127(t_col_127),
	.col_128(t_col_128),
	.col_129(t_col_129),
	.col_130(t_col_130),
	.col_131(t_col_131),
	.col_132(t_col_132),
	.col_133(t_col_133),
	.col_134(t_col_134),
	.col_135(t_col_135),
	.col_136(t_col_136),
	.col_137(t_col_137),
	.col_138(t_col_138),
	.col_139(t_col_139),
	.col_140(t_col_140),
	.col_141(t_col_141),
	.col_142(t_col_142),
	.col_143(t_col_143),
	.col_144(t_col_144),
	.col_145(t_col_145),
	.col_146(t_col_146),
	.col_147(t_col_147),
	.col_148(t_col_148),
	.col_149(t_col_149),
	.col_150(t_col_150),
	.col_151(t_col_151),
	.col_152(t_col_152),
	.col_153(t_col_153),
	.col_154(t_col_154),
	.col_155(t_col_155),
	.col_156(t_col_156),
	.col_157(t_col_157),
	.col_158(t_col_158),
	.col_159(t_col_159),
	.col_160(t_col_160),
	.col_161(t_col_161),
	.col_162(t_col_162),
	.col_163(t_col_163),
	.col_164(t_col_164),
	.col_165(t_col_165),
	.col_166(t_col_166),
	.col_167(t_col_167),
	.col_168(t_col_168),
	.col_169(t_col_169),
	.col_170(t_col_170),
	.col_171(t_col_171),
	.col_172(t_col_172),
	.col_173(t_col_173),
	.col_174(t_col_174),
	.col_175(t_col_175),
	.col_176(t_col_176),
	.col_177(t_col_177),
	.col_178(t_col_178),
	.col_179(t_col_179),
	.col_180(t_col_180),
	.col_181(t_col_181),
	.col_182(t_col_182),
	.col_183(t_col_183),
	.col_184(t_col_184),
	.col_185(t_col_185),
	.col_186(t_col_186),
	.col_187(t_col_187),
	.col_188(t_col_188),
	.col_189(t_col_189),
	.col_190(t_col_190),
	.col_191(t_col_191),
	.col_192(t_col_192),
	.col_193(t_col_193),
	.col_194(t_col_194),
	.col_195(t_col_195),
	.col_196(t_col_196),
	.col_197(t_col_197),
	.col_198(t_col_198),
	.col_199(t_col_199),
	.col_200(t_col_200),
	.col_201(t_col_201),
	.col_202(t_col_202),
	.col_203(t_col_203),
	.col_204(t_col_204),
	.col_205(t_col_205),
	.col_206(t_col_206),
	.col_207(t_col_207),
	.col_208(t_col_208),
	.col_209(t_col_209),
	.col_210(t_col_210),
	.col_211(t_col_211),
	.col_212(t_col_212),
	.col_213(t_col_213),
	.col_214(t_col_214),
	.col_215(t_col_215),
	.col_216(t_col_216),
	.col_217(t_col_217),
	.col_218(t_col_218),
	.col_219(t_col_219),
	.col_220(t_col_220),
	.col_221(t_col_221),
	.col_222(t_col_222),
	.col_223(t_col_223),
	.col_224(t_col_224),
	.col_225(t_col_225),
	.col_226(t_col_226),
	.col_227(t_col_227),
	.col_228(t_col_228),
	.col_229(t_col_229),
	.col_230(t_col_230),
	.col_231(t_col_231),
	.col_232(t_col_232),
	.col_233(t_col_233),
	.col_234(t_col_234),
	.col_235(t_col_235),
	.col_236(t_col_236),
	.col_237(t_col_237),
	.col_238(t_col_238),
	.col_239(t_col_239),
	.col_240(t_col_240),
	.col_241(t_col_241),
	.col_242(t_col_242),
	.col_243(t_col_243),
	.col_244(t_col_244),
	.col_245(t_col_245),
	.col_246(t_col_246),
	.col_247(t_col_247),
	.col_248(t_col_248),
	.col_249(t_col_249),
	.col_250(t_col_250),
	.col_251(t_col_251),
	.col_252(t_col_252),
	.col_253(t_col_253),
	.col_254(t_col_254),
	.col_255(t_col_255),
	.col_256(t_col_256),
	.col_257(t_col_257),
	.col_258(t_col_258),
	.col_259(t_col_259),
	.col_260(t_col_260),
	.col_261(t_col_261),
	.col_262(t_col_262),
	.col_263(t_col_263),
	.col_264(t_col_264),
	.col_265(t_col_265),
	.col_266(t_col_266),
	.col_267(t_col_267),
	.col_268(t_col_268),
	.col_269(t_col_269),
	.col_270(t_col_270),
	.col_271(t_col_271),
	.col_272(t_col_272),
	.col_273(t_col_273),
	.col_274(t_col_274),
	.col_275(t_col_275),
	.col_276(t_col_276),
	.col_277(t_col_277),
	.col_278(t_col_278),
	.col_279(t_col_279),
	.col_280(t_col_280),
	.col_281(t_col_281),
	.col_282(t_col_282),
	.col_283(t_col_283),
	.col_284(t_col_284),
	.col_285(t_col_285),
	.col_286(t_col_286),
	.col_287(t_col_287),
	.col_288(t_col_288),
	.col_289(t_col_289),
	.col_290(t_col_290),
	.col_291(t_col_291),
	.col_292(t_col_292),
	.col_293(t_col_293),
	.col_294(t_col_294),
	.col_295(t_col_295),
	.col_296(t_col_296),
	.col_297(t_col_297),
	.col_298(t_col_298),
	.col_299(t_col_299),
	.col_300(t_col_300),
	.col_301(t_col_301),
	.col_302(t_col_302),
	.col_303(t_col_303),
	.col_304(t_col_304),
	.col_305(t_col_305),
	.col_306(t_col_306),
	.col_307(t_col_307),
	.col_308(t_col_308),
	.col_309(t_col_309),
	.col_310(t_col_310),
	.col_311(t_col_311),
	.col_312(t_col_312),
	.col_313(t_col_313),
	.col_314(t_col_314),
	.col_315(t_col_315),
	.col_316(t_col_316),
	.col_317(t_col_317),
	.col_318(t_col_318),
	.col_319(t_col_319),
	.col_320(t_col_320),
	.col_321(t_col_321),
	.col_322(t_col_322),
	.col_323(t_col_323),
	.col_324(t_col_324),
	.col_325(t_col_325),
	.col_326(t_col_326),
	.col_327(t_col_327),
	.col_328(t_col_328),
	.col_329(t_col_329),
	.col_330(t_col_330),
	.col_331(t_col_331),
	.col_332(t_col_332),
	.col_333(t_col_333),
	.col_334(t_col_334),
	.col_335(t_col_335),
	.col_336(t_col_336),
	.col_337(t_col_337),
	.col_338(t_col_338),
	.col_339(t_col_339),
	.col_340(t_col_340),
	.col_341(t_col_341),
	.col_342(t_col_342),
	.col_343(t_col_343),
	.col_344(t_col_344),
	.col_345(t_col_345),
	.col_346(t_col_346),
	.col_347(t_col_347),
	.col_348(t_col_348),
	.col_349(t_col_349),
	.col_350(t_col_350),
	.col_351(t_col_351),
	.col_352(t_col_352),
	.col_353(t_col_353),
	.col_354(t_col_354),
	.col_355(t_col_355),
	.col_356(t_col_356),
	.col_357(t_col_357),
	.col_358(t_col_358),
	.col_359(t_col_359),
	.col_360(t_col_360),
	.col_361(t_col_361),
	.col_362(t_col_362),
	.col_363(t_col_363),
	.col_364(t_col_364),
	.col_365(t_col_365),
	.col_366(t_col_366),
	.col_367(t_col_367),
	.col_368(t_col_368),
	.col_369(t_col_369),
	.col_370(t_col_370),
	.col_371(t_col_371),
	.col_372(t_col_372),
	.col_373(t_col_373),
	.col_374(t_col_374),
	.col_375(t_col_375),
	.col_376(t_col_376),
	.col_377(t_col_377),
	.col_378(t_col_378),
	.col_379(t_col_379),
	.col_380(t_col_380),
	.col_381(t_col_381),
	.col_382(t_col_382),
	.col_383(t_col_383),
	.col_384(t_col_384),
	.col_385(t_col_385),
	.col_386(t_col_386),
	.col_387(t_col_387),
	.col_388(t_col_388),
	.col_389(t_col_389),
	.col_390(t_col_390),
	.col_391(t_col_391),
	.col_392(t_col_392),
	.col_393(t_col_393),
	.col_394(t_col_394),
	.col_395(t_col_395),
	.col_396(t_col_396),
	.col_397(t_col_397),
	.col_398(t_col_398),
	.col_399(t_col_399),
	.col_400(t_col_400),
	.col_401(t_col_401),
	.col_402(t_col_402),
	.col_403(t_col_403),
	.col_404(t_col_404),
	.col_405(t_col_405),
	.col_406(t_col_406),
	.col_407(t_col_407),
	.col_408(t_col_408),
	.col_409(t_col_409),
	.col_410(t_col_410),
	.col_411(t_col_411),
	.col_412(t_col_412),
	.col_413(t_col_413),
	.col_414(t_col_414),
	.col_415(t_col_415),
	.col_416(t_col_416),
	.col_417(t_col_417),
	.col_418(t_col_418),
	.col_419(t_col_419),
	.col_420(t_col_420),
	.col_421(t_col_421),
	.col_422(t_col_422),
	.col_423(t_col_423),
	.col_424(t_col_424),
	.col_425(t_col_425),
	.col_426(t_col_426),
	.col_427(t_col_427),
	.col_428(t_col_428),
	.col_429(t_col_429),
	.col_430(t_col_430),
	.col_431(t_col_431),
	.col_432(t_col_432),
	.col_433(t_col_433),
	.col_434(t_col_434),
	.col_435(t_col_435),
	.col_436(t_col_436),
	.col_437(t_col_437),
	.col_438(t_col_438),
	.col_439(t_col_439),
	.col_440(t_col_440),
	.col_441(t_col_441),
	.col_442(t_col_442),
	.col_443(t_col_443),
	.col_444(t_col_444),
	.col_445(t_col_445),
	.col_446(t_col_446),
	.col_447(t_col_447),
	.col_448(t_col_448),
	.col_449(t_col_449),
	.col_450(t_col_450),
	.col_451(t_col_451),
	.col_452(t_col_452),
	.col_453(t_col_453),
	.col_454(t_col_454),
	.col_455(t_col_455),
	.col_456(t_col_456),
	.col_457(t_col_457),
	.col_458(t_col_458),
	.col_459(t_col_459),
	.col_460(t_col_460),
	.col_461(t_col_461),
	.col_462(t_col_462),
	.col_463(t_col_463),
	.col_464(t_col_464),
	.col_465(t_col_465),
	.col_466(t_col_466),
	.col_467(t_col_467),
	.col_468(t_col_468),
	.col_469(t_col_469),
	.col_470(t_col_470),
	.col_471(t_col_471),
	.col_472(t_col_472),
	.col_473(t_col_473),
	.col_474(t_col_474),
	.col_475(t_col_475),
	.col_476(t_col_476),
	.col_477(t_col_477),
	.col_478(t_col_478),
	.col_479(t_col_479),
	.col_480(t_col_480),
	.col_481(t_col_481),
	.col_482(t_col_482),
	.col_483(t_col_483),
	.col_484(t_col_484),
	.col_485(t_col_485),
	.col_486(t_col_486),
	.col_487(t_col_487),
	.col_488(t_col_488),
	.col_489(t_col_489),
	.col_490(t_col_490),
	.col_491(t_col_491),
	.col_492(t_col_492),
	.col_493(t_col_493),
	.col_494(t_col_494),
	.col_495(t_col_495),
	.col_496(t_col_496),
	.col_497(t_col_497),
	.col_498(t_col_498),
	.col_499(t_col_499),
	.col_500(t_col_500),
	.col_501(t_col_501),
	.col_502(t_col_502),
	.col_503(t_col_503),
	.col_504(t_col_504),
	.col_505(t_col_505),
	.col_506(t_col_506),
	.col_507(t_col_507),
	.col_508(t_col_508),
	.col_509(t_col_509),
	.col_510(t_col_510),
	.col_511(t_col_511),
	.col_512(t_col_512),
	.col_513(t_col_513),
	.col_514(t_col_514),
	.col_515(t_col_515),
	.col_516(t_col_516),
	.col_517(t_col_517),
	.col_518(t_col_518),
	.col_519(t_col_519),
	.col_520(t_col_520),
	.col_521(t_col_521),
	.col_522(t_col_522),
	.col_523(t_col_523),
	.col_524(t_col_524),
	.col_525(t_col_525),
	.col_526(t_col_526),
	.col_527(t_col_527),
	.col_528(t_col_528),
	.col_529(t_col_529),
	.col_530(t_col_530),
	.col_531(t_col_531),
	.col_532(t_col_532),
	.col_533(t_col_533),
	.col_534(t_col_534),
	.col_535(t_col_535),
	.col_536(t_col_536),
	.col_537(t_col_537),
	.col_538(t_col_538),
	.col_539(t_col_539),
	.col_540(t_col_540),
	.col_541(t_col_541),
	.col_542(t_col_542),
	.col_543(t_col_543),
	.col_544(t_col_544),
	.col_545(t_col_545),
	.col_546(t_col_546),
	.col_547(t_col_547),
	.col_548(t_col_548),
	.col_549(t_col_549),
	.col_550(t_col_550),
	.col_551(t_col_551),
	.col_552(t_col_552),
	.col_553(t_col_553),
	.col_554(t_col_554),
	.col_555(t_col_555),
	.col_556(t_col_556),
	.col_557(t_col_557),
	.col_558(t_col_558),
	.col_559(t_col_559),
	.col_560(t_col_560),
	.col_561(t_col_561),
	.col_562(t_col_562),
	.col_563(t_col_563),
	.col_564(t_col_564),
	.col_565(t_col_565),
	.col_566(t_col_566),
	.col_567(t_col_567),
	.col_568(t_col_568),
	.col_569(t_col_569),
	.col_570(t_col_570),
	.col_571(t_col_571),
	.col_572(t_col_572),
	.col_573(t_col_573),
	.col_574(t_col_574),
	.col_575(t_col_575),
	.col_576(t_col_576),
	.col_577(t_col_577),
	.col_578(t_col_578),
	.col_579(t_col_579),
	.col_580(t_col_580),
	.col_581(t_col_581),
	.col_582(t_col_582),
	.col_583(t_col_583),
	.col_584(t_col_584),
	.col_585(t_col_585),
	.col_586(t_col_586),
	.col_587(t_col_587),
	.col_588(t_col_588),
	.col_589(t_col_589),
	.col_590(t_col_590),
	.col_591(t_col_591),
	.col_592(t_col_592),
	.col_593(t_col_593),
	.col_594(t_col_594),
	.col_595(t_col_595),
	.col_596(t_col_596),
	.col_597(t_col_597),
	.col_598(t_col_598),
	.col_599(t_col_599),
	.col_600(t_col_600),
	.col_601(t_col_601),
	.col_602(t_col_602),
	.col_603(t_col_603),
	.col_604(t_col_604),
	.col_605(t_col_605),
	.col_606(t_col_606),
	.col_607(t_col_607),
	.col_608(t_col_608),
	.col_609(t_col_609),
	.col_610(t_col_610),
	.col_611(t_col_611),
	.col_612(t_col_612),
	.col_613(t_col_613),
	.col_614(t_col_614),
	.col_615(t_col_615),
	.col_616(t_col_616),
	.col_617(t_col_617),
	.col_618(t_col_618),
	.col_619(t_col_619),
	.col_620(t_col_620),
	.col_621(t_col_621),
	.col_622(t_col_622),
	.col_623(t_col_623),
	.col_624(t_col_624),
	.col_625(t_col_625),
	.col_626(t_col_626),
	.col_627(t_col_627),
	.col_628(t_col_628),
	.col_629(t_col_629),
	.col_630(t_col_630),
	.col_631(t_col_631),
	.col_632(t_col_632),
	.col_633(t_col_633),
	.col_634(t_col_634),
	.col_635(t_col_635),
	.col_636(t_col_636),
	.col_637(t_col_637),
	.col_638(t_col_638),
	.col_639(t_col_639),
	.col_640(t_col_640),
	.col_641(t_col_641),
	.col_642(t_col_642),
	.col_643(t_col_643),
	.col_644(t_col_644),
	.col_645(t_col_645),
	.col_646(t_col_646),
	.col_647(t_col_647),
	.col_648(t_col_648),
	.col_649(t_col_649),
	.col_650(t_col_650),
	.col_651(t_col_651),
	.col_652(t_col_652),
	.col_653(t_col_653),
	.col_654(t_col_654),
	.col_655(t_col_655),
	.col_656(t_col_656),
	.col_657(t_col_657),
	.col_658(t_col_658),
	.col_659(t_col_659),
	.col_660(t_col_660),
	.col_661(t_col_661),
	.col_662(t_col_662),
	.col_663(t_col_663),
	.col_664(t_col_664),
	.col_665(t_col_665),
	.col_666(t_col_666),
	.col_667(t_col_667),
	.col_668(t_col_668),
	.col_669(t_col_669),
	.col_670(t_col_670),
	.col_671(t_col_671),
	.col_672(t_col_672),
	.col_673(t_col_673),
	.col_674(t_col_674),
	.col_675(t_col_675),
	.col_676(t_col_676),
	.col_677(t_col_677),
	.col_678(t_col_678),
	.col_679(t_col_679),
	.col_680(t_col_680),
	.col_681(t_col_681),
	.col_682(t_col_682),
	.col_683(t_col_683),
	.col_684(t_col_684),
	.col_685(t_col_685),
	.col_686(t_col_686),
	.col_687(t_col_687),
	.col_688(t_col_688),
	.col_689(t_col_689),
	.col_690(t_col_690),
	.col_691(t_col_691),
	.col_692(t_col_692),
	.col_693(t_col_693),
	.col_694(t_col_694),
	.col_695(t_col_695),
	.col_696(t_col_696),
	.col_697(t_col_697),
	.col_698(t_col_698),
	.col_699(t_col_699),
	.col_700(t_col_700),
	.col_701(t_col_701),
	.col_702(t_col_702),
	.col_703(t_col_703),
	.col_704(t_col_704),
	.col_705(t_col_705),
	.col_706(t_col_706),
	.col_707(t_col_707),
	.col_708(t_col_708),
	.col_709(t_col_709),
	.col_710(t_col_710),
	.col_711(t_col_711),
	.col_712(t_col_712),
	.col_713(t_col_713),
	.col_714(t_col_714),
	.col_715(t_col_715),
	.col_716(t_col_716),
	.col_717(t_col_717),
	.col_718(t_col_718),
	.col_719(t_col_719),
	.col_720(t_col_720),
	.col_721(t_col_721),
	.col_722(t_col_722),
	.col_723(t_col_723),
	.col_724(t_col_724),
	.col_725(t_col_725),
	.col_726(t_col_726),
	.col_727(t_col_727),
	.col_728(t_col_728),
	.col_729(t_col_729),
	.col_730(t_col_730),
	.col_731(t_col_731),
	.col_732(t_col_732),
	.col_733(t_col_733),
	.col_734(t_col_734),
	.col_735(t_col_735),
	.col_736(t_col_736),
	.col_737(t_col_737),
	.col_738(t_col_738),
	.col_739(t_col_739),
	.col_740(t_col_740),
	.col_741(t_col_741),
	.col_742(t_col_742),
	.col_743(t_col_743),
	.col_744(t_col_744),
	.col_745(t_col_745),
	.col_746(t_col_746),
	.col_747(t_col_747),
	.col_748(t_col_748),
	.col_749(t_col_749),
	.col_750(t_col_750),
	.col_751(t_col_751),
	.col_752(t_col_752),
	.col_753(t_col_753),
	.col_754(t_col_754),
	.col_755(t_col_755),
	.col_756(t_col_756),
	.col_757(t_col_757),
	.col_758(t_col_758),
	.col_759(t_col_759),
	.col_760(t_col_760),
	.col_761(t_col_761),
	.col_762(t_col_762),
	.col_763(t_col_763),
	.col_764(t_col_764),
	.col_765(t_col_765),
	.col_766(t_col_766),
	.col_767(t_col_767),
	.col_768(t_col_768),
	.col_769(t_col_769),
	.col_770(t_col_770),
	.col_771(t_col_771),
	.col_772(t_col_772),
	.col_773(t_col_773),
	.col_774(t_col_774),
	.col_775(t_col_775),
	.col_776(t_col_776),
	.col_777(t_col_777),
	.col_778(t_col_778),
	.col_779(t_col_779),
	.col_780(t_col_780),
	.col_781(t_col_781),
	.col_782(t_col_782),
	.col_783(t_col_783),
	.col_784(t_col_784),
	.col_785(t_col_785),
	.col_786(t_col_786),
	.col_787(t_col_787),
	.col_788(t_col_788),
	.col_789(t_col_789),
	.col_790(t_col_790),
	.col_791(t_col_791),
	.col_792(t_col_792),
	.col_793(t_col_793),
	.col_794(t_col_794),
	.col_795(t_col_795),
	.col_796(t_col_796),
	.col_797(t_col_797),
	.col_798(t_col_798),
	.col_799(t_col_799),
	.col_800(t_col_800),
	.col_801(t_col_801),
	.col_802(t_col_802),
	.col_803(t_col_803),
	.col_804(t_col_804),
	.col_805(t_col_805),
	.col_806(t_col_806),
	.col_807(t_col_807),
	.col_808(t_col_808),
	.col_809(t_col_809),
	.col_810(t_col_810),
	.col_811(t_col_811),
	.col_812(t_col_812),
	.col_813(t_col_813),
	.col_814(t_col_814),
	.col_815(t_col_815),
	.col_816(t_col_816),
	.col_817(t_col_817),
	.col_818(t_col_818),
	.col_819(t_col_819),
	.col_820(t_col_820),
	.col_821(t_col_821),
	.col_822(t_col_822),
	.col_823(t_col_823),
	.col_824(t_col_824),
	.col_825(t_col_825),
	.col_826(t_col_826),
	.col_827(t_col_827),
	.col_828(t_col_828),
	.col_829(t_col_829),
	.col_830(t_col_830),
	.col_831(t_col_831),
	.col_832(t_col_832),
	.col_833(t_col_833),
	.col_834(t_col_834),
	.col_835(t_col_835),
	.col_836(t_col_836),
	.col_837(t_col_837),
	.col_838(t_col_838),
	.col_839(t_col_839),
	.col_840(t_col_840),
	.col_841(t_col_841),
	.col_842(t_col_842),
	.col_843(t_col_843),
	.col_844(t_col_844),
	.col_845(t_col_845),
	.col_846(t_col_846),
	.col_847(t_col_847),
	.col_848(t_col_848),
	.col_849(t_col_849),
	.col_850(t_col_850),
	.col_851(t_col_851),
	.col_852(t_col_852),
	.col_853(t_col_853),
	.col_854(t_col_854),
	.col_855(t_col_855),
	.col_856(t_col_856),
	.col_857(t_col_857),
	.col_858(t_col_858),
	.col_859(t_col_859),
	.col_860(t_col_860),
	.col_861(t_col_861),
	.col_862(t_col_862),
	.col_863(t_col_863),
	.col_864(t_col_864),
	.col_865(t_col_865),
	.col_866(t_col_866),
	.col_867(t_col_867),
	.col_868(t_col_868),
	.col_869(t_col_869),
	.col_870(t_col_870),
	.col_871(t_col_871),
	.col_872(t_col_872),
	.col_873(t_col_873),
	.col_874(t_col_874),
	.col_875(t_col_875),
	.col_876(t_col_876),
	.col_877(t_col_877),
	.col_878(t_col_878),
	.col_879(t_col_879),
	.col_880(t_col_880),
	.col_881(t_col_881),
	.col_882(t_col_882),
	.col_883(t_col_883),
	.col_884(t_col_884),
	.col_885(t_col_885),
	.col_886(t_col_886),
	.col_887(t_col_887),
	.col_888(t_col_888),
	.col_889(t_col_889),
	.col_890(t_col_890),
	.col_891(t_col_891),
	.col_892(t_col_892),
	.col_893(t_col_893),
	.col_894(t_col_894),
	.col_895(t_col_895),
	.col_896(t_col_896),
	.col_897(t_col_897),
	.col_898(t_col_898),
	.col_899(t_col_899),
	.col_900(t_col_900),
	.col_901(t_col_901),
	.col_902(t_col_902),
	.col_903(t_col_903),
	.col_904(t_col_904),
	.col_905(t_col_905),
	.col_906(t_col_906),
	.col_907(t_col_907),
	.col_908(t_col_908),
	.col_909(t_col_909),
	.col_910(t_col_910),
	.col_911(t_col_911),
	.col_912(t_col_912),
	.col_913(t_col_913),
	.col_914(t_col_914),
	.col_915(t_col_915),
	.col_916(t_col_916),
	.col_917(t_col_917),
	.col_918(t_col_918),
	.col_919(t_col_919),
	.col_920(t_col_920),
	.col_921(t_col_921),
	.col_922(t_col_922),
	.col_923(t_col_923),
	.col_924(t_col_924),
	.col_925(t_col_925),
	.col_926(t_col_926),
	.col_927(t_col_927),
	.col_928(t_col_928),
	.col_929(t_col_929),
	.col_930(t_col_930),
	.col_931(t_col_931),
	.col_932(t_col_932),
	.col_933(t_col_933),
	.col_934(t_col_934),
	.col_935(t_col_935),
	.col_936(t_col_936),
	.col_937(t_col_937),
	.col_938(t_col_938),
	.col_939(t_col_939),
	.col_940(t_col_940),
	.col_941(t_col_941),
	.col_942(t_col_942),
	.col_943(t_col_943),
	.col_944(t_col_944),
	.col_945(t_col_945),
	.col_946(t_col_946),
	.col_947(t_col_947),
	.col_948(t_col_948),
	.col_949(t_col_949),
	.col_950(t_col_950),
	.col_951(t_col_951),
	.col_952(t_col_952),
	.col_953(t_col_953),
	.col_954(t_col_954),
	.col_955(t_col_955),
	.col_956(t_col_956),
	.col_957(t_col_957),
	.col_958(t_col_958),
	.col_959(t_col_959),
	.col_960(t_col_960),
	.col_961(t_col_961),
	.col_962(t_col_962),
	.col_963(t_col_963),
	.col_964(t_col_964),
	.col_965(t_col_965),
	.col_966(t_col_966),
	.col_967(t_col_967),
	.col_968(t_col_968),
	.col_969(t_col_969),
	.col_970(t_col_970),
	.col_971(t_col_971),
	.col_972(t_col_972),
	.col_973(t_col_973),
	.col_974(t_col_974),
	.col_975(t_col_975),
	.col_976(t_col_976),
	.col_977(t_col_977),
	.col_978(t_col_978),
	.col_979(t_col_979),
	.col_980(t_col_980),
	.col_981(t_col_981),
	.col_982(t_col_982),
	.col_983(t_col_983),
	.col_984(t_col_984),
	.col_985(t_col_985),
	.col_986(t_col_986),
	.col_987(t_col_987),
	.col_988(t_col_988),
	.col_989(t_col_989),
	.col_990(t_col_990),
	.col_991(t_col_991),
	.col_992(t_col_992),
	.col_993(t_col_993),
	.col_994(t_col_994),
	.col_995(t_col_995),
	.col_996(t_col_996),
	.col_997(t_col_997),
	.col_998(t_col_998),
	.col_999(t_col_999),
	.col_1000(t_col_1000),
	.col_1001(t_col_1001),
	.col_1002(t_col_1002),
	.col_1003(t_col_1003),
	.col_1004(t_col_1004),
	.col_1005(t_col_1005),
	.col_1006(t_col_1006),
	.col_1007(t_col_1007),
	.col_1008(t_col_1008),
	.col_1009(t_col_1009),
	.col_1010(t_col_1010),
	.col_1011(t_col_1011),
	.col_1012(t_col_1012),
	.col_1013(t_col_1013),
	.col_1014(t_col_1014),
	.col_1015(t_col_1015),
	.col_1016(t_col_1016),
	.col_1017(t_col_1017),
	.col_1018(t_col_1018),
	.col_1019(t_col_1019),
	.col_1020(t_col_1020),
	.col_1021(t_col_1021),
	.col_1022(t_col_1022),
	.col_1023(t_col_1023)
);

assign ta = sel ? {a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37], a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47], a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57], a[58], a[59], a[60], a[61], a[62], a[63], a[64], a[65], a[66], a[67], a[68], a[69], a[70], a[71], a[72], a[73], a[74], a[75], a[76], a[77], a[78], a[79], a[80], a[81], a[82], a[83], a[84], a[85], a[86], a[87], a[88], a[89], a[90], a[91], a[92], a[93], a[94], a[95], a[96], a[97], a[98], a[99], a[100], a[101], a[102], a[103], a[104], a[105], a[106], a[107], a[108], a[109], a[110], a[111], a[112], a[113], a[114], a[115], a[116], a[117], a[118], a[119], a[120], a[121], a[122], a[123], a[124], a[125], a[126], a[127], a[128], a[129], a[130], a[131], a[132], a[133], a[134], a[135], a[136], a[137], a[138], a[139], a[140], a[141], a[142], a[143], a[144], a[145], a[146], a[147], a[148], a[149], a[150], a[151], a[152], a[153], a[154], a[155], a[156], a[157], a[158], a[159], a[160], a[161], a[162], a[163], a[164], a[165], a[166], a[167], a[168], a[169], a[170], a[171], a[172], a[173], a[174], a[175], a[176], a[177], a[178], a[179], a[180], a[181], a[182], a[183], a[184], a[185], a[186], a[187], a[188], a[189], a[190], a[191], a[192], a[193], a[194], a[195], a[196], a[197], a[198], a[199], a[200], a[201], a[202], a[203], a[204], a[205], a[206], a[207], a[208], a[209], a[210], a[211], a[212], a[213], a[214], a[215], a[216], a[217], a[218], a[219], a[220], a[221], a[222], a[223], a[224], a[225], a[226], a[227], a[228], a[229], a[230], a[231], a[232], a[233], a[234], a[235], a[236], a[237], a[238], a[239], a[240], a[241], a[242], a[243], a[244], a[245], a[246], a[247], a[248], a[249], a[250], a[251], a[252], a[253], a[254], a[255], a[256], a[257], a[258], a[259], a[260], a[261], a[262], a[263], a[264], a[265], a[266], a[267], a[268], a[269], a[270], a[271], a[272], a[273], a[274], a[275], a[276], a[277], a[278], a[279], a[280], a[281], a[282], a[283], a[284], a[285], a[286], a[287], a[288], a[289], a[290], a[291], a[292], a[293], a[294], a[295], a[296], a[297], a[298], a[299], a[300], a[301], a[302], a[303], a[304], a[305], a[306], a[307], a[308], a[309], a[310], a[311], a[312], a[313], a[314], a[315], a[316], a[317], a[318], a[319], a[320], a[321], a[322], a[323], a[324], a[325], a[326], a[327], a[328], a[329], a[330], a[331], a[332], a[333], a[334], a[335], a[336], a[337], a[338], a[339], a[340], a[341], a[342], a[343], a[344], a[345], a[346], a[347], a[348], a[349], a[350], a[351], a[352], a[353], a[354], a[355], a[356], a[357], a[358], a[359], a[360], a[361], a[362], a[363], a[364], a[365], a[366], a[367], a[368], a[369], a[370], a[371], a[372], a[373], a[374], a[375], a[376], a[377], a[378], a[379], a[380], a[381], a[382], a[383], a[384], a[385], a[386], a[387], a[388], a[389], a[390], a[391], a[392], a[393], a[394], a[395], a[396], a[397], a[398], a[399], a[400], a[401], a[402], a[403], a[404], a[405], a[406], a[407], a[408], a[409], a[410], a[411], a[412], a[413], a[414], a[415], a[416], a[417], a[418], a[419], a[420], a[421], a[422], a[423], a[424], a[425], a[426], a[427], a[428], a[429], a[430], a[431], a[432], a[433], a[434], a[435], a[436], a[437], a[438], a[439], a[440], a[441], a[442], a[443], a[444], a[445], a[446], a[447], a[448], a[449], a[450], a[451], a[452], a[453], a[454], a[455], a[456], a[457], a[458], a[459], a[460], a[461], a[462], a[463], a[464], a[465], a[466], a[467], a[468], a[469], a[470], a[471], a[472], a[473], a[474], a[475], a[476], a[477], a[478], a[479], a[480], a[481], a[482], a[483], a[484], a[485], a[486], a[487], a[488], a[489], a[490], a[491], a[492], a[493], a[494], a[495], a[496], a[497], a[498], a[499], a[500], a[501], a[502], a[503], a[504], a[505], a[506], a[507], a[508], a[509], a[510], a[511], a[512], a[513], a[514], a[515], a[516], a[517], a[518], a[519], a[520], a[521], a[522], a[523], a[524], a[525], a[526], a[527], a[528], a[529], a[530], a[531], a[532], a[533], a[534], a[535], a[536], a[537], a[538], a[539], a[540], a[541], a[542], a[543], a[544], a[545], a[546], a[547], a[548], a[549], a[550], a[551], a[552], a[553], a[554], a[555], a[556], a[557], a[558], a[559], a[560], a[561], a[562], a[563], a[564], a[565], a[566], a[567], a[568], a[569], a[570], a[571], a[572], a[573], a[574], a[575], a[576], a[577], a[578], a[579], a[580], a[581], a[582], a[583], a[584], a[585], a[586], a[587], a[588], a[589], a[590], a[591], a[592], a[593], a[594], a[595], a[596], a[597], a[598], a[599], a[600], a[601], a[602], a[603], a[604], a[605], a[606], a[607], a[608], a[609], a[610], a[611], a[612], a[613], a[614], a[615], a[616], a[617], a[618], a[619], a[620], a[621], a[622], a[623], a[624], a[625], a[626], a[627], a[628], a[629], a[630], a[631], a[632], a[633], a[634], a[635], a[636], a[637], a[638], a[639], a[640], a[641], a[642], a[643], a[644], a[645], a[646], a[647], a[648], a[649], a[650], a[651], a[652], a[653], a[654], a[655], a[656], a[657], a[658], a[659], a[660], a[661], a[662], a[663], a[664], a[665], a[666], a[667], a[668], a[669], a[670], a[671], a[672], a[673], a[674], a[675], a[676], a[677], a[678], a[679], a[680], a[681], a[682], a[683], a[684], a[685], a[686], a[687], a[688], a[689], a[690], a[691], a[692], a[693], a[694], a[695], a[696], a[697], a[698], a[699], a[700], a[701], a[702], a[703], a[704], a[705], a[706], a[707], a[708], a[709], a[710], a[711], a[712], a[713], a[714], a[715], a[716], a[717], a[718], a[719], a[720], a[721], a[722], a[723], a[724], a[725], a[726], a[727], a[728], a[729], a[730], a[731], a[732], a[733], a[734], a[735], a[736], a[737], a[738], a[739], a[740], a[741], a[742], a[743], a[744], a[745], a[746], a[747], a[748], a[749], a[750], a[751], a[752], a[753], a[754], a[755], a[756], a[757], a[758], a[759], a[760], a[761], a[762], a[763], a[764], a[765], a[766], a[767], a[768], a[769], a[770], a[771], a[772], a[773], a[774], a[775], a[776], a[777], a[778], a[779], a[780], a[781], a[782], a[783], a[784], a[785], a[786], a[787], a[788], a[789], a[790], a[791], a[792], a[793], a[794], a[795], a[796], a[797], a[798], a[799], a[800], a[801], a[802], a[803], a[804], a[805], a[806], a[807], a[808], a[809], a[810], a[811], a[812], a[813], a[814], a[815], a[816], a[817], a[818], a[819], a[820], a[821], a[822], a[823], a[824], a[825], a[826], a[827], a[828], a[829], a[830], a[831], a[832], a[833], a[834], a[835], a[836], a[837], a[838], a[839], a[840], a[841], a[842], a[843], a[844], a[845], a[846], a[847], a[848], a[849], a[850], a[851], a[852], a[853], a[854], a[855], a[856], a[857], a[858], a[859], a[860], a[861], a[862], a[863], a[864], a[865], a[866], a[867], a[868], a[869], a[870], a[871], a[872], a[873], a[874], a[875], a[876], a[877], a[878], a[879], a[880], a[881], a[882], a[883], a[884], a[885], a[886], a[887], a[888], a[889], a[890], a[891], a[892], a[893], a[894], a[895], a[896], a[897], a[898], a[899], a[900], a[901], a[902], a[903], a[904], a[905], a[906], a[907], a[908], a[909], a[910], a[911], a[912], a[913], a[914], a[915], a[916], a[917], a[918], a[919], a[920], a[921], a[922], a[923], a[924], a[925], a[926], a[927], a[928], a[929], a[930], a[931], a[932], a[933], a[934], a[935], a[936], a[937], a[938], a[939], a[940], a[941], a[942], a[943], a[944], a[945], a[946], a[947], a[948], a[949], a[950], a[951], a[952], a[953], a[954], a[955], a[956], a[957], a[958], a[959], a[960], a[961], a[962], a[963], a[964], a[965], a[966], a[967], a[968], a[969], a[970], a[971], a[972], a[973], a[974], a[975], a[976], a[977], a[978], a[979], a[980], a[981], a[982], a[983], a[984], a[985], a[986], a[987], a[988], a[989], a[990], a[991], a[992], a[993], a[994], a[995], a[996], a[997], a[998], a[999], a[1000], a[1001], a[1002], a[1003], a[1004], a[1005], a[1006], a[1007], a[1008], a[1009], a[1010], a[1011], a[1012], a[1013], a[1014], a[1015], a[1016], a[1017], a[1018], a[1019], a[1020], a[1021], a[1022], a[1023]} : a;
assign col_0 = sel ? {a[1023] & a[0], a[1022] & a[1], a[1021] & a[2], a[1020] & a[3], a[1019] & a[4], a[1018] & a[5], a[1017] & a[6], a[1016] & a[7], a[1015] & a[8], a[1014] & a[9], a[1013] & a[10], a[1012] & a[11], a[1011] & a[12], a[1010] & a[13], a[1009] & a[14], a[1008] & a[15], a[1007] & a[16], a[1006] & a[17], a[1005] & a[18], a[1004] & a[19], a[1003] & a[20], a[1002] & a[21], a[1001] & a[22], a[1000] & a[23], a[999] & a[24], a[998] & a[25], a[997] & a[26], a[996] & a[27], a[995] & a[28], a[994] & a[29], a[993] & a[30], a[992] & a[31], a[991] & a[32], a[990] & a[33], a[989] & a[34], a[988] & a[35], a[987] & a[36], a[986] & a[37], a[985] & a[38], a[984] & a[39], a[983] & a[40], a[982] & a[41], a[981] & a[42], a[980] & a[43], a[979] & a[44], a[978] & a[45], a[977] & a[46], a[976] & a[47], a[975] & a[48], a[974] & a[49], a[973] & a[50], a[972] & a[51], a[971] & a[52], a[970] & a[53], a[969] & a[54], a[968] & a[55], a[967] & a[56], a[966] & a[57], a[965] & a[58], a[964] & a[59], a[963] & a[60], a[962] & a[61], a[961] & a[62], a[960] & a[63], a[959] & a[64], a[958] & a[65], a[957] & a[66], a[956] & a[67], a[955] & a[68], a[954] & a[69], a[953] & a[70], a[952] & a[71], a[951] & a[72], a[950] & a[73], a[949] & a[74], a[948] & a[75], a[947] & a[76], a[946] & a[77], a[945] & a[78], a[944] & a[79], a[943] & a[80], a[942] & a[81], a[941] & a[82], a[940] & a[83], a[939] & a[84], a[938] & a[85], a[937] & a[86], a[936] & a[87], a[935] & a[88], a[934] & a[89], a[933] & a[90], a[932] & a[91], a[931] & a[92], a[930] & a[93], a[929] & a[94], a[928] & a[95], a[927] & a[96], a[926] & a[97], a[925] & a[98], a[924] & a[99], a[923] & a[100], a[922] & a[101], a[921] & a[102], a[920] & a[103], a[919] & a[104], a[918] & a[105], a[917] & a[106], a[916] & a[107], a[915] & a[108], a[914] & a[109], a[913] & a[110], a[912] & a[111], a[911] & a[112], a[910] & a[113], a[909] & a[114], a[908] & a[115], a[907] & a[116], a[906] & a[117], a[905] & a[118], a[904] & a[119], a[903] & a[120], a[902] & a[121], a[901] & a[122], a[900] & a[123], a[899] & a[124], a[898] & a[125], a[897] & a[126], a[896] & a[127], a[895] & a[128], a[894] & a[129], a[893] & a[130], a[892] & a[131], a[891] & a[132], a[890] & a[133], a[889] & a[134], a[888] & a[135], a[887] & a[136], a[886] & a[137], a[885] & a[138], a[884] & a[139], a[883] & a[140], a[882] & a[141], a[881] & a[142], a[880] & a[143], a[879] & a[144], a[878] & a[145], a[877] & a[146], a[876] & a[147], a[875] & a[148], a[874] & a[149], a[873] & a[150], a[872] & a[151], a[871] & a[152], a[870] & a[153], a[869] & a[154], a[868] & a[155], a[867] & a[156], a[866] & a[157], a[865] & a[158], a[864] & a[159], a[863] & a[160], a[862] & a[161], a[861] & a[162], a[860] & a[163], a[859] & a[164], a[858] & a[165], a[857] & a[166], a[856] & a[167], a[855] & a[168], a[854] & a[169], a[853] & a[170], a[852] & a[171], a[851] & a[172], a[850] & a[173], a[849] & a[174], a[848] & a[175], a[847] & a[176], a[846] & a[177], a[845] & a[178], a[844] & a[179], a[843] & a[180], a[842] & a[181], a[841] & a[182], a[840] & a[183], a[839] & a[184], a[838] & a[185], a[837] & a[186], a[836] & a[187], a[835] & a[188], a[834] & a[189], a[833] & a[190], a[832] & a[191], a[831] & a[192], a[830] & a[193], a[829] & a[194], a[828] & a[195], a[827] & a[196], a[826] & a[197], a[825] & a[198], a[824] & a[199], a[823] & a[200], a[822] & a[201], a[821] & a[202], a[820] & a[203], a[819] & a[204], a[818] & a[205], a[817] & a[206], a[816] & a[207], a[815] & a[208], a[814] & a[209], a[813] & a[210], a[812] & a[211], a[811] & a[212], a[810] & a[213], a[809] & a[214], a[808] & a[215], a[807] & a[216], a[806] & a[217], a[805] & a[218], a[804] & a[219], a[803] & a[220], a[802] & a[221], a[801] & a[222], a[800] & a[223], a[799] & a[224], a[798] & a[225], a[797] & a[226], a[796] & a[227], a[795] & a[228], a[794] & a[229], a[793] & a[230], a[792] & a[231], a[791] & a[232], a[790] & a[233], a[789] & a[234], a[788] & a[235], a[787] & a[236], a[786] & a[237], a[785] & a[238], a[784] & a[239], a[783] & a[240], a[782] & a[241], a[781] & a[242], a[780] & a[243], a[779] & a[244], a[778] & a[245], a[777] & a[246], a[776] & a[247], a[775] & a[248], a[774] & a[249], a[773] & a[250], a[772] & a[251], a[771] & a[252], a[770] & a[253], a[769] & a[254], a[768] & a[255], a[767] & a[256], a[766] & a[257], a[765] & a[258], a[764] & a[259], a[763] & a[260], a[762] & a[261], a[761] & a[262], a[760] & a[263], a[759] & a[264], a[758] & a[265], a[757] & a[266], a[756] & a[267], a[755] & a[268], a[754] & a[269], a[753] & a[270], a[752] & a[271], a[751] & a[272], a[750] & a[273], a[749] & a[274], a[748] & a[275], a[747] & a[276], a[746] & a[277], a[745] & a[278], a[744] & a[279], a[743] & a[280], a[742] & a[281], a[741] & a[282], a[740] & a[283], a[739] & a[284], a[738] & a[285], a[737] & a[286], a[736] & a[287], a[735] & a[288], a[734] & a[289], a[733] & a[290], a[732] & a[291], a[731] & a[292], a[730] & a[293], a[729] & a[294], a[728] & a[295], a[727] & a[296], a[726] & a[297], a[725] & a[298], a[724] & a[299], a[723] & a[300], a[722] & a[301], a[721] & a[302], a[720] & a[303], a[719] & a[304], a[718] & a[305], a[717] & a[306], a[716] & a[307], a[715] & a[308], a[714] & a[309], a[713] & a[310], a[712] & a[311], a[711] & a[312], a[710] & a[313], a[709] & a[314], a[708] & a[315], a[707] & a[316], a[706] & a[317], a[705] & a[318], a[704] & a[319], a[703] & a[320], a[702] & a[321], a[701] & a[322], a[700] & a[323], a[699] & a[324], a[698] & a[325], a[697] & a[326], a[696] & a[327], a[695] & a[328], a[694] & a[329], a[693] & a[330], a[692] & a[331], a[691] & a[332], a[690] & a[333], a[689] & a[334], a[688] & a[335], a[687] & a[336], a[686] & a[337], a[685] & a[338], a[684] & a[339], a[683] & a[340], a[682] & a[341], a[681] & a[342], a[680] & a[343], a[679] & a[344], a[678] & a[345], a[677] & a[346], a[676] & a[347], a[675] & a[348], a[674] & a[349], a[673] & a[350], a[672] & a[351], a[671] & a[352], a[670] & a[353], a[669] & a[354], a[668] & a[355], a[667] & a[356], a[666] & a[357], a[665] & a[358], a[664] & a[359], a[663] & a[360], a[662] & a[361], a[661] & a[362], a[660] & a[363], a[659] & a[364], a[658] & a[365], a[657] & a[366], a[656] & a[367], a[655] & a[368], a[654] & a[369], a[653] & a[370], a[652] & a[371], a[651] & a[372], a[650] & a[373], a[649] & a[374], a[648] & a[375], a[647] & a[376], a[646] & a[377], a[645] & a[378], a[644] & a[379], a[643] & a[380], a[642] & a[381], a[641] & a[382], a[640] & a[383], a[639] & a[384], a[638] & a[385], a[637] & a[386], a[636] & a[387], a[635] & a[388], a[634] & a[389], a[633] & a[390], a[632] & a[391], a[631] & a[392], a[630] & a[393], a[629] & a[394], a[628] & a[395], a[627] & a[396], a[626] & a[397], a[625] & a[398], a[624] & a[399], a[623] & a[400], a[622] & a[401], a[621] & a[402], a[620] & a[403], a[619] & a[404], a[618] & a[405], a[617] & a[406], a[616] & a[407], a[615] & a[408], a[614] & a[409], a[613] & a[410], a[612] & a[411], a[611] & a[412], a[610] & a[413], a[609] & a[414], a[608] & a[415], a[607] & a[416], a[606] & a[417], a[605] & a[418], a[604] & a[419], a[603] & a[420], a[602] & a[421], a[601] & a[422], a[600] & a[423], a[599] & a[424], a[598] & a[425], a[597] & a[426], a[596] & a[427], a[595] & a[428], a[594] & a[429], a[593] & a[430], a[592] & a[431], a[591] & a[432], a[590] & a[433], a[589] & a[434], a[588] & a[435], a[587] & a[436], a[586] & a[437], a[585] & a[438], a[584] & a[439], a[583] & a[440], a[582] & a[441], a[581] & a[442], a[580] & a[443], a[579] & a[444], a[578] & a[445], a[577] & a[446], a[576] & a[447], a[575] & a[448], a[574] & a[449], a[573] & a[450], a[572] & a[451], a[571] & a[452], a[570] & a[453], a[569] & a[454], a[568] & a[455], a[567] & a[456], a[566] & a[457], a[565] & a[458], a[564] & a[459], a[563] & a[460], a[562] & a[461], a[561] & a[462], a[560] & a[463], a[559] & a[464], a[558] & a[465], a[557] & a[466], a[556] & a[467], a[555] & a[468], a[554] & a[469], a[553] & a[470], a[552] & a[471], a[551] & a[472], a[550] & a[473], a[549] & a[474], a[548] & a[475], a[547] & a[476], a[546] & a[477], a[545] & a[478], a[544] & a[479], a[543] & a[480], a[542] & a[481], a[541] & a[482], a[540] & a[483], a[539] & a[484], a[538] & a[485], a[537] & a[486], a[536] & a[487], a[535] & a[488], a[534] & a[489], a[533] & a[490], a[532] & a[491], a[531] & a[492], a[530] & a[493], a[529] & a[494], a[528] & a[495], a[527] & a[496], a[526] & a[497], a[525] & a[498], a[524] & a[499], a[523] & a[500], a[522] & a[501], a[521] & a[502], a[520] & a[503], a[519] & a[504], a[518] & a[505], a[517] & a[506], a[516] & a[507], a[515] & a[508], a[514] & a[509], a[513] & a[510], a[512] & ~a[511]} : {a[0], 511'b0};
assign col_1 = sel ? {t_col_1023, a[512] & a[511]} : 512'b0;
assign col_2 = sel ? {t_col_1022, ~a[512] & a[513]} : {t_col_2, ~a[0] & a[1]};
assign col_3 = sel ? {t_col_1021, a[513] & a[512]} : {t_col_3, a[0] & a[1]};
assign col_4 = sel ? {t_col_1020, ~a[513] & a[514]} : {t_col_4, ~a[1] & a[2]};
assign col_5 = sel ? {t_col_1019, a[514] & a[513]} : {t_col_5, a[1] & a[2]};
assign col_6 = sel ? {t_col_1018, ~a[514] & a[515]} : {t_col_6, ~a[2] & a[3]};
assign col_7 = sel ? {t_col_1017, a[515] & a[514]} : {t_col_7, a[2] & a[3]};
assign col_8 = sel ? {t_col_1016, ~a[515] & a[516]} : {t_col_8, ~a[3] & a[4]};
assign col_9 = sel ? {t_col_1015, a[516] & a[515]} : {t_col_9, a[3] & a[4]};
assign col_10 = sel ? {t_col_1014, ~a[516] & a[517]} : {t_col_10, ~a[4] & a[5]};
assign col_11 = sel ? {t_col_1013, a[517] & a[516]} : {t_col_11, a[4] & a[5]};
assign col_12 = sel ? {t_col_1012, ~a[517] & a[518]} : {t_col_12, ~a[5] & a[6]};
assign col_13 = sel ? {t_col_1011, a[518] & a[517]} : {t_col_13, a[5] & a[6]};
assign col_14 = sel ? {t_col_1010, ~a[518] & a[519]} : {t_col_14, ~a[6] & a[7]};
assign col_15 = sel ? {t_col_1009, a[519] & a[518]} : {t_col_15, a[6] & a[7]};
assign col_16 = sel ? {t_col_1008, ~a[519] & a[520]} : {t_col_16, ~a[7] & a[8]};
assign col_17 = sel ? {t_col_1007, a[520] & a[519]} : {t_col_17, a[7] & a[8]};
assign col_18 = sel ? {t_col_1006, ~a[520] & a[521]} : {t_col_18, ~a[8] & a[9]};
assign col_19 = sel ? {t_col_1005, a[521] & a[520]} : {t_col_19, a[8] & a[9]};
assign col_20 = sel ? {t_col_1004, ~a[521] & a[522]} : {t_col_20, ~a[9] & a[10]};
assign col_21 = sel ? {t_col_1003, a[522] & a[521]} : {t_col_21, a[9] & a[10]};
assign col_22 = sel ? {t_col_1002, ~a[522] & a[523]} : {t_col_22, ~a[10] & a[11]};
assign col_23 = sel ? {t_col_1001, a[523] & a[522]} : {t_col_23, a[10] & a[11]};
assign col_24 = sel ? {t_col_1000, ~a[523] & a[524]} : {t_col_24, ~a[11] & a[12]};
assign col_25 = sel ? {t_col_999, a[524] & a[523]} : {t_col_25, a[11] & a[12]};
assign col_26 = sel ? {t_col_998, ~a[524] & a[525]} : {t_col_26, ~a[12] & a[13]};
assign col_27 = sel ? {t_col_997, a[525] & a[524]} : {t_col_27, a[12] & a[13]};
assign col_28 = sel ? {t_col_996, ~a[525] & a[526]} : {t_col_28, ~a[13] & a[14]};
assign col_29 = sel ? {t_col_995, a[526] & a[525]} : {t_col_29, a[13] & a[14]};
assign col_30 = sel ? {t_col_994, ~a[526] & a[527]} : {t_col_30, ~a[14] & a[15]};
assign col_31 = sel ? {t_col_993, a[527] & a[526]} : {t_col_31, a[14] & a[15]};
assign col_32 = sel ? {t_col_992, ~a[527] & a[528]} : {t_col_32, ~a[15] & a[16]};
assign col_33 = sel ? {t_col_991, a[528] & a[527]} : {t_col_33, a[15] & a[16]};
assign col_34 = sel ? {t_col_990, ~a[528] & a[529]} : {t_col_34, ~a[16] & a[17]};
assign col_35 = sel ? {t_col_989, a[529] & a[528]} : {t_col_35, a[16] & a[17]};
assign col_36 = sel ? {t_col_988, ~a[529] & a[530]} : {t_col_36, ~a[17] & a[18]};
assign col_37 = sel ? {t_col_987, a[530] & a[529]} : {t_col_37, a[17] & a[18]};
assign col_38 = sel ? {t_col_986, ~a[530] & a[531]} : {t_col_38, ~a[18] & a[19]};
assign col_39 = sel ? {t_col_985, a[531] & a[530]} : {t_col_39, a[18] & a[19]};
assign col_40 = sel ? {t_col_984, ~a[531] & a[532]} : {t_col_40, ~a[19] & a[20]};
assign col_41 = sel ? {t_col_983, a[532] & a[531]} : {t_col_41, a[19] & a[20]};
assign col_42 = sel ? {t_col_982, ~a[532] & a[533]} : {t_col_42, ~a[20] & a[21]};
assign col_43 = sel ? {t_col_981, a[533] & a[532]} : {t_col_43, a[20] & a[21]};
assign col_44 = sel ? {t_col_980, ~a[533] & a[534]} : {t_col_44, ~a[21] & a[22]};
assign col_45 = sel ? {t_col_979, a[534] & a[533]} : {t_col_45, a[21] & a[22]};
assign col_46 = sel ? {t_col_978, ~a[534] & a[535]} : {t_col_46, ~a[22] & a[23]};
assign col_47 = sel ? {t_col_977, a[535] & a[534]} : {t_col_47, a[22] & a[23]};
assign col_48 = sel ? {t_col_976, ~a[535] & a[536]} : {t_col_48, ~a[23] & a[24]};
assign col_49 = sel ? {t_col_975, a[536] & a[535]} : {t_col_49, a[23] & a[24]};
assign col_50 = sel ? {t_col_974, ~a[536] & a[537]} : {t_col_50, ~a[24] & a[25]};
assign col_51 = sel ? {t_col_973, a[537] & a[536]} : {t_col_51, a[24] & a[25]};
assign col_52 = sel ? {t_col_972, ~a[537] & a[538]} : {t_col_52, ~a[25] & a[26]};
assign col_53 = sel ? {t_col_971, a[538] & a[537]} : {t_col_53, a[25] & a[26]};
assign col_54 = sel ? {t_col_970, ~a[538] & a[539]} : {t_col_54, ~a[26] & a[27]};
assign col_55 = sel ? {t_col_969, a[539] & a[538]} : {t_col_55, a[26] & a[27]};
assign col_56 = sel ? {t_col_968, ~a[539] & a[540]} : {t_col_56, ~a[27] & a[28]};
assign col_57 = sel ? {t_col_967, a[540] & a[539]} : {t_col_57, a[27] & a[28]};
assign col_58 = sel ? {t_col_966, ~a[540] & a[541]} : {t_col_58, ~a[28] & a[29]};
assign col_59 = sel ? {t_col_965, a[541] & a[540]} : {t_col_59, a[28] & a[29]};
assign col_60 = sel ? {t_col_964, ~a[541] & a[542]} : {t_col_60, ~a[29] & a[30]};
assign col_61 = sel ? {t_col_963, a[542] & a[541]} : {t_col_61, a[29] & a[30]};
assign col_62 = sel ? {t_col_962, ~a[542] & a[543]} : {t_col_62, ~a[30] & a[31]};
assign col_63 = sel ? {t_col_961, a[543] & a[542]} : {t_col_63, a[30] & a[31]};
assign col_64 = sel ? {t_col_960, ~a[543] & a[544]} : {t_col_64, ~a[31] & a[32]};
assign col_65 = sel ? {t_col_959, a[544] & a[543]} : {t_col_65, a[31] & a[32]};
assign col_66 = sel ? {t_col_958, ~a[544] & a[545]} : {t_col_66, ~a[32] & a[33]};
assign col_67 = sel ? {t_col_957, a[545] & a[544]} : {t_col_67, a[32] & a[33]};
assign col_68 = sel ? {t_col_956, ~a[545] & a[546]} : {t_col_68, ~a[33] & a[34]};
assign col_69 = sel ? {t_col_955, a[546] & a[545]} : {t_col_69, a[33] & a[34]};
assign col_70 = sel ? {t_col_954, ~a[546] & a[547]} : {t_col_70, ~a[34] & a[35]};
assign col_71 = sel ? {t_col_953, a[547] & a[546]} : {t_col_71, a[34] & a[35]};
assign col_72 = sel ? {t_col_952, ~a[547] & a[548]} : {t_col_72, ~a[35] & a[36]};
assign col_73 = sel ? {t_col_951, a[548] & a[547]} : {t_col_73, a[35] & a[36]};
assign col_74 = sel ? {t_col_950, ~a[548] & a[549]} : {t_col_74, ~a[36] & a[37]};
assign col_75 = sel ? {t_col_949, a[549] & a[548]} : {t_col_75, a[36] & a[37]};
assign col_76 = sel ? {t_col_948, ~a[549] & a[550]} : {t_col_76, ~a[37] & a[38]};
assign col_77 = sel ? {t_col_947, a[550] & a[549]} : {t_col_77, a[37] & a[38]};
assign col_78 = sel ? {t_col_946, ~a[550] & a[551]} : {t_col_78, ~a[38] & a[39]};
assign col_79 = sel ? {t_col_945, a[551] & a[550]} : {t_col_79, a[38] & a[39]};
assign col_80 = sel ? {t_col_944, ~a[551] & a[552]} : {t_col_80, ~a[39] & a[40]};
assign col_81 = sel ? {t_col_943, a[552] & a[551]} : {t_col_81, a[39] & a[40]};
assign col_82 = sel ? {t_col_942, ~a[552] & a[553]} : {t_col_82, ~a[40] & a[41]};
assign col_83 = sel ? {t_col_941, a[553] & a[552]} : {t_col_83, a[40] & a[41]};
assign col_84 = sel ? {t_col_940, ~a[553] & a[554]} : {t_col_84, ~a[41] & a[42]};
assign col_85 = sel ? {t_col_939, a[554] & a[553]} : {t_col_85, a[41] & a[42]};
assign col_86 = sel ? {t_col_938, ~a[554] & a[555]} : {t_col_86, ~a[42] & a[43]};
assign col_87 = sel ? {t_col_937, a[555] & a[554]} : {t_col_87, a[42] & a[43]};
assign col_88 = sel ? {t_col_936, ~a[555] & a[556]} : {t_col_88, ~a[43] & a[44]};
assign col_89 = sel ? {t_col_935, a[556] & a[555]} : {t_col_89, a[43] & a[44]};
assign col_90 = sel ? {t_col_934, ~a[556] & a[557]} : {t_col_90, ~a[44] & a[45]};
assign col_91 = sel ? {t_col_933, a[557] & a[556]} : {t_col_91, a[44] & a[45]};
assign col_92 = sel ? {t_col_932, ~a[557] & a[558]} : {t_col_92, ~a[45] & a[46]};
assign col_93 = sel ? {t_col_931, a[558] & a[557]} : {t_col_93, a[45] & a[46]};
assign col_94 = sel ? {t_col_930, ~a[558] & a[559]} : {t_col_94, ~a[46] & a[47]};
assign col_95 = sel ? {t_col_929, a[559] & a[558]} : {t_col_95, a[46] & a[47]};
assign col_96 = sel ? {t_col_928, ~a[559] & a[560]} : {t_col_96, ~a[47] & a[48]};
assign col_97 = sel ? {t_col_927, a[560] & a[559]} : {t_col_97, a[47] & a[48]};
assign col_98 = sel ? {t_col_926, ~a[560] & a[561]} : {t_col_98, ~a[48] & a[49]};
assign col_99 = sel ? {t_col_925, a[561] & a[560]} : {t_col_99, a[48] & a[49]};
assign col_100 = sel ? {t_col_924, ~a[561] & a[562]} : {t_col_100, ~a[49] & a[50]};
assign col_101 = sel ? {t_col_923, a[562] & a[561]} : {t_col_101, a[49] & a[50]};
assign col_102 = sel ? {t_col_922, ~a[562] & a[563]} : {t_col_102, ~a[50] & a[51]};
assign col_103 = sel ? {t_col_921, a[563] & a[562]} : {t_col_103, a[50] & a[51]};
assign col_104 = sel ? {t_col_920, ~a[563] & a[564]} : {t_col_104, ~a[51] & a[52]};
assign col_105 = sel ? {t_col_919, a[564] & a[563]} : {t_col_105, a[51] & a[52]};
assign col_106 = sel ? {t_col_918, ~a[564] & a[565]} : {t_col_106, ~a[52] & a[53]};
assign col_107 = sel ? {t_col_917, a[565] & a[564]} : {t_col_107, a[52] & a[53]};
assign col_108 = sel ? {t_col_916, ~a[565] & a[566]} : {t_col_108, ~a[53] & a[54]};
assign col_109 = sel ? {t_col_915, a[566] & a[565]} : {t_col_109, a[53] & a[54]};
assign col_110 = sel ? {t_col_914, ~a[566] & a[567]} : {t_col_110, ~a[54] & a[55]};
assign col_111 = sel ? {t_col_913, a[567] & a[566]} : {t_col_111, a[54] & a[55]};
assign col_112 = sel ? {t_col_912, ~a[567] & a[568]} : {t_col_112, ~a[55] & a[56]};
assign col_113 = sel ? {t_col_911, a[568] & a[567]} : {t_col_113, a[55] & a[56]};
assign col_114 = sel ? {t_col_910, ~a[568] & a[569]} : {t_col_114, ~a[56] & a[57]};
assign col_115 = sel ? {t_col_909, a[569] & a[568]} : {t_col_115, a[56] & a[57]};
assign col_116 = sel ? {t_col_908, ~a[569] & a[570]} : {t_col_116, ~a[57] & a[58]};
assign col_117 = sel ? {t_col_907, a[570] & a[569]} : {t_col_117, a[57] & a[58]};
assign col_118 = sel ? {t_col_906, ~a[570] & a[571]} : {t_col_118, ~a[58] & a[59]};
assign col_119 = sel ? {t_col_905, a[571] & a[570]} : {t_col_119, a[58] & a[59]};
assign col_120 = sel ? {t_col_904, ~a[571] & a[572]} : {t_col_120, ~a[59] & a[60]};
assign col_121 = sel ? {t_col_903, a[572] & a[571]} : {t_col_121, a[59] & a[60]};
assign col_122 = sel ? {t_col_902, ~a[572] & a[573]} : {t_col_122, ~a[60] & a[61]};
assign col_123 = sel ? {t_col_901, a[573] & a[572]} : {t_col_123, a[60] & a[61]};
assign col_124 = sel ? {t_col_900, ~a[573] & a[574]} : {t_col_124, ~a[61] & a[62]};
assign col_125 = sel ? {t_col_899, a[574] & a[573]} : {t_col_125, a[61] & a[62]};
assign col_126 = sel ? {t_col_898, ~a[574] & a[575]} : {t_col_126, ~a[62] & a[63]};
assign col_127 = sel ? {t_col_897, a[575] & a[574]} : {t_col_127, a[62] & a[63]};
assign col_128 = sel ? {t_col_896, ~a[575] & a[576]} : {t_col_128, ~a[63] & a[64]};
assign col_129 = sel ? {t_col_895, a[576] & a[575]} : {t_col_129, a[63] & a[64]};
assign col_130 = sel ? {t_col_894, ~a[576] & a[577]} : {t_col_130, ~a[64] & a[65]};
assign col_131 = sel ? {t_col_893, a[577] & a[576]} : {t_col_131, a[64] & a[65]};
assign col_132 = sel ? {t_col_892, ~a[577] & a[578]} : {t_col_132, ~a[65] & a[66]};
assign col_133 = sel ? {t_col_891, a[578] & a[577]} : {t_col_133, a[65] & a[66]};
assign col_134 = sel ? {t_col_890, ~a[578] & a[579]} : {t_col_134, ~a[66] & a[67]};
assign col_135 = sel ? {t_col_889, a[579] & a[578]} : {t_col_135, a[66] & a[67]};
assign col_136 = sel ? {t_col_888, ~a[579] & a[580]} : {t_col_136, ~a[67] & a[68]};
assign col_137 = sel ? {t_col_887, a[580] & a[579]} : {t_col_137, a[67] & a[68]};
assign col_138 = sel ? {t_col_886, ~a[580] & a[581]} : {t_col_138, ~a[68] & a[69]};
assign col_139 = sel ? {t_col_885, a[581] & a[580]} : {t_col_139, a[68] & a[69]};
assign col_140 = sel ? {t_col_884, ~a[581] & a[582]} : {t_col_140, ~a[69] & a[70]};
assign col_141 = sel ? {t_col_883, a[582] & a[581]} : {t_col_141, a[69] & a[70]};
assign col_142 = sel ? {t_col_882, ~a[582] & a[583]} : {t_col_142, ~a[70] & a[71]};
assign col_143 = sel ? {t_col_881, a[583] & a[582]} : {t_col_143, a[70] & a[71]};
assign col_144 = sel ? {t_col_880, ~a[583] & a[584]} : {t_col_144, ~a[71] & a[72]};
assign col_145 = sel ? {t_col_879, a[584] & a[583]} : {t_col_145, a[71] & a[72]};
assign col_146 = sel ? {t_col_878, ~a[584] & a[585]} : {t_col_146, ~a[72] & a[73]};
assign col_147 = sel ? {t_col_877, a[585] & a[584]} : {t_col_147, a[72] & a[73]};
assign col_148 = sel ? {t_col_876, ~a[585] & a[586]} : {t_col_148, ~a[73] & a[74]};
assign col_149 = sel ? {t_col_875, a[586] & a[585]} : {t_col_149, a[73] & a[74]};
assign col_150 = sel ? {t_col_874, ~a[586] & a[587]} : {t_col_150, ~a[74] & a[75]};
assign col_151 = sel ? {t_col_873, a[587] & a[586]} : {t_col_151, a[74] & a[75]};
assign col_152 = sel ? {t_col_872, ~a[587] & a[588]} : {t_col_152, ~a[75] & a[76]};
assign col_153 = sel ? {t_col_871, a[588] & a[587]} : {t_col_153, a[75] & a[76]};
assign col_154 = sel ? {t_col_870, ~a[588] & a[589]} : {t_col_154, ~a[76] & a[77]};
assign col_155 = sel ? {t_col_869, a[589] & a[588]} : {t_col_155, a[76] & a[77]};
assign col_156 = sel ? {t_col_868, ~a[589] & a[590]} : {t_col_156, ~a[77] & a[78]};
assign col_157 = sel ? {t_col_867, a[590] & a[589]} : {t_col_157, a[77] & a[78]};
assign col_158 = sel ? {t_col_866, ~a[590] & a[591]} : {t_col_158, ~a[78] & a[79]};
assign col_159 = sel ? {t_col_865, a[591] & a[590]} : {t_col_159, a[78] & a[79]};
assign col_160 = sel ? {t_col_864, ~a[591] & a[592]} : {t_col_160, ~a[79] & a[80]};
assign col_161 = sel ? {t_col_863, a[592] & a[591]} : {t_col_161, a[79] & a[80]};
assign col_162 = sel ? {t_col_862, ~a[592] & a[593]} : {t_col_162, ~a[80] & a[81]};
assign col_163 = sel ? {t_col_861, a[593] & a[592]} : {t_col_163, a[80] & a[81]};
assign col_164 = sel ? {t_col_860, ~a[593] & a[594]} : {t_col_164, ~a[81] & a[82]};
assign col_165 = sel ? {t_col_859, a[594] & a[593]} : {t_col_165, a[81] & a[82]};
assign col_166 = sel ? {t_col_858, ~a[594] & a[595]} : {t_col_166, ~a[82] & a[83]};
assign col_167 = sel ? {t_col_857, a[595] & a[594]} : {t_col_167, a[82] & a[83]};
assign col_168 = sel ? {t_col_856, ~a[595] & a[596]} : {t_col_168, ~a[83] & a[84]};
assign col_169 = sel ? {t_col_855, a[596] & a[595]} : {t_col_169, a[83] & a[84]};
assign col_170 = sel ? {t_col_854, ~a[596] & a[597]} : {t_col_170, ~a[84] & a[85]};
assign col_171 = sel ? {t_col_853, a[597] & a[596]} : {t_col_171, a[84] & a[85]};
assign col_172 = sel ? {t_col_852, ~a[597] & a[598]} : {t_col_172, ~a[85] & a[86]};
assign col_173 = sel ? {t_col_851, a[598] & a[597]} : {t_col_173, a[85] & a[86]};
assign col_174 = sel ? {t_col_850, ~a[598] & a[599]} : {t_col_174, ~a[86] & a[87]};
assign col_175 = sel ? {t_col_849, a[599] & a[598]} : {t_col_175, a[86] & a[87]};
assign col_176 = sel ? {t_col_848, ~a[599] & a[600]} : {t_col_176, ~a[87] & a[88]};
assign col_177 = sel ? {t_col_847, a[600] & a[599]} : {t_col_177, a[87] & a[88]};
assign col_178 = sel ? {t_col_846, ~a[600] & a[601]} : {t_col_178, ~a[88] & a[89]};
assign col_179 = sel ? {t_col_845, a[601] & a[600]} : {t_col_179, a[88] & a[89]};
assign col_180 = sel ? {t_col_844, ~a[601] & a[602]} : {t_col_180, ~a[89] & a[90]};
assign col_181 = sel ? {t_col_843, a[602] & a[601]} : {t_col_181, a[89] & a[90]};
assign col_182 = sel ? {t_col_842, ~a[602] & a[603]} : {t_col_182, ~a[90] & a[91]};
assign col_183 = sel ? {t_col_841, a[603] & a[602]} : {t_col_183, a[90] & a[91]};
assign col_184 = sel ? {t_col_840, ~a[603] & a[604]} : {t_col_184, ~a[91] & a[92]};
assign col_185 = sel ? {t_col_839, a[604] & a[603]} : {t_col_185, a[91] & a[92]};
assign col_186 = sel ? {t_col_838, ~a[604] & a[605]} : {t_col_186, ~a[92] & a[93]};
assign col_187 = sel ? {t_col_837, a[605] & a[604]} : {t_col_187, a[92] & a[93]};
assign col_188 = sel ? {t_col_836, ~a[605] & a[606]} : {t_col_188, ~a[93] & a[94]};
assign col_189 = sel ? {t_col_835, a[606] & a[605]} : {t_col_189, a[93] & a[94]};
assign col_190 = sel ? {t_col_834, ~a[606] & a[607]} : {t_col_190, ~a[94] & a[95]};
assign col_191 = sel ? {t_col_833, a[607] & a[606]} : {t_col_191, a[94] & a[95]};
assign col_192 = sel ? {t_col_832, ~a[607] & a[608]} : {t_col_192, ~a[95] & a[96]};
assign col_193 = sel ? {t_col_831, a[608] & a[607]} : {t_col_193, a[95] & a[96]};
assign col_194 = sel ? {t_col_830, ~a[608] & a[609]} : {t_col_194, ~a[96] & a[97]};
assign col_195 = sel ? {t_col_829, a[609] & a[608]} : {t_col_195, a[96] & a[97]};
assign col_196 = sel ? {t_col_828, ~a[609] & a[610]} : {t_col_196, ~a[97] & a[98]};
assign col_197 = sel ? {t_col_827, a[610] & a[609]} : {t_col_197, a[97] & a[98]};
assign col_198 = sel ? {t_col_826, ~a[610] & a[611]} : {t_col_198, ~a[98] & a[99]};
assign col_199 = sel ? {t_col_825, a[611] & a[610]} : {t_col_199, a[98] & a[99]};
assign col_200 = sel ? {t_col_824, ~a[611] & a[612]} : {t_col_200, ~a[99] & a[100]};
assign col_201 = sel ? {t_col_823, a[612] & a[611]} : {t_col_201, a[99] & a[100]};
assign col_202 = sel ? {t_col_822, ~a[612] & a[613]} : {t_col_202, ~a[100] & a[101]};
assign col_203 = sel ? {t_col_821, a[613] & a[612]} : {t_col_203, a[100] & a[101]};
assign col_204 = sel ? {t_col_820, ~a[613] & a[614]} : {t_col_204, ~a[101] & a[102]};
assign col_205 = sel ? {t_col_819, a[614] & a[613]} : {t_col_205, a[101] & a[102]};
assign col_206 = sel ? {t_col_818, ~a[614] & a[615]} : {t_col_206, ~a[102] & a[103]};
assign col_207 = sel ? {t_col_817, a[615] & a[614]} : {t_col_207, a[102] & a[103]};
assign col_208 = sel ? {t_col_816, ~a[615] & a[616]} : {t_col_208, ~a[103] & a[104]};
assign col_209 = sel ? {t_col_815, a[616] & a[615]} : {t_col_209, a[103] & a[104]};
assign col_210 = sel ? {t_col_814, ~a[616] & a[617]} : {t_col_210, ~a[104] & a[105]};
assign col_211 = sel ? {t_col_813, a[617] & a[616]} : {t_col_211, a[104] & a[105]};
assign col_212 = sel ? {t_col_812, ~a[617] & a[618]} : {t_col_212, ~a[105] & a[106]};
assign col_213 = sel ? {t_col_811, a[618] & a[617]} : {t_col_213, a[105] & a[106]};
assign col_214 = sel ? {t_col_810, ~a[618] & a[619]} : {t_col_214, ~a[106] & a[107]};
assign col_215 = sel ? {t_col_809, a[619] & a[618]} : {t_col_215, a[106] & a[107]};
assign col_216 = sel ? {t_col_808, ~a[619] & a[620]} : {t_col_216, ~a[107] & a[108]};
assign col_217 = sel ? {t_col_807, a[620] & a[619]} : {t_col_217, a[107] & a[108]};
assign col_218 = sel ? {t_col_806, ~a[620] & a[621]} : {t_col_218, ~a[108] & a[109]};
assign col_219 = sel ? {t_col_805, a[621] & a[620]} : {t_col_219, a[108] & a[109]};
assign col_220 = sel ? {t_col_804, ~a[621] & a[622]} : {t_col_220, ~a[109] & a[110]};
assign col_221 = sel ? {t_col_803, a[622] & a[621]} : {t_col_221, a[109] & a[110]};
assign col_222 = sel ? {t_col_802, ~a[622] & a[623]} : {t_col_222, ~a[110] & a[111]};
assign col_223 = sel ? {t_col_801, a[623] & a[622]} : {t_col_223, a[110] & a[111]};
assign col_224 = sel ? {t_col_800, ~a[623] & a[624]} : {t_col_224, ~a[111] & a[112]};
assign col_225 = sel ? {t_col_799, a[624] & a[623]} : {t_col_225, a[111] & a[112]};
assign col_226 = sel ? {t_col_798, ~a[624] & a[625]} : {t_col_226, ~a[112] & a[113]};
assign col_227 = sel ? {t_col_797, a[625] & a[624]} : {t_col_227, a[112] & a[113]};
assign col_228 = sel ? {t_col_796, ~a[625] & a[626]} : {t_col_228, ~a[113] & a[114]};
assign col_229 = sel ? {t_col_795, a[626] & a[625]} : {t_col_229, a[113] & a[114]};
assign col_230 = sel ? {t_col_794, ~a[626] & a[627]} : {t_col_230, ~a[114] & a[115]};
assign col_231 = sel ? {t_col_793, a[627] & a[626]} : {t_col_231, a[114] & a[115]};
assign col_232 = sel ? {t_col_792, ~a[627] & a[628]} : {t_col_232, ~a[115] & a[116]};
assign col_233 = sel ? {t_col_791, a[628] & a[627]} : {t_col_233, a[115] & a[116]};
assign col_234 = sel ? {t_col_790, ~a[628] & a[629]} : {t_col_234, ~a[116] & a[117]};
assign col_235 = sel ? {t_col_789, a[629] & a[628]} : {t_col_235, a[116] & a[117]};
assign col_236 = sel ? {t_col_788, ~a[629] & a[630]} : {t_col_236, ~a[117] & a[118]};
assign col_237 = sel ? {t_col_787, a[630] & a[629]} : {t_col_237, a[117] & a[118]};
assign col_238 = sel ? {t_col_786, ~a[630] & a[631]} : {t_col_238, ~a[118] & a[119]};
assign col_239 = sel ? {t_col_785, a[631] & a[630]} : {t_col_239, a[118] & a[119]};
assign col_240 = sel ? {t_col_784, ~a[631] & a[632]} : {t_col_240, ~a[119] & a[120]};
assign col_241 = sel ? {t_col_783, a[632] & a[631]} : {t_col_241, a[119] & a[120]};
assign col_242 = sel ? {t_col_782, ~a[632] & a[633]} : {t_col_242, ~a[120] & a[121]};
assign col_243 = sel ? {t_col_781, a[633] & a[632]} : {t_col_243, a[120] & a[121]};
assign col_244 = sel ? {t_col_780, ~a[633] & a[634]} : {t_col_244, ~a[121] & a[122]};
assign col_245 = sel ? {t_col_779, a[634] & a[633]} : {t_col_245, a[121] & a[122]};
assign col_246 = sel ? {t_col_778, ~a[634] & a[635]} : {t_col_246, ~a[122] & a[123]};
assign col_247 = sel ? {t_col_777, a[635] & a[634]} : {t_col_247, a[122] & a[123]};
assign col_248 = sel ? {t_col_776, ~a[635] & a[636]} : {t_col_248, ~a[123] & a[124]};
assign col_249 = sel ? {t_col_775, a[636] & a[635]} : {t_col_249, a[123] & a[124]};
assign col_250 = sel ? {t_col_774, ~a[636] & a[637]} : {t_col_250, ~a[124] & a[125]};
assign col_251 = sel ? {t_col_773, a[637] & a[636]} : {t_col_251, a[124] & a[125]};
assign col_252 = sel ? {t_col_772, ~a[637] & a[638]} : {t_col_252, ~a[125] & a[126]};
assign col_253 = sel ? {t_col_771, a[638] & a[637]} : {t_col_253, a[125] & a[126]};
assign col_254 = sel ? {t_col_770, ~a[638] & a[639]} : {t_col_254, ~a[126] & a[127]};
assign col_255 = sel ? {t_col_769, a[639] & a[638]} : {t_col_255, a[126] & a[127]};
assign col_256 = sel ? {t_col_768, ~a[639] & a[640]} : {t_col_256, ~a[127] & a[128]};
assign col_257 = sel ? {t_col_767, a[640] & a[639]} : {t_col_257, a[127] & a[128]};
assign col_258 = sel ? {t_col_766, ~a[640] & a[641]} : {t_col_258, ~a[128] & a[129]};
assign col_259 = sel ? {t_col_765, a[641] & a[640]} : {t_col_259, a[128] & a[129]};
assign col_260 = sel ? {t_col_764, ~a[641] & a[642]} : {t_col_260, ~a[129] & a[130]};
assign col_261 = sel ? {t_col_763, a[642] & a[641]} : {t_col_261, a[129] & a[130]};
assign col_262 = sel ? {t_col_762, ~a[642] & a[643]} : {t_col_262, ~a[130] & a[131]};
assign col_263 = sel ? {t_col_761, a[643] & a[642]} : {t_col_263, a[130] & a[131]};
assign col_264 = sel ? {t_col_760, ~a[643] & a[644]} : {t_col_264, ~a[131] & a[132]};
assign col_265 = sel ? {t_col_759, a[644] & a[643]} : {t_col_265, a[131] & a[132]};
assign col_266 = sel ? {t_col_758, ~a[644] & a[645]} : {t_col_266, ~a[132] & a[133]};
assign col_267 = sel ? {t_col_757, a[645] & a[644]} : {t_col_267, a[132] & a[133]};
assign col_268 = sel ? {t_col_756, ~a[645] & a[646]} : {t_col_268, ~a[133] & a[134]};
assign col_269 = sel ? {t_col_755, a[646] & a[645]} : {t_col_269, a[133] & a[134]};
assign col_270 = sel ? {t_col_754, ~a[646] & a[647]} : {t_col_270, ~a[134] & a[135]};
assign col_271 = sel ? {t_col_753, a[647] & a[646]} : {t_col_271, a[134] & a[135]};
assign col_272 = sel ? {t_col_752, ~a[647] & a[648]} : {t_col_272, ~a[135] & a[136]};
assign col_273 = sel ? {t_col_751, a[648] & a[647]} : {t_col_273, a[135] & a[136]};
assign col_274 = sel ? {t_col_750, ~a[648] & a[649]} : {t_col_274, ~a[136] & a[137]};
assign col_275 = sel ? {t_col_749, a[649] & a[648]} : {t_col_275, a[136] & a[137]};
assign col_276 = sel ? {t_col_748, ~a[649] & a[650]} : {t_col_276, ~a[137] & a[138]};
assign col_277 = sel ? {t_col_747, a[650] & a[649]} : {t_col_277, a[137] & a[138]};
assign col_278 = sel ? {t_col_746, ~a[650] & a[651]} : {t_col_278, ~a[138] & a[139]};
assign col_279 = sel ? {t_col_745, a[651] & a[650]} : {t_col_279, a[138] & a[139]};
assign col_280 = sel ? {t_col_744, ~a[651] & a[652]} : {t_col_280, ~a[139] & a[140]};
assign col_281 = sel ? {t_col_743, a[652] & a[651]} : {t_col_281, a[139] & a[140]};
assign col_282 = sel ? {t_col_742, ~a[652] & a[653]} : {t_col_282, ~a[140] & a[141]};
assign col_283 = sel ? {t_col_741, a[653] & a[652]} : {t_col_283, a[140] & a[141]};
assign col_284 = sel ? {t_col_740, ~a[653] & a[654]} : {t_col_284, ~a[141] & a[142]};
assign col_285 = sel ? {t_col_739, a[654] & a[653]} : {t_col_285, a[141] & a[142]};
assign col_286 = sel ? {t_col_738, ~a[654] & a[655]} : {t_col_286, ~a[142] & a[143]};
assign col_287 = sel ? {t_col_737, a[655] & a[654]} : {t_col_287, a[142] & a[143]};
assign col_288 = sel ? {t_col_736, ~a[655] & a[656]} : {t_col_288, ~a[143] & a[144]};
assign col_289 = sel ? {t_col_735, a[656] & a[655]} : {t_col_289, a[143] & a[144]};
assign col_290 = sel ? {t_col_734, ~a[656] & a[657]} : {t_col_290, ~a[144] & a[145]};
assign col_291 = sel ? {t_col_733, a[657] & a[656]} : {t_col_291, a[144] & a[145]};
assign col_292 = sel ? {t_col_732, ~a[657] & a[658]} : {t_col_292, ~a[145] & a[146]};
assign col_293 = sel ? {t_col_731, a[658] & a[657]} : {t_col_293, a[145] & a[146]};
assign col_294 = sel ? {t_col_730, ~a[658] & a[659]} : {t_col_294, ~a[146] & a[147]};
assign col_295 = sel ? {t_col_729, a[659] & a[658]} : {t_col_295, a[146] & a[147]};
assign col_296 = sel ? {t_col_728, ~a[659] & a[660]} : {t_col_296, ~a[147] & a[148]};
assign col_297 = sel ? {t_col_727, a[660] & a[659]} : {t_col_297, a[147] & a[148]};
assign col_298 = sel ? {t_col_726, ~a[660] & a[661]} : {t_col_298, ~a[148] & a[149]};
assign col_299 = sel ? {t_col_725, a[661] & a[660]} : {t_col_299, a[148] & a[149]};
assign col_300 = sel ? {t_col_724, ~a[661] & a[662]} : {t_col_300, ~a[149] & a[150]};
assign col_301 = sel ? {t_col_723, a[662] & a[661]} : {t_col_301, a[149] & a[150]};
assign col_302 = sel ? {t_col_722, ~a[662] & a[663]} : {t_col_302, ~a[150] & a[151]};
assign col_303 = sel ? {t_col_721, a[663] & a[662]} : {t_col_303, a[150] & a[151]};
assign col_304 = sel ? {t_col_720, ~a[663] & a[664]} : {t_col_304, ~a[151] & a[152]};
assign col_305 = sel ? {t_col_719, a[664] & a[663]} : {t_col_305, a[151] & a[152]};
assign col_306 = sel ? {t_col_718, ~a[664] & a[665]} : {t_col_306, ~a[152] & a[153]};
assign col_307 = sel ? {t_col_717, a[665] & a[664]} : {t_col_307, a[152] & a[153]};
assign col_308 = sel ? {t_col_716, ~a[665] & a[666]} : {t_col_308, ~a[153] & a[154]};
assign col_309 = sel ? {t_col_715, a[666] & a[665]} : {t_col_309, a[153] & a[154]};
assign col_310 = sel ? {t_col_714, ~a[666] & a[667]} : {t_col_310, ~a[154] & a[155]};
assign col_311 = sel ? {t_col_713, a[667] & a[666]} : {t_col_311, a[154] & a[155]};
assign col_312 = sel ? {t_col_712, ~a[667] & a[668]} : {t_col_312, ~a[155] & a[156]};
assign col_313 = sel ? {t_col_711, a[668] & a[667]} : {t_col_313, a[155] & a[156]};
assign col_314 = sel ? {t_col_710, ~a[668] & a[669]} : {t_col_314, ~a[156] & a[157]};
assign col_315 = sel ? {t_col_709, a[669] & a[668]} : {t_col_315, a[156] & a[157]};
assign col_316 = sel ? {t_col_708, ~a[669] & a[670]} : {t_col_316, ~a[157] & a[158]};
assign col_317 = sel ? {t_col_707, a[670] & a[669]} : {t_col_317, a[157] & a[158]};
assign col_318 = sel ? {t_col_706, ~a[670] & a[671]} : {t_col_318, ~a[158] & a[159]};
assign col_319 = sel ? {t_col_705, a[671] & a[670]} : {t_col_319, a[158] & a[159]};
assign col_320 = sel ? {t_col_704, ~a[671] & a[672]} : {t_col_320, ~a[159] & a[160]};
assign col_321 = sel ? {t_col_703, a[672] & a[671]} : {t_col_321, a[159] & a[160]};
assign col_322 = sel ? {t_col_702, ~a[672] & a[673]} : {t_col_322, ~a[160] & a[161]};
assign col_323 = sel ? {t_col_701, a[673] & a[672]} : {t_col_323, a[160] & a[161]};
assign col_324 = sel ? {t_col_700, ~a[673] & a[674]} : {t_col_324, ~a[161] & a[162]};
assign col_325 = sel ? {t_col_699, a[674] & a[673]} : {t_col_325, a[161] & a[162]};
assign col_326 = sel ? {t_col_698, ~a[674] & a[675]} : {t_col_326, ~a[162] & a[163]};
assign col_327 = sel ? {t_col_697, a[675] & a[674]} : {t_col_327, a[162] & a[163]};
assign col_328 = sel ? {t_col_696, ~a[675] & a[676]} : {t_col_328, ~a[163] & a[164]};
assign col_329 = sel ? {t_col_695, a[676] & a[675]} : {t_col_329, a[163] & a[164]};
assign col_330 = sel ? {t_col_694, ~a[676] & a[677]} : {t_col_330, ~a[164] & a[165]};
assign col_331 = sel ? {t_col_693, a[677] & a[676]} : {t_col_331, a[164] & a[165]};
assign col_332 = sel ? {t_col_692, ~a[677] & a[678]} : {t_col_332, ~a[165] & a[166]};
assign col_333 = sel ? {t_col_691, a[678] & a[677]} : {t_col_333, a[165] & a[166]};
assign col_334 = sel ? {t_col_690, ~a[678] & a[679]} : {t_col_334, ~a[166] & a[167]};
assign col_335 = sel ? {t_col_689, a[679] & a[678]} : {t_col_335, a[166] & a[167]};
assign col_336 = sel ? {t_col_688, ~a[679] & a[680]} : {t_col_336, ~a[167] & a[168]};
assign col_337 = sel ? {t_col_687, a[680] & a[679]} : {t_col_337, a[167] & a[168]};
assign col_338 = sel ? {t_col_686, ~a[680] & a[681]} : {t_col_338, ~a[168] & a[169]};
assign col_339 = sel ? {t_col_685, a[681] & a[680]} : {t_col_339, a[168] & a[169]};
assign col_340 = sel ? {t_col_684, ~a[681] & a[682]} : {t_col_340, ~a[169] & a[170]};
assign col_341 = sel ? {t_col_683, a[682] & a[681]} : {t_col_341, a[169] & a[170]};
assign col_342 = sel ? {t_col_682, ~a[682] & a[683]} : {t_col_342, ~a[170] & a[171]};
assign col_343 = sel ? {t_col_681, a[683] & a[682]} : {t_col_343, a[170] & a[171]};
assign col_344 = sel ? {t_col_680, ~a[683] & a[684]} : {t_col_344, ~a[171] & a[172]};
assign col_345 = sel ? {t_col_679, a[684] & a[683]} : {t_col_345, a[171] & a[172]};
assign col_346 = sel ? {t_col_678, ~a[684] & a[685]} : {t_col_346, ~a[172] & a[173]};
assign col_347 = sel ? {t_col_677, a[685] & a[684]} : {t_col_347, a[172] & a[173]};
assign col_348 = sel ? {t_col_676, ~a[685] & a[686]} : {t_col_348, ~a[173] & a[174]};
assign col_349 = sel ? {t_col_675, a[686] & a[685]} : {t_col_349, a[173] & a[174]};
assign col_350 = sel ? {t_col_674, ~a[686] & a[687]} : {t_col_350, ~a[174] & a[175]};
assign col_351 = sel ? {t_col_673, a[687] & a[686]} : {t_col_351, a[174] & a[175]};
assign col_352 = sel ? {t_col_672, ~a[687] & a[688]} : {t_col_352, ~a[175] & a[176]};
assign col_353 = sel ? {t_col_671, a[688] & a[687]} : {t_col_353, a[175] & a[176]};
assign col_354 = sel ? {t_col_670, ~a[688] & a[689]} : {t_col_354, ~a[176] & a[177]};
assign col_355 = sel ? {t_col_669, a[689] & a[688]} : {t_col_355, a[176] & a[177]};
assign col_356 = sel ? {t_col_668, ~a[689] & a[690]} : {t_col_356, ~a[177] & a[178]};
assign col_357 = sel ? {t_col_667, a[690] & a[689]} : {t_col_357, a[177] & a[178]};
assign col_358 = sel ? {t_col_666, ~a[690] & a[691]} : {t_col_358, ~a[178] & a[179]};
assign col_359 = sel ? {t_col_665, a[691] & a[690]} : {t_col_359, a[178] & a[179]};
assign col_360 = sel ? {t_col_664, ~a[691] & a[692]} : {t_col_360, ~a[179] & a[180]};
assign col_361 = sel ? {t_col_663, a[692] & a[691]} : {t_col_361, a[179] & a[180]};
assign col_362 = sel ? {t_col_662, ~a[692] & a[693]} : {t_col_362, ~a[180] & a[181]};
assign col_363 = sel ? {t_col_661, a[693] & a[692]} : {t_col_363, a[180] & a[181]};
assign col_364 = sel ? {t_col_660, ~a[693] & a[694]} : {t_col_364, ~a[181] & a[182]};
assign col_365 = sel ? {t_col_659, a[694] & a[693]} : {t_col_365, a[181] & a[182]};
assign col_366 = sel ? {t_col_658, ~a[694] & a[695]} : {t_col_366, ~a[182] & a[183]};
assign col_367 = sel ? {t_col_657, a[695] & a[694]} : {t_col_367, a[182] & a[183]};
assign col_368 = sel ? {t_col_656, ~a[695] & a[696]} : {t_col_368, ~a[183] & a[184]};
assign col_369 = sel ? {t_col_655, a[696] & a[695]} : {t_col_369, a[183] & a[184]};
assign col_370 = sel ? {t_col_654, ~a[696] & a[697]} : {t_col_370, ~a[184] & a[185]};
assign col_371 = sel ? {t_col_653, a[697] & a[696]} : {t_col_371, a[184] & a[185]};
assign col_372 = sel ? {t_col_652, ~a[697] & a[698]} : {t_col_372, ~a[185] & a[186]};
assign col_373 = sel ? {t_col_651, a[698] & a[697]} : {t_col_373, a[185] & a[186]};
assign col_374 = sel ? {t_col_650, ~a[698] & a[699]} : {t_col_374, ~a[186] & a[187]};
assign col_375 = sel ? {t_col_649, a[699] & a[698]} : {t_col_375, a[186] & a[187]};
assign col_376 = sel ? {t_col_648, ~a[699] & a[700]} : {t_col_376, ~a[187] & a[188]};
assign col_377 = sel ? {t_col_647, a[700] & a[699]} : {t_col_377, a[187] & a[188]};
assign col_378 = sel ? {t_col_646, ~a[700] & a[701]} : {t_col_378, ~a[188] & a[189]};
assign col_379 = sel ? {t_col_645, a[701] & a[700]} : {t_col_379, a[188] & a[189]};
assign col_380 = sel ? {t_col_644, ~a[701] & a[702]} : {t_col_380, ~a[189] & a[190]};
assign col_381 = sel ? {t_col_643, a[702] & a[701]} : {t_col_381, a[189] & a[190]};
assign col_382 = sel ? {t_col_642, ~a[702] & a[703]} : {t_col_382, ~a[190] & a[191]};
assign col_383 = sel ? {t_col_641, a[703] & a[702]} : {t_col_383, a[190] & a[191]};
assign col_384 = sel ? {t_col_640, ~a[703] & a[704]} : {t_col_384, ~a[191] & a[192]};
assign col_385 = sel ? {t_col_639, a[704] & a[703]} : {t_col_385, a[191] & a[192]};
assign col_386 = sel ? {t_col_638, ~a[704] & a[705]} : {t_col_386, ~a[192] & a[193]};
assign col_387 = sel ? {t_col_637, a[705] & a[704]} : {t_col_387, a[192] & a[193]};
assign col_388 = sel ? {t_col_636, ~a[705] & a[706]} : {t_col_388, ~a[193] & a[194]};
assign col_389 = sel ? {t_col_635, a[706] & a[705]} : {t_col_389, a[193] & a[194]};
assign col_390 = sel ? {t_col_634, ~a[706] & a[707]} : {t_col_390, ~a[194] & a[195]};
assign col_391 = sel ? {t_col_633, a[707] & a[706]} : {t_col_391, a[194] & a[195]};
assign col_392 = sel ? {t_col_632, ~a[707] & a[708]} : {t_col_392, ~a[195] & a[196]};
assign col_393 = sel ? {t_col_631, a[708] & a[707]} : {t_col_393, a[195] & a[196]};
assign col_394 = sel ? {t_col_630, ~a[708] & a[709]} : {t_col_394, ~a[196] & a[197]};
assign col_395 = sel ? {t_col_629, a[709] & a[708]} : {t_col_395, a[196] & a[197]};
assign col_396 = sel ? {t_col_628, ~a[709] & a[710]} : {t_col_396, ~a[197] & a[198]};
assign col_397 = sel ? {t_col_627, a[710] & a[709]} : {t_col_397, a[197] & a[198]};
assign col_398 = sel ? {t_col_626, ~a[710] & a[711]} : {t_col_398, ~a[198] & a[199]};
assign col_399 = sel ? {t_col_625, a[711] & a[710]} : {t_col_399, a[198] & a[199]};
assign col_400 = sel ? {t_col_624, ~a[711] & a[712]} : {t_col_400, ~a[199] & a[200]};
assign col_401 = sel ? {t_col_623, a[712] & a[711]} : {t_col_401, a[199] & a[200]};
assign col_402 = sel ? {t_col_622, ~a[712] & a[713]} : {t_col_402, ~a[200] & a[201]};
assign col_403 = sel ? {t_col_621, a[713] & a[712]} : {t_col_403, a[200] & a[201]};
assign col_404 = sel ? {t_col_620, ~a[713] & a[714]} : {t_col_404, ~a[201] & a[202]};
assign col_405 = sel ? {t_col_619, a[714] & a[713]} : {t_col_405, a[201] & a[202]};
assign col_406 = sel ? {t_col_618, ~a[714] & a[715]} : {t_col_406, ~a[202] & a[203]};
assign col_407 = sel ? {t_col_617, a[715] & a[714]} : {t_col_407, a[202] & a[203]};
assign col_408 = sel ? {t_col_616, ~a[715] & a[716]} : {t_col_408, ~a[203] & a[204]};
assign col_409 = sel ? {t_col_615, a[716] & a[715]} : {t_col_409, a[203] & a[204]};
assign col_410 = sel ? {t_col_614, ~a[716] & a[717]} : {t_col_410, ~a[204] & a[205]};
assign col_411 = sel ? {t_col_613, a[717] & a[716]} : {t_col_411, a[204] & a[205]};
assign col_412 = sel ? {t_col_612, ~a[717] & a[718]} : {t_col_412, ~a[205] & a[206]};
assign col_413 = sel ? {t_col_611, a[718] & a[717]} : {t_col_413, a[205] & a[206]};
assign col_414 = sel ? {t_col_610, ~a[718] & a[719]} : {t_col_414, ~a[206] & a[207]};
assign col_415 = sel ? {t_col_609, a[719] & a[718]} : {t_col_415, a[206] & a[207]};
assign col_416 = sel ? {t_col_608, ~a[719] & a[720]} : {t_col_416, ~a[207] & a[208]};
assign col_417 = sel ? {t_col_607, a[720] & a[719]} : {t_col_417, a[207] & a[208]};
assign col_418 = sel ? {t_col_606, ~a[720] & a[721]} : {t_col_418, ~a[208] & a[209]};
assign col_419 = sel ? {t_col_605, a[721] & a[720]} : {t_col_419, a[208] & a[209]};
assign col_420 = sel ? {t_col_604, ~a[721] & a[722]} : {t_col_420, ~a[209] & a[210]};
assign col_421 = sel ? {t_col_603, a[722] & a[721]} : {t_col_421, a[209] & a[210]};
assign col_422 = sel ? {t_col_602, ~a[722] & a[723]} : {t_col_422, ~a[210] & a[211]};
assign col_423 = sel ? {t_col_601, a[723] & a[722]} : {t_col_423, a[210] & a[211]};
assign col_424 = sel ? {t_col_600, ~a[723] & a[724]} : {t_col_424, ~a[211] & a[212]};
assign col_425 = sel ? {t_col_599, a[724] & a[723]} : {t_col_425, a[211] & a[212]};
assign col_426 = sel ? {t_col_598, ~a[724] & a[725]} : {t_col_426, ~a[212] & a[213]};
assign col_427 = sel ? {t_col_597, a[725] & a[724]} : {t_col_427, a[212] & a[213]};
assign col_428 = sel ? {t_col_596, ~a[725] & a[726]} : {t_col_428, ~a[213] & a[214]};
assign col_429 = sel ? {t_col_595, a[726] & a[725]} : {t_col_429, a[213] & a[214]};
assign col_430 = sel ? {t_col_594, ~a[726] & a[727]} : {t_col_430, ~a[214] & a[215]};
assign col_431 = sel ? {t_col_593, a[727] & a[726]} : {t_col_431, a[214] & a[215]};
assign col_432 = sel ? {t_col_592, ~a[727] & a[728]} : {t_col_432, ~a[215] & a[216]};
assign col_433 = sel ? {t_col_591, a[728] & a[727]} : {t_col_433, a[215] & a[216]};
assign col_434 = sel ? {t_col_590, ~a[728] & a[729]} : {t_col_434, ~a[216] & a[217]};
assign col_435 = sel ? {t_col_589, a[729] & a[728]} : {t_col_435, a[216] & a[217]};
assign col_436 = sel ? {t_col_588, ~a[729] & a[730]} : {t_col_436, ~a[217] & a[218]};
assign col_437 = sel ? {t_col_587, a[730] & a[729]} : {t_col_437, a[217] & a[218]};
assign col_438 = sel ? {t_col_586, ~a[730] & a[731]} : {t_col_438, ~a[218] & a[219]};
assign col_439 = sel ? {t_col_585, a[731] & a[730]} : {t_col_439, a[218] & a[219]};
assign col_440 = sel ? {t_col_584, ~a[731] & a[732]} : {t_col_440, ~a[219] & a[220]};
assign col_441 = sel ? {t_col_583, a[732] & a[731]} : {t_col_441, a[219] & a[220]};
assign col_442 = sel ? {t_col_582, ~a[732] & a[733]} : {t_col_442, ~a[220] & a[221]};
assign col_443 = sel ? {t_col_581, a[733] & a[732]} : {t_col_443, a[220] & a[221]};
assign col_444 = sel ? {t_col_580, ~a[733] & a[734]} : {t_col_444, ~a[221] & a[222]};
assign col_445 = sel ? {t_col_579, a[734] & a[733]} : {t_col_445, a[221] & a[222]};
assign col_446 = sel ? {t_col_578, ~a[734] & a[735]} : {t_col_446, ~a[222] & a[223]};
assign col_447 = sel ? {t_col_577, a[735] & a[734]} : {t_col_447, a[222] & a[223]};
assign col_448 = sel ? {t_col_576, ~a[735] & a[736]} : {t_col_448, ~a[223] & a[224]};
assign col_449 = sel ? {t_col_575, a[736] & a[735]} : {t_col_449, a[223] & a[224]};
assign col_450 = sel ? {t_col_574, ~a[736] & a[737]} : {t_col_450, ~a[224] & a[225]};
assign col_451 = sel ? {t_col_573, a[737] & a[736]} : {t_col_451, a[224] & a[225]};
assign col_452 = sel ? {t_col_572, ~a[737] & a[738]} : {t_col_452, ~a[225] & a[226]};
assign col_453 = sel ? {t_col_571, a[738] & a[737]} : {t_col_453, a[225] & a[226]};
assign col_454 = sel ? {t_col_570, ~a[738] & a[739]} : {t_col_454, ~a[226] & a[227]};
assign col_455 = sel ? {t_col_569, a[739] & a[738]} : {t_col_455, a[226] & a[227]};
assign col_456 = sel ? {t_col_568, ~a[739] & a[740]} : {t_col_456, ~a[227] & a[228]};
assign col_457 = sel ? {t_col_567, a[740] & a[739]} : {t_col_457, a[227] & a[228]};
assign col_458 = sel ? {t_col_566, ~a[740] & a[741]} : {t_col_458, ~a[228] & a[229]};
assign col_459 = sel ? {t_col_565, a[741] & a[740]} : {t_col_459, a[228] & a[229]};
assign col_460 = sel ? {t_col_564, ~a[741] & a[742]} : {t_col_460, ~a[229] & a[230]};
assign col_461 = sel ? {t_col_563, a[742] & a[741]} : {t_col_461, a[229] & a[230]};
assign col_462 = sel ? {t_col_562, ~a[742] & a[743]} : {t_col_462, ~a[230] & a[231]};
assign col_463 = sel ? {t_col_561, a[743] & a[742]} : {t_col_463, a[230] & a[231]};
assign col_464 = sel ? {t_col_560, ~a[743] & a[744]} : {t_col_464, ~a[231] & a[232]};
assign col_465 = sel ? {t_col_559, a[744] & a[743]} : {t_col_465, a[231] & a[232]};
assign col_466 = sel ? {t_col_558, ~a[744] & a[745]} : {t_col_466, ~a[232] & a[233]};
assign col_467 = sel ? {t_col_557, a[745] & a[744]} : {t_col_467, a[232] & a[233]};
assign col_468 = sel ? {t_col_556, ~a[745] & a[746]} : {t_col_468, ~a[233] & a[234]};
assign col_469 = sel ? {t_col_555, a[746] & a[745]} : {t_col_469, a[233] & a[234]};
assign col_470 = sel ? {t_col_554, ~a[746] & a[747]} : {t_col_470, ~a[234] & a[235]};
assign col_471 = sel ? {t_col_553, a[747] & a[746]} : {t_col_471, a[234] & a[235]};
assign col_472 = sel ? {t_col_552, ~a[747] & a[748]} : {t_col_472, ~a[235] & a[236]};
assign col_473 = sel ? {t_col_551, a[748] & a[747]} : {t_col_473, a[235] & a[236]};
assign col_474 = sel ? {t_col_550, ~a[748] & a[749]} : {t_col_474, ~a[236] & a[237]};
assign col_475 = sel ? {t_col_549, a[749] & a[748]} : {t_col_475, a[236] & a[237]};
assign col_476 = sel ? {t_col_548, ~a[749] & a[750]} : {t_col_476, ~a[237] & a[238]};
assign col_477 = sel ? {t_col_547, a[750] & a[749]} : {t_col_477, a[237] & a[238]};
assign col_478 = sel ? {t_col_546, ~a[750] & a[751]} : {t_col_478, ~a[238] & a[239]};
assign col_479 = sel ? {t_col_545, a[751] & a[750]} : {t_col_479, a[238] & a[239]};
assign col_480 = sel ? {t_col_544, ~a[751] & a[752]} : {t_col_480, ~a[239] & a[240]};
assign col_481 = sel ? {t_col_543, a[752] & a[751]} : {t_col_481, a[239] & a[240]};
assign col_482 = sel ? {t_col_542, ~a[752] & a[753]} : {t_col_482, ~a[240] & a[241]};
assign col_483 = sel ? {t_col_541, a[753] & a[752]} : {t_col_483, a[240] & a[241]};
assign col_484 = sel ? {t_col_540, ~a[753] & a[754]} : {t_col_484, ~a[241] & a[242]};
assign col_485 = sel ? {t_col_539, a[754] & a[753]} : {t_col_485, a[241] & a[242]};
assign col_486 = sel ? {t_col_538, ~a[754] & a[755]} : {t_col_486, ~a[242] & a[243]};
assign col_487 = sel ? {t_col_537, a[755] & a[754]} : {t_col_487, a[242] & a[243]};
assign col_488 = sel ? {t_col_536, ~a[755] & a[756]} : {t_col_488, ~a[243] & a[244]};
assign col_489 = sel ? {t_col_535, a[756] & a[755]} : {t_col_489, a[243] & a[244]};
assign col_490 = sel ? {t_col_534, ~a[756] & a[757]} : {t_col_490, ~a[244] & a[245]};
assign col_491 = sel ? {t_col_533, a[757] & a[756]} : {t_col_491, a[244] & a[245]};
assign col_492 = sel ? {t_col_532, ~a[757] & a[758]} : {t_col_492, ~a[245] & a[246]};
assign col_493 = sel ? {t_col_531, a[758] & a[757]} : {t_col_493, a[245] & a[246]};
assign col_494 = sel ? {t_col_530, ~a[758] & a[759]} : {t_col_494, ~a[246] & a[247]};
assign col_495 = sel ? {t_col_529, a[759] & a[758]} : {t_col_495, a[246] & a[247]};
assign col_496 = sel ? {t_col_528, ~a[759] & a[760]} : {t_col_496, ~a[247] & a[248]};
assign col_497 = sel ? {t_col_527, a[760] & a[759]} : {t_col_497, a[247] & a[248]};
assign col_498 = sel ? {t_col_526, ~a[760] & a[761]} : {t_col_498, ~a[248] & a[249]};
assign col_499 = sel ? {t_col_525, a[761] & a[760]} : {t_col_499, a[248] & a[249]};
assign col_500 = sel ? {t_col_524, ~a[761] & a[762]} : {t_col_500, ~a[249] & a[250]};
assign col_501 = sel ? {t_col_523, a[762] & a[761]} : {t_col_501, a[249] & a[250]};
assign col_502 = sel ? {t_col_522, ~a[762] & a[763]} : {t_col_502, ~a[250] & a[251]};
assign col_503 = sel ? {t_col_521, a[763] & a[762]} : {t_col_503, a[250] & a[251]};
assign col_504 = sel ? {t_col_520, ~a[763] & a[764]} : {t_col_504, ~a[251] & a[252]};
assign col_505 = sel ? {t_col_519, a[764] & a[763]} : {t_col_505, a[251] & a[252]};
assign col_506 = sel ? {t_col_518, ~a[764] & a[765]} : {t_col_506, ~a[252] & a[253]};
assign col_507 = sel ? {t_col_517, a[765] & a[764]} : {t_col_507, a[252] & a[253]};
assign col_508 = sel ? {t_col_516, ~a[765] & a[766]} : {t_col_508, ~a[253] & a[254]};
assign col_509 = sel ? {t_col_515, a[766] & a[765]} : {t_col_509, a[253] & a[254]};
assign col_510 = sel ? {t_col_514, ~a[766] & a[767]} : {t_col_510, ~a[254] & a[255]};
assign col_511 = sel ? {t_col_513, a[767] & a[766]} : {t_col_511, a[254] & a[255]};
assign col_512 = sel ? {t_col_512, ~a[767] & a[768]} : {t_col_512, ~a[255] & a[256]};
assign col_513 = sel ? {t_col_511, a[768] & a[767]} : {t_col_513, a[255] & a[256]};
assign col_514 = sel ? {t_col_510, ~a[768] & a[769]} : {t_col_514, ~a[256] & a[257]};
assign col_515 = sel ? {t_col_509, a[769] & a[768]} : {t_col_515, a[256] & a[257]};
assign col_516 = sel ? {t_col_508, ~a[769] & a[770]} : {t_col_516, ~a[257] & a[258]};
assign col_517 = sel ? {t_col_507, a[770] & a[769]} : {t_col_517, a[257] & a[258]};
assign col_518 = sel ? {t_col_506, ~a[770] & a[771]} : {t_col_518, ~a[258] & a[259]};
assign col_519 = sel ? {t_col_505, a[771] & a[770]} : {t_col_519, a[258] & a[259]};
assign col_520 = sel ? {t_col_504, ~a[771] & a[772]} : {t_col_520, ~a[259] & a[260]};
assign col_521 = sel ? {t_col_503, a[772] & a[771]} : {t_col_521, a[259] & a[260]};
assign col_522 = sel ? {t_col_502, ~a[772] & a[773]} : {t_col_522, ~a[260] & a[261]};
assign col_523 = sel ? {t_col_501, a[773] & a[772]} : {t_col_523, a[260] & a[261]};
assign col_524 = sel ? {t_col_500, ~a[773] & a[774]} : {t_col_524, ~a[261] & a[262]};
assign col_525 = sel ? {t_col_499, a[774] & a[773]} : {t_col_525, a[261] & a[262]};
assign col_526 = sel ? {t_col_498, ~a[774] & a[775]} : {t_col_526, ~a[262] & a[263]};
assign col_527 = sel ? {t_col_497, a[775] & a[774]} : {t_col_527, a[262] & a[263]};
assign col_528 = sel ? {t_col_496, ~a[775] & a[776]} : {t_col_528, ~a[263] & a[264]};
assign col_529 = sel ? {t_col_495, a[776] & a[775]} : {t_col_529, a[263] & a[264]};
assign col_530 = sel ? {t_col_494, ~a[776] & a[777]} : {t_col_530, ~a[264] & a[265]};
assign col_531 = sel ? {t_col_493, a[777] & a[776]} : {t_col_531, a[264] & a[265]};
assign col_532 = sel ? {t_col_492, ~a[777] & a[778]} : {t_col_532, ~a[265] & a[266]};
assign col_533 = sel ? {t_col_491, a[778] & a[777]} : {t_col_533, a[265] & a[266]};
assign col_534 = sel ? {t_col_490, ~a[778] & a[779]} : {t_col_534, ~a[266] & a[267]};
assign col_535 = sel ? {t_col_489, a[779] & a[778]} : {t_col_535, a[266] & a[267]};
assign col_536 = sel ? {t_col_488, ~a[779] & a[780]} : {t_col_536, ~a[267] & a[268]};
assign col_537 = sel ? {t_col_487, a[780] & a[779]} : {t_col_537, a[267] & a[268]};
assign col_538 = sel ? {t_col_486, ~a[780] & a[781]} : {t_col_538, ~a[268] & a[269]};
assign col_539 = sel ? {t_col_485, a[781] & a[780]} : {t_col_539, a[268] & a[269]};
assign col_540 = sel ? {t_col_484, ~a[781] & a[782]} : {t_col_540, ~a[269] & a[270]};
assign col_541 = sel ? {t_col_483, a[782] & a[781]} : {t_col_541, a[269] & a[270]};
assign col_542 = sel ? {t_col_482, ~a[782] & a[783]} : {t_col_542, ~a[270] & a[271]};
assign col_543 = sel ? {t_col_481, a[783] & a[782]} : {t_col_543, a[270] & a[271]};
assign col_544 = sel ? {t_col_480, ~a[783] & a[784]} : {t_col_544, ~a[271] & a[272]};
assign col_545 = sel ? {t_col_479, a[784] & a[783]} : {t_col_545, a[271] & a[272]};
assign col_546 = sel ? {t_col_478, ~a[784] & a[785]} : {t_col_546, ~a[272] & a[273]};
assign col_547 = sel ? {t_col_477, a[785] & a[784]} : {t_col_547, a[272] & a[273]};
assign col_548 = sel ? {t_col_476, ~a[785] & a[786]} : {t_col_548, ~a[273] & a[274]};
assign col_549 = sel ? {t_col_475, a[786] & a[785]} : {t_col_549, a[273] & a[274]};
assign col_550 = sel ? {t_col_474, ~a[786] & a[787]} : {t_col_550, ~a[274] & a[275]};
assign col_551 = sel ? {t_col_473, a[787] & a[786]} : {t_col_551, a[274] & a[275]};
assign col_552 = sel ? {t_col_472, ~a[787] & a[788]} : {t_col_552, ~a[275] & a[276]};
assign col_553 = sel ? {t_col_471, a[788] & a[787]} : {t_col_553, a[275] & a[276]};
assign col_554 = sel ? {t_col_470, ~a[788] & a[789]} : {t_col_554, ~a[276] & a[277]};
assign col_555 = sel ? {t_col_469, a[789] & a[788]} : {t_col_555, a[276] & a[277]};
assign col_556 = sel ? {t_col_468, ~a[789] & a[790]} : {t_col_556, ~a[277] & a[278]};
assign col_557 = sel ? {t_col_467, a[790] & a[789]} : {t_col_557, a[277] & a[278]};
assign col_558 = sel ? {t_col_466, ~a[790] & a[791]} : {t_col_558, ~a[278] & a[279]};
assign col_559 = sel ? {t_col_465, a[791] & a[790]} : {t_col_559, a[278] & a[279]};
assign col_560 = sel ? {t_col_464, ~a[791] & a[792]} : {t_col_560, ~a[279] & a[280]};
assign col_561 = sel ? {t_col_463, a[792] & a[791]} : {t_col_561, a[279] & a[280]};
assign col_562 = sel ? {t_col_462, ~a[792] & a[793]} : {t_col_562, ~a[280] & a[281]};
assign col_563 = sel ? {t_col_461, a[793] & a[792]} : {t_col_563, a[280] & a[281]};
assign col_564 = sel ? {t_col_460, ~a[793] & a[794]} : {t_col_564, ~a[281] & a[282]};
assign col_565 = sel ? {t_col_459, a[794] & a[793]} : {t_col_565, a[281] & a[282]};
assign col_566 = sel ? {t_col_458, ~a[794] & a[795]} : {t_col_566, ~a[282] & a[283]};
assign col_567 = sel ? {t_col_457, a[795] & a[794]} : {t_col_567, a[282] & a[283]};
assign col_568 = sel ? {t_col_456, ~a[795] & a[796]} : {t_col_568, ~a[283] & a[284]};
assign col_569 = sel ? {t_col_455, a[796] & a[795]} : {t_col_569, a[283] & a[284]};
assign col_570 = sel ? {t_col_454, ~a[796] & a[797]} : {t_col_570, ~a[284] & a[285]};
assign col_571 = sel ? {t_col_453, a[797] & a[796]} : {t_col_571, a[284] & a[285]};
assign col_572 = sel ? {t_col_452, ~a[797] & a[798]} : {t_col_572, ~a[285] & a[286]};
assign col_573 = sel ? {t_col_451, a[798] & a[797]} : {t_col_573, a[285] & a[286]};
assign col_574 = sel ? {t_col_450, ~a[798] & a[799]} : {t_col_574, ~a[286] & a[287]};
assign col_575 = sel ? {t_col_449, a[799] & a[798]} : {t_col_575, a[286] & a[287]};
assign col_576 = sel ? {t_col_448, ~a[799] & a[800]} : {t_col_576, ~a[287] & a[288]};
assign col_577 = sel ? {t_col_447, a[800] & a[799]} : {t_col_577, a[287] & a[288]};
assign col_578 = sel ? {t_col_446, ~a[800] & a[801]} : {t_col_578, ~a[288] & a[289]};
assign col_579 = sel ? {t_col_445, a[801] & a[800]} : {t_col_579, a[288] & a[289]};
assign col_580 = sel ? {t_col_444, ~a[801] & a[802]} : {t_col_580, ~a[289] & a[290]};
assign col_581 = sel ? {t_col_443, a[802] & a[801]} : {t_col_581, a[289] & a[290]};
assign col_582 = sel ? {t_col_442, ~a[802] & a[803]} : {t_col_582, ~a[290] & a[291]};
assign col_583 = sel ? {t_col_441, a[803] & a[802]} : {t_col_583, a[290] & a[291]};
assign col_584 = sel ? {t_col_440, ~a[803] & a[804]} : {t_col_584, ~a[291] & a[292]};
assign col_585 = sel ? {t_col_439, a[804] & a[803]} : {t_col_585, a[291] & a[292]};
assign col_586 = sel ? {t_col_438, ~a[804] & a[805]} : {t_col_586, ~a[292] & a[293]};
assign col_587 = sel ? {t_col_437, a[805] & a[804]} : {t_col_587, a[292] & a[293]};
assign col_588 = sel ? {t_col_436, ~a[805] & a[806]} : {t_col_588, ~a[293] & a[294]};
assign col_589 = sel ? {t_col_435, a[806] & a[805]} : {t_col_589, a[293] & a[294]};
assign col_590 = sel ? {t_col_434, ~a[806] & a[807]} : {t_col_590, ~a[294] & a[295]};
assign col_591 = sel ? {t_col_433, a[807] & a[806]} : {t_col_591, a[294] & a[295]};
assign col_592 = sel ? {t_col_432, ~a[807] & a[808]} : {t_col_592, ~a[295] & a[296]};
assign col_593 = sel ? {t_col_431, a[808] & a[807]} : {t_col_593, a[295] & a[296]};
assign col_594 = sel ? {t_col_430, ~a[808] & a[809]} : {t_col_594, ~a[296] & a[297]};
assign col_595 = sel ? {t_col_429, a[809] & a[808]} : {t_col_595, a[296] & a[297]};
assign col_596 = sel ? {t_col_428, ~a[809] & a[810]} : {t_col_596, ~a[297] & a[298]};
assign col_597 = sel ? {t_col_427, a[810] & a[809]} : {t_col_597, a[297] & a[298]};
assign col_598 = sel ? {t_col_426, ~a[810] & a[811]} : {t_col_598, ~a[298] & a[299]};
assign col_599 = sel ? {t_col_425, a[811] & a[810]} : {t_col_599, a[298] & a[299]};
assign col_600 = sel ? {t_col_424, ~a[811] & a[812]} : {t_col_600, ~a[299] & a[300]};
assign col_601 = sel ? {t_col_423, a[812] & a[811]} : {t_col_601, a[299] & a[300]};
assign col_602 = sel ? {t_col_422, ~a[812] & a[813]} : {t_col_602, ~a[300] & a[301]};
assign col_603 = sel ? {t_col_421, a[813] & a[812]} : {t_col_603, a[300] & a[301]};
assign col_604 = sel ? {t_col_420, ~a[813] & a[814]} : {t_col_604, ~a[301] & a[302]};
assign col_605 = sel ? {t_col_419, a[814] & a[813]} : {t_col_605, a[301] & a[302]};
assign col_606 = sel ? {t_col_418, ~a[814] & a[815]} : {t_col_606, ~a[302] & a[303]};
assign col_607 = sel ? {t_col_417, a[815] & a[814]} : {t_col_607, a[302] & a[303]};
assign col_608 = sel ? {t_col_416, ~a[815] & a[816]} : {t_col_608, ~a[303] & a[304]};
assign col_609 = sel ? {t_col_415, a[816] & a[815]} : {t_col_609, a[303] & a[304]};
assign col_610 = sel ? {t_col_414, ~a[816] & a[817]} : {t_col_610, ~a[304] & a[305]};
assign col_611 = sel ? {t_col_413, a[817] & a[816]} : {t_col_611, a[304] & a[305]};
assign col_612 = sel ? {t_col_412, ~a[817] & a[818]} : {t_col_612, ~a[305] & a[306]};
assign col_613 = sel ? {t_col_411, a[818] & a[817]} : {t_col_613, a[305] & a[306]};
assign col_614 = sel ? {t_col_410, ~a[818] & a[819]} : {t_col_614, ~a[306] & a[307]};
assign col_615 = sel ? {t_col_409, a[819] & a[818]} : {t_col_615, a[306] & a[307]};
assign col_616 = sel ? {t_col_408, ~a[819] & a[820]} : {t_col_616, ~a[307] & a[308]};
assign col_617 = sel ? {t_col_407, a[820] & a[819]} : {t_col_617, a[307] & a[308]};
assign col_618 = sel ? {t_col_406, ~a[820] & a[821]} : {t_col_618, ~a[308] & a[309]};
assign col_619 = sel ? {t_col_405, a[821] & a[820]} : {t_col_619, a[308] & a[309]};
assign col_620 = sel ? {t_col_404, ~a[821] & a[822]} : {t_col_620, ~a[309] & a[310]};
assign col_621 = sel ? {t_col_403, a[822] & a[821]} : {t_col_621, a[309] & a[310]};
assign col_622 = sel ? {t_col_402, ~a[822] & a[823]} : {t_col_622, ~a[310] & a[311]};
assign col_623 = sel ? {t_col_401, a[823] & a[822]} : {t_col_623, a[310] & a[311]};
assign col_624 = sel ? {t_col_400, ~a[823] & a[824]} : {t_col_624, ~a[311] & a[312]};
assign col_625 = sel ? {t_col_399, a[824] & a[823]} : {t_col_625, a[311] & a[312]};
assign col_626 = sel ? {t_col_398, ~a[824] & a[825]} : {t_col_626, ~a[312] & a[313]};
assign col_627 = sel ? {t_col_397, a[825] & a[824]} : {t_col_627, a[312] & a[313]};
assign col_628 = sel ? {t_col_396, ~a[825] & a[826]} : {t_col_628, ~a[313] & a[314]};
assign col_629 = sel ? {t_col_395, a[826] & a[825]} : {t_col_629, a[313] & a[314]};
assign col_630 = sel ? {t_col_394, ~a[826] & a[827]} : {t_col_630, ~a[314] & a[315]};
assign col_631 = sel ? {t_col_393, a[827] & a[826]} : {t_col_631, a[314] & a[315]};
assign col_632 = sel ? {t_col_392, ~a[827] & a[828]} : {t_col_632, ~a[315] & a[316]};
assign col_633 = sel ? {t_col_391, a[828] & a[827]} : {t_col_633, a[315] & a[316]};
assign col_634 = sel ? {t_col_390, ~a[828] & a[829]} : {t_col_634, ~a[316] & a[317]};
assign col_635 = sel ? {t_col_389, a[829] & a[828]} : {t_col_635, a[316] & a[317]};
assign col_636 = sel ? {t_col_388, ~a[829] & a[830]} : {t_col_636, ~a[317] & a[318]};
assign col_637 = sel ? {t_col_387, a[830] & a[829]} : {t_col_637, a[317] & a[318]};
assign col_638 = sel ? {t_col_386, ~a[830] & a[831]} : {t_col_638, ~a[318] & a[319]};
assign col_639 = sel ? {t_col_385, a[831] & a[830]} : {t_col_639, a[318] & a[319]};
assign col_640 = sel ? {t_col_384, ~a[831] & a[832]} : {t_col_640, ~a[319] & a[320]};
assign col_641 = sel ? {t_col_383, a[832] & a[831]} : {t_col_641, a[319] & a[320]};
assign col_642 = sel ? {t_col_382, ~a[832] & a[833]} : {t_col_642, ~a[320] & a[321]};
assign col_643 = sel ? {t_col_381, a[833] & a[832]} : {t_col_643, a[320] & a[321]};
assign col_644 = sel ? {t_col_380, ~a[833] & a[834]} : {t_col_644, ~a[321] & a[322]};
assign col_645 = sel ? {t_col_379, a[834] & a[833]} : {t_col_645, a[321] & a[322]};
assign col_646 = sel ? {t_col_378, ~a[834] & a[835]} : {t_col_646, ~a[322] & a[323]};
assign col_647 = sel ? {t_col_377, a[835] & a[834]} : {t_col_647, a[322] & a[323]};
assign col_648 = sel ? {t_col_376, ~a[835] & a[836]} : {t_col_648, ~a[323] & a[324]};
assign col_649 = sel ? {t_col_375, a[836] & a[835]} : {t_col_649, a[323] & a[324]};
assign col_650 = sel ? {t_col_374, ~a[836] & a[837]} : {t_col_650, ~a[324] & a[325]};
assign col_651 = sel ? {t_col_373, a[837] & a[836]} : {t_col_651, a[324] & a[325]};
assign col_652 = sel ? {t_col_372, ~a[837] & a[838]} : {t_col_652, ~a[325] & a[326]};
assign col_653 = sel ? {t_col_371, a[838] & a[837]} : {t_col_653, a[325] & a[326]};
assign col_654 = sel ? {t_col_370, ~a[838] & a[839]} : {t_col_654, ~a[326] & a[327]};
assign col_655 = sel ? {t_col_369, a[839] & a[838]} : {t_col_655, a[326] & a[327]};
assign col_656 = sel ? {t_col_368, ~a[839] & a[840]} : {t_col_656, ~a[327] & a[328]};
assign col_657 = sel ? {t_col_367, a[840] & a[839]} : {t_col_657, a[327] & a[328]};
assign col_658 = sel ? {t_col_366, ~a[840] & a[841]} : {t_col_658, ~a[328] & a[329]};
assign col_659 = sel ? {t_col_365, a[841] & a[840]} : {t_col_659, a[328] & a[329]};
assign col_660 = sel ? {t_col_364, ~a[841] & a[842]} : {t_col_660, ~a[329] & a[330]};
assign col_661 = sel ? {t_col_363, a[842] & a[841]} : {t_col_661, a[329] & a[330]};
assign col_662 = sel ? {t_col_362, ~a[842] & a[843]} : {t_col_662, ~a[330] & a[331]};
assign col_663 = sel ? {t_col_361, a[843] & a[842]} : {t_col_663, a[330] & a[331]};
assign col_664 = sel ? {t_col_360, ~a[843] & a[844]} : {t_col_664, ~a[331] & a[332]};
assign col_665 = sel ? {t_col_359, a[844] & a[843]} : {t_col_665, a[331] & a[332]};
assign col_666 = sel ? {t_col_358, ~a[844] & a[845]} : {t_col_666, ~a[332] & a[333]};
assign col_667 = sel ? {t_col_357, a[845] & a[844]} : {t_col_667, a[332] & a[333]};
assign col_668 = sel ? {t_col_356, ~a[845] & a[846]} : {t_col_668, ~a[333] & a[334]};
assign col_669 = sel ? {t_col_355, a[846] & a[845]} : {t_col_669, a[333] & a[334]};
assign col_670 = sel ? {t_col_354, ~a[846] & a[847]} : {t_col_670, ~a[334] & a[335]};
assign col_671 = sel ? {t_col_353, a[847] & a[846]} : {t_col_671, a[334] & a[335]};
assign col_672 = sel ? {t_col_352, ~a[847] & a[848]} : {t_col_672, ~a[335] & a[336]};
assign col_673 = sel ? {t_col_351, a[848] & a[847]} : {t_col_673, a[335] & a[336]};
assign col_674 = sel ? {t_col_350, ~a[848] & a[849]} : {t_col_674, ~a[336] & a[337]};
assign col_675 = sel ? {t_col_349, a[849] & a[848]} : {t_col_675, a[336] & a[337]};
assign col_676 = sel ? {t_col_348, ~a[849] & a[850]} : {t_col_676, ~a[337] & a[338]};
assign col_677 = sel ? {t_col_347, a[850] & a[849]} : {t_col_677, a[337] & a[338]};
assign col_678 = sel ? {t_col_346, ~a[850] & a[851]} : {t_col_678, ~a[338] & a[339]};
assign col_679 = sel ? {t_col_345, a[851] & a[850]} : {t_col_679, a[338] & a[339]};
assign col_680 = sel ? {t_col_344, ~a[851] & a[852]} : {t_col_680, ~a[339] & a[340]};
assign col_681 = sel ? {t_col_343, a[852] & a[851]} : {t_col_681, a[339] & a[340]};
assign col_682 = sel ? {t_col_342, ~a[852] & a[853]} : {t_col_682, ~a[340] & a[341]};
assign col_683 = sel ? {t_col_341, a[853] & a[852]} : {t_col_683, a[340] & a[341]};
assign col_684 = sel ? {t_col_340, ~a[853] & a[854]} : {t_col_684, ~a[341] & a[342]};
assign col_685 = sel ? {t_col_339, a[854] & a[853]} : {t_col_685, a[341] & a[342]};
assign col_686 = sel ? {t_col_338, ~a[854] & a[855]} : {t_col_686, ~a[342] & a[343]};
assign col_687 = sel ? {t_col_337, a[855] & a[854]} : {t_col_687, a[342] & a[343]};
assign col_688 = sel ? {t_col_336, ~a[855] & a[856]} : {t_col_688, ~a[343] & a[344]};
assign col_689 = sel ? {t_col_335, a[856] & a[855]} : {t_col_689, a[343] & a[344]};
assign col_690 = sel ? {t_col_334, ~a[856] & a[857]} : {t_col_690, ~a[344] & a[345]};
assign col_691 = sel ? {t_col_333, a[857] & a[856]} : {t_col_691, a[344] & a[345]};
assign col_692 = sel ? {t_col_332, ~a[857] & a[858]} : {t_col_692, ~a[345] & a[346]};
assign col_693 = sel ? {t_col_331, a[858] & a[857]} : {t_col_693, a[345] & a[346]};
assign col_694 = sel ? {t_col_330, ~a[858] & a[859]} : {t_col_694, ~a[346] & a[347]};
assign col_695 = sel ? {t_col_329, a[859] & a[858]} : {t_col_695, a[346] & a[347]};
assign col_696 = sel ? {t_col_328, ~a[859] & a[860]} : {t_col_696, ~a[347] & a[348]};
assign col_697 = sel ? {t_col_327, a[860] & a[859]} : {t_col_697, a[347] & a[348]};
assign col_698 = sel ? {t_col_326, ~a[860] & a[861]} : {t_col_698, ~a[348] & a[349]};
assign col_699 = sel ? {t_col_325, a[861] & a[860]} : {t_col_699, a[348] & a[349]};
assign col_700 = sel ? {t_col_324, ~a[861] & a[862]} : {t_col_700, ~a[349] & a[350]};
assign col_701 = sel ? {t_col_323, a[862] & a[861]} : {t_col_701, a[349] & a[350]};
assign col_702 = sel ? {t_col_322, ~a[862] & a[863]} : {t_col_702, ~a[350] & a[351]};
assign col_703 = sel ? {t_col_321, a[863] & a[862]} : {t_col_703, a[350] & a[351]};
assign col_704 = sel ? {t_col_320, ~a[863] & a[864]} : {t_col_704, ~a[351] & a[352]};
assign col_705 = sel ? {t_col_319, a[864] & a[863]} : {t_col_705, a[351] & a[352]};
assign col_706 = sel ? {t_col_318, ~a[864] & a[865]} : {t_col_706, ~a[352] & a[353]};
assign col_707 = sel ? {t_col_317, a[865] & a[864]} : {t_col_707, a[352] & a[353]};
assign col_708 = sel ? {t_col_316, ~a[865] & a[866]} : {t_col_708, ~a[353] & a[354]};
assign col_709 = sel ? {t_col_315, a[866] & a[865]} : {t_col_709, a[353] & a[354]};
assign col_710 = sel ? {t_col_314, ~a[866] & a[867]} : {t_col_710, ~a[354] & a[355]};
assign col_711 = sel ? {t_col_313, a[867] & a[866]} : {t_col_711, a[354] & a[355]};
assign col_712 = sel ? {t_col_312, ~a[867] & a[868]} : {t_col_712, ~a[355] & a[356]};
assign col_713 = sel ? {t_col_311, a[868] & a[867]} : {t_col_713, a[355] & a[356]};
assign col_714 = sel ? {t_col_310, ~a[868] & a[869]} : {t_col_714, ~a[356] & a[357]};
assign col_715 = sel ? {t_col_309, a[869] & a[868]} : {t_col_715, a[356] & a[357]};
assign col_716 = sel ? {t_col_308, ~a[869] & a[870]} : {t_col_716, ~a[357] & a[358]};
assign col_717 = sel ? {t_col_307, a[870] & a[869]} : {t_col_717, a[357] & a[358]};
assign col_718 = sel ? {t_col_306, ~a[870] & a[871]} : {t_col_718, ~a[358] & a[359]};
assign col_719 = sel ? {t_col_305, a[871] & a[870]} : {t_col_719, a[358] & a[359]};
assign col_720 = sel ? {t_col_304, ~a[871] & a[872]} : {t_col_720, ~a[359] & a[360]};
assign col_721 = sel ? {t_col_303, a[872] & a[871]} : {t_col_721, a[359] & a[360]};
assign col_722 = sel ? {t_col_302, ~a[872] & a[873]} : {t_col_722, ~a[360] & a[361]};
assign col_723 = sel ? {t_col_301, a[873] & a[872]} : {t_col_723, a[360] & a[361]};
assign col_724 = sel ? {t_col_300, ~a[873] & a[874]} : {t_col_724, ~a[361] & a[362]};
assign col_725 = sel ? {t_col_299, a[874] & a[873]} : {t_col_725, a[361] & a[362]};
assign col_726 = sel ? {t_col_298, ~a[874] & a[875]} : {t_col_726, ~a[362] & a[363]};
assign col_727 = sel ? {t_col_297, a[875] & a[874]} : {t_col_727, a[362] & a[363]};
assign col_728 = sel ? {t_col_296, ~a[875] & a[876]} : {t_col_728, ~a[363] & a[364]};
assign col_729 = sel ? {t_col_295, a[876] & a[875]} : {t_col_729, a[363] & a[364]};
assign col_730 = sel ? {t_col_294, ~a[876] & a[877]} : {t_col_730, ~a[364] & a[365]};
assign col_731 = sel ? {t_col_293, a[877] & a[876]} : {t_col_731, a[364] & a[365]};
assign col_732 = sel ? {t_col_292, ~a[877] & a[878]} : {t_col_732, ~a[365] & a[366]};
assign col_733 = sel ? {t_col_291, a[878] & a[877]} : {t_col_733, a[365] & a[366]};
assign col_734 = sel ? {t_col_290, ~a[878] & a[879]} : {t_col_734, ~a[366] & a[367]};
assign col_735 = sel ? {t_col_289, a[879] & a[878]} : {t_col_735, a[366] & a[367]};
assign col_736 = sel ? {t_col_288, ~a[879] & a[880]} : {t_col_736, ~a[367] & a[368]};
assign col_737 = sel ? {t_col_287, a[880] & a[879]} : {t_col_737, a[367] & a[368]};
assign col_738 = sel ? {t_col_286, ~a[880] & a[881]} : {t_col_738, ~a[368] & a[369]};
assign col_739 = sel ? {t_col_285, a[881] & a[880]} : {t_col_739, a[368] & a[369]};
assign col_740 = sel ? {t_col_284, ~a[881] & a[882]} : {t_col_740, ~a[369] & a[370]};
assign col_741 = sel ? {t_col_283, a[882] & a[881]} : {t_col_741, a[369] & a[370]};
assign col_742 = sel ? {t_col_282, ~a[882] & a[883]} : {t_col_742, ~a[370] & a[371]};
assign col_743 = sel ? {t_col_281, a[883] & a[882]} : {t_col_743, a[370] & a[371]};
assign col_744 = sel ? {t_col_280, ~a[883] & a[884]} : {t_col_744, ~a[371] & a[372]};
assign col_745 = sel ? {t_col_279, a[884] & a[883]} : {t_col_745, a[371] & a[372]};
assign col_746 = sel ? {t_col_278, ~a[884] & a[885]} : {t_col_746, ~a[372] & a[373]};
assign col_747 = sel ? {t_col_277, a[885] & a[884]} : {t_col_747, a[372] & a[373]};
assign col_748 = sel ? {t_col_276, ~a[885] & a[886]} : {t_col_748, ~a[373] & a[374]};
assign col_749 = sel ? {t_col_275, a[886] & a[885]} : {t_col_749, a[373] & a[374]};
assign col_750 = sel ? {t_col_274, ~a[886] & a[887]} : {t_col_750, ~a[374] & a[375]};
assign col_751 = sel ? {t_col_273, a[887] & a[886]} : {t_col_751, a[374] & a[375]};
assign col_752 = sel ? {t_col_272, ~a[887] & a[888]} : {t_col_752, ~a[375] & a[376]};
assign col_753 = sel ? {t_col_271, a[888] & a[887]} : {t_col_753, a[375] & a[376]};
assign col_754 = sel ? {t_col_270, ~a[888] & a[889]} : {t_col_754, ~a[376] & a[377]};
assign col_755 = sel ? {t_col_269, a[889] & a[888]} : {t_col_755, a[376] & a[377]};
assign col_756 = sel ? {t_col_268, ~a[889] & a[890]} : {t_col_756, ~a[377] & a[378]};
assign col_757 = sel ? {t_col_267, a[890] & a[889]} : {t_col_757, a[377] & a[378]};
assign col_758 = sel ? {t_col_266, ~a[890] & a[891]} : {t_col_758, ~a[378] & a[379]};
assign col_759 = sel ? {t_col_265, a[891] & a[890]} : {t_col_759, a[378] & a[379]};
assign col_760 = sel ? {t_col_264, ~a[891] & a[892]} : {t_col_760, ~a[379] & a[380]};
assign col_761 = sel ? {t_col_263, a[892] & a[891]} : {t_col_761, a[379] & a[380]};
assign col_762 = sel ? {t_col_262, ~a[892] & a[893]} : {t_col_762, ~a[380] & a[381]};
assign col_763 = sel ? {t_col_261, a[893] & a[892]} : {t_col_763, a[380] & a[381]};
assign col_764 = sel ? {t_col_260, ~a[893] & a[894]} : {t_col_764, ~a[381] & a[382]};
assign col_765 = sel ? {t_col_259, a[894] & a[893]} : {t_col_765, a[381] & a[382]};
assign col_766 = sel ? {t_col_258, ~a[894] & a[895]} : {t_col_766, ~a[382] & a[383]};
assign col_767 = sel ? {t_col_257, a[895] & a[894]} : {t_col_767, a[382] & a[383]};
assign col_768 = sel ? {t_col_256, ~a[895] & a[896]} : {t_col_768, ~a[383] & a[384]};
assign col_769 = sel ? {t_col_255, a[896] & a[895]} : {t_col_769, a[383] & a[384]};
assign col_770 = sel ? {t_col_254, ~a[896] & a[897]} : {t_col_770, ~a[384] & a[385]};
assign col_771 = sel ? {t_col_253, a[897] & a[896]} : {t_col_771, a[384] & a[385]};
assign col_772 = sel ? {t_col_252, ~a[897] & a[898]} : {t_col_772, ~a[385] & a[386]};
assign col_773 = sel ? {t_col_251, a[898] & a[897]} : {t_col_773, a[385] & a[386]};
assign col_774 = sel ? {t_col_250, ~a[898] & a[899]} : {t_col_774, ~a[386] & a[387]};
assign col_775 = sel ? {t_col_249, a[899] & a[898]} : {t_col_775, a[386] & a[387]};
assign col_776 = sel ? {t_col_248, ~a[899] & a[900]} : {t_col_776, ~a[387] & a[388]};
assign col_777 = sel ? {t_col_247, a[900] & a[899]} : {t_col_777, a[387] & a[388]};
assign col_778 = sel ? {t_col_246, ~a[900] & a[901]} : {t_col_778, ~a[388] & a[389]};
assign col_779 = sel ? {t_col_245, a[901] & a[900]} : {t_col_779, a[388] & a[389]};
assign col_780 = sel ? {t_col_244, ~a[901] & a[902]} : {t_col_780, ~a[389] & a[390]};
assign col_781 = sel ? {t_col_243, a[902] & a[901]} : {t_col_781, a[389] & a[390]};
assign col_782 = sel ? {t_col_242, ~a[902] & a[903]} : {t_col_782, ~a[390] & a[391]};
assign col_783 = sel ? {t_col_241, a[903] & a[902]} : {t_col_783, a[390] & a[391]};
assign col_784 = sel ? {t_col_240, ~a[903] & a[904]} : {t_col_784, ~a[391] & a[392]};
assign col_785 = sel ? {t_col_239, a[904] & a[903]} : {t_col_785, a[391] & a[392]};
assign col_786 = sel ? {t_col_238, ~a[904] & a[905]} : {t_col_786, ~a[392] & a[393]};
assign col_787 = sel ? {t_col_237, a[905] & a[904]} : {t_col_787, a[392] & a[393]};
assign col_788 = sel ? {t_col_236, ~a[905] & a[906]} : {t_col_788, ~a[393] & a[394]};
assign col_789 = sel ? {t_col_235, a[906] & a[905]} : {t_col_789, a[393] & a[394]};
assign col_790 = sel ? {t_col_234, ~a[906] & a[907]} : {t_col_790, ~a[394] & a[395]};
assign col_791 = sel ? {t_col_233, a[907] & a[906]} : {t_col_791, a[394] & a[395]};
assign col_792 = sel ? {t_col_232, ~a[907] & a[908]} : {t_col_792, ~a[395] & a[396]};
assign col_793 = sel ? {t_col_231, a[908] & a[907]} : {t_col_793, a[395] & a[396]};
assign col_794 = sel ? {t_col_230, ~a[908] & a[909]} : {t_col_794, ~a[396] & a[397]};
assign col_795 = sel ? {t_col_229, a[909] & a[908]} : {t_col_795, a[396] & a[397]};
assign col_796 = sel ? {t_col_228, ~a[909] & a[910]} : {t_col_796, ~a[397] & a[398]};
assign col_797 = sel ? {t_col_227, a[910] & a[909]} : {t_col_797, a[397] & a[398]};
assign col_798 = sel ? {t_col_226, ~a[910] & a[911]} : {t_col_798, ~a[398] & a[399]};
assign col_799 = sel ? {t_col_225, a[911] & a[910]} : {t_col_799, a[398] & a[399]};
assign col_800 = sel ? {t_col_224, ~a[911] & a[912]} : {t_col_800, ~a[399] & a[400]};
assign col_801 = sel ? {t_col_223, a[912] & a[911]} : {t_col_801, a[399] & a[400]};
assign col_802 = sel ? {t_col_222, ~a[912] & a[913]} : {t_col_802, ~a[400] & a[401]};
assign col_803 = sel ? {t_col_221, a[913] & a[912]} : {t_col_803, a[400] & a[401]};
assign col_804 = sel ? {t_col_220, ~a[913] & a[914]} : {t_col_804, ~a[401] & a[402]};
assign col_805 = sel ? {t_col_219, a[914] & a[913]} : {t_col_805, a[401] & a[402]};
assign col_806 = sel ? {t_col_218, ~a[914] & a[915]} : {t_col_806, ~a[402] & a[403]};
assign col_807 = sel ? {t_col_217, a[915] & a[914]} : {t_col_807, a[402] & a[403]};
assign col_808 = sel ? {t_col_216, ~a[915] & a[916]} : {t_col_808, ~a[403] & a[404]};
assign col_809 = sel ? {t_col_215, a[916] & a[915]} : {t_col_809, a[403] & a[404]};
assign col_810 = sel ? {t_col_214, ~a[916] & a[917]} : {t_col_810, ~a[404] & a[405]};
assign col_811 = sel ? {t_col_213, a[917] & a[916]} : {t_col_811, a[404] & a[405]};
assign col_812 = sel ? {t_col_212, ~a[917] & a[918]} : {t_col_812, ~a[405] & a[406]};
assign col_813 = sel ? {t_col_211, a[918] & a[917]} : {t_col_813, a[405] & a[406]};
assign col_814 = sel ? {t_col_210, ~a[918] & a[919]} : {t_col_814, ~a[406] & a[407]};
assign col_815 = sel ? {t_col_209, a[919] & a[918]} : {t_col_815, a[406] & a[407]};
assign col_816 = sel ? {t_col_208, ~a[919] & a[920]} : {t_col_816, ~a[407] & a[408]};
assign col_817 = sel ? {t_col_207, a[920] & a[919]} : {t_col_817, a[407] & a[408]};
assign col_818 = sel ? {t_col_206, ~a[920] & a[921]} : {t_col_818, ~a[408] & a[409]};
assign col_819 = sel ? {t_col_205, a[921] & a[920]} : {t_col_819, a[408] & a[409]};
assign col_820 = sel ? {t_col_204, ~a[921] & a[922]} : {t_col_820, ~a[409] & a[410]};
assign col_821 = sel ? {t_col_203, a[922] & a[921]} : {t_col_821, a[409] & a[410]};
assign col_822 = sel ? {t_col_202, ~a[922] & a[923]} : {t_col_822, ~a[410] & a[411]};
assign col_823 = sel ? {t_col_201, a[923] & a[922]} : {t_col_823, a[410] & a[411]};
assign col_824 = sel ? {t_col_200, ~a[923] & a[924]} : {t_col_824, ~a[411] & a[412]};
assign col_825 = sel ? {t_col_199, a[924] & a[923]} : {t_col_825, a[411] & a[412]};
assign col_826 = sel ? {t_col_198, ~a[924] & a[925]} : {t_col_826, ~a[412] & a[413]};
assign col_827 = sel ? {t_col_197, a[925] & a[924]} : {t_col_827, a[412] & a[413]};
assign col_828 = sel ? {t_col_196, ~a[925] & a[926]} : {t_col_828, ~a[413] & a[414]};
assign col_829 = sel ? {t_col_195, a[926] & a[925]} : {t_col_829, a[413] & a[414]};
assign col_830 = sel ? {t_col_194, ~a[926] & a[927]} : {t_col_830, ~a[414] & a[415]};
assign col_831 = sel ? {t_col_193, a[927] & a[926]} : {t_col_831, a[414] & a[415]};
assign col_832 = sel ? {t_col_192, ~a[927] & a[928]} : {t_col_832, ~a[415] & a[416]};
assign col_833 = sel ? {t_col_191, a[928] & a[927]} : {t_col_833, a[415] & a[416]};
assign col_834 = sel ? {t_col_190, ~a[928] & a[929]} : {t_col_834, ~a[416] & a[417]};
assign col_835 = sel ? {t_col_189, a[929] & a[928]} : {t_col_835, a[416] & a[417]};
assign col_836 = sel ? {t_col_188, ~a[929] & a[930]} : {t_col_836, ~a[417] & a[418]};
assign col_837 = sel ? {t_col_187, a[930] & a[929]} : {t_col_837, a[417] & a[418]};
assign col_838 = sel ? {t_col_186, ~a[930] & a[931]} : {t_col_838, ~a[418] & a[419]};
assign col_839 = sel ? {t_col_185, a[931] & a[930]} : {t_col_839, a[418] & a[419]};
assign col_840 = sel ? {t_col_184, ~a[931] & a[932]} : {t_col_840, ~a[419] & a[420]};
assign col_841 = sel ? {t_col_183, a[932] & a[931]} : {t_col_841, a[419] & a[420]};
assign col_842 = sel ? {t_col_182, ~a[932] & a[933]} : {t_col_842, ~a[420] & a[421]};
assign col_843 = sel ? {t_col_181, a[933] & a[932]} : {t_col_843, a[420] & a[421]};
assign col_844 = sel ? {t_col_180, ~a[933] & a[934]} : {t_col_844, ~a[421] & a[422]};
assign col_845 = sel ? {t_col_179, a[934] & a[933]} : {t_col_845, a[421] & a[422]};
assign col_846 = sel ? {t_col_178, ~a[934] & a[935]} : {t_col_846, ~a[422] & a[423]};
assign col_847 = sel ? {t_col_177, a[935] & a[934]} : {t_col_847, a[422] & a[423]};
assign col_848 = sel ? {t_col_176, ~a[935] & a[936]} : {t_col_848, ~a[423] & a[424]};
assign col_849 = sel ? {t_col_175, a[936] & a[935]} : {t_col_849, a[423] & a[424]};
assign col_850 = sel ? {t_col_174, ~a[936] & a[937]} : {t_col_850, ~a[424] & a[425]};
assign col_851 = sel ? {t_col_173, a[937] & a[936]} : {t_col_851, a[424] & a[425]};
assign col_852 = sel ? {t_col_172, ~a[937] & a[938]} : {t_col_852, ~a[425] & a[426]};
assign col_853 = sel ? {t_col_171, a[938] & a[937]} : {t_col_853, a[425] & a[426]};
assign col_854 = sel ? {t_col_170, ~a[938] & a[939]} : {t_col_854, ~a[426] & a[427]};
assign col_855 = sel ? {t_col_169, a[939] & a[938]} : {t_col_855, a[426] & a[427]};
assign col_856 = sel ? {t_col_168, ~a[939] & a[940]} : {t_col_856, ~a[427] & a[428]};
assign col_857 = sel ? {t_col_167, a[940] & a[939]} : {t_col_857, a[427] & a[428]};
assign col_858 = sel ? {t_col_166, ~a[940] & a[941]} : {t_col_858, ~a[428] & a[429]};
assign col_859 = sel ? {t_col_165, a[941] & a[940]} : {t_col_859, a[428] & a[429]};
assign col_860 = sel ? {t_col_164, ~a[941] & a[942]} : {t_col_860, ~a[429] & a[430]};
assign col_861 = sel ? {t_col_163, a[942] & a[941]} : {t_col_861, a[429] & a[430]};
assign col_862 = sel ? {t_col_162, ~a[942] & a[943]} : {t_col_862, ~a[430] & a[431]};
assign col_863 = sel ? {t_col_161, a[943] & a[942]} : {t_col_863, a[430] & a[431]};
assign col_864 = sel ? {t_col_160, ~a[943] & a[944]} : {t_col_864, ~a[431] & a[432]};
assign col_865 = sel ? {t_col_159, a[944] & a[943]} : {t_col_865, a[431] & a[432]};
assign col_866 = sel ? {t_col_158, ~a[944] & a[945]} : {t_col_866, ~a[432] & a[433]};
assign col_867 = sel ? {t_col_157, a[945] & a[944]} : {t_col_867, a[432] & a[433]};
assign col_868 = sel ? {t_col_156, ~a[945] & a[946]} : {t_col_868, ~a[433] & a[434]};
assign col_869 = sel ? {t_col_155, a[946] & a[945]} : {t_col_869, a[433] & a[434]};
assign col_870 = sel ? {t_col_154, ~a[946] & a[947]} : {t_col_870, ~a[434] & a[435]};
assign col_871 = sel ? {t_col_153, a[947] & a[946]} : {t_col_871, a[434] & a[435]};
assign col_872 = sel ? {t_col_152, ~a[947] & a[948]} : {t_col_872, ~a[435] & a[436]};
assign col_873 = sel ? {t_col_151, a[948] & a[947]} : {t_col_873, a[435] & a[436]};
assign col_874 = sel ? {t_col_150, ~a[948] & a[949]} : {t_col_874, ~a[436] & a[437]};
assign col_875 = sel ? {t_col_149, a[949] & a[948]} : {t_col_875, a[436] & a[437]};
assign col_876 = sel ? {t_col_148, ~a[949] & a[950]} : {t_col_876, ~a[437] & a[438]};
assign col_877 = sel ? {t_col_147, a[950] & a[949]} : {t_col_877, a[437] & a[438]};
assign col_878 = sel ? {t_col_146, ~a[950] & a[951]} : {t_col_878, ~a[438] & a[439]};
assign col_879 = sel ? {t_col_145, a[951] & a[950]} : {t_col_879, a[438] & a[439]};
assign col_880 = sel ? {t_col_144, ~a[951] & a[952]} : {t_col_880, ~a[439] & a[440]};
assign col_881 = sel ? {t_col_143, a[952] & a[951]} : {t_col_881, a[439] & a[440]};
assign col_882 = sel ? {t_col_142, ~a[952] & a[953]} : {t_col_882, ~a[440] & a[441]};
assign col_883 = sel ? {t_col_141, a[953] & a[952]} : {t_col_883, a[440] & a[441]};
assign col_884 = sel ? {t_col_140, ~a[953] & a[954]} : {t_col_884, ~a[441] & a[442]};
assign col_885 = sel ? {t_col_139, a[954] & a[953]} : {t_col_885, a[441] & a[442]};
assign col_886 = sel ? {t_col_138, ~a[954] & a[955]} : {t_col_886, ~a[442] & a[443]};
assign col_887 = sel ? {t_col_137, a[955] & a[954]} : {t_col_887, a[442] & a[443]};
assign col_888 = sel ? {t_col_136, ~a[955] & a[956]} : {t_col_888, ~a[443] & a[444]};
assign col_889 = sel ? {t_col_135, a[956] & a[955]} : {t_col_889, a[443] & a[444]};
assign col_890 = sel ? {t_col_134, ~a[956] & a[957]} : {t_col_890, ~a[444] & a[445]};
assign col_891 = sel ? {t_col_133, a[957] & a[956]} : {t_col_891, a[444] & a[445]};
assign col_892 = sel ? {t_col_132, ~a[957] & a[958]} : {t_col_892, ~a[445] & a[446]};
assign col_893 = sel ? {t_col_131, a[958] & a[957]} : {t_col_893, a[445] & a[446]};
assign col_894 = sel ? {t_col_130, ~a[958] & a[959]} : {t_col_894, ~a[446] & a[447]};
assign col_895 = sel ? {t_col_129, a[959] & a[958]} : {t_col_895, a[446] & a[447]};
assign col_896 = sel ? {t_col_128, ~a[959] & a[960]} : {t_col_896, ~a[447] & a[448]};
assign col_897 = sel ? {t_col_127, a[960] & a[959]} : {t_col_897, a[447] & a[448]};
assign col_898 = sel ? {t_col_126, ~a[960] & a[961]} : {t_col_898, ~a[448] & a[449]};
assign col_899 = sel ? {t_col_125, a[961] & a[960]} : {t_col_899, a[448] & a[449]};
assign col_900 = sel ? {t_col_124, ~a[961] & a[962]} : {t_col_900, ~a[449] & a[450]};
assign col_901 = sel ? {t_col_123, a[962] & a[961]} : {t_col_901, a[449] & a[450]};
assign col_902 = sel ? {t_col_122, ~a[962] & a[963]} : {t_col_902, ~a[450] & a[451]};
assign col_903 = sel ? {t_col_121, a[963] & a[962]} : {t_col_903, a[450] & a[451]};
assign col_904 = sel ? {t_col_120, ~a[963] & a[964]} : {t_col_904, ~a[451] & a[452]};
assign col_905 = sel ? {t_col_119, a[964] & a[963]} : {t_col_905, a[451] & a[452]};
assign col_906 = sel ? {t_col_118, ~a[964] & a[965]} : {t_col_906, ~a[452] & a[453]};
assign col_907 = sel ? {t_col_117, a[965] & a[964]} : {t_col_907, a[452] & a[453]};
assign col_908 = sel ? {t_col_116, ~a[965] & a[966]} : {t_col_908, ~a[453] & a[454]};
assign col_909 = sel ? {t_col_115, a[966] & a[965]} : {t_col_909, a[453] & a[454]};
assign col_910 = sel ? {t_col_114, ~a[966] & a[967]} : {t_col_910, ~a[454] & a[455]};
assign col_911 = sel ? {t_col_113, a[967] & a[966]} : {t_col_911, a[454] & a[455]};
assign col_912 = sel ? {t_col_112, ~a[967] & a[968]} : {t_col_912, ~a[455] & a[456]};
assign col_913 = sel ? {t_col_111, a[968] & a[967]} : {t_col_913, a[455] & a[456]};
assign col_914 = sel ? {t_col_110, ~a[968] & a[969]} : {t_col_914, ~a[456] & a[457]};
assign col_915 = sel ? {t_col_109, a[969] & a[968]} : {t_col_915, a[456] & a[457]};
assign col_916 = sel ? {t_col_108, ~a[969] & a[970]} : {t_col_916, ~a[457] & a[458]};
assign col_917 = sel ? {t_col_107, a[970] & a[969]} : {t_col_917, a[457] & a[458]};
assign col_918 = sel ? {t_col_106, ~a[970] & a[971]} : {t_col_918, ~a[458] & a[459]};
assign col_919 = sel ? {t_col_105, a[971] & a[970]} : {t_col_919, a[458] & a[459]};
assign col_920 = sel ? {t_col_104, ~a[971] & a[972]} : {t_col_920, ~a[459] & a[460]};
assign col_921 = sel ? {t_col_103, a[972] & a[971]} : {t_col_921, a[459] & a[460]};
assign col_922 = sel ? {t_col_102, ~a[972] & a[973]} : {t_col_922, ~a[460] & a[461]};
assign col_923 = sel ? {t_col_101, a[973] & a[972]} : {t_col_923, a[460] & a[461]};
assign col_924 = sel ? {t_col_100, ~a[973] & a[974]} : {t_col_924, ~a[461] & a[462]};
assign col_925 = sel ? {t_col_99, a[974] & a[973]} : {t_col_925, a[461] & a[462]};
assign col_926 = sel ? {t_col_98, ~a[974] & a[975]} : {t_col_926, ~a[462] & a[463]};
assign col_927 = sel ? {t_col_97, a[975] & a[974]} : {t_col_927, a[462] & a[463]};
assign col_928 = sel ? {t_col_96, ~a[975] & a[976]} : {t_col_928, ~a[463] & a[464]};
assign col_929 = sel ? {t_col_95, a[976] & a[975]} : {t_col_929, a[463] & a[464]};
assign col_930 = sel ? {t_col_94, ~a[976] & a[977]} : {t_col_930, ~a[464] & a[465]};
assign col_931 = sel ? {t_col_93, a[977] & a[976]} : {t_col_931, a[464] & a[465]};
assign col_932 = sel ? {t_col_92, ~a[977] & a[978]} : {t_col_932, ~a[465] & a[466]};
assign col_933 = sel ? {t_col_91, a[978] & a[977]} : {t_col_933, a[465] & a[466]};
assign col_934 = sel ? {t_col_90, ~a[978] & a[979]} : {t_col_934, ~a[466] & a[467]};
assign col_935 = sel ? {t_col_89, a[979] & a[978]} : {t_col_935, a[466] & a[467]};
assign col_936 = sel ? {t_col_88, ~a[979] & a[980]} : {t_col_936, ~a[467] & a[468]};
assign col_937 = sel ? {t_col_87, a[980] & a[979]} : {t_col_937, a[467] & a[468]};
assign col_938 = sel ? {t_col_86, ~a[980] & a[981]} : {t_col_938, ~a[468] & a[469]};
assign col_939 = sel ? {t_col_85, a[981] & a[980]} : {t_col_939, a[468] & a[469]};
assign col_940 = sel ? {t_col_84, ~a[981] & a[982]} : {t_col_940, ~a[469] & a[470]};
assign col_941 = sel ? {t_col_83, a[982] & a[981]} : {t_col_941, a[469] & a[470]};
assign col_942 = sel ? {t_col_82, ~a[982] & a[983]} : {t_col_942, ~a[470] & a[471]};
assign col_943 = sel ? {t_col_81, a[983] & a[982]} : {t_col_943, a[470] & a[471]};
assign col_944 = sel ? {t_col_80, ~a[983] & a[984]} : {t_col_944, ~a[471] & a[472]};
assign col_945 = sel ? {t_col_79, a[984] & a[983]} : {t_col_945, a[471] & a[472]};
assign col_946 = sel ? {t_col_78, ~a[984] & a[985]} : {t_col_946, ~a[472] & a[473]};
assign col_947 = sel ? {t_col_77, a[985] & a[984]} : {t_col_947, a[472] & a[473]};
assign col_948 = sel ? {t_col_76, ~a[985] & a[986]} : {t_col_948, ~a[473] & a[474]};
assign col_949 = sel ? {t_col_75, a[986] & a[985]} : {t_col_949, a[473] & a[474]};
assign col_950 = sel ? {t_col_74, ~a[986] & a[987]} : {t_col_950, ~a[474] & a[475]};
assign col_951 = sel ? {t_col_73, a[987] & a[986]} : {t_col_951, a[474] & a[475]};
assign col_952 = sel ? {t_col_72, ~a[987] & a[988]} : {t_col_952, ~a[475] & a[476]};
assign col_953 = sel ? {t_col_71, a[988] & a[987]} : {t_col_953, a[475] & a[476]};
assign col_954 = sel ? {t_col_70, ~a[988] & a[989]} : {t_col_954, ~a[476] & a[477]};
assign col_955 = sel ? {t_col_69, a[989] & a[988]} : {t_col_955, a[476] & a[477]};
assign col_956 = sel ? {t_col_68, ~a[989] & a[990]} : {t_col_956, ~a[477] & a[478]};
assign col_957 = sel ? {t_col_67, a[990] & a[989]} : {t_col_957, a[477] & a[478]};
assign col_958 = sel ? {t_col_66, ~a[990] & a[991]} : {t_col_958, ~a[478] & a[479]};
assign col_959 = sel ? {t_col_65, a[991] & a[990]} : {t_col_959, a[478] & a[479]};
assign col_960 = sel ? {t_col_64, ~a[991] & a[992]} : {t_col_960, ~a[479] & a[480]};
assign col_961 = sel ? {t_col_63, a[992] & a[991]} : {t_col_961, a[479] & a[480]};
assign col_962 = sel ? {t_col_62, ~a[992] & a[993]} : {t_col_962, ~a[480] & a[481]};
assign col_963 = sel ? {t_col_61, a[993] & a[992]} : {t_col_963, a[480] & a[481]};
assign col_964 = sel ? {t_col_60, ~a[993] & a[994]} : {t_col_964, ~a[481] & a[482]};
assign col_965 = sel ? {t_col_59, a[994] & a[993]} : {t_col_965, a[481] & a[482]};
assign col_966 = sel ? {t_col_58, ~a[994] & a[995]} : {t_col_966, ~a[482] & a[483]};
assign col_967 = sel ? {t_col_57, a[995] & a[994]} : {t_col_967, a[482] & a[483]};
assign col_968 = sel ? {t_col_56, ~a[995] & a[996]} : {t_col_968, ~a[483] & a[484]};
assign col_969 = sel ? {t_col_55, a[996] & a[995]} : {t_col_969, a[483] & a[484]};
assign col_970 = sel ? {t_col_54, ~a[996] & a[997]} : {t_col_970, ~a[484] & a[485]};
assign col_971 = sel ? {t_col_53, a[997] & a[996]} : {t_col_971, a[484] & a[485]};
assign col_972 = sel ? {t_col_52, ~a[997] & a[998]} : {t_col_972, ~a[485] & a[486]};
assign col_973 = sel ? {t_col_51, a[998] & a[997]} : {t_col_973, a[485] & a[486]};
assign col_974 = sel ? {t_col_50, ~a[998] & a[999]} : {t_col_974, ~a[486] & a[487]};
assign col_975 = sel ? {t_col_49, a[999] & a[998]} : {t_col_975, a[486] & a[487]};
assign col_976 = sel ? {t_col_48, ~a[999] & a[1000]} : {t_col_976, ~a[487] & a[488]};
assign col_977 = sel ? {t_col_47, a[1000] & a[999]} : {t_col_977, a[487] & a[488]};
assign col_978 = sel ? {t_col_46, ~a[1000] & a[1001]} : {t_col_978, ~a[488] & a[489]};
assign col_979 = sel ? {t_col_45, a[1001] & a[1000]} : {t_col_979, a[488] & a[489]};
assign col_980 = sel ? {t_col_44, ~a[1001] & a[1002]} : {t_col_980, ~a[489] & a[490]};
assign col_981 = sel ? {t_col_43, a[1002] & a[1001]} : {t_col_981, a[489] & a[490]};
assign col_982 = sel ? {t_col_42, ~a[1002] & a[1003]} : {t_col_982, ~a[490] & a[491]};
assign col_983 = sel ? {t_col_41, a[1003] & a[1002]} : {t_col_983, a[490] & a[491]};
assign col_984 = sel ? {t_col_40, ~a[1003] & a[1004]} : {t_col_984, ~a[491] & a[492]};
assign col_985 = sel ? {t_col_39, a[1004] & a[1003]} : {t_col_985, a[491] & a[492]};
assign col_986 = sel ? {t_col_38, ~a[1004] & a[1005]} : {t_col_986, ~a[492] & a[493]};
assign col_987 = sel ? {t_col_37, a[1005] & a[1004]} : {t_col_987, a[492] & a[493]};
assign col_988 = sel ? {t_col_36, ~a[1005] & a[1006]} : {t_col_988, ~a[493] & a[494]};
assign col_989 = sel ? {t_col_35, a[1006] & a[1005]} : {t_col_989, a[493] & a[494]};
assign col_990 = sel ? {t_col_34, ~a[1006] & a[1007]} : {t_col_990, ~a[494] & a[495]};
assign col_991 = sel ? {t_col_33, a[1007] & a[1006]} : {t_col_991, a[494] & a[495]};
assign col_992 = sel ? {t_col_32, ~a[1007] & a[1008]} : {t_col_992, ~a[495] & a[496]};
assign col_993 = sel ? {t_col_31, a[1008] & a[1007]} : {t_col_993, a[495] & a[496]};
assign col_994 = sel ? {t_col_30, ~a[1008] & a[1009]} : {t_col_994, ~a[496] & a[497]};
assign col_995 = sel ? {t_col_29, a[1009] & a[1008]} : {t_col_995, a[496] & a[497]};
assign col_996 = sel ? {t_col_28, ~a[1009] & a[1010]} : {t_col_996, ~a[497] & a[498]};
assign col_997 = sel ? {t_col_27, a[1010] & a[1009]} : {t_col_997, a[497] & a[498]};
assign col_998 = sel ? {t_col_26, ~a[1010] & a[1011]} : {t_col_998, ~a[498] & a[499]};
assign col_999 = sel ? {t_col_25, a[1011] & a[1010]} : {t_col_999, a[498] & a[499]};
assign col_1000 = sel ? {t_col_24, ~a[1011] & a[1012]} : {t_col_1000, ~a[499] & a[500]};
assign col_1001 = sel ? {t_col_23, a[1012] & a[1011]} : {t_col_1001, a[499] & a[500]};
assign col_1002 = sel ? {t_col_22, ~a[1012] & a[1013]} : {t_col_1002, ~a[500] & a[501]};
assign col_1003 = sel ? {t_col_21, a[1013] & a[1012]} : {t_col_1003, a[500] & a[501]};
assign col_1004 = sel ? {t_col_20, ~a[1013] & a[1014]} : {t_col_1004, ~a[501] & a[502]};
assign col_1005 = sel ? {t_col_19, a[1014] & a[1013]} : {t_col_1005, a[501] & a[502]};
assign col_1006 = sel ? {t_col_18, ~a[1014] & a[1015]} : {t_col_1006, ~a[502] & a[503]};
assign col_1007 = sel ? {t_col_17, a[1015] & a[1014]} : {t_col_1007, a[502] & a[503]};
assign col_1008 = sel ? {t_col_16, ~a[1015] & a[1016]} : {t_col_1008, ~a[503] & a[504]};
assign col_1009 = sel ? {t_col_15, a[1016] & a[1015]} : {t_col_1009, a[503] & a[504]};
assign col_1010 = sel ? {t_col_14, ~a[1016] & a[1017]} : {t_col_1010, ~a[504] & a[505]};
assign col_1011 = sel ? {t_col_13, a[1017] & a[1016]} : {t_col_1011, a[504] & a[505]};
assign col_1012 = sel ? {t_col_12, ~a[1017] & a[1018]} : {t_col_1012, ~a[505] & a[506]};
assign col_1013 = sel ? {t_col_11, a[1018] & a[1017]} : {t_col_1013, a[505] & a[506]};
assign col_1014 = sel ? {t_col_10, ~a[1018] & a[1019]} : {t_col_1014, ~a[506] & a[507]};
assign col_1015 = sel ? {t_col_9, a[1019] & a[1018]} : {t_col_1015, a[506] & a[507]};
assign col_1016 = sel ? {t_col_8, ~a[1019] & a[1020]} : {t_col_1016, ~a[507] & a[508]};
assign col_1017 = sel ? {t_col_7, a[1020] & a[1019]} : {t_col_1017, a[507] & a[508]};
assign col_1018 = sel ? {t_col_6, ~a[1020] & a[1021]} : {t_col_1018, ~a[508] & a[509]};
assign col_1019 = sel ? {t_col_5, a[1021] & a[1020]} : {t_col_1019, a[508] & a[509]};
assign col_1020 = sel ? {t_col_4, ~a[1021] & a[1022]} : {t_col_1020, ~a[509] & a[510]};
assign col_1021 = sel ? {t_col_3, a[1022] & a[1021]} : {t_col_1021, a[509] & a[510]};
assign col_1022 = sel ? {t_col_2, ~a[1022] & a[1023]} : {t_col_1022, ~a[510] & a[511]};
assign col_1023 = sel ? {a[1023] & a[1022], 511'b0} : {t_col_1023, a[510] & a[511]};

endmodule

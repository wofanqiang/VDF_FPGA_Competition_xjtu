module xpb_5_285
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hab20270b9e27c248930ec5cfb7452fcb1011c43c6dd3628da23a0ac964a0f4b4b73c4236e1191b56dfc7f950a9991b5dd277f2890d3dd76a16deff0465d0f10fe5b7f2bc1533dec9eda11766f360d49b045e993cf731d762aa20a368f7f0043e34330b8a4c9b441777ddc07c043f821bc77b219e2d85c012c8b71cefcaa7a4c5;
    5'b00010 : xpb = 1024'ha59308c17a614fc85b1813c85e301844aead8548062f24a3c6975c3d163f3c616b3006f4f80bb81f2031b35a6fd425f140d5bd2bf7c8de887d1ebeaa90cf6d6e5720b0c97ad6c04ec8a82c2b4de5e50514b838e161dd81b49eb4b4d735b565ea395e84eae86d8fa168fb9a1910aede0e401c645a0ac022f54afebedb0c6ce31f;
    5'b00011 : xpb = 1024'ha005ea77569add48232161c1051b00be4d4946539e8ae6b9eaf4adb0c7dd840e1f23cbb30efe54e7609b6d64360f3084af3387cee253e5a6e35e7e50bbcde9ccc8896ed6e079a1d3a3af40efa86af56f2511d885cc892c069348c645737ac7963e89fe4b843fdb2b5a1973b61d1e3a00b8bda715e7fa85d7cd4660c64e322179;
    5'b00100 : xpb = 1024'h9a78cc2d32d46ac7eb2aafb9ac05e937ebe5075f36e6a8d00f51ff24797bcbbad317907125f0f1afa105276dfc4a3b181d915271ccdeecc5499e3df6e6cc662b39f22ce4461c83587eb655b402f005d9356b782a3734d65887dcd7b3b140294243b577ac201226b54b374d53298d95f3315ee9d1c534e8ba4f8e02b18ff75fd3;
    5'b00101 : xpb = 1024'h94ebade30f0df847b333fdb252f0d1b18a80c86acf426ae633af50982b1a1367870b552f3ce38e77e16ee177c28545ab8bef1d14b769f3e3afddfd9d11cae289ab5aeaf1abbf64dd59bd6a785d75164345c517cea1e080aa7c70e921ef058aee48e0f10cbbe4723f3c5526f035fcf1e5aa002c8da26f4b9cd1d5a49cd1bc9e2d;
    5'b00110 : xpb = 1024'h8f5e8f98eb4785c77b3d4baaf9dbba2b291c8976679e2cfc580ca20bdcb85b143aff19ed53d62b4021d89b8188c0503efa4ce7b7a1f4fb02161dbd433cc95ee81cc3a8ff1162466234c47f3cb7fa26ad561eb7730c8c2afc7104fa902ccaec9a4e0c6a6d57b6bdc92d73008d426c4dd822a16f497fa9ae7f541d46881381dc87;
    5'b00111 : xpb = 1024'h89d1714ec7811347434699a3a0c6a2a4c7b84a81fff9ef127c69f37f8e56a2c0eef2deab6ac8c8086242558b4efb5ad268aab25a8c8002207c5d7ce967c7db468e2c670c770527e70fcb9401127f3717667857177737d54e65990bfe6a904e465337e3cdf38909531e90da2a4edba9ca9b42b2055ce41161d664e87355471ae1;
    5'b01000 : xpb = 1024'h84445304a3baa0c70b4fe79c47b18b1e66540b8d9855b128a0c744f33ff4ea6da2e6a36981bb64d0a2ac0f9515366565d7087cfd770b093ee29d3c8f92c657a4ff952519dca8096bead2a8c56d04478176d1f6bbe1e37fa05a2d1d6ca855aff258635d2e8f5b54dd0faeb3c75b4b05bd13e3f4c13a1e744458ac8a5e970c593b;
    5'b01001 : xpb = 1024'h7eb734ba7ff42e46d3593594ee9c739804efcc9930b1733ec5249666f193321a56da682798ae0198e315c99edb716ff9456647a06196105d48dcfc35bdc4d40370fde327424aeaf0c5d9bd89c78957eb872b96604c8f29f24ec12edae61b119e5d8ed68f2b2da06700cc8d6467ba61af8c85377d1758d726daf42c49d8d19795;
    5'b01010 : xpb = 1024'h792a16705c2dbbc69b62838d95875c11a38b8da4c90d3554e981e7daa33179c70ace2ce5afa09e61237f83a8a1ac7a8cb3c412434c21177baf1cbbdbe8c35061e266a134a7edcc75a0e0d24e220e685597853604b73ad4444355404923e0734a62ba4fefc6ffebf0f1ea67017429bda205267a38f4933a095d3bce351a96d5ef;
    5'b01011 : xpb = 1024'h739cf82638674946636bd1863c72448b42274eb06168f76b0ddf394e54cfc173bec1f1a3c6933b2963e93db267e785202221dce636ac1e9a155c7b8213c1ccc053cf5f420d90adfa7be7e7127c9378bfa7ded5a921e67e9637e951b761a5d4f667e5c95062d2377ae308409e809919947dc7bcf4d1cd9cebdf8370205c5c1449;
    5'b01100 : xpb = 1024'h6e0fd9dc14a0d6c62b751f7ee35d2d04e0c30fbbf9c4b981323c8ac2066e092072b5b661dd85d7f1a452f7bc2e228fb3907fa789213725b87b9c3b283ec0491ec5381d4f73338f7f56eefbd6d7188929b838754d8c9228e82c7d63259f6b36a26d1142b0fea48304d4261a3b8d087586f668ffb0af07ffce61cb120b9e2152a3;
    5'b01101 : xpb = 1024'h6882bb91f0da6445f37e6d778a48157e7f5ed0c792207b975699dc35b80c50cd26a97b1ff47874b9e4bcb1c5f45d9a46fedd722c0bc22cd6e1dbface69bec57d36a0db5cd8d6710431f6109b319d9993c89214f1f73dd33a21117493dd30984e723cbc119a76ce8ec543f3d89977d1796f0a426c8c4262b0e412b3f6dfe690fd;
    5'b01110 : xpb = 1024'h62f59d47cd13f1c5bb87bb703132fdf81dfa91d32a7c3dad7af72da969aa9879da9d3fde0b6b118225266bcfba98a4da6d3b3ccef64d33f5481bba7494bd41dba809996a3e7952890cfd255f8c22a9fdd8ebb49661e97d8c15a586021af5f9fa7768357236491a18b661cd75a5e72d6be7ab8528697cc593665a55e221abcf57;
    5'b01111 : xpb = 1024'h5d687efda94d7f4583910968d81de671bc9652dec2d7ffc39f547f1d1b48e0268e91049c225dae4a659025d980d3af6ddb990771e0d83b13ae5b7a1abfbbbe3a19725777a41c340de8043a23e6a7ba67e945543acc9527de0a39977058bb5ba67c93aed2d21b65a2a77fa712b256895e604cc7e446b72875e8a1f7cd63710db1;
    5'b10000 : xpb = 1024'h57db60b385870cc54b9a57617f08ceeb5b3213ea5b33c1d9c3b1d090cce727d34284c95a39504b12a5f9dfe3470eba0149f6d214cb634232149b39c0eaba3a988adb158509bf1592c30b4ee8412ccad1f99ef3df3740d22ffecda8de9680bd5281bf28336dedb12c989d80afbec5e550d8ee0aa023f18b586ae999b8a5364c0b;
    5'b10001 : xpb = 1024'h524e426961c09a4513a3a55a25f3b764f9cdd4f5f38f83efe80f22047e856f7ff6788e185042e7dae66399ed0d49c494b8549cb7b5ee49507adaf96715b8b6f6fc43d3926f61f7179e1263ac9bb1db3c09f89383a1ec7c81f361ba4cd4461efe86eaa19409bffcb689bb5a4ccb354143518f4d5c012bee3aed313ba3e6fb8a65;
    5'b10010 : xpb = 1024'h4cc1241f3dfa27c4dbacf352ccde9fde986996018beb46060c6c73783023b72caa6c52d6673584a326cd53f6d384cf2826b2675aa079506ee11ab90d40b733556dac919fd504d89c79197870f636eba61a5233280c9826d3e7f5cbbb120b80aa8c161af4a59248407ad933e9d7a49d35ca309017de66511d6f78dd8f28c0c8bf;
    5'b10011 : xpb = 1024'h473405d51a33b544a3b6414b73c988583705570d2447081c30c9c4ebe1c1fed95e6017947e28216b67370e0099bfd9bb951031fd8b04578d475a78b36bb5afb3df154fad3aa7ba2154208d3550bbfc102aabd2cc7743d125dc89dd294fd0e25691419455416493ca6bf70d86e413f92842d1d2d3bba0b3fff1c07f7a6a860719;
    5'b10100 : xpb = 1024'h41a6e78af66d42c46bbf8f441ab470d1d5a11818bca2ca325527165f936046861253dc52951abe33a7a0c80a5ffae44f036dfca0758f5eabad9a385996b42c12507e0dbaa04a9ba62f27a1f9ab410c7a3b057270e1ef7b77d11dee978d964402966d0db5dd36df545d14e723f083551abb73158f98db16e274082165ac4b4573;
    5'b10101 : xpb = 1024'h3c19c940d2a6d04433c8dd3cc19f594b743cd92454fe8c48798467d344fe8e32c647a110ac0d5afbe80a82142635eee271cbc743601a65ca13d9f7ffc1b2a870c1e6cbc805ed7d2b0a2eb6be05c61ce44b5f12154c9b25c9c5b20005cb5ba5ae9b98871679092ade4e32c0c0fcf2b10d3414584b761579c4f64fc350ee1083cd;
    5'b10110 : xpb = 1024'h368caaf6aee05dc3fbd22b35688a41c512d89a2fed5a4e5e9de1b946f69cd5df7a3b65cec2fff7c428743c1dec70f975e02991e64aa56ce87a19b7a5ecb124cf334f89d56b905eafe535cb82604b2d4e5bb8b1b9b746d01bba4611740921075aa0c4007714db76683f509a5e09620cffacb59b07534fdca77897653c2fd5c227;
    5'b10111 : xpb = 1024'h30ff8cac8b19eb43c3db792e0f752a3eb1745b3b85b61074c23f0abaa83b1d8c2e2f2a8cd9f2948c68ddf627b2ac04094e875c8935307406e059774c17afa12da4b847e2d1334034c03ce046bad03db86c12515e21f27a6daeda22e246e66906a5ef79d7b0adc1f2306e73fb15d168f22556ddc3308a3f89fadf0727719b0081;
    5'b11000 : xpb = 1024'h2b726e62675378c38be4c726b66012b850101c471e11d28ae69c5c2e59d96538e222ef4af0e53154a947b03178e70e9cbce5272c1fbb7b25469936f242ae1d8c162105f036d621b99b43f50b15554e227c6bf1028c9e24bfa36e345084abcab2ab1af3384c800d7c218c4d982240c4e49df8207f0dc4a26c7d26a912b3603edb;
    5'b11001 : xpb = 1024'h25e55018438d064353ee151f5d4afb31eeabdd52b66d94a10af9ada20b77ace59616b40907d7ce1ce9b16a3b3f2219302b42f1cf0a468243acd8f6986dac99ea8789c3fd9c79033e764b09cf6fda5e8c8cc590a6f749cf11980245bec2712c5eb0466c98e852590612aa27352eb020d71699633aeaff054eff6e4afdf5257d35;
    5'b11010 : xpb = 1024'h205831ce1fc693c31bf763180435e3ab8d479e5e4ec956b72f56ff15bd15f4924a0a78c71eca6ae52a1b2445055d23c399a0bc71f4d189621318b63e98ab1648f8f2820b021be4c351521e93ca5f6ef69d1f304b61f579638c96572d00368e0ab571e5f98424a49003c800d23b1f7cc98f3aa5f6c839683181b5ece936eabb8f;
    5'b11011 : xpb = 1024'h1acb1383fc002142e400b110ab20cc252be35f69e72518cd53b450896eb43c3efdfe3d8535bd07ad6a84de4ecb982e5707fe8714df5c9080795875e4c3a992a76a5b401867bec6482c59335824e47f60ad78cfefcca123b5812a689b3dfbefb6ba9d5f5a1ff6f019f4e5da6f478ed8bc07dbe8b2a573cb1403fd8ed478aff9e9;
    5'b11100 : xpb = 1024'h153df539d839aec2ac09ff09520bb49eca7f20757f80dae37811a1fd205283ebb1f202434cafa475aaee985891d338ea765c51b7c9e7979edf98358aeea80f05dbc3fe25cd61a7cd0760481c7f698fcabdd26f94374cce0775be7a097bc15162bfc8d8babbc93ba3e603b40c53fe34ae807d2b6e82ae2df6864530bfba753843;
    5'b11101 : xpb = 1024'hfb0d6efb4733c4274134d01f8f69d18691ae18117dc9cf99c6ef370d1f0cb9865e5c70163a2413deb585262580e437de4ba1c5ab4729ebd45d7f53119a68b644d2cbc3333048951e2675ce0d9eea034ce2c0f38a1f878596a528b77b986b30ec4f4521b579b872dd7218da9606d90a0f91e6e2a5fe890d9088cd2aafc3a769d;
    5'b11110 : xpb = 1024'ha23b8a590acc9c23c1c9afa9fe1859207b6a28cb0385f0fc0cc44e4838f134519d98bbf7a94de062bc20c6c1e494e115317e6fd9efda5dbac17b4d744a507c2be957a4098a76ad6bd6e71a53473b09ede85aedd0ca422ab5ee69ce5f74c14baca1fcb7bf36dd2b7c83f67466cdcec9371bfb0e63d22f3bb8ad474963dffb4f7;
    5'b11111 : xpb = 1024'h4969a5b6ce657420425e8f346cc6e0ba652639848942125e5299658352d5af1cdcd507d91877ace6c2bc675e48458a4c175b1a08988acfa1257747d6fa384212ffe384dfe4a4c5b987586698ef8c108eedf4e81774fccfd537aae5435117666cf4b44dc8f401e41b95d40e3794c4885ea60f3a21a5d569e0d1c16817fc4f351;
    endcase
end

endmodule

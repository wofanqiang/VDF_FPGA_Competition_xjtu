module xpb_5_100
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h79ba968c4955054dbbf38b86b80267766e0862bf8ebbdecdee44b6050aeba77b8ae57421ef64d505974897b7107345cad73d2d690e18dc1438126a973b89ea7821efb64fd743e1a2d418452175c3f80fa7ed40cc21f78a045ed532a7d07b1b3398649c0e90ff0436bef33017772fc88225691e4959421f40d79d5b2b39038d7c;
    5'b00010 : xpb = 1024'h42c7e7c2d0bbd5d2ace19f365faa879b6a9ac24e48001d245eacb2b462d4a1ef12826acb14a32b7c8f32f0273d887acb4a6032ebf97ee7dcbf8595d03c41603ecf9037f0fef6c600959687a052ac2bee5bd587ffb768e6f8081dd354e6cb93d501c1a5f371350fdff726794ff68f6adafbf85db06238e15168cb3b51e924b48d;
    5'b00011 : xpb = 1024'hbd538f95822a6579dcfb2e60752a7c0672d21dd01445b7acf14af63babd9c629a1f617439e181f3871d48976a9dafcbbd83386ee4e4f3a546f8c1093cf8d6057d30b99226a9aa5e5714ca1f2f945fcd0fbdcf334cda43ebb1667401fd1c0c766b1eafd8516b1b892f59c28875ef0d33d2879d176b2fa361f9f91b789945db9e;
    5'b00100 : xpb = 1024'h858fcf85a177aba559c33e6cbf550f36d535849c90003a48bd596568c5a943de2504d596294656f91e65e04e7b10f59694c065d7f2fdcfb97f0b2ba07882c07d9f206fe1fded8c012b2d0f40a55857dcb7ab0fff6ed1cdf0103ba6a9cd9727aa03834be6e26a1fbfee4cf29fed1ed5b5f7f0bb60c471c2a2d19676a3d249691a;
    5'b00101 : xpb = 1024'h4e9d20bc28de7c2a4ab1521c66fd2f5bd1c7e42b4944789f2dc162181d923e51aca1cc3f4e84ad70165038bea8262a9707e36b5ade63db82067e56d9793a36444cc0f18325a0705eecab51bf82408bbb6b93573304432ae3b9844756e3e7a04b6ce055cbc2a02b6926803bd86c7e780ece7ffac7cd6884b362c456ca826a902b;
    5'b00110 : xpb = 1024'h17aa71f2b0454caf3b9f65cc0ea54f80ce5a43ba0288b6f59e295ec7757b38c5343ec2e873c303e70e3a912ed53b5f977b0670ddc9c9e74a8df1821279f1ac0afa6173244d5354bcae29943e5f28bf9a1f7b9e6699b487d762cce803fa3818ecd63d5fb0a2d637125eb38510ebde1a67a50f3a2ed65f46c3f3f236f1328bb73c;
    5'b00111 : xpb = 1024'h9165087ef99a51fcf792f152c6a7b6f73c62a679914495c38c6e14cc8066e040bf24370a6327d8eca58328e5e5aea56252439e46d7e2c35ec603eca9b57b96831c5129742497365f8241d95fd4ecb7a9c768df32bbac11dbc1a21aabcab334206ea1fbbf33d53b491da6b528630de2e9ca7858782fa16604cb8f921c6b8f44b8;
    5'b01000 : xpb = 1024'h5a7259b581012281e88105026e4fd71c38f506084a88d419fcd6117bd84fdab446c12db388662f639d6d815612c3da62c566a3c9c348cf274d7717e2b6330c49c9f1ab154c4a1abd43c01bdeb1d4eb887b512666511d6ecf6aeabb58e103acc1d7ff05a4140b46f255d9fe60e26d8542a10797df389828155cbd72431bb06bc9;
    5'b01001 : xpb = 1024'h237faaec0867f306d96f18b215f7f7413587659703cd12706d3e0e2b3038d527ce5e245cada485da9557d9c63fd90f633889a94caeaedaefd4ea431bb6ea821077922cb673fcff1b053e5e5d8ebd1f672f396d99e68ecbc314335c05f7542563415c0f88f441529b8e0d479961cd279b7796d746418eea25edeb5269cbd192da;
    5'b01010 : xpb = 1024'h9d3a417851bcf8549562a438cdfa5eb7a38fc8569288f13e5b82c4303b247ca35943987e9d095ae02ca0717d504c552e0fc6d6b5bcc7b7040cfcadb2f2746c889981e3064b40e0bdd956a37f04811776d726ae66088655c773088eadc7cf4096d9c0ab97854056d24d0077b0d8fcf01d9cfff58f9ad10966c588ad9504d52056;
    5'b01011 : xpb = 1024'h664792aed923c8d98650b7e875a27edca02227e54bcd2f94cbeac0df930d7716e0e08f27c247b157248ac9ed7d618a2e82e9dc38a82dc2cc946fd8ebf32be24f472264a772f3c51b9ad4e5fde1694b558b0ef5999df7b2bb1c512f5ade1fb938431db57c6576627b8533c0e9585c9276738f34f6a3c7cb7756b68dbbb4f64767;
    5'b01100 : xpb = 1024'h2f54e3e5608a995e773ecb981d4a9f019cb4877405116deb3c52bd8eeaf6718a687d85d0e78607ce1c75225daa76bf2ef60ce1bb9393ce951be30424f3e35815f4c2e6489aa6a9795c53287cbe517f343ef73ccd33690faec599d007f47031d9ac7abf6145ac6e24bd670a21d7bc34cf4a1e745dacbe8d87e7e46de265176e78;
    5'b01101 : xpb = 1024'ha90f7a71a9df9eac3332571ed54d06780abcea3393cd4cb92a977393f5e21905f362f9f2d6eadcd3b3bdba14baea04f9cd4a0f24a1acaaa953f56ebc2f6d428e16b29c9871ea8b1c306b6d9e34157743e6e47d99556099b3246f02afc4eb4d0d44df5b6fd6ab725b7c5a3a394eebfd516f8792a70600acc8bf81c90d9e1afbf4;
    5'b01110 : xpb = 1024'h721ccba831466f3124206ace7cf5269d074f49c24d118b0f9aff70434dcb13797afff09bfc29334aaba81284e7ff39fa406d14a78d12b671db6899f53024b854c4531e39999d6f79f1e9b01d10fdab229accc4ccead1f6a6cdb7a35cdb3bc5aeae3c6554b6e17e04b48d8371ce4b9faa4616d20e0ef76ed950afa9344e3c2305;
    5'b01111 : xpb = 1024'h3b2a1cdeb8ad3fb6150e7e7e249d46c203e1a9510655c9660b676cf2a5b40ded029ce745216789c1a3926af515146efab3901a2a7878c23a62dbc52e30dc2e1b71f39fdac15053d7b367f29bede5df014eb50c008043539a77004409f18c3e5017996f39971789adecc0ccaa4dab42031ca6117517ee30e9e1dd895afe5d4a16;
    5'b10000 : xpb = 1024'h4376e154014103b05fc922dcc4566e7007408dfbf9a07bc7bcf69a1fd9d08608a39ddee46a5e0389b7cc3654229a3fb26b31fad63dece02ea4ef0673193a3e21f94217be903383574e6351acace12e0029d533415b4b08e2048e4b707dcb6f180f6791e774d955724f415e2cd0ae45bf33550dc20e4f2fa730b6981ae7e7127;
    5'b10001 : xpb = 1024'h7df204a189691588c1f01db48447ce5d6e7c6b9f4e55e68a6a141fa70888afdc151f5210360ab53e32c55b1c529ce9c5fdf04d1671f7aa1722615afe6d1d8e5a4183d7cbc04719d848fe7a3c40920aefaa8a940037ac3a927f1e175ed857d225195b152d084c998de3e745fa443aacde189e6f257a27123b4aa8c4ace781fea3;
    5'b10010 : xpb = 1024'h46ff55d810cfe60db2de31642befee826b0ecb2e079a24e0da7c1c566071aa4f9cbc48b95b490bb52aafb38c7fb21ec6711352995d5db5dfa9d486376dd50420ef24596ce7f9fe360a7cbcbb1d7a3ece5e72db33cd1d97862866b80beea84ac682b81f11e882a5371c1a8f32c39a4f36ef2dae8c831dd44bdbd6a4d397a325b4;
    5'b10011 : xpb = 1024'h100ca70e9836b692a3cc4513d3980ea767a12abcc0de63374ae41905b85aa4c324593f628087622c229a0bfcacc753c6e436581c48c3c1a83147b1706e8c79e79cc4db0e0face293cbfaff39fa6272ad125b2267628ef479d1af58b904f8c367ec1528f6c8b8b0e0544dd86b42f9f18fc5bcedf38c14965c6d0484fa47c44cc5;
    5'b10100 : xpb = 1024'h89c73d9ae18bbbe05fbfd09a8b9a761dd5a98d7c4f9a42053928cf0ac3464c3eaf3eb3846fec3731b9e2a3b3bd3a9991bb73858556dc9dbc695a1c07aa16645fbeb4915de6f0c436a013445b70266abcba48633384867e7e30848b60d573de9b8479c50559b7b51713410882ba29ba11eb260c3ce556b59d44a1e02580c7da41;
    5'b10101 : xpb = 1024'h52d48ed168f28c6550ade44a33429642d23bed0b08de805ba990cbba1b2f46b236dbaa2d952a8da8b1ccfc23ea4fce922e968b084242a984f0cd4740aacdda266c5512ff0ea3a894619186da4d0e9e9b6e30aa6719f7db71d9cd2c0debc4573cedd6ceea39edc0c04b7451bb39895c6ac1b54ba3ee4d77add5cfc04c30e90152;
    5'b10110 : xpb = 1024'h1be1e007f0595cea419bf7f9daeab667cece4c99c222beb219f8c86973184125be78a0d6ba68e41fa9b7549417650392a1b9908b2da8b54d78407279ab854fed19f594a036568cf2230fc95929f6d27a2218f19aaf6938658315ccbb0214cfde5733d8cf1a23cc6983a79af3b8e8fec398448b0af74439be66fda072e10a2863;
    5'b10111 : xpb = 1024'h959c769439ae6237fd8f838092ed1dde3cd6af5950de9d80083d7e6e7e03e8a1495e14f8a9cdb92540ffec4b27d8495d78f6bdf43bc19161b052dd10e70f3a653be54af00d9a6e94f7280e7a9fbaca89ca063266d160c269e1eaff62d28feb11ef9874ddab22d0a0429acb0b3018c745bdada954508658ff3e9afb9e1a0db5df;
    5'b11000 : xpb = 1024'h5ea9c7cac11532bcee7d97303a953e0339690ee80a22dbd678a57b1dd5ece314d0fb0ba1cf0c0f9c38ea44bb54ed7e5dec19c37727279d2a37c60849e7c6b02be985cc91354d52f2b8a650f97ca2fe687dee799a66d21f5d8b33a00fe8e063b358f57ec28b58dc497ace1443af78699e943ce8bb597d1b0fcfc8dbc4ca2edcf0;
    5'b11001 : xpb = 1024'h27b71901487c0341df6baadfe23d5e2835fb6e76c3671a2ce90d77cd2dd5dd885898024af44a661330d49d2b8202b35e5f3cc8fa128da8f2bf393382e87e25f297264e325d0037507a249378598b324731d6c0cdfc437c51347c40bcff30dc54c25288a76b8ee7f2b3015d7c2ed80bf76acc28226273dd2060f6bbeb7a500401;
    5'b11010 : xpb = 1024'ha171af8d91d1088f9b5f36669a3fc59ea403d1365222f8fad7522dd238c18503e37d766ce3af3b18c81d34e29275f9293679f66320a68506f74b9e1a2408106ab9160482344418f34e3cd899cf4f2a56d9c4019a1e3b065593517364cfabf7885ab724b5fc8dec2971f48d93a607d4799035466bbbb5fc6138941716b353917d;
    5'b11011 : xpb = 1024'h6a7f00c41937d9148c4d4a1641e7e5c3a09630c50b67375147ba2a8190aa7f776b1a6d1608ed918fc0078d52bf8b2e29a99cfbe60c0c90cf7ebec95324bf863166b686235bf6fd510fbb1b18ac375e358dac48cdb3ac63493c9a1411e5fc7029c4142e9adcc3f7d2aa27d6cc256776d266c485d2c4acbe71c9c1f73d6374b88e;
    5'b11100 : xpb = 1024'h338c51faa09ea9997d3b5dc5e99005e89d289053c4ab75a7b8222730e89379eaf2b763bf2e2be806b7f1e5c2eca0632a1cc00168f7729c980631f48c2576fbf8145707c483a9e1aed1395d97891f921441949001491dc03ce5e2b4befc4ce8cb2d71387fbcfa037be25b2004a4c7192b3d53c539cda380825aefd7641395df9f;
    5'b11101 : xpb = 1024'had46e886e9f3aee7392ee94ca1926d5f0b30f31353675475a666dd35f37f21667d9cd7e11d90bd0c4f3a7d79fd13a8f4f3fd2ed2058b78ac3e445f236100e6703646be145aedc351a551a2b8fee38a23e981d0cd6b154a4144b7e766ccc803fec5d5d48e4df907b2a14e501c1bf6e1ad62bce38326e59fc3328d328f4c996d1b;
    5'b11110 : xpb = 1024'h765439bd715a7f6c2a1cfcfc493a8d8407c352a20cab92cc16ced9e54b681bda0539ce8a42cf13834724d5ea2a28ddf567203454f0f18474c5b78a5c61b85c36e3e73fb582a0a7af66cfe537dbcbbe029d6a18010086a734ee008813e3187ca02f32de732e2f135bd98199549b568406394c22ea2fdc61d3c3bb12b5fcba942c;
    5'b11111 : xpb = 1024'h3f618af3f8c14ff11b0b10abf0e2ada90455b230c5efd1228736d694a351164d8cd6c533680d69fa3f0f2e5a573e12f5da4339d7dc57903d4d2ab595626fd1fd9187c156aa538c0d284e27b6b8b3f1e151525f3495f80428974928c0f968f541988fe8580e651f0511b4e28d1ab6265f0fdb625138d323e454e8f2dcacdbbb3d;
    endcase
end

endmodule

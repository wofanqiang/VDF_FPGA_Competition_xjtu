module xpb_5_850
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h73089ebab524ed1e6960eb25faad4c1d827598adcee0b7a325325b6e8437cf755a91de91c191f5f07e19b2bd05013a68437d4b7993d7a40e2d67d3151dc6abde795a228c8c5d5820ae648e4e7dd6e09afa2f999304b0eaced657763c39586f167567cd154759b6faf238837e18d3418b99532f4d7e54d0d3b508f63b85c2afb6;
    5'b00010 : xpb = 1024'h3563f81fa85ba57407bc5e74e50050e993752e2ac849cececc87fd87556cf1e2b1db3faab8fd6d525cd5263326a4640622e06f0d04fc77d0aa3066cc00bae30b7e65106a6929b2fc4a2f19fa62d1fd05005a398d7cdba88cf7225a7db8863b9abbc80800ddea75685db1201d39d65cede3cc7fb8ac5e447723a2717282a2f901;
    5'b00011 : xpb = 1024'ha86c96da5d809292711d499adfad9d0715eac6d8972a8671f1ba58f5d9a4c1580c6d1e3c7a8f6342daeed8f02ba59e6e665dba8698d41bded79839e11e818ee9f7bf32f6f5870b1cf893a848e0a8dd9ffa89d320818c935bcd79d0b9f1deaab1312fd51625442c634fe9a39b52a99e797d1faf062ab3154ad8ab67ae0865a8b7;
    5'b00100 : xpb = 1024'h6ac7f03f50b74ae80f78bce9ca00a1d326ea5c5590939d9d990ffb0eaad9e3c563b67f5571fadaa4b9aa4c664d48c80c45c0de1a09f8efa15460cd980175c616fcca20d4d25365f8945e33f4c5a3fa0a00b4731af9b75119ee44b4fb710c773577901001bbd4ead0bb62403a73acb9dbc798ff7158bc88ee4744e2e50545f202;
    5'b00101 : xpb = 1024'h2d2349a443ee033dadd43038b453a69f37e9f1d289fcb4c940659d277c0f0632baffe06e696652069865bfdc6eebf1aa252401ad7b1dc363d129614ee469fd4401d50eb2af1fc0d43028bfa0aa9f167406df131571e20ed80f0f993cf03a43b9bdf04aed5265a93e26dadcd994afd53e12124fdc86c5fc91b5de5e1c02263b4d;
    5'b00110 : xpb = 1024'ha02be85ef912f05c17351b5eaf00f2bcba5f8a8058dd6c6c6597f8960046d5a81591bf002af847f7167f729973ed2c1268a14d270ef56771fe9134640230a9227b2f313f3b7d18f4de8d4def2875f70f010eaca87692f9a6e5670f792992b2d03358180299bf603919136057ad8316c9ab657f2a051acd656ae7545787e8eb03;
    5'b00111 : xpb = 1024'h628741c3ec49a8b1b5908ead9953f788cb5f1ffd524683980ced9aaed17bf8156cdb20192263bf58f53ae60f959055b0480470ba801a3b347b59c81ae524e04f803a1f1d184973d07a57d99b0d71137907394ca2eebdb7650631f3baa8c07f5479b852ee30501ea6848bfcf6ce86322bf5decf9533244108d980cf8e84c9344e;
    5'b01000 : xpb = 1024'h24e29b28df80610753ec01fc83a6fc54dc5eb57a4baf9ac3b4433cc7a2b11a82c424813219cf36bad3f65985b7337f4e2767944df13f0ef6f8225bd1c819177c85450cfaf515ceac16226546f26c2fe30d63ec9d66e8752326fcd7fc27ee4bd8c0188dd9c6e0dd13f0049995ef894d8e40582000612db4ac481a4ac581a97d99;
    5'b01001 : xpb = 1024'h97eb39e394a54e25bd4ced227e5448725ed44e281a905266d975983626e8e9f81eb65fc3db612cab52100c42bc34b9b66ae4dfc78516b305258a2ee6e5dfc35afe9f2f87817326ccc486f3957043107e079386306b995ff1fd544e386146baef35805aef0e3a940ee23d1d14085c8f19d9ab4f4ddf82857ffd234101076c2d4f;
    5'b01010 : xpb = 1024'h5a46934887dc067b5ba8607168a74d3e6fd3e3a513f9699280cb3a4ef81e0c6575ffc0dcd2cca40d30cb7fb8ddd7e3544a48035af63b86c7a252c29dc8d3fa8803aa1d655e3f81a860517f41553e2ce80dbe262ae3c41db01e1f3279e07487737be095daa4cb527c4db5b9b3295faa7c24249fb90d8bf9236bbcbc38044c769a;
    5'b01011 : xpb = 1024'h1ca1ecad7b12bed0fa03d3c052fa520a80d379220d6280be2820dc67c9532ed2cd4921f5ca381b6f0f86f32eff7b0cf229ab26ee67605a8a1f1b5654abc831b508b50b433b0bdc83fc1c0aed3a39495213e8c6255beedb6e3eea16bb5fa253f7c240d0c63b5c10e9b92e56524a62c5de6e9df0243b956cc6da56376f012cbfe5;
    5'b01100 : xpb = 1024'h8faa8b683037abef6364bee64da79e28034911cfdc4338614d5337d64d8afe4827db00878bca115f8da0a5ec047c475a6d287267fb37fe984c832969c98edd93820f2dcfc76934a4aa80993bb81029ed0e185fb8609fc63d15418cf798fac30e37a89ddb82b5c7e4ab66d9d06336076a07f11f71b9ea3d9a8f5f2daa86ef6f9b;
    5'b01101 : xpb = 1024'h5205e4cd236e644501c0323537faa2f41448a74cd5ac4f8cf4a8d9ef1ec020b57f2461a0833588c16c5c1962261f70f84c8b95fb6c5cd25ac94bbd20ac8314c0871a1bada4358f80464b24e79d0b46571442ffb2d8ca83fb360c713918288f927e08d8c71946865216df766f843922cc526a6fdce7f3b13dfdf8a8e183cfb8e6;
    5'b01110 : xpb = 1024'h14613e3216a51c9aa01ba584224da7c025483cc9cf1566b89bfe7c07eff54322d66dc2b97aa100234b178cd847c29a962beeb98edd81a61d461450d78f774bed8c25098b8101ea5be215b093820662c11a6d9fad50f541b956d7557a97565c16c46913b2afd744bf8258130ea53c3e2e9ce3c04815fd24e16c92241880b00231;
    5'b01111 : xpb = 1024'h8769dceccbca09b9097c90aa1cfaf3dda7bdd5779df61e5bc130d776742d129830ffa14b3c32f613c9313f954cc3d4fe6f6c050871594a2b737c23ecad3df7cc057f2c180d5f427c907a3ee1ffdd435c149d394055a62c882d2ecbb6d0aecb2d39d0e0c7f730fbba7490968cbe0f7fba3636ef959451f5b5219b1a540672b1e7;
    5'b10000 : xpb = 1024'h49c53651bf00c20ea7d803f9074df8a9b8bd6af4975f35876886798f4562350588490264339e6d75a7ecb30b6e66fe9c4ecf289be27e1dedf044b7a390322ef90a8a19f5ea2b9d582c44ca8de4d85fc61ac7d93acdd0ea464df9aff84fdc97b180311bb38dc1ba27e009332bdf129b1c80b04000c25b69589034958b0352fb32;
    5'b10001 : xpb = 1024'hc208fb6b2377a6446337747f1a0fd75c9bd007190c84cb30fdc1ba816975772df92637d2b09e4d786a82681900a283a2e324c2f53a2f1b06d0d4b5a732666260f9507d3c6f7f833c80f5639c9d37c3020f2793545fba8046ec49439cf0a6435c691569f245278954b81cfcb0015b67ecb29906bf064dcfbfece10c20033447d;
    5'b10010 : xpb = 1024'h7f292e71675c6782af94626dec4e49934c32991f5fa90456350e77169acf26e83a24420eec9bdac804c1d93e950b62a271af97a8e77a95be9a751e6f90ed120488ef2a60535550547673e48847aa5ccb1b2212c84aac92d3451c0a760862d34c3bf923b46bac2f903dba534918e8f80a647cbfb96eb9adcfb3d706fd85f5f433;
    5'b10011 : xpb = 1024'h418487d65a931fd84defd5bcd6a14e5f5d322e9c59121b81dc64192f6c044955916da327e4075229e37d4cb4b6ae8c405112bb3c589f6981173db22673e149318dfa183e3021ab30123e70342ca57935214cb2c2c2d7509165e6eeb787909fd082595ea0023cedfda932efe839ec136caef610249cc321732270823482d63d7e;
    5'b10100 : xpb = 1024'h3dfe13b4dc9d82dec4b490bc0f4532b6e31c419527b32ad83b9bb483d396bc2e8b70440db72c98bc238c02ad851b5de3075decfc9c43d43940645dd56d5805e9305061c0cee060bae08fbe011a0959f277752bd3b020e4f86b1d2f906be6c54c8b9998b98cdac6b14ab8c875aef2ecef96f608fcacc95169109fd6b7fb686c9;
    5'b10101 : xpb = 1024'h76e87ff602eec54c55ac3431bba19f48f0a75cc7215bea50a8ec16b6c1713b384348e2d29d04bf7c405272e7dd52f04673f32a495d9be151c16e18f2749c2c3d0c5f28a8994b5e2c5c6d8a2e8f77763a21a6ec503fb2f91e5d0949354016db6b3e2166a0e027636606e4100573c2705a92c28fdd492165ea4612f3a70579367f;
    5'b10110 : xpb = 1024'h3943d95af6257da1f407a780a5f4a41501a6f2441ac5017c5041b8cf92a65da59a9243eb947036de1f0de65dfef619e453564ddccec0b5143e36aca95790636a116a16867617b907f83815da747292a427d18c4ab7ddb6dc7dd42d76bf44a7ef8481a18c76b821d3725caca494c58bbcdd3be048772ad98db4ac6ede02597fca;
    5'b10111 : xpb = 1024'hac4c7815ab4a6ac05d6892a6a0a1f032841c8af1e9a5b91f7574143e16de2d1af524227d56022cce9d27991b03f7544c96d39956629859226b9e7fbe75570f488ac4391302751128a69ca428f249733f220125ddbc8ea1ab542ba3b2f89d1705f9e96ea1be11d8ce64953022ad98cd48768f0f95f57faa6169b56519881c2f80;
    5'b11000 : xpb = 1024'h6ea7d17a9e812315fbc405f58af4f4fe951c206ee30ed04b1cc9b656e8134f884c6d83964d6da4307be30c91259a7dea7636bce9d3bd2ce4e8671375584b46758fcf26f0df416c0442672fd4d7448fa9282bc5d834b95f6974f687f477cae38a4049a98d54a2973bd00dccc1ce9be8aac108600123891e04d84ee05084fc78cb;
    5'b11001 : xpb = 1024'h31032adf91b7db6b9a1f79447547f9caa61bb5ebdc77e776c41f586fb94871f5a3b6e4af44d91b925a9e8007473da7885599e07d44e200a7652fa72c3b3f7da294da14cebc0dc6dfde31bb80bc3fac132e5665d2ace41d2795c16c35f6f8b00e86a9e478eb3355a93b866960ef9f040d0b81b06c519291a846e85b8781dcc216;
    5'b11010 : xpb = 1024'ha40bc99a46dcc88a0380646a6ff545e828914e99ab589f19e951b3de3d80416afe48c341066b1182d8b832c44c3ee1f099172bf6d8b9a4b592977a41590629810e34375b486b1f008c9649cf3a168cae2885ff65b19507f66c18e27230511f24fc11b18e328d0ca42dbeecdf08724598a4d4dfb9cfe7627bfbf151c3079f71cc;
    5'b11011 : xpb = 1024'h666722ff3a1380dfa1dbd7b95a484ab43990e416a4c1b64590a755f70eb563d855922459fdd688e4b773a63a6de20b8e787a4f8a49de78780f600df83bfa60ae133f2539253779dc2860d57b1f11a9182eb09f6029bfc5b48ce3c6b3af7eeba94271ec79c91dcb119937897e297560faef4e3024fdf0d61f6a8accfa047fbb17;
    5'b11100 : xpb = 1024'h28c27c642d4a393540374b08449b4f804a9079939e2acd7137fcf80fdfea8645acdb8572f5420046962f19b08f85352c57dd731dbb034c3a8c28a1af1eee97db184a13170203d4b7c42b6127040cc58234db3f5aa1ea8372adaeaaf52eacb82d88d227655fae897f04b0261d4a787c5d39c780902bfa49c2d924483101600462;
    5'b11101 : xpb = 1024'h9bcb1b1ee26f2653a998362e3f489b9dcd0612416d0b85145d2f537e642255bb076d6404b6d3f6371448cc6d94866f949b5abe974edaf048b99074c43cb543b991a435a38e612cd8728fef7581e3a61d2f0ad8eda69b6e418406213168052743fe39f47aa7084079f6e8a99b634bbde8d31aafddaa4f1a968e2d3e6c8722b418;
    5'b11110 : xpb = 1024'h5e267483d5a5dea947f3a97d299ba069de05a7be66749c400484f597355778285eb6c51dae3f6d98f3043fe3b62999327abde22abfffc40b3659087b1fa97ae696af23816b2d87b40e5a7b2166dec287353578e81ec62bffa4d10572e732f3c8449a2f663d98fee76261463a844ed94b1d940048d8588e39fcc6b9a38402fd63;
    5'b11111 : xpb = 1024'h2081cde8c8dc96fee64f1ccc13eea535ef053d3b5fddb36babda97b0068c9a95b6002636a5aae4fad1bfb359d7ccc2d05a2105be312497cdb3219c32029db2139bba115f47f9e28faa2506cd4bd9def13b6018e296f0e9bdc59be9b46660c04c8afa6a51d429bd54cdd9e2d9a551f4ad680d50b4066201dd6b6034da80e346ae;
    endcase
end

endmodule

module xpb_5_105
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h86edc2a802820760bf9245b988acdce00e811bf7f340f78f79ed343fb3a10c11473bbdc8d4bc07136f986ca845347f64d663f5ac7bd9c05d49de0ce632747c43f2842f7d206706ae9cc6a35959c25c0053aa6682b69611c4091c96e0fb96de301ecf23cee9b2aae49e82bc59a15c8b7e66aa1b841c9e5f4e616d3035cfce24e;
    5'b00010 : xpb = 1024'h10ddb855005040ec17f248b731159b9c01d0237efe681ef1ef3da687f674218228e777b91a9780e26df30d9508a68fec9acc7eb58f7b380ba93bc19cc64e8f887e5085efa40ce0d5d398d46b2b384b800a754cd056d2c238812392dc1f72dbc603d9e479dd36555c93d0578b342b916fccd543708393cbe9cc2da606b9f9c49c;
    5'b00011 : xpb = 1024'h194c947f8078616223eb6d12c9a0696a02b8353e7d9c2e6ae6dc79cbf1ae32433d5b3395a7e34153a4ec945f8cf9d7e2e832be105738d4117dd9a26b2975d74cbd78c8e776135140bd653ea0c0d471400faff338823c2354c1b55c4a2f2c49a905c6d6b6cbd1800addb88350ce415a27b33fe528c55db1deb244790a16f6a6ea;
    5'b00100 : xpb = 1024'h21bb70aa00a081d82fe4916e622b373803a046fdfcd03de3de7b4d0fece8430451ceef72352f01c4dbe61b2a114d1fd93598fd6b1ef67017527783398c9d1f10fca10bdf4819c1aba731a8d65670970014ea99a0ada58471024725b83ee5b78c07b3c8f3ba6caab927a0af16685722df99aa86e1072797d3985b4c0d73f38938;
    5'b00101 : xpb = 1024'h2a2a4cd480c8a24e3bddb5c9fab60506048858bd7c044d5cd61a2053e82253c56642ab4ec27ac23612dfa1f495a067cf82ff3cc5e6b40c1d27156407efc466d53bc94ed71a20321690fe130bec0cbcc01a254008d90ee58d42d8ef264e9f256f09a0bb30a907d5677188dadc026ceb978015289948f17dc87e721f10d0f06b86;
    5'b00110 : xpb = 1024'h329928ff00f0c2c447d6da259340d2d405706a7cfb385cd5cdb8f397e35c64867ab6672b4fc682a749d928bf19f3afc5d0657c20ae71a822fbb344d652ebae997af191ceec26a2817aca7d4181a8e2801f5fe671047846a9836ab8945e5893520b8dad6d97a30015bb7106a19c82b44f667fca518abb63bd6488f2142ded4dd4;
    5'b00111 : xpb = 1024'h3b0805298118e33a53cffe812bcba0a206587c3c7a6c6c4ec557c6dbde9675478f2a2307dd12431880d2af899e46f7bc1dcbbb7b762f4428d05125a4b612f65dba19d4c6be2d12ec6496e77717450840249a8cd92fe1a7c5c3fc82026e1201350d7a9faa863e2ac40559326736987d074cea6c09cc8549b24a9fc5178aea3022;
    5'b01000 : xpb = 1024'h4376e154014103b05fc922dcc4566e7007408dfbf9a07bc7bcf69a1fd9d08608a39ddee46a5e0389b7cc3654229a3fb26b31fad63dece02ea4ef0673193a3e21f94217be903383574e6351acace12e0029d533415b4b08e2048e4b707dcb6f180f6791e774d955724f415e2cd0ae45bf33550dc20e4f2fa730b6981ae7e71270;
    5'b01001 : xpb = 1024'h4be5bd7e816924266bc247385ce13c3e08289fbb78d48b40b4956d63d50a96c9b8119ac0f7a9c3faeec5bd1ea6ed87a8b8983a3105aa7c34798ce7417c6185e6386a5ab66239f3c2382fbbe2427d53c02f0fd9a986b469fe452014de8d84dcfb1154842463748020992989f26ac40e7719bfaf7a5019159c16cd6b1e44e3f4be;
    5'b01010 : xpb = 1024'h545499a90191449c77bb6b93f56c0a0c0910b17af8089ab9ac3440a7d044a78acc85569d84f5846c25bf43e92b40cf9f05fe798bcd68183a4e2ac80fdf88cdaa77929dae3440642d21fc2617d8197980344a8011b21dcb1a85b1de4c9d3e4ade13417661520faacee311b5b804d9d72f002a513291e2fb90fce43e21a1e0d70c;
    5'b01011 : xpb = 1024'h5cc375d381b9651283b48fef8df6d7da09f8c33a773caa32a3d313ebcb7eb84be0f9127a124144dd5cb8cab3af9417955364b8e69525b44022c8a8de42b0156eb6bae0a60646d4980bc8904d6db59f4039852679dd872c36c643a7baacf7b8c1152e689e40aad57d2cf9e17d9eef9fe6e694f2ead3ace185e2fb1124feddb95a;
    5'b01100 : xpb = 1024'h653251fe01e185888fadb44b2681a5a80ae0d4f9f670b9ab9b71e72fc6b8c90cf56cce569f8d054e93b2517e33e75f8ba0caf8415ce35045f76689aca5d75d32f5e3239dd84d4502f594fa830351c5003ebfcce208f08d5306d57128bcb126a4171b5adb2f46002b76e20d433905689eccff94a31576c77ac911e4285bda9ba8;
    5'b01101 : xpb = 1024'h6da12e288209a5fe9ba6d8a6bf0c73760bc8e6b975a4c9249310ba73c1f2d9ce09e08a332cd8c5bfcaabd848b83aa781ee31379c24a0ec4bcc046a7b08fea4f7350b6695aa53b56ddf6164b898edeac043fa734a3459ee6f47673a96cc6a948719084d181de12ad9c0ca3908d31b3156b36a365b5740ad6faf28b72bb8d77df6;
    5'b01110 : xpb = 1024'h76100a530231c674a79ffd02579741440cb0f878f4d8d89d8aaf8db7bd2cea8f1e54460fba24863101a55f133c8def783b9776f6ec5e8851a0a24b496c25ecbb7433a98d7c5a25d8c92dceee2e8a1080493519b25fc34f8b87f90404dc24026a1af53f550c7c55880ab264ce6d30fa0e99d4d813990a9364953f8a2f15d46044;
    5'b01111 : xpb = 1024'h7e7ee67d8259e6eab399215df0220f120d990a38740ce816824e60fbb866fb5032c801ec477046a2389ee5ddc0e1376e88fdb651b41c245775402c17cf4d347fb35bec854e609643b2fa3923c42636404e6fc01a8b2cb0a7c88acd72ebdd704d1ce23191fb178036549a90940746c2c6803f79cbdad479597b565d3272d14292;
    5'b10000 : xpb = 1024'h86edc2a802820760bf9245b988acdce00e811bf7f340f78f79ed343fb3a10c11473bbdc8d4bc07136f986ca845347f64d663f5ac7bd9c05d49de0ce632747c43f2842f7d206706ae9cc6a35959c25c0053aa6682b69611c4091c96e0fb96de301ecf23cee9b2aae49e82bc59a15c8b7e66aa1b841c9e5f4e616d3035cfce24e0;
    5'b10001 : xpb = 1024'h8f5c9ed282aa27d6cb8b6a152137aaae0f692db772750708718c0783aedb1cd25baf79a56207c784a691f372c987c75b23ca350743975c631e7bedb4959bc40831ac7274f26d771986930d8eef5e81c058e50ceae1ff72e049ae604f0b504c1320bc160bd84dd592e86ae81f3b7254364d14bd3c5e684543478403392ccb072e;
    5'b10010 : xpb = 1024'h97cb7afd02d2484cd7848e70b9c2787c10513f76f1a91681692adac7aa152d9370233581ef5387f5dd8b7a3d4ddb0f51713074620b54f868f319ce82f8c30bcc70d4b56cc473e784705f77c484faa7805e1fb3530d68d3fc8a4029bd1b09b9f622a90848c6e90041325313e4d5881cee337f5ef4a0322b382d9ad63c89c7e97c;
    5'b10011 : xpb = 1024'ha03a572782fa68c2e37db2cc524d464a1139513670dd25fa60c9ae0ba54f3e548496f15e7c9f486714850107d22e5747be96b3bcd312946ec7b7af515bea5390affcf864967a57ef5a2be1fa1a96cd40635a59bb38d23518cad1f32b2ac327d92495fa85b5842aef7c3b3faa6f9de5a619ea00ace1fc112d13b1a93fe6c4cbca;
    5'b10100 : xpb = 1024'ha8a9335203228938ef76d727ead81418122162f5f01135735868814fa0894f15990aad3b09eb08d84b7e87d256819f3e0bfcf3179ad030749c55901fbf119b54ef253b5c6880c85a43f84c2fb032f30068950023643b96350b63bc993a7c95bc2682ecc2a41f559dc6236b7009b3ae5e0054a26523c5f721f9c87c4343c1ae18;
    5'b10101 : xpb = 1024'h6aca26c15c74e6306a83ac73089a94a193718499cda474d22a9b3de8c0b2ceaa35eb9ecd104abae319cf55f776d669f5490a8c3fdafc2ec054318fe7666e67b9fe49a58af63b801b2ab3c2acf3548f79caacf3031eca409668f40c900b610cf9684cd5e1f187be894bb056abf950ec97e5653b15447fe6996fd44217dc29fb;
    5'b10110 : xpb = 1024'h8d9a6514184955c3c63a8080b936862a27b83441901b3edc9c96e81e3fac38fbea9a77b5a5c0b2c1a1356207bca1e6042af49e70798983494f2125e4a8db62bf9268c9d5cfcabeb04f71df8428f7a4f7f05535b2e882b5cd6fabd7a9fc4ceeffb553f12d08cb26cd333dc1c460f19a47e5006f3570e65db7f86a74574d90c49;
    5'b10111 : xpb = 1024'h1148827bc1acb5d2485ccc63a41e3630a36395039835c366c16841c5df34d450d31d6357e7a7cb9d510cdceb001d665690158941cf56343a698ff32cadb4fdf0384ecf952f031c55eec3882dd82ba00f843ff9c359f18c79178c86e8af7e3cd2fd42314fbf27dd1b1d1c07e1e024e25c64baa8ab98d84bd0659d7a48d1d5ee97;
    5'b11000 : xpb = 1024'h19b75ea641d4d6485455f0bf3ca903fea44ba6c31769d2dfb9071509da6ee511e7911f3474f38c0e880663b58470ae4cdd7bc89c9713d0403e2dd3fb10dc45b47777128d01098cc0d88ff2636dc7c5cf897aa02b855aed95581e5056bf37aab5ff2f238cadc307c9670433a77a3aab144b254a63daa231c54bb44d4c2ed2d0e5;
    5'b11001 : xpb = 1024'h22263ad0c1fcf6be604f151ad533d1cca533b882969de258b0a5e84dd5a8f5d2fc04db11023f4c7fbeffea8008c3f6432ae207f75ed16c4612cbb4c974038d78b69f5584d30ffd2bc25c5c990363eb8f8eb54693b0c44eb198b019c4cef11899011c15c99c5e3277b0ec5f6d145073cc318fec1c1c6c17ba31cb204f8bcfb333;
    5'b11010 : xpb = 1024'h2a9516fb422517346c4839766dbe9f9aa61bca4215d1f1d1a844bb91d0e30694107896ed8f8b0cf0f5f9714a8d173e3978484752268f084be7699597d72ad53cf5c7987ca5166d96ac28c6ce9900114f93efecfbdc2dafcdd941e332deaa867c030908068af95d25fad48b32ae663c8417fa8dd45e35fdaf17e1f352e8cc9581;
    5'b11011 : xpb = 1024'h3303f325c24d37aa78415dd206496d68a703dc019506014a9fe38ed5cc1d175524ec52ca1cd6cd622cf2f815116a862fc5ae86acee4ca451bc0776663a521d0134efdb74771cde0195f531042e9c370f992a9364079710ea19d3aca0ee63f45f04f5fa43799487d444bcb6f8487c053bfe652f8c9fffe3a3fdf8c65645c977cf;
    5'b11100 : xpb = 1024'h3b72cf5042755820843a822d9ed43b36a7ebedc1143a10c397826219c757281639600ea6aa228dd363ec7edf95bdce261314c607b60a405790a557349d7964c574181e6c49234e6c7fc19b39c4385ccf9e6539cc330072065a65760efe1d624206e2ec80682fb2828ea4e2bde291cdf3e4cfd144e1c9c998e40f9959a2c65a1d;
    5'b11101 : xpb = 1024'h43e1ab7ac29d78969033a689375f0904a8d3ff80936e203c8f21355dc29138d74dd3ca83376e4e449ae605aa1a11161c607b05627dc7dc5d6543380300a0ac89b34061641b29bed7698e056f59d4828fa39fe0345e69d3229af73f7d0dd6d02508cfdebd56cadd30d88d0e837ca796abcb3a72fd2393af8dca266c5cffc33c6b;
    5'b11110 : xpb = 1024'h4c5087a542c5990c9c2ccae4cfe9d6d2a9bc114012a22fb586c008a1bdcb49986247865fc4ba0eb5d1df8c749e645e12ade144bd4585786339e118d163c7f44df268a45bed302f42535a6fa4ef70a84fa8da869c89d3343edb8908eb1d903e080abcd0fa456607df22753a4916bd5f63b1a514b5655d9582b03d3f605cc01eb9;
    5'b11111 : xpb = 1024'h54bf63cfc2edb982a825ef406874a4a0aaa422ff91d63f2e7e5edbe5b9055a5976bb423c5205cf2708d9133f22b7a608fb4784180d4314690e7ef99fc6ef3c123190e753bf369fad3d26d9da850cce0fae152d04b53c955b1c1ad2592d49abeb0ca9c3373401328d6c5d660eb0d3281b980fb66da7277b7796541263b9bd0107;
    endcase
end

endmodule

module xpb_5_155
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h16f54fa08ac47c3bc62eb3e4111fb4e9009c586e6f0327894f65b2be6bb06e5cf3eee2c5f5b3ec7b3d8128c9f911c3797ce6cd1e9c7ef695e74ebe27d9dc9cb917d54f965f806850c02c7bd5153b622ac15d4881478a9384b2287bf15183c8b9f5c9b9b029af4cf4d675f34523db2e7e69ceb9c2b279ce51a9920986e1f1757e;
    5'b00010 : xpb = 1024'h2dea9f411588f8778c5d67c8223f69d20138b0dcde064f129ecb657cd760dcb9e7ddc58beb67d8f67b025193f22386f2f9cd9a3d38fded2bce9d7c4fb3b939722faa9f2cbf00d0a18058f7aa2a76c45582ba91028f1527096450f7e2a3079173eb937360535e99e9acebe68a47b65cfcd39d738564f39ca35324130dc3e2eafc;
    5'b00011 : xpb = 1024'h44dfeee1a04d74b3528c1bac335f1ebb01d5094b4d09769bee31183b43114b16dbcca851e11bc571b8837a5deb354a6c76b4675bd57ce3c1b5ec3a778d95d62b477feec31e8138f24085737f3fb226804417d983d69fba8e167973d3f48b5a2de15d2d107d0de6de8361d9cf6b918b7b3d6c2d48176d6af4fcb61c94a5d4607a;
    5'b00100 : xpb = 1024'h5bd53e822b11f0ef18bacf90447ed3a4027161b9bc0c9e253d96caf9aec1b973cfbb8b17d6cfb1ecf604a327e4470de5f39b347a71fbda579d3af89f677272e45f553e597e01a14300b1ef5454ed88ab057522051e2a4e12c8a1efc5460f22e7d726e6c0a6bd33d359d7cd148f6cb9f9a73ae70ac9e73946a648261b87c5d5f8;
    5'b00101 : xpb = 1024'h72ca8e22b5d66d2adee98374559e888d030dba282b0fc5ae8cfc7db81a7227d0c3aa6dddcc839e683385cbf1dd58d15f708201990e7ad0ed8489b6c7414f0f9d772a8defdd820993c0de6b296a28ead5c6d26a8665b4e1977aca6bb69792eba1ccf0a070d06c80c8304dc059b347e8781109a0cd7c6107984fda2fa269b74b76;
    5'b00110 : xpb = 1024'h89bfddc3409ae966a518375866be3d7603aa12969a12ed37dc6230768622962db79950a3c2378ae37106f4bbd66a94d8ed68ceb7aaf9c7836bd874ef1b2bac568effdd863d0271e4810ae6fe7f644d00882fb307ad3f751c2cf2e7a7e916b45bc2ba5a20fa1bcdbd06c3b39ed72316f67ad85a902edad5e9f96c39294ba8c0f4;
    5'b00111 : xpb = 1024'ha0b52d63cb5f65a26b46eb3c77ddf25f04466b05091614c12bc7e334f1d3048aab883369b7eb775eae881d85cf7c58526a4f9bd64778be1953273316f508490fa6d52d1c9c82da35413762d3949faf2b498cfb88f4ca08a0df1b63993a9a7d15b88413d123cb1ab1dd39a6e3fafe4574e4a71452e154a43ba2fe42b02d9a3672;
    5'b01000 : xpb = 1024'h6fd37ae9435ad156670274978a35ff6936cc042a2a19bd2fd50dc9daa80c5df9c2e98b6e378e54b4cab0708e5300b01831c410ec144e46389d6b1e0941271174a5b48044c724540eec9dc0610ff4d2516e54a71afce6f14dbb74d8fd1f3a33d7f463b579cb16f192cefb34a27094dc9ff9bef334383155d0620d13286a94585;
    5'b01001 : xpb = 1024'h1df2874f1efa29512c9edb2d89c314df940918b111a4c35c4cb68f5c1631343c901d7b7cd92cd1c68a2c2fd2de41ce7b00030e2d5dc3daf9712570086def0dd06230979aabf2ad91aef657db263aaf4fd84292f2f75902998ddfc98123776bf7750ff507c660bc0e0365a68f4ae47c48696aa8f5f5fce3aeafb2dab9689abb03;
    5'b01010 : xpb = 1024'h34e7d6efa9bea58cf2cd8f119ae2c9c894a5711f80a7eae59c1c421a81e1a299840c5e42cee0be41c7ad589cd75391f47ce9db4bfa42d18f58742e3047cbaa897a05e7310b7315e26f22d3b03b76117a999fdb743ee3961e4008457274fb34b16ad9aeb7f0100902d9db99d46ebfaac6d33962b8a876b2005944e4404a8c3081;
    5'b01011 : xpb = 1024'h4bdd2690348321c8b8fc42f5ac027eb19541c98defab126eeb81f4d8ed9210f677fb4108c494aabd052e8166d065556df9d0a86a96c1c8253fc2ec5821a8474291db36c76af37e332f4f4f8550b173a55afd23f5866e29a2f230c163c67efd6b60a3686819bf55f7b0518d19929ad9453d081c7b5af0805202d6edc72c7da5ff;
    5'b01100 : xpb = 1024'h62d27630bf479e047f2af6d9bd22339a95de21fc5eae39f83ae7a79759427f536bea23ceba48973842afaa30c97718e776b775893340bebb2711aa7ffb84e3fba9b0865dca73e683ef7bcb5a65ecd5d01c5a6c76cdf8bd27a4593d551802c625566d2218436ea2ec86c7805eb67607c3a6d6d63e0d6a4ea3ac68f74e0e6f1b7d;
    5'b01101 : xpb = 1024'h79c7c5d14a0c1a404559aabdce41e883967a7a6acdb161818a4d5a55c4f2edb05fd90694affc83b38030d2fac288dc60f39e42a7cfbfb5510e6068a7d56180b4c185d5f429f44ed4afa8472f7b2837faddb7b4f8158350ac5681b94669868edf4c36dbc86d1defe15d3d73a3da51364210a59000bfe41cf555fb00d4f06090fb;
    5'b01110 : xpb = 1024'h90bd1571d4d0967c0b885ea1df619d6c9716d2d93cb4890ad9b30d1430a35c0d53c7e95aa5b0702ebdb1fbc4bb9a9fda70850fc66c3eabe6f5af26cfaf3e1d6dd95b258a8974b7256fd4c30490639a259f14fd795d0de43108aa3537bb0a57994200957896cd3cd633b366e8fe2c64c07a7449c3725deb46ff8d0a5bd2520679;
    5'b01111 : xpb = 1024'ha7b265125f9512b7d1b71285f081525597b32b47abb7b0942918bfd29c53ca6a47b6cc209b645ca9fb33248eb4ac6353ed6bdce508bda27cdcfde4f7891aba26f1307520e8f51f7630013ed9a59efc50607245faa49877b5bad2b1290c8e205337ca4f28c07c89cb0a295a2e2207933ee443038624d7b998a91f13e2b4437bf7;
    5'b10000 : xpb = 1024'hdfa6f5d286b5a2acce04e92f146bfed26d98085454337a5faa1b93b55018bbf385d316dc6f1ca9699560e11ca6016030638821d8289c8c713ad63c12824e22e94b6900898e48a81dd93b80c21fe9a4a2dca94e35f9cde29b76e9b1fa3e7467afe8c76af3962de3259df66944e129b93ff37de6687062aba0c41a2650d528b0a;
    5'b10001 : xpb = 1024'h24efbefdb32fd666930f0277026674d62775d8f3b4465f2f4a076bf9c0b1fa1c2c4c1433bca5b711d6d736dbc371d97c831f4f3c1f08bf5cfafc21e902017ee7ac8bdf9ef864f2d29dc033e13739fc74ef27dd64a72771ae69971710f56b0f34f456305f63122b27305559d971edca1269069829397ff90bb5d3abebef440088;
    5'b10010 : xpb = 1024'h3be50e9e3df452a2593db65b138629bf28123162234986b8996d1eb82c626879203af6f9b259a38d14585fa5bc839cf600061c5abb87b5f2e24ae010dbde1ba0c4612f3557e55b235decafb64c755e9fb08525e5eeb205331bbf930246eed7eeea1fea0f8cc1781c06cb4d1e95c8f890d2d551ebebf9c75d5f65b572d1357606;
    5'b10011 : xpb = 1024'h52da5e3ec8b8cede1f6c6a3f24a5dea828ae89d0924cae41e8d2d1769812d6d61429d9bfa80d900851d9886fb595606f7cece9795806ac88c9999e38b5bab859dc367ecbb765c3741e192b8b61b0c0ca71e26e67363c98b7cde80ef39872a0a8dfe9a3bfb670c510dd414063b9a4270f3ca40bae9e7395af08f7bef9b326eb84;
    5'b10100 : xpb = 1024'h69cfaddf537d4b19e59b1e2335c59391294ae23f014fd5cb3838843503c345330818bc859dc17c838f5ab139aea723e8f9d3b697f485a31eb0e85c608f975512f40bce6216e62bc4de45a76076ec22f5333fb6e87dc72c3c80108ae4e9f66962d5b35d6fe0201205b3b733a8dd7f558da672c57150ed6400b289c88095186102;
    5'b10101 : xpb = 1024'h80c4fd7fde41c755abc9d20746e5487a29e73aad7052fd54879e36f36f73b38ffc079f4b937568feccdbda03a7b8e76276ba83b6910499b498371a886973f1cc0be11df8766694159e7223358c27851ff49cff69c551bfc1323906d63b7a321ccb7d172009cf5efa8a2d26ee015a840c10417f34036732525c1bd2077709d680;
    5'b10110 : xpb = 1024'h97ba4d206906439171f885eb5804fd632a83931bdf5624ddd703e9b1db2421eceff682118929557a0a5d02cda0caaadbf3a150d52d83904a7f85d8b043508e8523b66d8ed5e6fc665e9e9f0aa162e74ab5fa47eb0cdc5345e46182c78cfdfad6c146d0d0337eabef60a31a332535b28a7a1038f6b5e100a405addb8e58fb4bfe;
    5'b10111 : xpb = 1024'haeaf9cc0f3cabfcd382739cf6924b24c2b1feb8a4e594c6726699c7046d49049e3e564d77edd41f547de2b9799dc6e5570881df3ca0286e066d496d81d2d2b3e3b8bbd25356764b71ecb1adfb69e49757757906c5466e6ca9689feb8de81c390b7108a805d2df8e437190d784910e108e3def2b9685acef5af3fe5153aecc17c;
    5'b11000 : xpb = 1024'h14f7a70bbca10740335075dc69ea1fe3ba4640c7e7e4d378f7f295d8ff82519ed48bca24aa6aafe1e601151aaf9021048954c32c43cead2a9d8415a1bc375345df11d80ce556cfc2cc5d941232fde76f44afdf550f6b4d3e9325e8af75dae9b87dd2b206d6144d4b86cf19de751be95dfed3cd99ca8940171262739793fbd08f;
    5'b11001 : xpb = 1024'h2becf6ac4765837bf97f29c07b09d4ccbae2993656e7fb02475848976b32bffbc87aaceaa01e9c5d23823de4a8a1e47e063b904ae04da3c084d2d3c99613effef6e727a344d738138c8a0fe74839499a060d27d656f5e0c3454e64a0c75eb272739c6bb6ffc39a405d450d2398f717dc68a2875c7d030e68bbf47d1e75ed460d;
    5'b11010 : xpb = 1024'h42e2464cd229ffb7bfaddda48c2989b5bb7ef1a4c5eb228b96bdfb55d6e32e58bc698fb095d288d8610366aea1b3a7f783225d697ccc9a566c2191f16ff08cb80ebc7739a457a0644cb68bbc5d74abc4c76a70579e807447f776e09218e27b2c696625672972e73533bb0068bcd2465ad271411f2f7cdcba658686a557debb8b;
    5'b11011 : xpb = 1024'h59d795ed5cee7bf385dc91889d493e9ebc1b4a1334ee4a14e623ae1442939cb5b05872768b8675539e848f789ac56b7100092a88194b90ec5370501949cd29712691c6d003d808b50ce3079172b00def88c7b8d8e60b07cca99f5c836a6643e65f2fdf175322342a0a30f3ade0ad74d93c3ffae1e1f6ab0c0f18902c39d03109;
    5'b11100 : xpb = 1024'h70cce58de7b2f82f4c0b456cae68f387bcb7a281a3f1719e358960d2ae440b12a447553c813a61cedc05b84293d72eea7ceff7a6b5ca87823abf0e4123a9c62a3e67166663587105cd0f836687eb701a4a25015a2d959b515bc7d874bbea0ca054f998c77cd1811ee0a6e6f30488a357a60eb4a49470795db8aa99b31bc1a687;
    5'b11101 : xpb = 1024'h87c2352e7277746b1239f950bf88a870bd53faf012f4992784ef139119f4796f9836380276ee4e4a1986e10c8ce8f263f9d6c4c552497e18220dcc68fd8662e3563c65fcc2d8d9568d3bff3b9d26d2450b8249db75202ed60df054660d6dd55a4ac35277a680ce13b71cda382863d1d60fdd6e6746ea47af623ca339fdb31c05;
    5'b11110 : xpb = 1024'h9eb784cefd3bf0a6d868ad34d0a85d59bdf0535e81f7c0b0d454c64f85a4e7cc8c251ac86ca23ac5570809d685fab5dd76bd91e3eec874ae095c8a90d762ff9c6e11b593225941a74d687b10b262346fccdf925cbcaac25ac018d0575ef19e14408d0c27d0301b088d92cd7d4c3f005479ac2829f96416010bceacc0dfa49183;
    5'b11111 : xpb = 1024'h4ff8f19c6123819d391e941d16dcaf14d16a89c1b8347c2a5ddbfb83e52a9217ccb8015982fa8b1f52af3599bae688c8f8a371c68949af8400c095a766d27a41197d07ad248acb2fafaf4432ec1d2699a37e14577af28cebcb4ba4df64ac43c074f33ae49166f6fdd48d9e3784a08a994a1030a5b9287226ef13b4338b3a096;
    endcase
end

endmodule

module xpb_5_90
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h18461f205c95e678c730bc4548ea585a001ea4885d1309e809b0be8438bc1891f755a2848c1f1c82c12fb4cc9ed9f91d1e6562bfd101f8b15e33ca4487d9a86ee0ef502175f6a398da40146d83437cd0b546a9700e3ed60bc9e9ed41f167f300c9542222b6cfb9bc671bf95c81bf4129c65123c083509e4569d72528698534e4;
    5'b00010 : xpb = 1024'h308c3e40b92bccf18e61788a91d4b0b4003d4910ba2613d013617d0871783123eeab4509183e3905825f69993db3f23a3ccac57fa203f162bc6794890fb350ddc1dea042ebed4731b48028db0686f9a16a8d52e01c7dac1793d3da83e2cfe60192a844456d9f7378ce37f2b9037e82538ca2478106a13c8ad3ae4a50d30a69c8;
    5'b00011 : xpb = 1024'h48d25d6115c1b36a559234cfdabf090e005bed9917391db81d123b8caa3449b5e600e78da45d5588438f1e65dc8deb575b30283f7305ea141a9b5ecd978cf94ca2cdf06461e3eaca8ec03d4889ca76721fd3fc502abc82235dbdc7c5d437d9025bfc6668246f2d353553ec15853dc37d52f36b4189f1dad03d856f793c8f9eac;
    5'b00100 : xpb = 1024'h61187c81725799e31cc2f11523a96168007a9221744c27a026c2fa10e2f06247dd568a12307c720b04bed3327b67e47479958aff4407e2c578cf29121f66a1bb83bd4085d7da8e63690051b60d0df342d51aa5c038fb582f27a7b507c59fcc032550888adb3ee6f19c6fe57206fd04a719448f020d427915a75c94a1a614d390;
    5'b00101 : xpb = 1024'h795e9ba1ceed805be3f3ad5a6c93b9c2009936a9d15f31883073b8951bac7ad9d4ac2c96bc9b8e8dc5ee87ff1a41dd9197faedbf1509db76d702f356a7404a2a64ac90a74dd131fc43406623905170138a614f30473a2e3af191a249b707bf03eea4aaad920ea0ae038bdece88bc45d0df95b2c29093175b1133b9ca0f9a0874;
    5'b00110 : xpb = 1024'h91a4bac22b8366d4ab24699fb57e121c00b7db322e723b703a2477195468936bcc01cf1b48baab10871e3ccbb91bd6aeb660507ee60bd4283536bd9b2f19f299459be0c8c3c7d5951d807a911394ece43fa7f8a055790446bb7b8f8ba86fb204b7f8ccd048de5a6a6aa7d82b0a7b86faa5e6d68313e3b5a07b0adef2791f3d58;
    5'b00111 : xpb = 1024'ha9ead9e288194d4d725525e4fe686a7600d67fba8b85455843d5359d8d24abfdc357719fd4d9c793484df19857f5cfcbd4c5b33eb70dccd9936a87dfb6f39b08268b30ea39be792df7c08efe96d869b4f4eea21063b7da5285657ccd99d7a505814ceef2ffae1426d1c3d1878c3ac8246c37fa43973453e5e4e2041ae2a4723c;
    5'b01000 : xpb = 1024'h1183b3ad22c0fefd6e806a5336f87b7e8f7f21121320aec8cfa93acc12de1787b76496ab96d265876a1f671e1371b81e8f10ee18655cf53f40ff12c603facec5932b4c5d00241f81bf66a0c981402254b63051e7e570834d99c2d814d114f5741b997eec05b4d555b21fe4051629e324e3af3f21ca3994fb0849ae3ec34740b5;
    5'b01001 : xpb = 1024'h29c9d2cd7f56e57635b126987fe2d3d88f9dc59a7033b8b0d959f9504b9a3019aeba393022f1820a2b4f1beab24bb13bad7650d8365eedf09f32dd0a8bd47734741a9c7e761ac31a99a6b53704839f256b76fb57f3af595963acc556c27ce874e4eda10ebc848f12193bdd6197e9244eaa0062e24d8a33407220d3672ccc7599;
    5'b01010 : xpb = 1024'h420ff1eddbeccbeefce1e2ddc8cd2c328fbc6a22cd46c298e30ab7d4845648aba60fdbb4af109e8cec7ed0b75125aa58cbdbb3980760e6a1fd66a74f13ae1fa35509ec9fec1166b373e6c9a487c71bf620bda4c801ee2f652d96b298b3e4db75ae41c331735448ce8057d6be19a86578705186a2d0dad185dbf7f88f9651aa7d;
    5'b01011 : xpb = 1024'h5a56110e3882b267c4129f2311b7848c8fdb0eab2a59cc80ecbb7658bd12613d9d657e393b2fbb0fadae8583efffa375ea411657d862df535b9a71939b87c81235f93cc162080a4c4e26de120b0a98c6d6044e38102d0570f7809fdaa54cce767795e5542a24028ae773d01a9b67a6a236a2aa63542b6fcb45cf1db7ffd6df61;
    5'b01100 : xpb = 1024'h729c302e951898e08b435b685aa1dce68ff9b333876cd668f66c34dcf5ce79cf94bb20bdc74ed7926ede3a508ed99c9308a67917a964d804b9ce3bd82361708116e88ce2d7feade52866f27f8e4e15978b4af7a81e6bdb7cc16a8d1c96b4c17740ea0776e0f3bc474e8fc9771d26e7cbfcf3ce23d77c0e10afa642e0695c1445;
    5'b01101 : xpb = 1024'h8ae24f4ef1ae7f59527417ada38c3540901857bbe47fe051001cf3612e8a92618c10c342536df415300def1d2db395b0270bdbd77a66d0b61802061cab3b18eff7d7dd044df5517e02a706ed119192684091a1182caab1888b547a5e881cb4780a3e299997c37603b5abc2d39ee628f5c344f1e45accac56197d6808d2e14929;
    5'b01110 : xpb = 1024'ha3286e6f4e4465d219a4d3f2ec768d9a9036fc444192ea3909cdb1e56746aaf3836665c6df8d1097f13da3e9cc8d8ecd45713e974b68c9677635d0613314c15ed8c72d25c3ebf516dce71b5a94d50f38f5d84a883ae98794553e67a07984a778d3924bbc4e932fc01cc7bc3020a56a1f899615a4de1d4a9b83548d313c667e0d;
    5'b01111 : xpb = 1024'hac14839e8ec178215d0186125069ea31edf9d9bc92e53a995a1b713ed00167d77738ad2a185ae8c130f196f8809771fffbc7970f9b7f1cd23ca5b47801bf51c456748988a519b6aa48d2d257f3cc7d8b719fa5fbca2308f699bc2e7b0c1f7e76ddedbb55499f0eefd23ceadaa948520010d5a8311228bb0a6bc37551d094c86;
    5'b10000 : xpb = 1024'h2307675a4581fdfadd00d4a66df0f6fd1efe422426415d919f52759825bc2f0f6ec92d572da4cb0ed43ece3c26e3703d1e21dc30cab9ea7e81fe258c07f59d8b265698ba00483f037ecd4193028044a96c60a3cfcae1069b3385b029a229eae83732fdd80b69aaab643fc80a2c53c649c75e7e43947329f610935c7d868e816a;
    5'b10001 : xpb = 1024'h3b4d867aa217e473a43190ebb6db4f571f1ce6ac83546779a903341c5e7847a1661ecfdbb9c3e791956e8308c5bd695a3c873ef09bbbe32fe031efd08fcf45fa0745e8db763ee29c590d560085c3c17a21a74d3fd91fdca6fd6f9d6b9391dde900871ffac2396467cb5bc166ae1307738dafa20417c3c83b7a6a81a5f013b64e;
    5'b10010 : xpb = 1024'h5393a59afeadcaec6b624d30ffc5a7b11f3b8b34e0677161b2b3f2a0973460335d74726045e30414569e37d5649762775aeca1b06cbddbe13e65ba1517a8ee68e83538fcec358635334d6a6e09073e4ad6edf6afe75eb2b2c7598aad84f9d0e9c9db421d79091e243277bac32fd2489d5400c5c49b146680e441a6ce5998eb32;
    5'b10011 : xpb = 1024'h6bd9c4bb5b43b1653293097648b0000b1f5a2fbd3d7a7b49bc64b124cff078c554ca14e4d202209717cdeca203715b94795204703dbfd4929c9984599f8296d7c924891e622c29ce0d8d7edb8c4abb1b8c34a01ff59d88be914377ef7661c3ea932f64402fd8d7e09993b41fb19189c71a51e9851e6504c64e18cbf6c31e2016;
    5'b10100 : xpb = 1024'h841fe3dbb7d997ddf9c3c5bb919a58651f78d4459a8d8531c6156fa908ac91574c1fb7695e213d19d8fda16ea24b54b197b767300ec1cd43facd4e9e275c3f46aa13d93fd822cd66e7cd93490f8e37ec417b499003dc5eca5b2d653167c9b6eb5c838662e6a8919d00afad7c3350caf0e0a30d45a1b5a30bb7eff11f2ca354fa;
    5'b10101 : xpb = 1024'h9c6602fc146f7e56c0f48200da84b0bf1f9778cdf7a08f19cfc62e2d4168a9e9437559edea40599c9a2d563b41254dceb61cc9efdfc3c5f5590118e2af35e7b58b0329614e1970ffc20da7b692d1b4bcf6c1f300121b34d6251752735931a9ec25d7a8859d784b5967cba6d8b5100c1aa6f431062506415121c71647962889de;
    5'b10110 : xpb = 1024'h3fedcc6af173006bd1fc66f1314c1c7ae401a257f3bf88a5b9a335bc722157337827ef9ac38f790bbfecbc0fca13621706804c98e12ee5b0695a3c8fc3d1b72f7a344d4147f175389b3b9817d396d5cb803a2d793d3ddd13974adba906efa5ac024387ea37f0c884827b9563eff271b1e6b75e4580b8266452ec06b76cb5857;
    5'b10111 : xpb = 1024'h1c44fbe70bad167f845082b45bff1a21ae5ebeaddc4f0272654af1dfffde2e052ed8217e385814137d2e808d9b7b2f3e8ecd67895f14e70c64c96e0d8416c3e1d89294f58a75baec63f3cdef007cea2d6d4a4c47a212b3dd035e9afc81d6ed5b89785aa15a4ec644af43b2b2c0be6844e4bc99a4db5c20abaf05e593e0508d3b;
    5'b11000 : xpb = 1024'h348b1b076842fcf84b813ef9a4e9727bae7d633639620c5a6efbb064389a4697262dc402c47730963e5e355a3a55285bad32ca493016dfbdc2fd38520bf06c50b981e517006c5e853e33e25c83c066fe2290f5b7b05189e8cd48883e733ee05c52cc7cc4111e8001165fac0f427da96eab0dbd655eacbef118dd0abc49d5c21f;
    5'b11001 : xpb = 1024'h4cd13a27c4d8e37112b1fb3eedd3cad5ae9c07be9675164278ac6ee871565f291d83668750964d18ff8dea26d92f2178cb982d090118d86f2131029693ca14bf9a7135387663021e1873f6ca0703e3ced7d79f27be905ff49732758064a6d35d1c209ee6c7ee39bd7d7ba56bc43cea98715ee125e1fd5d3682b42fe4b35af703;
    5'b11010 : xpb = 1024'h65175948216ec9e9d9e2b78436be232faebaac46f388202a825d2d6caa1277bb14d9090bdcb5699bc0bd9ef378091a95e9fd8fc8d21ad1207f64ccdb1ba3bd2e7b608559ec59a5b6f2b40b378a47609f8d1e4897cccf3600611c62c2560ec65de574c1097ebdf379e4979ec845fc2bc237b004e6654dfb7bec8b550d1ce02be7;
    5'b11011 : xpb = 1024'h7d5d78687e04b062a11373c97fa87b89aed950cf509b2a128c0debf0e2ce904d0c2eab9068d4861e81ed53c016e313b30862f288a31cc9d1dd98971fa37d659d5c4fd57b6250494fccf41fa50d8add704264f207db0e0c0c2b0650044776b95eaec8e32c358dad364bb39824c7bb6cebfe0128a6e89e99c156627a35866560cb;
    5'b11100 : xpb = 1024'h95a39788da9a96db6844300ec892d3e3aef7f557adae33fa95beaa751b8aa8df03844e14f4f3a2a1431d088cb5bd0cd026c85548741ec2833bcc61642b570e0c3d3f259cd846ece8a734341290ce5a40f7ab9b77e94ce217f4f03d4638deac5f781d054eec5d66f2b2cf9181497aae15c4524c676bef3806c0399f5defea95af;
    5'b11101 : xpb = 1024'hade9b6a937307d542f74ec54117d2c3daf1699e00ac13de29f6f68f95446c170fad9f0998112bf24044cbd59549705ed452db8084520bb349a002ba8b330b67b1e2e75be4e3d9081817448801411d711acf244e7f78bb823beda2a882a469f6041712771a32d20af19eb8addcb39ef3f8aa37027ef3fd64c2a10c486596fca93;
    5'b11110 : xpb = 1024'h15829073d1d82f042ba030c24a0d3d463dbf3b37925ca7532b436e27da002cfaeee715a5430b5d18261e32df1012ee3fff78f2e1f36fe39a4794b68f0037ea388ace913114a336d5491a5a4afe798fb16e33f4bf7944611ed33785cf6183efcedbbdb76aa933e1ddfa479d5b55290a40021ab506224517614d786eaa3a12990c;
    5'b11111 : xpb = 1024'h2dc8af942e6e157cf2d0ed0792f795a03ddddfbfef6fb13b34f42cac12bc458ce63cb829cf2a799ae74de7abaeece75d1dde55a1c471dc4ba5c880d3881192a76bbde1528a99da6e235a6eb881bd0c82237a9e2f8783372a9d21731152ebe2cfa511d98d60039b9a616396b7d6e84b69c86bd8c6a595b5a6b74f93d2a397cdf0;
    endcase
end

endmodule

module compressor_array_48_16_1030
(
    input  [47:0] col_in_0,
    input  [47:0] col_in_1,
    input  [47:0] col_in_2,
    input  [47:0] col_in_3,
    input  [47:0] col_in_4,
    input  [47:0] col_in_5,
    input  [47:0] col_in_6,
    input  [47:0] col_in_7,
    input  [47:0] col_in_8,
    input  [47:0] col_in_9,
    input  [47:0] col_in_10,
    input  [47:0] col_in_11,
    input  [47:0] col_in_12,
    input  [47:0] col_in_13,
    input  [47:0] col_in_14,
    input  [47:0] col_in_15,
    input  [47:0] col_in_16,
    input  [47:0] col_in_17,
    input  [47:0] col_in_18,
    input  [47:0] col_in_19,
    input  [47:0] col_in_20,
    input  [47:0] col_in_21,
    input  [47:0] col_in_22,
    input  [47:0] col_in_23,
    input  [47:0] col_in_24,
    input  [47:0] col_in_25,
    input  [47:0] col_in_26,
    input  [47:0] col_in_27,
    input  [47:0] col_in_28,
    input  [47:0] col_in_29,
    input  [47:0] col_in_30,
    input  [47:0] col_in_31,
    input  [47:0] col_in_32,
    input  [47:0] col_in_33,
    input  [47:0] col_in_34,
    input  [47:0] col_in_35,
    input  [47:0] col_in_36,
    input  [47:0] col_in_37,
    input  [47:0] col_in_38,
    input  [47:0] col_in_39,
    input  [47:0] col_in_40,
    input  [47:0] col_in_41,
    input  [47:0] col_in_42,
    input  [47:0] col_in_43,
    input  [47:0] col_in_44,
    input  [47:0] col_in_45,
    input  [47:0] col_in_46,
    input  [47:0] col_in_47,
    input  [47:0] col_in_48,
    input  [47:0] col_in_49,
    input  [47:0] col_in_50,
    input  [47:0] col_in_51,
    input  [47:0] col_in_52,
    input  [47:0] col_in_53,
    input  [47:0] col_in_54,
    input  [47:0] col_in_55,
    input  [47:0] col_in_56,
    input  [47:0] col_in_57,
    input  [47:0] col_in_58,
    input  [47:0] col_in_59,
    input  [47:0] col_in_60,
    input  [47:0] col_in_61,
    input  [47:0] col_in_62,
    input  [47:0] col_in_63,
    input  [47:0] col_in_64,
    input  [47:0] col_in_65,
    input  [47:0] col_in_66,
    input  [47:0] col_in_67,
    input  [47:0] col_in_68,
    input  [47:0] col_in_69,
    input  [47:0] col_in_70,
    input  [47:0] col_in_71,
    input  [47:0] col_in_72,
    input  [47:0] col_in_73,
    input  [47:0] col_in_74,
    input  [47:0] col_in_75,
    input  [47:0] col_in_76,
    input  [47:0] col_in_77,
    input  [47:0] col_in_78,
    input  [47:0] col_in_79,
    input  [47:0] col_in_80,
    input  [47:0] col_in_81,
    input  [47:0] col_in_82,
    input  [47:0] col_in_83,
    input  [47:0] col_in_84,
    input  [47:0] col_in_85,
    input  [47:0] col_in_86,
    input  [47:0] col_in_87,
    input  [47:0] col_in_88,
    input  [47:0] col_in_89,
    input  [47:0] col_in_90,
    input  [47:0] col_in_91,
    input  [47:0] col_in_92,
    input  [47:0] col_in_93,
    input  [47:0] col_in_94,
    input  [47:0] col_in_95,
    input  [47:0] col_in_96,
    input  [47:0] col_in_97,
    input  [47:0] col_in_98,
    input  [47:0] col_in_99,
    input  [47:0] col_in_100,
    input  [47:0] col_in_101,
    input  [47:0] col_in_102,
    input  [47:0] col_in_103,
    input  [47:0] col_in_104,
    input  [47:0] col_in_105,
    input  [47:0] col_in_106,
    input  [47:0] col_in_107,
    input  [47:0] col_in_108,
    input  [47:0] col_in_109,
    input  [47:0] col_in_110,
    input  [47:0] col_in_111,
    input  [47:0] col_in_112,
    input  [47:0] col_in_113,
    input  [47:0] col_in_114,
    input  [47:0] col_in_115,
    input  [47:0] col_in_116,
    input  [47:0] col_in_117,
    input  [47:0] col_in_118,
    input  [47:0] col_in_119,
    input  [47:0] col_in_120,
    input  [47:0] col_in_121,
    input  [47:0] col_in_122,
    input  [47:0] col_in_123,
    input  [47:0] col_in_124,
    input  [47:0] col_in_125,
    input  [47:0] col_in_126,
    input  [47:0] col_in_127,
    input  [47:0] col_in_128,
    input  [47:0] col_in_129,
    input  [47:0] col_in_130,
    input  [47:0] col_in_131,
    input  [47:0] col_in_132,
    input  [47:0] col_in_133,
    input  [47:0] col_in_134,
    input  [47:0] col_in_135,
    input  [47:0] col_in_136,
    input  [47:0] col_in_137,
    input  [47:0] col_in_138,
    input  [47:0] col_in_139,
    input  [47:0] col_in_140,
    input  [47:0] col_in_141,
    input  [47:0] col_in_142,
    input  [47:0] col_in_143,
    input  [47:0] col_in_144,
    input  [47:0] col_in_145,
    input  [47:0] col_in_146,
    input  [47:0] col_in_147,
    input  [47:0] col_in_148,
    input  [47:0] col_in_149,
    input  [47:0] col_in_150,
    input  [47:0] col_in_151,
    input  [47:0] col_in_152,
    input  [47:0] col_in_153,
    input  [47:0] col_in_154,
    input  [47:0] col_in_155,
    input  [47:0] col_in_156,
    input  [47:0] col_in_157,
    input  [47:0] col_in_158,
    input  [47:0] col_in_159,
    input  [47:0] col_in_160,
    input  [47:0] col_in_161,
    input  [47:0] col_in_162,
    input  [47:0] col_in_163,
    input  [47:0] col_in_164,
    input  [47:0] col_in_165,
    input  [47:0] col_in_166,
    input  [47:0] col_in_167,
    input  [47:0] col_in_168,
    input  [47:0] col_in_169,
    input  [47:0] col_in_170,
    input  [47:0] col_in_171,
    input  [47:0] col_in_172,
    input  [47:0] col_in_173,
    input  [47:0] col_in_174,
    input  [47:0] col_in_175,
    input  [47:0] col_in_176,
    input  [47:0] col_in_177,
    input  [47:0] col_in_178,
    input  [47:0] col_in_179,
    input  [47:0] col_in_180,
    input  [47:0] col_in_181,
    input  [47:0] col_in_182,
    input  [47:0] col_in_183,
    input  [47:0] col_in_184,
    input  [47:0] col_in_185,
    input  [47:0] col_in_186,
    input  [47:0] col_in_187,
    input  [47:0] col_in_188,
    input  [47:0] col_in_189,
    input  [47:0] col_in_190,
    input  [47:0] col_in_191,
    input  [47:0] col_in_192,
    input  [47:0] col_in_193,
    input  [47:0] col_in_194,
    input  [47:0] col_in_195,
    input  [47:0] col_in_196,
    input  [47:0] col_in_197,
    input  [47:0] col_in_198,
    input  [47:0] col_in_199,
    input  [47:0] col_in_200,
    input  [47:0] col_in_201,
    input  [47:0] col_in_202,
    input  [47:0] col_in_203,
    input  [47:0] col_in_204,
    input  [47:0] col_in_205,
    input  [47:0] col_in_206,
    input  [47:0] col_in_207,
    input  [47:0] col_in_208,
    input  [47:0] col_in_209,
    input  [47:0] col_in_210,
    input  [47:0] col_in_211,
    input  [47:0] col_in_212,
    input  [47:0] col_in_213,
    input  [47:0] col_in_214,
    input  [47:0] col_in_215,
    input  [47:0] col_in_216,
    input  [47:0] col_in_217,
    input  [47:0] col_in_218,
    input  [47:0] col_in_219,
    input  [47:0] col_in_220,
    input  [47:0] col_in_221,
    input  [47:0] col_in_222,
    input  [47:0] col_in_223,
    input  [47:0] col_in_224,
    input  [47:0] col_in_225,
    input  [47:0] col_in_226,
    input  [47:0] col_in_227,
    input  [47:0] col_in_228,
    input  [47:0] col_in_229,
    input  [47:0] col_in_230,
    input  [47:0] col_in_231,
    input  [47:0] col_in_232,
    input  [47:0] col_in_233,
    input  [47:0] col_in_234,
    input  [47:0] col_in_235,
    input  [47:0] col_in_236,
    input  [47:0] col_in_237,
    input  [47:0] col_in_238,
    input  [47:0] col_in_239,
    input  [47:0] col_in_240,
    input  [47:0] col_in_241,
    input  [47:0] col_in_242,
    input  [47:0] col_in_243,
    input  [47:0] col_in_244,
    input  [47:0] col_in_245,
    input  [47:0] col_in_246,
    input  [47:0] col_in_247,
    input  [47:0] col_in_248,
    input  [47:0] col_in_249,
    input  [47:0] col_in_250,
    input  [47:0] col_in_251,
    input  [47:0] col_in_252,
    input  [47:0] col_in_253,
    input  [47:0] col_in_254,
    input  [47:0] col_in_255,
    input  [47:0] col_in_256,
    input  [47:0] col_in_257,
    input  [47:0] col_in_258,
    input  [47:0] col_in_259,
    input  [47:0] col_in_260,
    input  [47:0] col_in_261,
    input  [47:0] col_in_262,
    input  [47:0] col_in_263,
    input  [47:0] col_in_264,
    input  [47:0] col_in_265,
    input  [47:0] col_in_266,
    input  [47:0] col_in_267,
    input  [47:0] col_in_268,
    input  [47:0] col_in_269,
    input  [47:0] col_in_270,
    input  [47:0] col_in_271,
    input  [47:0] col_in_272,
    input  [47:0] col_in_273,
    input  [47:0] col_in_274,
    input  [47:0] col_in_275,
    input  [47:0] col_in_276,
    input  [47:0] col_in_277,
    input  [47:0] col_in_278,
    input  [47:0] col_in_279,
    input  [47:0] col_in_280,
    input  [47:0] col_in_281,
    input  [47:0] col_in_282,
    input  [47:0] col_in_283,
    input  [47:0] col_in_284,
    input  [47:0] col_in_285,
    input  [47:0] col_in_286,
    input  [47:0] col_in_287,
    input  [47:0] col_in_288,
    input  [47:0] col_in_289,
    input  [47:0] col_in_290,
    input  [47:0] col_in_291,
    input  [47:0] col_in_292,
    input  [47:0] col_in_293,
    input  [47:0] col_in_294,
    input  [47:0] col_in_295,
    input  [47:0] col_in_296,
    input  [47:0] col_in_297,
    input  [47:0] col_in_298,
    input  [47:0] col_in_299,
    input  [47:0] col_in_300,
    input  [47:0] col_in_301,
    input  [47:0] col_in_302,
    input  [47:0] col_in_303,
    input  [47:0] col_in_304,
    input  [47:0] col_in_305,
    input  [47:0] col_in_306,
    input  [47:0] col_in_307,
    input  [47:0] col_in_308,
    input  [47:0] col_in_309,
    input  [47:0] col_in_310,
    input  [47:0] col_in_311,
    input  [47:0] col_in_312,
    input  [47:0] col_in_313,
    input  [47:0] col_in_314,
    input  [47:0] col_in_315,
    input  [47:0] col_in_316,
    input  [47:0] col_in_317,
    input  [47:0] col_in_318,
    input  [47:0] col_in_319,
    input  [47:0] col_in_320,
    input  [47:0] col_in_321,
    input  [47:0] col_in_322,
    input  [47:0] col_in_323,
    input  [47:0] col_in_324,
    input  [47:0] col_in_325,
    input  [47:0] col_in_326,
    input  [47:0] col_in_327,
    input  [47:0] col_in_328,
    input  [47:0] col_in_329,
    input  [47:0] col_in_330,
    input  [47:0] col_in_331,
    input  [47:0] col_in_332,
    input  [47:0] col_in_333,
    input  [47:0] col_in_334,
    input  [47:0] col_in_335,
    input  [47:0] col_in_336,
    input  [47:0] col_in_337,
    input  [47:0] col_in_338,
    input  [47:0] col_in_339,
    input  [47:0] col_in_340,
    input  [47:0] col_in_341,
    input  [47:0] col_in_342,
    input  [47:0] col_in_343,
    input  [47:0] col_in_344,
    input  [47:0] col_in_345,
    input  [47:0] col_in_346,
    input  [47:0] col_in_347,
    input  [47:0] col_in_348,
    input  [47:0] col_in_349,
    input  [47:0] col_in_350,
    input  [47:0] col_in_351,
    input  [47:0] col_in_352,
    input  [47:0] col_in_353,
    input  [47:0] col_in_354,
    input  [47:0] col_in_355,
    input  [47:0] col_in_356,
    input  [47:0] col_in_357,
    input  [47:0] col_in_358,
    input  [47:0] col_in_359,
    input  [47:0] col_in_360,
    input  [47:0] col_in_361,
    input  [47:0] col_in_362,
    input  [47:0] col_in_363,
    input  [47:0] col_in_364,
    input  [47:0] col_in_365,
    input  [47:0] col_in_366,
    input  [47:0] col_in_367,
    input  [47:0] col_in_368,
    input  [47:0] col_in_369,
    input  [47:0] col_in_370,
    input  [47:0] col_in_371,
    input  [47:0] col_in_372,
    input  [47:0] col_in_373,
    input  [47:0] col_in_374,
    input  [47:0] col_in_375,
    input  [47:0] col_in_376,
    input  [47:0] col_in_377,
    input  [47:0] col_in_378,
    input  [47:0] col_in_379,
    input  [47:0] col_in_380,
    input  [47:0] col_in_381,
    input  [47:0] col_in_382,
    input  [47:0] col_in_383,
    input  [47:0] col_in_384,
    input  [47:0] col_in_385,
    input  [47:0] col_in_386,
    input  [47:0] col_in_387,
    input  [47:0] col_in_388,
    input  [47:0] col_in_389,
    input  [47:0] col_in_390,
    input  [47:0] col_in_391,
    input  [47:0] col_in_392,
    input  [47:0] col_in_393,
    input  [47:0] col_in_394,
    input  [47:0] col_in_395,
    input  [47:0] col_in_396,
    input  [47:0] col_in_397,
    input  [47:0] col_in_398,
    input  [47:0] col_in_399,
    input  [47:0] col_in_400,
    input  [47:0] col_in_401,
    input  [47:0] col_in_402,
    input  [47:0] col_in_403,
    input  [47:0] col_in_404,
    input  [47:0] col_in_405,
    input  [47:0] col_in_406,
    input  [47:0] col_in_407,
    input  [47:0] col_in_408,
    input  [47:0] col_in_409,
    input  [47:0] col_in_410,
    input  [47:0] col_in_411,
    input  [47:0] col_in_412,
    input  [47:0] col_in_413,
    input  [47:0] col_in_414,
    input  [47:0] col_in_415,
    input  [47:0] col_in_416,
    input  [47:0] col_in_417,
    input  [47:0] col_in_418,
    input  [47:0] col_in_419,
    input  [47:0] col_in_420,
    input  [47:0] col_in_421,
    input  [47:0] col_in_422,
    input  [47:0] col_in_423,
    input  [47:0] col_in_424,
    input  [47:0] col_in_425,
    input  [47:0] col_in_426,
    input  [47:0] col_in_427,
    input  [47:0] col_in_428,
    input  [47:0] col_in_429,
    input  [47:0] col_in_430,
    input  [47:0] col_in_431,
    input  [47:0] col_in_432,
    input  [47:0] col_in_433,
    input  [47:0] col_in_434,
    input  [47:0] col_in_435,
    input  [47:0] col_in_436,
    input  [47:0] col_in_437,
    input  [47:0] col_in_438,
    input  [47:0] col_in_439,
    input  [47:0] col_in_440,
    input  [47:0] col_in_441,
    input  [47:0] col_in_442,
    input  [47:0] col_in_443,
    input  [47:0] col_in_444,
    input  [47:0] col_in_445,
    input  [47:0] col_in_446,
    input  [47:0] col_in_447,
    input  [47:0] col_in_448,
    input  [47:0] col_in_449,
    input  [47:0] col_in_450,
    input  [47:0] col_in_451,
    input  [47:0] col_in_452,
    input  [47:0] col_in_453,
    input  [47:0] col_in_454,
    input  [47:0] col_in_455,
    input  [47:0] col_in_456,
    input  [47:0] col_in_457,
    input  [47:0] col_in_458,
    input  [47:0] col_in_459,
    input  [47:0] col_in_460,
    input  [47:0] col_in_461,
    input  [47:0] col_in_462,
    input  [47:0] col_in_463,
    input  [47:0] col_in_464,
    input  [47:0] col_in_465,
    input  [47:0] col_in_466,
    input  [47:0] col_in_467,
    input  [47:0] col_in_468,
    input  [47:0] col_in_469,
    input  [47:0] col_in_470,
    input  [47:0] col_in_471,
    input  [47:0] col_in_472,
    input  [47:0] col_in_473,
    input  [47:0] col_in_474,
    input  [47:0] col_in_475,
    input  [47:0] col_in_476,
    input  [47:0] col_in_477,
    input  [47:0] col_in_478,
    input  [47:0] col_in_479,
    input  [47:0] col_in_480,
    input  [47:0] col_in_481,
    input  [47:0] col_in_482,
    input  [47:0] col_in_483,
    input  [47:0] col_in_484,
    input  [47:0] col_in_485,
    input  [47:0] col_in_486,
    input  [47:0] col_in_487,
    input  [47:0] col_in_488,
    input  [47:0] col_in_489,
    input  [47:0] col_in_490,
    input  [47:0] col_in_491,
    input  [47:0] col_in_492,
    input  [47:0] col_in_493,
    input  [47:0] col_in_494,
    input  [47:0] col_in_495,
    input  [47:0] col_in_496,
    input  [47:0] col_in_497,
    input  [47:0] col_in_498,
    input  [47:0] col_in_499,
    input  [47:0] col_in_500,
    input  [47:0] col_in_501,
    input  [47:0] col_in_502,
    input  [47:0] col_in_503,
    input  [47:0] col_in_504,
    input  [47:0] col_in_505,
    input  [47:0] col_in_506,
    input  [47:0] col_in_507,
    input  [47:0] col_in_508,
    input  [47:0] col_in_509,
    input  [47:0] col_in_510,
    input  [47:0] col_in_511,
    input  [47:0] col_in_512,
    input  [47:0] col_in_513,
    input  [47:0] col_in_514,
    input  [47:0] col_in_515,
    input  [47:0] col_in_516,
    input  [47:0] col_in_517,
    input  [47:0] col_in_518,
    input  [47:0] col_in_519,
    input  [47:0] col_in_520,
    input  [47:0] col_in_521,
    input  [47:0] col_in_522,
    input  [47:0] col_in_523,
    input  [47:0] col_in_524,
    input  [47:0] col_in_525,
    input  [47:0] col_in_526,
    input  [47:0] col_in_527,
    input  [47:0] col_in_528,
    input  [47:0] col_in_529,
    input  [47:0] col_in_530,
    input  [47:0] col_in_531,
    input  [47:0] col_in_532,
    input  [47:0] col_in_533,
    input  [47:0] col_in_534,
    input  [47:0] col_in_535,
    input  [47:0] col_in_536,
    input  [47:0] col_in_537,
    input  [47:0] col_in_538,
    input  [47:0] col_in_539,
    input  [47:0] col_in_540,
    input  [47:0] col_in_541,
    input  [47:0] col_in_542,
    input  [47:0] col_in_543,
    input  [47:0] col_in_544,
    input  [47:0] col_in_545,
    input  [47:0] col_in_546,
    input  [47:0] col_in_547,
    input  [47:0] col_in_548,
    input  [47:0] col_in_549,
    input  [47:0] col_in_550,
    input  [47:0] col_in_551,
    input  [47:0] col_in_552,
    input  [47:0] col_in_553,
    input  [47:0] col_in_554,
    input  [47:0] col_in_555,
    input  [47:0] col_in_556,
    input  [47:0] col_in_557,
    input  [47:0] col_in_558,
    input  [47:0] col_in_559,
    input  [47:0] col_in_560,
    input  [47:0] col_in_561,
    input  [47:0] col_in_562,
    input  [47:0] col_in_563,
    input  [47:0] col_in_564,
    input  [47:0] col_in_565,
    input  [47:0] col_in_566,
    input  [47:0] col_in_567,
    input  [47:0] col_in_568,
    input  [47:0] col_in_569,
    input  [47:0] col_in_570,
    input  [47:0] col_in_571,
    input  [47:0] col_in_572,
    input  [47:0] col_in_573,
    input  [47:0] col_in_574,
    input  [47:0] col_in_575,
    input  [47:0] col_in_576,
    input  [47:0] col_in_577,
    input  [47:0] col_in_578,
    input  [47:0] col_in_579,
    input  [47:0] col_in_580,
    input  [47:0] col_in_581,
    input  [47:0] col_in_582,
    input  [47:0] col_in_583,
    input  [47:0] col_in_584,
    input  [47:0] col_in_585,
    input  [47:0] col_in_586,
    input  [47:0] col_in_587,
    input  [47:0] col_in_588,
    input  [47:0] col_in_589,
    input  [47:0] col_in_590,
    input  [47:0] col_in_591,
    input  [47:0] col_in_592,
    input  [47:0] col_in_593,
    input  [47:0] col_in_594,
    input  [47:0] col_in_595,
    input  [47:0] col_in_596,
    input  [47:0] col_in_597,
    input  [47:0] col_in_598,
    input  [47:0] col_in_599,
    input  [47:0] col_in_600,
    input  [47:0] col_in_601,
    input  [47:0] col_in_602,
    input  [47:0] col_in_603,
    input  [47:0] col_in_604,
    input  [47:0] col_in_605,
    input  [47:0] col_in_606,
    input  [47:0] col_in_607,
    input  [47:0] col_in_608,
    input  [47:0] col_in_609,
    input  [47:0] col_in_610,
    input  [47:0] col_in_611,
    input  [47:0] col_in_612,
    input  [47:0] col_in_613,
    input  [47:0] col_in_614,
    input  [47:0] col_in_615,
    input  [47:0] col_in_616,
    input  [47:0] col_in_617,
    input  [47:0] col_in_618,
    input  [47:0] col_in_619,
    input  [47:0] col_in_620,
    input  [47:0] col_in_621,
    input  [47:0] col_in_622,
    input  [47:0] col_in_623,
    input  [47:0] col_in_624,
    input  [47:0] col_in_625,
    input  [47:0] col_in_626,
    input  [47:0] col_in_627,
    input  [47:0] col_in_628,
    input  [47:0] col_in_629,
    input  [47:0] col_in_630,
    input  [47:0] col_in_631,
    input  [47:0] col_in_632,
    input  [47:0] col_in_633,
    input  [47:0] col_in_634,
    input  [47:0] col_in_635,
    input  [47:0] col_in_636,
    input  [47:0] col_in_637,
    input  [47:0] col_in_638,
    input  [47:0] col_in_639,
    input  [47:0] col_in_640,
    input  [47:0] col_in_641,
    input  [47:0] col_in_642,
    input  [47:0] col_in_643,
    input  [47:0] col_in_644,
    input  [47:0] col_in_645,
    input  [47:0] col_in_646,
    input  [47:0] col_in_647,
    input  [47:0] col_in_648,
    input  [47:0] col_in_649,
    input  [47:0] col_in_650,
    input  [47:0] col_in_651,
    input  [47:0] col_in_652,
    input  [47:0] col_in_653,
    input  [47:0] col_in_654,
    input  [47:0] col_in_655,
    input  [47:0] col_in_656,
    input  [47:0] col_in_657,
    input  [47:0] col_in_658,
    input  [47:0] col_in_659,
    input  [47:0] col_in_660,
    input  [47:0] col_in_661,
    input  [47:0] col_in_662,
    input  [47:0] col_in_663,
    input  [47:0] col_in_664,
    input  [47:0] col_in_665,
    input  [47:0] col_in_666,
    input  [47:0] col_in_667,
    input  [47:0] col_in_668,
    input  [47:0] col_in_669,
    input  [47:0] col_in_670,
    input  [47:0] col_in_671,
    input  [47:0] col_in_672,
    input  [47:0] col_in_673,
    input  [47:0] col_in_674,
    input  [47:0] col_in_675,
    input  [47:0] col_in_676,
    input  [47:0] col_in_677,
    input  [47:0] col_in_678,
    input  [47:0] col_in_679,
    input  [47:0] col_in_680,
    input  [47:0] col_in_681,
    input  [47:0] col_in_682,
    input  [47:0] col_in_683,
    input  [47:0] col_in_684,
    input  [47:0] col_in_685,
    input  [47:0] col_in_686,
    input  [47:0] col_in_687,
    input  [47:0] col_in_688,
    input  [47:0] col_in_689,
    input  [47:0] col_in_690,
    input  [47:0] col_in_691,
    input  [47:0] col_in_692,
    input  [47:0] col_in_693,
    input  [47:0] col_in_694,
    input  [47:0] col_in_695,
    input  [47:0] col_in_696,
    input  [47:0] col_in_697,
    input  [47:0] col_in_698,
    input  [47:0] col_in_699,
    input  [47:0] col_in_700,
    input  [47:0] col_in_701,
    input  [47:0] col_in_702,
    input  [47:0] col_in_703,
    input  [47:0] col_in_704,
    input  [47:0] col_in_705,
    input  [47:0] col_in_706,
    input  [47:0] col_in_707,
    input  [47:0] col_in_708,
    input  [47:0] col_in_709,
    input  [47:0] col_in_710,
    input  [47:0] col_in_711,
    input  [47:0] col_in_712,
    input  [47:0] col_in_713,
    input  [47:0] col_in_714,
    input  [47:0] col_in_715,
    input  [47:0] col_in_716,
    input  [47:0] col_in_717,
    input  [47:0] col_in_718,
    input  [47:0] col_in_719,
    input  [47:0] col_in_720,
    input  [47:0] col_in_721,
    input  [47:0] col_in_722,
    input  [47:0] col_in_723,
    input  [47:0] col_in_724,
    input  [47:0] col_in_725,
    input  [47:0] col_in_726,
    input  [47:0] col_in_727,
    input  [47:0] col_in_728,
    input  [47:0] col_in_729,
    input  [47:0] col_in_730,
    input  [47:0] col_in_731,
    input  [47:0] col_in_732,
    input  [47:0] col_in_733,
    input  [47:0] col_in_734,
    input  [47:0] col_in_735,
    input  [47:0] col_in_736,
    input  [47:0] col_in_737,
    input  [47:0] col_in_738,
    input  [47:0] col_in_739,
    input  [47:0] col_in_740,
    input  [47:0] col_in_741,
    input  [47:0] col_in_742,
    input  [47:0] col_in_743,
    input  [47:0] col_in_744,
    input  [47:0] col_in_745,
    input  [47:0] col_in_746,
    input  [47:0] col_in_747,
    input  [47:0] col_in_748,
    input  [47:0] col_in_749,
    input  [47:0] col_in_750,
    input  [47:0] col_in_751,
    input  [47:0] col_in_752,
    input  [47:0] col_in_753,
    input  [47:0] col_in_754,
    input  [47:0] col_in_755,
    input  [47:0] col_in_756,
    input  [47:0] col_in_757,
    input  [47:0] col_in_758,
    input  [47:0] col_in_759,
    input  [47:0] col_in_760,
    input  [47:0] col_in_761,
    input  [47:0] col_in_762,
    input  [47:0] col_in_763,
    input  [47:0] col_in_764,
    input  [47:0] col_in_765,
    input  [47:0] col_in_766,
    input  [47:0] col_in_767,
    input  [47:0] col_in_768,
    input  [47:0] col_in_769,
    input  [47:0] col_in_770,
    input  [47:0] col_in_771,
    input  [47:0] col_in_772,
    input  [47:0] col_in_773,
    input  [47:0] col_in_774,
    input  [47:0] col_in_775,
    input  [47:0] col_in_776,
    input  [47:0] col_in_777,
    input  [47:0] col_in_778,
    input  [47:0] col_in_779,
    input  [47:0] col_in_780,
    input  [47:0] col_in_781,
    input  [47:0] col_in_782,
    input  [47:0] col_in_783,
    input  [47:0] col_in_784,
    input  [47:0] col_in_785,
    input  [47:0] col_in_786,
    input  [47:0] col_in_787,
    input  [47:0] col_in_788,
    input  [47:0] col_in_789,
    input  [47:0] col_in_790,
    input  [47:0] col_in_791,
    input  [47:0] col_in_792,
    input  [47:0] col_in_793,
    input  [47:0] col_in_794,
    input  [47:0] col_in_795,
    input  [47:0] col_in_796,
    input  [47:0] col_in_797,
    input  [47:0] col_in_798,
    input  [47:0] col_in_799,
    input  [47:0] col_in_800,
    input  [47:0] col_in_801,
    input  [47:0] col_in_802,
    input  [47:0] col_in_803,
    input  [47:0] col_in_804,
    input  [47:0] col_in_805,
    input  [47:0] col_in_806,
    input  [47:0] col_in_807,
    input  [47:0] col_in_808,
    input  [47:0] col_in_809,
    input  [47:0] col_in_810,
    input  [47:0] col_in_811,
    input  [47:0] col_in_812,
    input  [47:0] col_in_813,
    input  [47:0] col_in_814,
    input  [47:0] col_in_815,
    input  [47:0] col_in_816,
    input  [47:0] col_in_817,
    input  [47:0] col_in_818,
    input  [47:0] col_in_819,
    input  [47:0] col_in_820,
    input  [47:0] col_in_821,
    input  [47:0] col_in_822,
    input  [47:0] col_in_823,
    input  [47:0] col_in_824,
    input  [47:0] col_in_825,
    input  [47:0] col_in_826,
    input  [47:0] col_in_827,
    input  [47:0] col_in_828,
    input  [47:0] col_in_829,
    input  [47:0] col_in_830,
    input  [47:0] col_in_831,
    input  [47:0] col_in_832,
    input  [47:0] col_in_833,
    input  [47:0] col_in_834,
    input  [47:0] col_in_835,
    input  [47:0] col_in_836,
    input  [47:0] col_in_837,
    input  [47:0] col_in_838,
    input  [47:0] col_in_839,
    input  [47:0] col_in_840,
    input  [47:0] col_in_841,
    input  [47:0] col_in_842,
    input  [47:0] col_in_843,
    input  [47:0] col_in_844,
    input  [47:0] col_in_845,
    input  [47:0] col_in_846,
    input  [47:0] col_in_847,
    input  [47:0] col_in_848,
    input  [47:0] col_in_849,
    input  [47:0] col_in_850,
    input  [47:0] col_in_851,
    input  [47:0] col_in_852,
    input  [47:0] col_in_853,
    input  [47:0] col_in_854,
    input  [47:0] col_in_855,
    input  [47:0] col_in_856,
    input  [47:0] col_in_857,
    input  [47:0] col_in_858,
    input  [47:0] col_in_859,
    input  [47:0] col_in_860,
    input  [47:0] col_in_861,
    input  [47:0] col_in_862,
    input  [47:0] col_in_863,
    input  [47:0] col_in_864,
    input  [47:0] col_in_865,
    input  [47:0] col_in_866,
    input  [47:0] col_in_867,
    input  [47:0] col_in_868,
    input  [47:0] col_in_869,
    input  [47:0] col_in_870,
    input  [47:0] col_in_871,
    input  [47:0] col_in_872,
    input  [47:0] col_in_873,
    input  [47:0] col_in_874,
    input  [47:0] col_in_875,
    input  [47:0] col_in_876,
    input  [47:0] col_in_877,
    input  [47:0] col_in_878,
    input  [47:0] col_in_879,
    input  [47:0] col_in_880,
    input  [47:0] col_in_881,
    input  [47:0] col_in_882,
    input  [47:0] col_in_883,
    input  [47:0] col_in_884,
    input  [47:0] col_in_885,
    input  [47:0] col_in_886,
    input  [47:0] col_in_887,
    input  [47:0] col_in_888,
    input  [47:0] col_in_889,
    input  [47:0] col_in_890,
    input  [47:0] col_in_891,
    input  [47:0] col_in_892,
    input  [47:0] col_in_893,
    input  [47:0] col_in_894,
    input  [47:0] col_in_895,
    input  [47:0] col_in_896,
    input  [47:0] col_in_897,
    input  [47:0] col_in_898,
    input  [47:0] col_in_899,
    input  [47:0] col_in_900,
    input  [47:0] col_in_901,
    input  [47:0] col_in_902,
    input  [47:0] col_in_903,
    input  [47:0] col_in_904,
    input  [47:0] col_in_905,
    input  [47:0] col_in_906,
    input  [47:0] col_in_907,
    input  [47:0] col_in_908,
    input  [47:0] col_in_909,
    input  [47:0] col_in_910,
    input  [47:0] col_in_911,
    input  [47:0] col_in_912,
    input  [47:0] col_in_913,
    input  [47:0] col_in_914,
    input  [47:0] col_in_915,
    input  [47:0] col_in_916,
    input  [47:0] col_in_917,
    input  [47:0] col_in_918,
    input  [47:0] col_in_919,
    input  [47:0] col_in_920,
    input  [47:0] col_in_921,
    input  [47:0] col_in_922,
    input  [47:0] col_in_923,
    input  [47:0] col_in_924,
    input  [47:0] col_in_925,
    input  [47:0] col_in_926,
    input  [47:0] col_in_927,
    input  [47:0] col_in_928,
    input  [47:0] col_in_929,
    input  [47:0] col_in_930,
    input  [47:0] col_in_931,
    input  [47:0] col_in_932,
    input  [47:0] col_in_933,
    input  [47:0] col_in_934,
    input  [47:0] col_in_935,
    input  [47:0] col_in_936,
    input  [47:0] col_in_937,
    input  [47:0] col_in_938,
    input  [47:0] col_in_939,
    input  [47:0] col_in_940,
    input  [47:0] col_in_941,
    input  [47:0] col_in_942,
    input  [47:0] col_in_943,
    input  [47:0] col_in_944,
    input  [47:0] col_in_945,
    input  [47:0] col_in_946,
    input  [47:0] col_in_947,
    input  [47:0] col_in_948,
    input  [47:0] col_in_949,
    input  [47:0] col_in_950,
    input  [47:0] col_in_951,
    input  [47:0] col_in_952,
    input  [47:0] col_in_953,
    input  [47:0] col_in_954,
    input  [47:0] col_in_955,
    input  [47:0] col_in_956,
    input  [47:0] col_in_957,
    input  [47:0] col_in_958,
    input  [47:0] col_in_959,
    input  [47:0] col_in_960,
    input  [47:0] col_in_961,
    input  [47:0] col_in_962,
    input  [47:0] col_in_963,
    input  [47:0] col_in_964,
    input  [47:0] col_in_965,
    input  [47:0] col_in_966,
    input  [47:0] col_in_967,
    input  [47:0] col_in_968,
    input  [47:0] col_in_969,
    input  [47:0] col_in_970,
    input  [47:0] col_in_971,
    input  [47:0] col_in_972,
    input  [47:0] col_in_973,
    input  [47:0] col_in_974,
    input  [47:0] col_in_975,
    input  [47:0] col_in_976,
    input  [47:0] col_in_977,
    input  [47:0] col_in_978,
    input  [47:0] col_in_979,
    input  [47:0] col_in_980,
    input  [47:0] col_in_981,
    input  [47:0] col_in_982,
    input  [47:0] col_in_983,
    input  [47:0] col_in_984,
    input  [47:0] col_in_985,
    input  [47:0] col_in_986,
    input  [47:0] col_in_987,
    input  [47:0] col_in_988,
    input  [47:0] col_in_989,
    input  [47:0] col_in_990,
    input  [47:0] col_in_991,
    input  [47:0] col_in_992,
    input  [47:0] col_in_993,
    input  [47:0] col_in_994,
    input  [47:0] col_in_995,
    input  [47:0] col_in_996,
    input  [47:0] col_in_997,
    input  [47:0] col_in_998,
    input  [47:0] col_in_999,
    input  [47:0] col_in_1000,
    input  [47:0] col_in_1001,
    input  [47:0] col_in_1002,
    input  [47:0] col_in_1003,
    input  [47:0] col_in_1004,
    input  [47:0] col_in_1005,
    input  [47:0] col_in_1006,
    input  [47:0] col_in_1007,
    input  [47:0] col_in_1008,
    input  [47:0] col_in_1009,
    input  [47:0] col_in_1010,
    input  [47:0] col_in_1011,
    input  [47:0] col_in_1012,
    input  [47:0] col_in_1013,
    input  [47:0] col_in_1014,
    input  [47:0] col_in_1015,
    input  [47:0] col_in_1016,
    input  [47:0] col_in_1017,
    input  [47:0] col_in_1018,
    input  [47:0] col_in_1019,
    input  [47:0] col_in_1020,
    input  [47:0] col_in_1021,
    input  [47:0] col_in_1022,
    input  [47:0] col_in_1023,
    input  [47:0] col_in_1024,
    input  [47:0] col_in_1025,
    input  [47:0] col_in_1026,
    input  [47:0] col_in_1027,
    input  [47:0] col_in_1028,
    input  [47:0] col_in_1029,

    output [15:0] col_out_0,
    output [15:0] col_out_1,
    output [15:0] col_out_2,
    output [15:0] col_out_3,
    output [15:0] col_out_4,
    output [15:0] col_out_5,
    output [15:0] col_out_6,
    output [15:0] col_out_7,
    output [15:0] col_out_8,
    output [15:0] col_out_9,
    output [15:0] col_out_10,
    output [15:0] col_out_11,
    output [15:0] col_out_12,
    output [15:0] col_out_13,
    output [15:0] col_out_14,
    output [15:0] col_out_15,
    output [15:0] col_out_16,
    output [15:0] col_out_17,
    output [15:0] col_out_18,
    output [15:0] col_out_19,
    output [15:0] col_out_20,
    output [15:0] col_out_21,
    output [15:0] col_out_22,
    output [15:0] col_out_23,
    output [15:0] col_out_24,
    output [15:0] col_out_25,
    output [15:0] col_out_26,
    output [15:0] col_out_27,
    output [15:0] col_out_28,
    output [15:0] col_out_29,
    output [15:0] col_out_30,
    output [15:0] col_out_31,
    output [15:0] col_out_32,
    output [15:0] col_out_33,
    output [15:0] col_out_34,
    output [15:0] col_out_35,
    output [15:0] col_out_36,
    output [15:0] col_out_37,
    output [15:0] col_out_38,
    output [15:0] col_out_39,
    output [15:0] col_out_40,
    output [15:0] col_out_41,
    output [15:0] col_out_42,
    output [15:0] col_out_43,
    output [15:0] col_out_44,
    output [15:0] col_out_45,
    output [15:0] col_out_46,
    output [15:0] col_out_47,
    output [15:0] col_out_48,
    output [15:0] col_out_49,
    output [15:0] col_out_50,
    output [15:0] col_out_51,
    output [15:0] col_out_52,
    output [15:0] col_out_53,
    output [15:0] col_out_54,
    output [15:0] col_out_55,
    output [15:0] col_out_56,
    output [15:0] col_out_57,
    output [15:0] col_out_58,
    output [15:0] col_out_59,
    output [15:0] col_out_60,
    output [15:0] col_out_61,
    output [15:0] col_out_62,
    output [15:0] col_out_63,
    output [15:0] col_out_64,
    output [15:0] col_out_65,
    output [15:0] col_out_66,
    output [15:0] col_out_67,
    output [15:0] col_out_68,
    output [15:0] col_out_69,
    output [15:0] col_out_70,
    output [15:0] col_out_71,
    output [15:0] col_out_72,
    output [15:0] col_out_73,
    output [15:0] col_out_74,
    output [15:0] col_out_75,
    output [15:0] col_out_76,
    output [15:0] col_out_77,
    output [15:0] col_out_78,
    output [15:0] col_out_79,
    output [15:0] col_out_80,
    output [15:0] col_out_81,
    output [15:0] col_out_82,
    output [15:0] col_out_83,
    output [15:0] col_out_84,
    output [15:0] col_out_85,
    output [15:0] col_out_86,
    output [15:0] col_out_87,
    output [15:0] col_out_88,
    output [15:0] col_out_89,
    output [15:0] col_out_90,
    output [15:0] col_out_91,
    output [15:0] col_out_92,
    output [15:0] col_out_93,
    output [15:0] col_out_94,
    output [15:0] col_out_95,
    output [15:0] col_out_96,
    output [15:0] col_out_97,
    output [15:0] col_out_98,
    output [15:0] col_out_99,
    output [15:0] col_out_100,
    output [15:0] col_out_101,
    output [15:0] col_out_102,
    output [15:0] col_out_103,
    output [15:0] col_out_104,
    output [15:0] col_out_105,
    output [15:0] col_out_106,
    output [15:0] col_out_107,
    output [15:0] col_out_108,
    output [15:0] col_out_109,
    output [15:0] col_out_110,
    output [15:0] col_out_111,
    output [15:0] col_out_112,
    output [15:0] col_out_113,
    output [15:0] col_out_114,
    output [15:0] col_out_115,
    output [15:0] col_out_116,
    output [15:0] col_out_117,
    output [15:0] col_out_118,
    output [15:0] col_out_119,
    output [15:0] col_out_120,
    output [15:0] col_out_121,
    output [15:0] col_out_122,
    output [15:0] col_out_123,
    output [15:0] col_out_124,
    output [15:0] col_out_125,
    output [15:0] col_out_126,
    output [15:0] col_out_127,
    output [15:0] col_out_128,
    output [15:0] col_out_129,
    output [15:0] col_out_130,
    output [15:0] col_out_131,
    output [15:0] col_out_132,
    output [15:0] col_out_133,
    output [15:0] col_out_134,
    output [15:0] col_out_135,
    output [15:0] col_out_136,
    output [15:0] col_out_137,
    output [15:0] col_out_138,
    output [15:0] col_out_139,
    output [15:0] col_out_140,
    output [15:0] col_out_141,
    output [15:0] col_out_142,
    output [15:0] col_out_143,
    output [15:0] col_out_144,
    output [15:0] col_out_145,
    output [15:0] col_out_146,
    output [15:0] col_out_147,
    output [15:0] col_out_148,
    output [15:0] col_out_149,
    output [15:0] col_out_150,
    output [15:0] col_out_151,
    output [15:0] col_out_152,
    output [15:0] col_out_153,
    output [15:0] col_out_154,
    output [15:0] col_out_155,
    output [15:0] col_out_156,
    output [15:0] col_out_157,
    output [15:0] col_out_158,
    output [15:0] col_out_159,
    output [15:0] col_out_160,
    output [15:0] col_out_161,
    output [15:0] col_out_162,
    output [15:0] col_out_163,
    output [15:0] col_out_164,
    output [15:0] col_out_165,
    output [15:0] col_out_166,
    output [15:0] col_out_167,
    output [15:0] col_out_168,
    output [15:0] col_out_169,
    output [15:0] col_out_170,
    output [15:0] col_out_171,
    output [15:0] col_out_172,
    output [15:0] col_out_173,
    output [15:0] col_out_174,
    output [15:0] col_out_175,
    output [15:0] col_out_176,
    output [15:0] col_out_177,
    output [15:0] col_out_178,
    output [15:0] col_out_179,
    output [15:0] col_out_180,
    output [15:0] col_out_181,
    output [15:0] col_out_182,
    output [15:0] col_out_183,
    output [15:0] col_out_184,
    output [15:0] col_out_185,
    output [15:0] col_out_186,
    output [15:0] col_out_187,
    output [15:0] col_out_188,
    output [15:0] col_out_189,
    output [15:0] col_out_190,
    output [15:0] col_out_191,
    output [15:0] col_out_192,
    output [15:0] col_out_193,
    output [15:0] col_out_194,
    output [15:0] col_out_195,
    output [15:0] col_out_196,
    output [15:0] col_out_197,
    output [15:0] col_out_198,
    output [15:0] col_out_199,
    output [15:0] col_out_200,
    output [15:0] col_out_201,
    output [15:0] col_out_202,
    output [15:0] col_out_203,
    output [15:0] col_out_204,
    output [15:0] col_out_205,
    output [15:0] col_out_206,
    output [15:0] col_out_207,
    output [15:0] col_out_208,
    output [15:0] col_out_209,
    output [15:0] col_out_210,
    output [15:0] col_out_211,
    output [15:0] col_out_212,
    output [15:0] col_out_213,
    output [15:0] col_out_214,
    output [15:0] col_out_215,
    output [15:0] col_out_216,
    output [15:0] col_out_217,
    output [15:0] col_out_218,
    output [15:0] col_out_219,
    output [15:0] col_out_220,
    output [15:0] col_out_221,
    output [15:0] col_out_222,
    output [15:0] col_out_223,
    output [15:0] col_out_224,
    output [15:0] col_out_225,
    output [15:0] col_out_226,
    output [15:0] col_out_227,
    output [15:0] col_out_228,
    output [15:0] col_out_229,
    output [15:0] col_out_230,
    output [15:0] col_out_231,
    output [15:0] col_out_232,
    output [15:0] col_out_233,
    output [15:0] col_out_234,
    output [15:0] col_out_235,
    output [15:0] col_out_236,
    output [15:0] col_out_237,
    output [15:0] col_out_238,
    output [15:0] col_out_239,
    output [15:0] col_out_240,
    output [15:0] col_out_241,
    output [15:0] col_out_242,
    output [15:0] col_out_243,
    output [15:0] col_out_244,
    output [15:0] col_out_245,
    output [15:0] col_out_246,
    output [15:0] col_out_247,
    output [15:0] col_out_248,
    output [15:0] col_out_249,
    output [15:0] col_out_250,
    output [15:0] col_out_251,
    output [15:0] col_out_252,
    output [15:0] col_out_253,
    output [15:0] col_out_254,
    output [15:0] col_out_255,
    output [15:0] col_out_256,
    output [15:0] col_out_257,
    output [15:0] col_out_258,
    output [15:0] col_out_259,
    output [15:0] col_out_260,
    output [15:0] col_out_261,
    output [15:0] col_out_262,
    output [15:0] col_out_263,
    output [15:0] col_out_264,
    output [15:0] col_out_265,
    output [15:0] col_out_266,
    output [15:0] col_out_267,
    output [15:0] col_out_268,
    output [15:0] col_out_269,
    output [15:0] col_out_270,
    output [15:0] col_out_271,
    output [15:0] col_out_272,
    output [15:0] col_out_273,
    output [15:0] col_out_274,
    output [15:0] col_out_275,
    output [15:0] col_out_276,
    output [15:0] col_out_277,
    output [15:0] col_out_278,
    output [15:0] col_out_279,
    output [15:0] col_out_280,
    output [15:0] col_out_281,
    output [15:0] col_out_282,
    output [15:0] col_out_283,
    output [15:0] col_out_284,
    output [15:0] col_out_285,
    output [15:0] col_out_286,
    output [15:0] col_out_287,
    output [15:0] col_out_288,
    output [15:0] col_out_289,
    output [15:0] col_out_290,
    output [15:0] col_out_291,
    output [15:0] col_out_292,
    output [15:0] col_out_293,
    output [15:0] col_out_294,
    output [15:0] col_out_295,
    output [15:0] col_out_296,
    output [15:0] col_out_297,
    output [15:0] col_out_298,
    output [15:0] col_out_299,
    output [15:0] col_out_300,
    output [15:0] col_out_301,
    output [15:0] col_out_302,
    output [15:0] col_out_303,
    output [15:0] col_out_304,
    output [15:0] col_out_305,
    output [15:0] col_out_306,
    output [15:0] col_out_307,
    output [15:0] col_out_308,
    output [15:0] col_out_309,
    output [15:0] col_out_310,
    output [15:0] col_out_311,
    output [15:0] col_out_312,
    output [15:0] col_out_313,
    output [15:0] col_out_314,
    output [15:0] col_out_315,
    output [15:0] col_out_316,
    output [15:0] col_out_317,
    output [15:0] col_out_318,
    output [15:0] col_out_319,
    output [15:0] col_out_320,
    output [15:0] col_out_321,
    output [15:0] col_out_322,
    output [15:0] col_out_323,
    output [15:0] col_out_324,
    output [15:0] col_out_325,
    output [15:0] col_out_326,
    output [15:0] col_out_327,
    output [15:0] col_out_328,
    output [15:0] col_out_329,
    output [15:0] col_out_330,
    output [15:0] col_out_331,
    output [15:0] col_out_332,
    output [15:0] col_out_333,
    output [15:0] col_out_334,
    output [15:0] col_out_335,
    output [15:0] col_out_336,
    output [15:0] col_out_337,
    output [15:0] col_out_338,
    output [15:0] col_out_339,
    output [15:0] col_out_340,
    output [15:0] col_out_341,
    output [15:0] col_out_342,
    output [15:0] col_out_343,
    output [15:0] col_out_344,
    output [15:0] col_out_345,
    output [15:0] col_out_346,
    output [15:0] col_out_347,
    output [15:0] col_out_348,
    output [15:0] col_out_349,
    output [15:0] col_out_350,
    output [15:0] col_out_351,
    output [15:0] col_out_352,
    output [15:0] col_out_353,
    output [15:0] col_out_354,
    output [15:0] col_out_355,
    output [15:0] col_out_356,
    output [15:0] col_out_357,
    output [15:0] col_out_358,
    output [15:0] col_out_359,
    output [15:0] col_out_360,
    output [15:0] col_out_361,
    output [15:0] col_out_362,
    output [15:0] col_out_363,
    output [15:0] col_out_364,
    output [15:0] col_out_365,
    output [15:0] col_out_366,
    output [15:0] col_out_367,
    output [15:0] col_out_368,
    output [15:0] col_out_369,
    output [15:0] col_out_370,
    output [15:0] col_out_371,
    output [15:0] col_out_372,
    output [15:0] col_out_373,
    output [15:0] col_out_374,
    output [15:0] col_out_375,
    output [15:0] col_out_376,
    output [15:0] col_out_377,
    output [15:0] col_out_378,
    output [15:0] col_out_379,
    output [15:0] col_out_380,
    output [15:0] col_out_381,
    output [15:0] col_out_382,
    output [15:0] col_out_383,
    output [15:0] col_out_384,
    output [15:0] col_out_385,
    output [15:0] col_out_386,
    output [15:0] col_out_387,
    output [15:0] col_out_388,
    output [15:0] col_out_389,
    output [15:0] col_out_390,
    output [15:0] col_out_391,
    output [15:0] col_out_392,
    output [15:0] col_out_393,
    output [15:0] col_out_394,
    output [15:0] col_out_395,
    output [15:0] col_out_396,
    output [15:0] col_out_397,
    output [15:0] col_out_398,
    output [15:0] col_out_399,
    output [15:0] col_out_400,
    output [15:0] col_out_401,
    output [15:0] col_out_402,
    output [15:0] col_out_403,
    output [15:0] col_out_404,
    output [15:0] col_out_405,
    output [15:0] col_out_406,
    output [15:0] col_out_407,
    output [15:0] col_out_408,
    output [15:0] col_out_409,
    output [15:0] col_out_410,
    output [15:0] col_out_411,
    output [15:0] col_out_412,
    output [15:0] col_out_413,
    output [15:0] col_out_414,
    output [15:0] col_out_415,
    output [15:0] col_out_416,
    output [15:0] col_out_417,
    output [15:0] col_out_418,
    output [15:0] col_out_419,
    output [15:0] col_out_420,
    output [15:0] col_out_421,
    output [15:0] col_out_422,
    output [15:0] col_out_423,
    output [15:0] col_out_424,
    output [15:0] col_out_425,
    output [15:0] col_out_426,
    output [15:0] col_out_427,
    output [15:0] col_out_428,
    output [15:0] col_out_429,
    output [15:0] col_out_430,
    output [15:0] col_out_431,
    output [15:0] col_out_432,
    output [15:0] col_out_433,
    output [15:0] col_out_434,
    output [15:0] col_out_435,
    output [15:0] col_out_436,
    output [15:0] col_out_437,
    output [15:0] col_out_438,
    output [15:0] col_out_439,
    output [15:0] col_out_440,
    output [15:0] col_out_441,
    output [15:0] col_out_442,
    output [15:0] col_out_443,
    output [15:0] col_out_444,
    output [15:0] col_out_445,
    output [15:0] col_out_446,
    output [15:0] col_out_447,
    output [15:0] col_out_448,
    output [15:0] col_out_449,
    output [15:0] col_out_450,
    output [15:0] col_out_451,
    output [15:0] col_out_452,
    output [15:0] col_out_453,
    output [15:0] col_out_454,
    output [15:0] col_out_455,
    output [15:0] col_out_456,
    output [15:0] col_out_457,
    output [15:0] col_out_458,
    output [15:0] col_out_459,
    output [15:0] col_out_460,
    output [15:0] col_out_461,
    output [15:0] col_out_462,
    output [15:0] col_out_463,
    output [15:0] col_out_464,
    output [15:0] col_out_465,
    output [15:0] col_out_466,
    output [15:0] col_out_467,
    output [15:0] col_out_468,
    output [15:0] col_out_469,
    output [15:0] col_out_470,
    output [15:0] col_out_471,
    output [15:0] col_out_472,
    output [15:0] col_out_473,
    output [15:0] col_out_474,
    output [15:0] col_out_475,
    output [15:0] col_out_476,
    output [15:0] col_out_477,
    output [15:0] col_out_478,
    output [15:0] col_out_479,
    output [15:0] col_out_480,
    output [15:0] col_out_481,
    output [15:0] col_out_482,
    output [15:0] col_out_483,
    output [15:0] col_out_484,
    output [15:0] col_out_485,
    output [15:0] col_out_486,
    output [15:0] col_out_487,
    output [15:0] col_out_488,
    output [15:0] col_out_489,
    output [15:0] col_out_490,
    output [15:0] col_out_491,
    output [15:0] col_out_492,
    output [15:0] col_out_493,
    output [15:0] col_out_494,
    output [15:0] col_out_495,
    output [15:0] col_out_496,
    output [15:0] col_out_497,
    output [15:0] col_out_498,
    output [15:0] col_out_499,
    output [15:0] col_out_500,
    output [15:0] col_out_501,
    output [15:0] col_out_502,
    output [15:0] col_out_503,
    output [15:0] col_out_504,
    output [15:0] col_out_505,
    output [15:0] col_out_506,
    output [15:0] col_out_507,
    output [15:0] col_out_508,
    output [15:0] col_out_509,
    output [15:0] col_out_510,
    output [15:0] col_out_511,
    output [15:0] col_out_512,
    output [15:0] col_out_513,
    output [15:0] col_out_514,
    output [15:0] col_out_515,
    output [15:0] col_out_516,
    output [15:0] col_out_517,
    output [15:0] col_out_518,
    output [15:0] col_out_519,
    output [15:0] col_out_520,
    output [15:0] col_out_521,
    output [15:0] col_out_522,
    output [15:0] col_out_523,
    output [15:0] col_out_524,
    output [15:0] col_out_525,
    output [15:0] col_out_526,
    output [15:0] col_out_527,
    output [15:0] col_out_528,
    output [15:0] col_out_529,
    output [15:0] col_out_530,
    output [15:0] col_out_531,
    output [15:0] col_out_532,
    output [15:0] col_out_533,
    output [15:0] col_out_534,
    output [15:0] col_out_535,
    output [15:0] col_out_536,
    output [15:0] col_out_537,
    output [15:0] col_out_538,
    output [15:0] col_out_539,
    output [15:0] col_out_540,
    output [15:0] col_out_541,
    output [15:0] col_out_542,
    output [15:0] col_out_543,
    output [15:0] col_out_544,
    output [15:0] col_out_545,
    output [15:0] col_out_546,
    output [15:0] col_out_547,
    output [15:0] col_out_548,
    output [15:0] col_out_549,
    output [15:0] col_out_550,
    output [15:0] col_out_551,
    output [15:0] col_out_552,
    output [15:0] col_out_553,
    output [15:0] col_out_554,
    output [15:0] col_out_555,
    output [15:0] col_out_556,
    output [15:0] col_out_557,
    output [15:0] col_out_558,
    output [15:0] col_out_559,
    output [15:0] col_out_560,
    output [15:0] col_out_561,
    output [15:0] col_out_562,
    output [15:0] col_out_563,
    output [15:0] col_out_564,
    output [15:0] col_out_565,
    output [15:0] col_out_566,
    output [15:0] col_out_567,
    output [15:0] col_out_568,
    output [15:0] col_out_569,
    output [15:0] col_out_570,
    output [15:0] col_out_571,
    output [15:0] col_out_572,
    output [15:0] col_out_573,
    output [15:0] col_out_574,
    output [15:0] col_out_575,
    output [15:0] col_out_576,
    output [15:0] col_out_577,
    output [15:0] col_out_578,
    output [15:0] col_out_579,
    output [15:0] col_out_580,
    output [15:0] col_out_581,
    output [15:0] col_out_582,
    output [15:0] col_out_583,
    output [15:0] col_out_584,
    output [15:0] col_out_585,
    output [15:0] col_out_586,
    output [15:0] col_out_587,
    output [15:0] col_out_588,
    output [15:0] col_out_589,
    output [15:0] col_out_590,
    output [15:0] col_out_591,
    output [15:0] col_out_592,
    output [15:0] col_out_593,
    output [15:0] col_out_594,
    output [15:0] col_out_595,
    output [15:0] col_out_596,
    output [15:0] col_out_597,
    output [15:0] col_out_598,
    output [15:0] col_out_599,
    output [15:0] col_out_600,
    output [15:0] col_out_601,
    output [15:0] col_out_602,
    output [15:0] col_out_603,
    output [15:0] col_out_604,
    output [15:0] col_out_605,
    output [15:0] col_out_606,
    output [15:0] col_out_607,
    output [15:0] col_out_608,
    output [15:0] col_out_609,
    output [15:0] col_out_610,
    output [15:0] col_out_611,
    output [15:0] col_out_612,
    output [15:0] col_out_613,
    output [15:0] col_out_614,
    output [15:0] col_out_615,
    output [15:0] col_out_616,
    output [15:0] col_out_617,
    output [15:0] col_out_618,
    output [15:0] col_out_619,
    output [15:0] col_out_620,
    output [15:0] col_out_621,
    output [15:0] col_out_622,
    output [15:0] col_out_623,
    output [15:0] col_out_624,
    output [15:0] col_out_625,
    output [15:0] col_out_626,
    output [15:0] col_out_627,
    output [15:0] col_out_628,
    output [15:0] col_out_629,
    output [15:0] col_out_630,
    output [15:0] col_out_631,
    output [15:0] col_out_632,
    output [15:0] col_out_633,
    output [15:0] col_out_634,
    output [15:0] col_out_635,
    output [15:0] col_out_636,
    output [15:0] col_out_637,
    output [15:0] col_out_638,
    output [15:0] col_out_639,
    output [15:0] col_out_640,
    output [15:0] col_out_641,
    output [15:0] col_out_642,
    output [15:0] col_out_643,
    output [15:0] col_out_644,
    output [15:0] col_out_645,
    output [15:0] col_out_646,
    output [15:0] col_out_647,
    output [15:0] col_out_648,
    output [15:0] col_out_649,
    output [15:0] col_out_650,
    output [15:0] col_out_651,
    output [15:0] col_out_652,
    output [15:0] col_out_653,
    output [15:0] col_out_654,
    output [15:0] col_out_655,
    output [15:0] col_out_656,
    output [15:0] col_out_657,
    output [15:0] col_out_658,
    output [15:0] col_out_659,
    output [15:0] col_out_660,
    output [15:0] col_out_661,
    output [15:0] col_out_662,
    output [15:0] col_out_663,
    output [15:0] col_out_664,
    output [15:0] col_out_665,
    output [15:0] col_out_666,
    output [15:0] col_out_667,
    output [15:0] col_out_668,
    output [15:0] col_out_669,
    output [15:0] col_out_670,
    output [15:0] col_out_671,
    output [15:0] col_out_672,
    output [15:0] col_out_673,
    output [15:0] col_out_674,
    output [15:0] col_out_675,
    output [15:0] col_out_676,
    output [15:0] col_out_677,
    output [15:0] col_out_678,
    output [15:0] col_out_679,
    output [15:0] col_out_680,
    output [15:0] col_out_681,
    output [15:0] col_out_682,
    output [15:0] col_out_683,
    output [15:0] col_out_684,
    output [15:0] col_out_685,
    output [15:0] col_out_686,
    output [15:0] col_out_687,
    output [15:0] col_out_688,
    output [15:0] col_out_689,
    output [15:0] col_out_690,
    output [15:0] col_out_691,
    output [15:0] col_out_692,
    output [15:0] col_out_693,
    output [15:0] col_out_694,
    output [15:0] col_out_695,
    output [15:0] col_out_696,
    output [15:0] col_out_697,
    output [15:0] col_out_698,
    output [15:0] col_out_699,
    output [15:0] col_out_700,
    output [15:0] col_out_701,
    output [15:0] col_out_702,
    output [15:0] col_out_703,
    output [15:0] col_out_704,
    output [15:0] col_out_705,
    output [15:0] col_out_706,
    output [15:0] col_out_707,
    output [15:0] col_out_708,
    output [15:0] col_out_709,
    output [15:0] col_out_710,
    output [15:0] col_out_711,
    output [15:0] col_out_712,
    output [15:0] col_out_713,
    output [15:0] col_out_714,
    output [15:0] col_out_715,
    output [15:0] col_out_716,
    output [15:0] col_out_717,
    output [15:0] col_out_718,
    output [15:0] col_out_719,
    output [15:0] col_out_720,
    output [15:0] col_out_721,
    output [15:0] col_out_722,
    output [15:0] col_out_723,
    output [15:0] col_out_724,
    output [15:0] col_out_725,
    output [15:0] col_out_726,
    output [15:0] col_out_727,
    output [15:0] col_out_728,
    output [15:0] col_out_729,
    output [15:0] col_out_730,
    output [15:0] col_out_731,
    output [15:0] col_out_732,
    output [15:0] col_out_733,
    output [15:0] col_out_734,
    output [15:0] col_out_735,
    output [15:0] col_out_736,
    output [15:0] col_out_737,
    output [15:0] col_out_738,
    output [15:0] col_out_739,
    output [15:0] col_out_740,
    output [15:0] col_out_741,
    output [15:0] col_out_742,
    output [15:0] col_out_743,
    output [15:0] col_out_744,
    output [15:0] col_out_745,
    output [15:0] col_out_746,
    output [15:0] col_out_747,
    output [15:0] col_out_748,
    output [15:0] col_out_749,
    output [15:0] col_out_750,
    output [15:0] col_out_751,
    output [15:0] col_out_752,
    output [15:0] col_out_753,
    output [15:0] col_out_754,
    output [15:0] col_out_755,
    output [15:0] col_out_756,
    output [15:0] col_out_757,
    output [15:0] col_out_758,
    output [15:0] col_out_759,
    output [15:0] col_out_760,
    output [15:0] col_out_761,
    output [15:0] col_out_762,
    output [15:0] col_out_763,
    output [15:0] col_out_764,
    output [15:0] col_out_765,
    output [15:0] col_out_766,
    output [15:0] col_out_767,
    output [15:0] col_out_768,
    output [15:0] col_out_769,
    output [15:0] col_out_770,
    output [15:0] col_out_771,
    output [15:0] col_out_772,
    output [15:0] col_out_773,
    output [15:0] col_out_774,
    output [15:0] col_out_775,
    output [15:0] col_out_776,
    output [15:0] col_out_777,
    output [15:0] col_out_778,
    output [15:0] col_out_779,
    output [15:0] col_out_780,
    output [15:0] col_out_781,
    output [15:0] col_out_782,
    output [15:0] col_out_783,
    output [15:0] col_out_784,
    output [15:0] col_out_785,
    output [15:0] col_out_786,
    output [15:0] col_out_787,
    output [15:0] col_out_788,
    output [15:0] col_out_789,
    output [15:0] col_out_790,
    output [15:0] col_out_791,
    output [15:0] col_out_792,
    output [15:0] col_out_793,
    output [15:0] col_out_794,
    output [15:0] col_out_795,
    output [15:0] col_out_796,
    output [15:0] col_out_797,
    output [15:0] col_out_798,
    output [15:0] col_out_799,
    output [15:0] col_out_800,
    output [15:0] col_out_801,
    output [15:0] col_out_802,
    output [15:0] col_out_803,
    output [15:0] col_out_804,
    output [15:0] col_out_805,
    output [15:0] col_out_806,
    output [15:0] col_out_807,
    output [15:0] col_out_808,
    output [15:0] col_out_809,
    output [15:0] col_out_810,
    output [15:0] col_out_811,
    output [15:0] col_out_812,
    output [15:0] col_out_813,
    output [15:0] col_out_814,
    output [15:0] col_out_815,
    output [15:0] col_out_816,
    output [15:0] col_out_817,
    output [15:0] col_out_818,
    output [15:0] col_out_819,
    output [15:0] col_out_820,
    output [15:0] col_out_821,
    output [15:0] col_out_822,
    output [15:0] col_out_823,
    output [15:0] col_out_824,
    output [15:0] col_out_825,
    output [15:0] col_out_826,
    output [15:0] col_out_827,
    output [15:0] col_out_828,
    output [15:0] col_out_829,
    output [15:0] col_out_830,
    output [15:0] col_out_831,
    output [15:0] col_out_832,
    output [15:0] col_out_833,
    output [15:0] col_out_834,
    output [15:0] col_out_835,
    output [15:0] col_out_836,
    output [15:0] col_out_837,
    output [15:0] col_out_838,
    output [15:0] col_out_839,
    output [15:0] col_out_840,
    output [15:0] col_out_841,
    output [15:0] col_out_842,
    output [15:0] col_out_843,
    output [15:0] col_out_844,
    output [15:0] col_out_845,
    output [15:0] col_out_846,
    output [15:0] col_out_847,
    output [15:0] col_out_848,
    output [15:0] col_out_849,
    output [15:0] col_out_850,
    output [15:0] col_out_851,
    output [15:0] col_out_852,
    output [15:0] col_out_853,
    output [15:0] col_out_854,
    output [15:0] col_out_855,
    output [15:0] col_out_856,
    output [15:0] col_out_857,
    output [15:0] col_out_858,
    output [15:0] col_out_859,
    output [15:0] col_out_860,
    output [15:0] col_out_861,
    output [15:0] col_out_862,
    output [15:0] col_out_863,
    output [15:0] col_out_864,
    output [15:0] col_out_865,
    output [15:0] col_out_866,
    output [15:0] col_out_867,
    output [15:0] col_out_868,
    output [15:0] col_out_869,
    output [15:0] col_out_870,
    output [15:0] col_out_871,
    output [15:0] col_out_872,
    output [15:0] col_out_873,
    output [15:0] col_out_874,
    output [15:0] col_out_875,
    output [15:0] col_out_876,
    output [15:0] col_out_877,
    output [15:0] col_out_878,
    output [15:0] col_out_879,
    output [15:0] col_out_880,
    output [15:0] col_out_881,
    output [15:0] col_out_882,
    output [15:0] col_out_883,
    output [15:0] col_out_884,
    output [15:0] col_out_885,
    output [15:0] col_out_886,
    output [15:0] col_out_887,
    output [15:0] col_out_888,
    output [15:0] col_out_889,
    output [15:0] col_out_890,
    output [15:0] col_out_891,
    output [15:0] col_out_892,
    output [15:0] col_out_893,
    output [15:0] col_out_894,
    output [15:0] col_out_895,
    output [15:0] col_out_896,
    output [15:0] col_out_897,
    output [15:0] col_out_898,
    output [15:0] col_out_899,
    output [15:0] col_out_900,
    output [15:0] col_out_901,
    output [15:0] col_out_902,
    output [15:0] col_out_903,
    output [15:0] col_out_904,
    output [15:0] col_out_905,
    output [15:0] col_out_906,
    output [15:0] col_out_907,
    output [15:0] col_out_908,
    output [15:0] col_out_909,
    output [15:0] col_out_910,
    output [15:0] col_out_911,
    output [15:0] col_out_912,
    output [15:0] col_out_913,
    output [15:0] col_out_914,
    output [15:0] col_out_915,
    output [15:0] col_out_916,
    output [15:0] col_out_917,
    output [15:0] col_out_918,
    output [15:0] col_out_919,
    output [15:0] col_out_920,
    output [15:0] col_out_921,
    output [15:0] col_out_922,
    output [15:0] col_out_923,
    output [15:0] col_out_924,
    output [15:0] col_out_925,
    output [15:0] col_out_926,
    output [15:0] col_out_927,
    output [15:0] col_out_928,
    output [15:0] col_out_929,
    output [15:0] col_out_930,
    output [15:0] col_out_931,
    output [15:0] col_out_932,
    output [15:0] col_out_933,
    output [15:0] col_out_934,
    output [15:0] col_out_935,
    output [15:0] col_out_936,
    output [15:0] col_out_937,
    output [15:0] col_out_938,
    output [15:0] col_out_939,
    output [15:0] col_out_940,
    output [15:0] col_out_941,
    output [15:0] col_out_942,
    output [15:0] col_out_943,
    output [15:0] col_out_944,
    output [15:0] col_out_945,
    output [15:0] col_out_946,
    output [15:0] col_out_947,
    output [15:0] col_out_948,
    output [15:0] col_out_949,
    output [15:0] col_out_950,
    output [15:0] col_out_951,
    output [15:0] col_out_952,
    output [15:0] col_out_953,
    output [15:0] col_out_954,
    output [15:0] col_out_955,
    output [15:0] col_out_956,
    output [15:0] col_out_957,
    output [15:0] col_out_958,
    output [15:0] col_out_959,
    output [15:0] col_out_960,
    output [15:0] col_out_961,
    output [15:0] col_out_962,
    output [15:0] col_out_963,
    output [15:0] col_out_964,
    output [15:0] col_out_965,
    output [15:0] col_out_966,
    output [15:0] col_out_967,
    output [15:0] col_out_968,
    output [15:0] col_out_969,
    output [15:0] col_out_970,
    output [15:0] col_out_971,
    output [15:0] col_out_972,
    output [15:0] col_out_973,
    output [15:0] col_out_974,
    output [15:0] col_out_975,
    output [15:0] col_out_976,
    output [15:0] col_out_977,
    output [15:0] col_out_978,
    output [15:0] col_out_979,
    output [15:0] col_out_980,
    output [15:0] col_out_981,
    output [15:0] col_out_982,
    output [15:0] col_out_983,
    output [15:0] col_out_984,
    output [15:0] col_out_985,
    output [15:0] col_out_986,
    output [15:0] col_out_987,
    output [15:0] col_out_988,
    output [15:0] col_out_989,
    output [15:0] col_out_990,
    output [15:0] col_out_991,
    output [15:0] col_out_992,
    output [15:0] col_out_993,
    output [15:0] col_out_994,
    output [15:0] col_out_995,
    output [15:0] col_out_996,
    output [15:0] col_out_997,
    output [15:0] col_out_998,
    output [15:0] col_out_999,
    output [15:0] col_out_1000,
    output [15:0] col_out_1001,
    output [15:0] col_out_1002,
    output [15:0] col_out_1003,
    output [15:0] col_out_1004,
    output [15:0] col_out_1005,
    output [15:0] col_out_1006,
    output [15:0] col_out_1007,
    output [15:0] col_out_1008,
    output [15:0] col_out_1009,
    output [15:0] col_out_1010,
    output [15:0] col_out_1011,
    output [15:0] col_out_1012,
    output [15:0] col_out_1013,
    output [15:0] col_out_1014,
    output [15:0] col_out_1015,
    output [15:0] col_out_1016,
    output [15:0] col_out_1017,
    output [15:0] col_out_1018,
    output [15:0] col_out_1019,
    output [15:0] col_out_1020,
    output [15:0] col_out_1021,
    output [15:0] col_out_1022,
    output [15:0] col_out_1023,
    output [15:0] col_out_1024,
    output [15:0] col_out_1025,
    output [15:0] col_out_1026,
    output [15:0] col_out_1027,
    output [15:0] col_out_1028,
    output [15:0] col_out_1029,
    output [15:0] col_out_1030,
    output [15:0] col_out_1031,
    output [15:0] col_out_1032
);



//--compressor_array input and output----------------------

wire [53:0] u_ca_in_0;
wire [53:0] u_ca_in_1;
wire [53:0] u_ca_in_2;
wire [53:0] u_ca_in_3;
wire [53:0] u_ca_in_4;
wire [53:0] u_ca_in_5;
wire [53:0] u_ca_in_6;
wire [53:0] u_ca_in_7;
wire [53:0] u_ca_in_8;
wire [53:0] u_ca_in_9;
wire [53:0] u_ca_in_10;
wire [53:0] u_ca_in_11;
wire [53:0] u_ca_in_12;
wire [53:0] u_ca_in_13;
wire [53:0] u_ca_in_14;
wire [53:0] u_ca_in_15;
wire [53:0] u_ca_in_16;
wire [53:0] u_ca_in_17;
wire [53:0] u_ca_in_18;
wire [53:0] u_ca_in_19;
wire [53:0] u_ca_in_20;
wire [53:0] u_ca_in_21;
wire [53:0] u_ca_in_22;
wire [53:0] u_ca_in_23;
wire [53:0] u_ca_in_24;
wire [53:0] u_ca_in_25;
wire [53:0] u_ca_in_26;
wire [53:0] u_ca_in_27;
wire [53:0] u_ca_in_28;
wire [53:0] u_ca_in_29;
wire [53:0] u_ca_in_30;
wire [53:0] u_ca_in_31;
wire [53:0] u_ca_in_32;
wire [53:0] u_ca_in_33;
wire [53:0] u_ca_in_34;
wire [53:0] u_ca_in_35;
wire [53:0] u_ca_in_36;
wire [53:0] u_ca_in_37;
wire [53:0] u_ca_in_38;
wire [53:0] u_ca_in_39;
wire [53:0] u_ca_in_40;
wire [53:0] u_ca_in_41;
wire [53:0] u_ca_in_42;
wire [53:0] u_ca_in_43;
wire [53:0] u_ca_in_44;
wire [53:0] u_ca_in_45;
wire [53:0] u_ca_in_46;
wire [53:0] u_ca_in_47;
wire [53:0] u_ca_in_48;
wire [53:0] u_ca_in_49;
wire [53:0] u_ca_in_50;
wire [53:0] u_ca_in_51;
wire [53:0] u_ca_in_52;
wire [53:0] u_ca_in_53;
wire [53:0] u_ca_in_54;
wire [53:0] u_ca_in_55;
wire [53:0] u_ca_in_56;
wire [53:0] u_ca_in_57;
wire [53:0] u_ca_in_58;
wire [53:0] u_ca_in_59;
wire [53:0] u_ca_in_60;
wire [53:0] u_ca_in_61;
wire [53:0] u_ca_in_62;
wire [53:0] u_ca_in_63;
wire [53:0] u_ca_in_64;
wire [53:0] u_ca_in_65;
wire [53:0] u_ca_in_66;
wire [53:0] u_ca_in_67;
wire [53:0] u_ca_in_68;
wire [53:0] u_ca_in_69;
wire [53:0] u_ca_in_70;
wire [53:0] u_ca_in_71;
wire [53:0] u_ca_in_72;
wire [53:0] u_ca_in_73;
wire [53:0] u_ca_in_74;
wire [53:0] u_ca_in_75;
wire [53:0] u_ca_in_76;
wire [53:0] u_ca_in_77;
wire [53:0] u_ca_in_78;
wire [53:0] u_ca_in_79;
wire [53:0] u_ca_in_80;
wire [53:0] u_ca_in_81;
wire [53:0] u_ca_in_82;
wire [53:0] u_ca_in_83;
wire [53:0] u_ca_in_84;
wire [53:0] u_ca_in_85;
wire [53:0] u_ca_in_86;
wire [53:0] u_ca_in_87;
wire [53:0] u_ca_in_88;
wire [53:0] u_ca_in_89;
wire [53:0] u_ca_in_90;
wire [53:0] u_ca_in_91;
wire [53:0] u_ca_in_92;
wire [53:0] u_ca_in_93;
wire [53:0] u_ca_in_94;
wire [53:0] u_ca_in_95;
wire [53:0] u_ca_in_96;
wire [53:0] u_ca_in_97;
wire [53:0] u_ca_in_98;
wire [53:0] u_ca_in_99;
wire [53:0] u_ca_in_100;
wire [53:0] u_ca_in_101;
wire [53:0] u_ca_in_102;
wire [53:0] u_ca_in_103;
wire [53:0] u_ca_in_104;
wire [53:0] u_ca_in_105;
wire [53:0] u_ca_in_106;
wire [53:0] u_ca_in_107;
wire [53:0] u_ca_in_108;
wire [53:0] u_ca_in_109;
wire [53:0] u_ca_in_110;
wire [53:0] u_ca_in_111;
wire [53:0] u_ca_in_112;
wire [53:0] u_ca_in_113;
wire [53:0] u_ca_in_114;
wire [53:0] u_ca_in_115;
wire [53:0] u_ca_in_116;
wire [53:0] u_ca_in_117;
wire [53:0] u_ca_in_118;
wire [53:0] u_ca_in_119;
wire [53:0] u_ca_in_120;
wire [53:0] u_ca_in_121;
wire [53:0] u_ca_in_122;
wire [53:0] u_ca_in_123;
wire [53:0] u_ca_in_124;
wire [53:0] u_ca_in_125;
wire [53:0] u_ca_in_126;
wire [53:0] u_ca_in_127;
wire [53:0] u_ca_in_128;
wire [53:0] u_ca_in_129;
wire [53:0] u_ca_in_130;
wire [53:0] u_ca_in_131;
wire [53:0] u_ca_in_132;
wire [53:0] u_ca_in_133;
wire [53:0] u_ca_in_134;
wire [53:0] u_ca_in_135;
wire [53:0] u_ca_in_136;
wire [53:0] u_ca_in_137;
wire [53:0] u_ca_in_138;
wire [53:0] u_ca_in_139;
wire [53:0] u_ca_in_140;
wire [53:0] u_ca_in_141;
wire [53:0] u_ca_in_142;
wire [53:0] u_ca_in_143;
wire [53:0] u_ca_in_144;
wire [53:0] u_ca_in_145;
wire [53:0] u_ca_in_146;
wire [53:0] u_ca_in_147;
wire [53:0] u_ca_in_148;
wire [53:0] u_ca_in_149;
wire [53:0] u_ca_in_150;
wire [53:0] u_ca_in_151;
wire [53:0] u_ca_in_152;
wire [53:0] u_ca_in_153;
wire [53:0] u_ca_in_154;
wire [53:0] u_ca_in_155;
wire [53:0] u_ca_in_156;
wire [53:0] u_ca_in_157;
wire [53:0] u_ca_in_158;
wire [53:0] u_ca_in_159;
wire [53:0] u_ca_in_160;
wire [53:0] u_ca_in_161;
wire [53:0] u_ca_in_162;
wire [53:0] u_ca_in_163;
wire [53:0] u_ca_in_164;
wire [53:0] u_ca_in_165;
wire [53:0] u_ca_in_166;
wire [53:0] u_ca_in_167;
wire [53:0] u_ca_in_168;
wire [53:0] u_ca_in_169;
wire [53:0] u_ca_in_170;
wire [53:0] u_ca_in_171;
wire [53:0] u_ca_in_172;
wire [53:0] u_ca_in_173;
wire [53:0] u_ca_in_174;
wire [53:0] u_ca_in_175;
wire [53:0] u_ca_in_176;
wire [53:0] u_ca_in_177;
wire [53:0] u_ca_in_178;
wire [53:0] u_ca_in_179;
wire [53:0] u_ca_in_180;
wire [53:0] u_ca_in_181;
wire [53:0] u_ca_in_182;
wire [53:0] u_ca_in_183;
wire [53:0] u_ca_in_184;
wire [53:0] u_ca_in_185;
wire [53:0] u_ca_in_186;
wire [53:0] u_ca_in_187;
wire [53:0] u_ca_in_188;
wire [53:0] u_ca_in_189;
wire [53:0] u_ca_in_190;
wire [53:0] u_ca_in_191;
wire [53:0] u_ca_in_192;
wire [53:0] u_ca_in_193;
wire [53:0] u_ca_in_194;
wire [53:0] u_ca_in_195;
wire [53:0] u_ca_in_196;
wire [53:0] u_ca_in_197;
wire [53:0] u_ca_in_198;
wire [53:0] u_ca_in_199;
wire [53:0] u_ca_in_200;
wire [53:0] u_ca_in_201;
wire [53:0] u_ca_in_202;
wire [53:0] u_ca_in_203;
wire [53:0] u_ca_in_204;
wire [53:0] u_ca_in_205;
wire [53:0] u_ca_in_206;
wire [53:0] u_ca_in_207;
wire [53:0] u_ca_in_208;
wire [53:0] u_ca_in_209;
wire [53:0] u_ca_in_210;
wire [53:0] u_ca_in_211;
wire [53:0] u_ca_in_212;
wire [53:0] u_ca_in_213;
wire [53:0] u_ca_in_214;
wire [53:0] u_ca_in_215;
wire [53:0] u_ca_in_216;
wire [53:0] u_ca_in_217;
wire [53:0] u_ca_in_218;
wire [53:0] u_ca_in_219;
wire [53:0] u_ca_in_220;
wire [53:0] u_ca_in_221;
wire [53:0] u_ca_in_222;
wire [53:0] u_ca_in_223;
wire [53:0] u_ca_in_224;
wire [53:0] u_ca_in_225;
wire [53:0] u_ca_in_226;
wire [53:0] u_ca_in_227;
wire [53:0] u_ca_in_228;
wire [53:0] u_ca_in_229;
wire [53:0] u_ca_in_230;
wire [53:0] u_ca_in_231;
wire [53:0] u_ca_in_232;
wire [53:0] u_ca_in_233;
wire [53:0] u_ca_in_234;
wire [53:0] u_ca_in_235;
wire [53:0] u_ca_in_236;
wire [53:0] u_ca_in_237;
wire [53:0] u_ca_in_238;
wire [53:0] u_ca_in_239;
wire [53:0] u_ca_in_240;
wire [53:0] u_ca_in_241;
wire [53:0] u_ca_in_242;
wire [53:0] u_ca_in_243;
wire [53:0] u_ca_in_244;
wire [53:0] u_ca_in_245;
wire [53:0] u_ca_in_246;
wire [53:0] u_ca_in_247;
wire [53:0] u_ca_in_248;
wire [53:0] u_ca_in_249;
wire [53:0] u_ca_in_250;
wire [53:0] u_ca_in_251;
wire [53:0] u_ca_in_252;
wire [53:0] u_ca_in_253;
wire [53:0] u_ca_in_254;
wire [53:0] u_ca_in_255;
wire [53:0] u_ca_in_256;
wire [53:0] u_ca_in_257;
wire [53:0] u_ca_in_258;
wire [53:0] u_ca_in_259;
wire [53:0] u_ca_in_260;
wire [53:0] u_ca_in_261;
wire [53:0] u_ca_in_262;
wire [53:0] u_ca_in_263;
wire [53:0] u_ca_in_264;
wire [53:0] u_ca_in_265;
wire [53:0] u_ca_in_266;
wire [53:0] u_ca_in_267;
wire [53:0] u_ca_in_268;
wire [53:0] u_ca_in_269;
wire [53:0] u_ca_in_270;
wire [53:0] u_ca_in_271;
wire [53:0] u_ca_in_272;
wire [53:0] u_ca_in_273;
wire [53:0] u_ca_in_274;
wire [53:0] u_ca_in_275;
wire [53:0] u_ca_in_276;
wire [53:0] u_ca_in_277;
wire [53:0] u_ca_in_278;
wire [53:0] u_ca_in_279;
wire [53:0] u_ca_in_280;
wire [53:0] u_ca_in_281;
wire [53:0] u_ca_in_282;
wire [53:0] u_ca_in_283;
wire [53:0] u_ca_in_284;
wire [53:0] u_ca_in_285;
wire [53:0] u_ca_in_286;
wire [53:0] u_ca_in_287;
wire [53:0] u_ca_in_288;
wire [53:0] u_ca_in_289;
wire [53:0] u_ca_in_290;
wire [53:0] u_ca_in_291;
wire [53:0] u_ca_in_292;
wire [53:0] u_ca_in_293;
wire [53:0] u_ca_in_294;
wire [53:0] u_ca_in_295;
wire [53:0] u_ca_in_296;
wire [53:0] u_ca_in_297;
wire [53:0] u_ca_in_298;
wire [53:0] u_ca_in_299;
wire [53:0] u_ca_in_300;
wire [53:0] u_ca_in_301;
wire [53:0] u_ca_in_302;
wire [53:0] u_ca_in_303;
wire [53:0] u_ca_in_304;
wire [53:0] u_ca_in_305;
wire [53:0] u_ca_in_306;
wire [53:0] u_ca_in_307;
wire [53:0] u_ca_in_308;
wire [53:0] u_ca_in_309;
wire [53:0] u_ca_in_310;
wire [53:0] u_ca_in_311;
wire [53:0] u_ca_in_312;
wire [53:0] u_ca_in_313;
wire [53:0] u_ca_in_314;
wire [53:0] u_ca_in_315;
wire [53:0] u_ca_in_316;
wire [53:0] u_ca_in_317;
wire [53:0] u_ca_in_318;
wire [53:0] u_ca_in_319;
wire [53:0] u_ca_in_320;
wire [53:0] u_ca_in_321;
wire [53:0] u_ca_in_322;
wire [53:0] u_ca_in_323;
wire [53:0] u_ca_in_324;
wire [53:0] u_ca_in_325;
wire [53:0] u_ca_in_326;
wire [53:0] u_ca_in_327;
wire [53:0] u_ca_in_328;
wire [53:0] u_ca_in_329;
wire [53:0] u_ca_in_330;
wire [53:0] u_ca_in_331;
wire [53:0] u_ca_in_332;
wire [53:0] u_ca_in_333;
wire [53:0] u_ca_in_334;
wire [53:0] u_ca_in_335;
wire [53:0] u_ca_in_336;
wire [53:0] u_ca_in_337;
wire [53:0] u_ca_in_338;
wire [53:0] u_ca_in_339;
wire [53:0] u_ca_in_340;
wire [53:0] u_ca_in_341;
wire [53:0] u_ca_in_342;
wire [53:0] u_ca_in_343;
wire [53:0] u_ca_in_344;
wire [53:0] u_ca_in_345;
wire [53:0] u_ca_in_346;
wire [53:0] u_ca_in_347;
wire [53:0] u_ca_in_348;
wire [53:0] u_ca_in_349;
wire [53:0] u_ca_in_350;
wire [53:0] u_ca_in_351;
wire [53:0] u_ca_in_352;
wire [53:0] u_ca_in_353;
wire [53:0] u_ca_in_354;
wire [53:0] u_ca_in_355;
wire [53:0] u_ca_in_356;
wire [53:0] u_ca_in_357;
wire [53:0] u_ca_in_358;
wire [53:0] u_ca_in_359;
wire [53:0] u_ca_in_360;
wire [53:0] u_ca_in_361;
wire [53:0] u_ca_in_362;
wire [53:0] u_ca_in_363;
wire [53:0] u_ca_in_364;
wire [53:0] u_ca_in_365;
wire [53:0] u_ca_in_366;
wire [53:0] u_ca_in_367;
wire [53:0] u_ca_in_368;
wire [53:0] u_ca_in_369;
wire [53:0] u_ca_in_370;
wire [53:0] u_ca_in_371;
wire [53:0] u_ca_in_372;
wire [53:0] u_ca_in_373;
wire [53:0] u_ca_in_374;
wire [53:0] u_ca_in_375;
wire [53:0] u_ca_in_376;
wire [53:0] u_ca_in_377;
wire [53:0] u_ca_in_378;
wire [53:0] u_ca_in_379;
wire [53:0] u_ca_in_380;
wire [53:0] u_ca_in_381;
wire [53:0] u_ca_in_382;
wire [53:0] u_ca_in_383;
wire [53:0] u_ca_in_384;
wire [53:0] u_ca_in_385;
wire [53:0] u_ca_in_386;
wire [53:0] u_ca_in_387;
wire [53:0] u_ca_in_388;
wire [53:0] u_ca_in_389;
wire [53:0] u_ca_in_390;
wire [53:0] u_ca_in_391;
wire [53:0] u_ca_in_392;
wire [53:0] u_ca_in_393;
wire [53:0] u_ca_in_394;
wire [53:0] u_ca_in_395;
wire [53:0] u_ca_in_396;
wire [53:0] u_ca_in_397;
wire [53:0] u_ca_in_398;
wire [53:0] u_ca_in_399;
wire [53:0] u_ca_in_400;
wire [53:0] u_ca_in_401;
wire [53:0] u_ca_in_402;
wire [53:0] u_ca_in_403;
wire [53:0] u_ca_in_404;
wire [53:0] u_ca_in_405;
wire [53:0] u_ca_in_406;
wire [53:0] u_ca_in_407;
wire [53:0] u_ca_in_408;
wire [53:0] u_ca_in_409;
wire [53:0] u_ca_in_410;
wire [53:0] u_ca_in_411;
wire [53:0] u_ca_in_412;
wire [53:0] u_ca_in_413;
wire [53:0] u_ca_in_414;
wire [53:0] u_ca_in_415;
wire [53:0] u_ca_in_416;
wire [53:0] u_ca_in_417;
wire [53:0] u_ca_in_418;
wire [53:0] u_ca_in_419;
wire [53:0] u_ca_in_420;
wire [53:0] u_ca_in_421;
wire [53:0] u_ca_in_422;
wire [53:0] u_ca_in_423;
wire [53:0] u_ca_in_424;
wire [53:0] u_ca_in_425;
wire [53:0] u_ca_in_426;
wire [53:0] u_ca_in_427;
wire [53:0] u_ca_in_428;
wire [53:0] u_ca_in_429;
wire [53:0] u_ca_in_430;
wire [53:0] u_ca_in_431;
wire [53:0] u_ca_in_432;
wire [53:0] u_ca_in_433;
wire [53:0] u_ca_in_434;
wire [53:0] u_ca_in_435;
wire [53:0] u_ca_in_436;
wire [53:0] u_ca_in_437;
wire [53:0] u_ca_in_438;
wire [53:0] u_ca_in_439;
wire [53:0] u_ca_in_440;
wire [53:0] u_ca_in_441;
wire [53:0] u_ca_in_442;
wire [53:0] u_ca_in_443;
wire [53:0] u_ca_in_444;
wire [53:0] u_ca_in_445;
wire [53:0] u_ca_in_446;
wire [53:0] u_ca_in_447;
wire [53:0] u_ca_in_448;
wire [53:0] u_ca_in_449;
wire [53:0] u_ca_in_450;
wire [53:0] u_ca_in_451;
wire [53:0] u_ca_in_452;
wire [53:0] u_ca_in_453;
wire [53:0] u_ca_in_454;
wire [53:0] u_ca_in_455;
wire [53:0] u_ca_in_456;
wire [53:0] u_ca_in_457;
wire [53:0] u_ca_in_458;
wire [53:0] u_ca_in_459;
wire [53:0] u_ca_in_460;
wire [53:0] u_ca_in_461;
wire [53:0] u_ca_in_462;
wire [53:0] u_ca_in_463;
wire [53:0] u_ca_in_464;
wire [53:0] u_ca_in_465;
wire [53:0] u_ca_in_466;
wire [53:0] u_ca_in_467;
wire [53:0] u_ca_in_468;
wire [53:0] u_ca_in_469;
wire [53:0] u_ca_in_470;
wire [53:0] u_ca_in_471;
wire [53:0] u_ca_in_472;
wire [53:0] u_ca_in_473;
wire [53:0] u_ca_in_474;
wire [53:0] u_ca_in_475;
wire [53:0] u_ca_in_476;
wire [53:0] u_ca_in_477;
wire [53:0] u_ca_in_478;
wire [53:0] u_ca_in_479;
wire [53:0] u_ca_in_480;
wire [53:0] u_ca_in_481;
wire [53:0] u_ca_in_482;
wire [53:0] u_ca_in_483;
wire [53:0] u_ca_in_484;
wire [53:0] u_ca_in_485;
wire [53:0] u_ca_in_486;
wire [53:0] u_ca_in_487;
wire [53:0] u_ca_in_488;
wire [53:0] u_ca_in_489;
wire [53:0] u_ca_in_490;
wire [53:0] u_ca_in_491;
wire [53:0] u_ca_in_492;
wire [53:0] u_ca_in_493;
wire [53:0] u_ca_in_494;
wire [53:0] u_ca_in_495;
wire [53:0] u_ca_in_496;
wire [53:0] u_ca_in_497;
wire [53:0] u_ca_in_498;
wire [53:0] u_ca_in_499;
wire [53:0] u_ca_in_500;
wire [53:0] u_ca_in_501;
wire [53:0] u_ca_in_502;
wire [53:0] u_ca_in_503;
wire [53:0] u_ca_in_504;
wire [53:0] u_ca_in_505;
wire [53:0] u_ca_in_506;
wire [53:0] u_ca_in_507;
wire [53:0] u_ca_in_508;
wire [53:0] u_ca_in_509;
wire [53:0] u_ca_in_510;
wire [53:0] u_ca_in_511;
wire [53:0] u_ca_in_512;
wire [53:0] u_ca_in_513;
wire [53:0] u_ca_in_514;
wire [53:0] u_ca_in_515;
wire [53:0] u_ca_in_516;
wire [53:0] u_ca_in_517;
wire [53:0] u_ca_in_518;
wire [53:0] u_ca_in_519;
wire [53:0] u_ca_in_520;
wire [53:0] u_ca_in_521;
wire [53:0] u_ca_in_522;
wire [53:0] u_ca_in_523;
wire [53:0] u_ca_in_524;
wire [53:0] u_ca_in_525;
wire [53:0] u_ca_in_526;
wire [53:0] u_ca_in_527;
wire [53:0] u_ca_in_528;
wire [53:0] u_ca_in_529;
wire [53:0] u_ca_in_530;
wire [53:0] u_ca_in_531;
wire [53:0] u_ca_in_532;
wire [53:0] u_ca_in_533;
wire [53:0] u_ca_in_534;
wire [53:0] u_ca_in_535;
wire [53:0] u_ca_in_536;
wire [53:0] u_ca_in_537;
wire [53:0] u_ca_in_538;
wire [53:0] u_ca_in_539;
wire [53:0] u_ca_in_540;
wire [53:0] u_ca_in_541;
wire [53:0] u_ca_in_542;
wire [53:0] u_ca_in_543;
wire [53:0] u_ca_in_544;
wire [53:0] u_ca_in_545;
wire [53:0] u_ca_in_546;
wire [53:0] u_ca_in_547;
wire [53:0] u_ca_in_548;
wire [53:0] u_ca_in_549;
wire [53:0] u_ca_in_550;
wire [53:0] u_ca_in_551;
wire [53:0] u_ca_in_552;
wire [53:0] u_ca_in_553;
wire [53:0] u_ca_in_554;
wire [53:0] u_ca_in_555;
wire [53:0] u_ca_in_556;
wire [53:0] u_ca_in_557;
wire [53:0] u_ca_in_558;
wire [53:0] u_ca_in_559;
wire [53:0] u_ca_in_560;
wire [53:0] u_ca_in_561;
wire [53:0] u_ca_in_562;
wire [53:0] u_ca_in_563;
wire [53:0] u_ca_in_564;
wire [53:0] u_ca_in_565;
wire [53:0] u_ca_in_566;
wire [53:0] u_ca_in_567;
wire [53:0] u_ca_in_568;
wire [53:0] u_ca_in_569;
wire [53:0] u_ca_in_570;
wire [53:0] u_ca_in_571;
wire [53:0] u_ca_in_572;
wire [53:0] u_ca_in_573;
wire [53:0] u_ca_in_574;
wire [53:0] u_ca_in_575;
wire [53:0] u_ca_in_576;
wire [53:0] u_ca_in_577;
wire [53:0] u_ca_in_578;
wire [53:0] u_ca_in_579;
wire [53:0] u_ca_in_580;
wire [53:0] u_ca_in_581;
wire [53:0] u_ca_in_582;
wire [53:0] u_ca_in_583;
wire [53:0] u_ca_in_584;
wire [53:0] u_ca_in_585;
wire [53:0] u_ca_in_586;
wire [53:0] u_ca_in_587;
wire [53:0] u_ca_in_588;
wire [53:0] u_ca_in_589;
wire [53:0] u_ca_in_590;
wire [53:0] u_ca_in_591;
wire [53:0] u_ca_in_592;
wire [53:0] u_ca_in_593;
wire [53:0] u_ca_in_594;
wire [53:0] u_ca_in_595;
wire [53:0] u_ca_in_596;
wire [53:0] u_ca_in_597;
wire [53:0] u_ca_in_598;
wire [53:0] u_ca_in_599;
wire [53:0] u_ca_in_600;
wire [53:0] u_ca_in_601;
wire [53:0] u_ca_in_602;
wire [53:0] u_ca_in_603;
wire [53:0] u_ca_in_604;
wire [53:0] u_ca_in_605;
wire [53:0] u_ca_in_606;
wire [53:0] u_ca_in_607;
wire [53:0] u_ca_in_608;
wire [53:0] u_ca_in_609;
wire [53:0] u_ca_in_610;
wire [53:0] u_ca_in_611;
wire [53:0] u_ca_in_612;
wire [53:0] u_ca_in_613;
wire [53:0] u_ca_in_614;
wire [53:0] u_ca_in_615;
wire [53:0] u_ca_in_616;
wire [53:0] u_ca_in_617;
wire [53:0] u_ca_in_618;
wire [53:0] u_ca_in_619;
wire [53:0] u_ca_in_620;
wire [53:0] u_ca_in_621;
wire [53:0] u_ca_in_622;
wire [53:0] u_ca_in_623;
wire [53:0] u_ca_in_624;
wire [53:0] u_ca_in_625;
wire [53:0] u_ca_in_626;
wire [53:0] u_ca_in_627;
wire [53:0] u_ca_in_628;
wire [53:0] u_ca_in_629;
wire [53:0] u_ca_in_630;
wire [53:0] u_ca_in_631;
wire [53:0] u_ca_in_632;
wire [53:0] u_ca_in_633;
wire [53:0] u_ca_in_634;
wire [53:0] u_ca_in_635;
wire [53:0] u_ca_in_636;
wire [53:0] u_ca_in_637;
wire [53:0] u_ca_in_638;
wire [53:0] u_ca_in_639;
wire [53:0] u_ca_in_640;
wire [53:0] u_ca_in_641;
wire [53:0] u_ca_in_642;
wire [53:0] u_ca_in_643;
wire [53:0] u_ca_in_644;
wire [53:0] u_ca_in_645;
wire [53:0] u_ca_in_646;
wire [53:0] u_ca_in_647;
wire [53:0] u_ca_in_648;
wire [53:0] u_ca_in_649;
wire [53:0] u_ca_in_650;
wire [53:0] u_ca_in_651;
wire [53:0] u_ca_in_652;
wire [53:0] u_ca_in_653;
wire [53:0] u_ca_in_654;
wire [53:0] u_ca_in_655;
wire [53:0] u_ca_in_656;
wire [53:0] u_ca_in_657;
wire [53:0] u_ca_in_658;
wire [53:0] u_ca_in_659;
wire [53:0] u_ca_in_660;
wire [53:0] u_ca_in_661;
wire [53:0] u_ca_in_662;
wire [53:0] u_ca_in_663;
wire [53:0] u_ca_in_664;
wire [53:0] u_ca_in_665;
wire [53:0] u_ca_in_666;
wire [53:0] u_ca_in_667;
wire [53:0] u_ca_in_668;
wire [53:0] u_ca_in_669;
wire [53:0] u_ca_in_670;
wire [53:0] u_ca_in_671;
wire [53:0] u_ca_in_672;
wire [53:0] u_ca_in_673;
wire [53:0] u_ca_in_674;
wire [53:0] u_ca_in_675;
wire [53:0] u_ca_in_676;
wire [53:0] u_ca_in_677;
wire [53:0] u_ca_in_678;
wire [53:0] u_ca_in_679;
wire [53:0] u_ca_in_680;
wire [53:0] u_ca_in_681;
wire [53:0] u_ca_in_682;
wire [53:0] u_ca_in_683;
wire [53:0] u_ca_in_684;
wire [53:0] u_ca_in_685;
wire [53:0] u_ca_in_686;
wire [53:0] u_ca_in_687;
wire [53:0] u_ca_in_688;
wire [53:0] u_ca_in_689;
wire [53:0] u_ca_in_690;
wire [53:0] u_ca_in_691;
wire [53:0] u_ca_in_692;
wire [53:0] u_ca_in_693;
wire [53:0] u_ca_in_694;
wire [53:0] u_ca_in_695;
wire [53:0] u_ca_in_696;
wire [53:0] u_ca_in_697;
wire [53:0] u_ca_in_698;
wire [53:0] u_ca_in_699;
wire [53:0] u_ca_in_700;
wire [53:0] u_ca_in_701;
wire [53:0] u_ca_in_702;
wire [53:0] u_ca_in_703;
wire [53:0] u_ca_in_704;
wire [53:0] u_ca_in_705;
wire [53:0] u_ca_in_706;
wire [53:0] u_ca_in_707;
wire [53:0] u_ca_in_708;
wire [53:0] u_ca_in_709;
wire [53:0] u_ca_in_710;
wire [53:0] u_ca_in_711;
wire [53:0] u_ca_in_712;
wire [53:0] u_ca_in_713;
wire [53:0] u_ca_in_714;
wire [53:0] u_ca_in_715;
wire [53:0] u_ca_in_716;
wire [53:0] u_ca_in_717;
wire [53:0] u_ca_in_718;
wire [53:0] u_ca_in_719;
wire [53:0] u_ca_in_720;
wire [53:0] u_ca_in_721;
wire [53:0] u_ca_in_722;
wire [53:0] u_ca_in_723;
wire [53:0] u_ca_in_724;
wire [53:0] u_ca_in_725;
wire [53:0] u_ca_in_726;
wire [53:0] u_ca_in_727;
wire [53:0] u_ca_in_728;
wire [53:0] u_ca_in_729;
wire [53:0] u_ca_in_730;
wire [53:0] u_ca_in_731;
wire [53:0] u_ca_in_732;
wire [53:0] u_ca_in_733;
wire [53:0] u_ca_in_734;
wire [53:0] u_ca_in_735;
wire [53:0] u_ca_in_736;
wire [53:0] u_ca_in_737;
wire [53:0] u_ca_in_738;
wire [53:0] u_ca_in_739;
wire [53:0] u_ca_in_740;
wire [53:0] u_ca_in_741;
wire [53:0] u_ca_in_742;
wire [53:0] u_ca_in_743;
wire [53:0] u_ca_in_744;
wire [53:0] u_ca_in_745;
wire [53:0] u_ca_in_746;
wire [53:0] u_ca_in_747;
wire [53:0] u_ca_in_748;
wire [53:0] u_ca_in_749;
wire [53:0] u_ca_in_750;
wire [53:0] u_ca_in_751;
wire [53:0] u_ca_in_752;
wire [53:0] u_ca_in_753;
wire [53:0] u_ca_in_754;
wire [53:0] u_ca_in_755;
wire [53:0] u_ca_in_756;
wire [53:0] u_ca_in_757;
wire [53:0] u_ca_in_758;
wire [53:0] u_ca_in_759;
wire [53:0] u_ca_in_760;
wire [53:0] u_ca_in_761;
wire [53:0] u_ca_in_762;
wire [53:0] u_ca_in_763;
wire [53:0] u_ca_in_764;
wire [53:0] u_ca_in_765;
wire [53:0] u_ca_in_766;
wire [53:0] u_ca_in_767;
wire [53:0] u_ca_in_768;
wire [53:0] u_ca_in_769;
wire [53:0] u_ca_in_770;
wire [53:0] u_ca_in_771;
wire [53:0] u_ca_in_772;
wire [53:0] u_ca_in_773;
wire [53:0] u_ca_in_774;
wire [53:0] u_ca_in_775;
wire [53:0] u_ca_in_776;
wire [53:0] u_ca_in_777;
wire [53:0] u_ca_in_778;
wire [53:0] u_ca_in_779;
wire [53:0] u_ca_in_780;
wire [53:0] u_ca_in_781;
wire [53:0] u_ca_in_782;
wire [53:0] u_ca_in_783;
wire [53:0] u_ca_in_784;
wire [53:0] u_ca_in_785;
wire [53:0] u_ca_in_786;
wire [53:0] u_ca_in_787;
wire [53:0] u_ca_in_788;
wire [53:0] u_ca_in_789;
wire [53:0] u_ca_in_790;
wire [53:0] u_ca_in_791;
wire [53:0] u_ca_in_792;
wire [53:0] u_ca_in_793;
wire [53:0] u_ca_in_794;
wire [53:0] u_ca_in_795;
wire [53:0] u_ca_in_796;
wire [53:0] u_ca_in_797;
wire [53:0] u_ca_in_798;
wire [53:0] u_ca_in_799;
wire [53:0] u_ca_in_800;
wire [53:0] u_ca_in_801;
wire [53:0] u_ca_in_802;
wire [53:0] u_ca_in_803;
wire [53:0] u_ca_in_804;
wire [53:0] u_ca_in_805;
wire [53:0] u_ca_in_806;
wire [53:0] u_ca_in_807;
wire [53:0] u_ca_in_808;
wire [53:0] u_ca_in_809;
wire [53:0] u_ca_in_810;
wire [53:0] u_ca_in_811;
wire [53:0] u_ca_in_812;
wire [53:0] u_ca_in_813;
wire [53:0] u_ca_in_814;
wire [53:0] u_ca_in_815;
wire [53:0] u_ca_in_816;
wire [53:0] u_ca_in_817;
wire [53:0] u_ca_in_818;
wire [53:0] u_ca_in_819;
wire [53:0] u_ca_in_820;
wire [53:0] u_ca_in_821;
wire [53:0] u_ca_in_822;
wire [53:0] u_ca_in_823;
wire [53:0] u_ca_in_824;
wire [53:0] u_ca_in_825;
wire [53:0] u_ca_in_826;
wire [53:0] u_ca_in_827;
wire [53:0] u_ca_in_828;
wire [53:0] u_ca_in_829;
wire [53:0] u_ca_in_830;
wire [53:0] u_ca_in_831;
wire [53:0] u_ca_in_832;
wire [53:0] u_ca_in_833;
wire [53:0] u_ca_in_834;
wire [53:0] u_ca_in_835;
wire [53:0] u_ca_in_836;
wire [53:0] u_ca_in_837;
wire [53:0] u_ca_in_838;
wire [53:0] u_ca_in_839;
wire [53:0] u_ca_in_840;
wire [53:0] u_ca_in_841;
wire [53:0] u_ca_in_842;
wire [53:0] u_ca_in_843;
wire [53:0] u_ca_in_844;
wire [53:0] u_ca_in_845;
wire [53:0] u_ca_in_846;
wire [53:0] u_ca_in_847;
wire [53:0] u_ca_in_848;
wire [53:0] u_ca_in_849;
wire [53:0] u_ca_in_850;
wire [53:0] u_ca_in_851;
wire [53:0] u_ca_in_852;
wire [53:0] u_ca_in_853;
wire [53:0] u_ca_in_854;
wire [53:0] u_ca_in_855;
wire [53:0] u_ca_in_856;
wire [53:0] u_ca_in_857;
wire [53:0] u_ca_in_858;
wire [53:0] u_ca_in_859;
wire [53:0] u_ca_in_860;
wire [53:0] u_ca_in_861;
wire [53:0] u_ca_in_862;
wire [53:0] u_ca_in_863;
wire [53:0] u_ca_in_864;
wire [53:0] u_ca_in_865;
wire [53:0] u_ca_in_866;
wire [53:0] u_ca_in_867;
wire [53:0] u_ca_in_868;
wire [53:0] u_ca_in_869;
wire [53:0] u_ca_in_870;
wire [53:0] u_ca_in_871;
wire [53:0] u_ca_in_872;
wire [53:0] u_ca_in_873;
wire [53:0] u_ca_in_874;
wire [53:0] u_ca_in_875;
wire [53:0] u_ca_in_876;
wire [53:0] u_ca_in_877;
wire [53:0] u_ca_in_878;
wire [53:0] u_ca_in_879;
wire [53:0] u_ca_in_880;
wire [53:0] u_ca_in_881;
wire [53:0] u_ca_in_882;
wire [53:0] u_ca_in_883;
wire [53:0] u_ca_in_884;
wire [53:0] u_ca_in_885;
wire [53:0] u_ca_in_886;
wire [53:0] u_ca_in_887;
wire [53:0] u_ca_in_888;
wire [53:0] u_ca_in_889;
wire [53:0] u_ca_in_890;
wire [53:0] u_ca_in_891;
wire [53:0] u_ca_in_892;
wire [53:0] u_ca_in_893;
wire [53:0] u_ca_in_894;
wire [53:0] u_ca_in_895;
wire [53:0] u_ca_in_896;
wire [53:0] u_ca_in_897;
wire [53:0] u_ca_in_898;
wire [53:0] u_ca_in_899;
wire [53:0] u_ca_in_900;
wire [53:0] u_ca_in_901;
wire [53:0] u_ca_in_902;
wire [53:0] u_ca_in_903;
wire [53:0] u_ca_in_904;
wire [53:0] u_ca_in_905;
wire [53:0] u_ca_in_906;
wire [53:0] u_ca_in_907;
wire [53:0] u_ca_in_908;
wire [53:0] u_ca_in_909;
wire [53:0] u_ca_in_910;
wire [53:0] u_ca_in_911;
wire [53:0] u_ca_in_912;
wire [53:0] u_ca_in_913;
wire [53:0] u_ca_in_914;
wire [53:0] u_ca_in_915;
wire [53:0] u_ca_in_916;
wire [53:0] u_ca_in_917;
wire [53:0] u_ca_in_918;
wire [53:0] u_ca_in_919;
wire [53:0] u_ca_in_920;
wire [53:0] u_ca_in_921;
wire [53:0] u_ca_in_922;
wire [53:0] u_ca_in_923;
wire [53:0] u_ca_in_924;
wire [53:0] u_ca_in_925;
wire [53:0] u_ca_in_926;
wire [53:0] u_ca_in_927;
wire [53:0] u_ca_in_928;
wire [53:0] u_ca_in_929;
wire [53:0] u_ca_in_930;
wire [53:0] u_ca_in_931;
wire [53:0] u_ca_in_932;
wire [53:0] u_ca_in_933;
wire [53:0] u_ca_in_934;
wire [53:0] u_ca_in_935;
wire [53:0] u_ca_in_936;
wire [53:0] u_ca_in_937;
wire [53:0] u_ca_in_938;
wire [53:0] u_ca_in_939;
wire [53:0] u_ca_in_940;
wire [53:0] u_ca_in_941;
wire [53:0] u_ca_in_942;
wire [53:0] u_ca_in_943;
wire [53:0] u_ca_in_944;
wire [53:0] u_ca_in_945;
wire [53:0] u_ca_in_946;
wire [53:0] u_ca_in_947;
wire [53:0] u_ca_in_948;
wire [53:0] u_ca_in_949;
wire [53:0] u_ca_in_950;
wire [53:0] u_ca_in_951;
wire [53:0] u_ca_in_952;
wire [53:0] u_ca_in_953;
wire [53:0] u_ca_in_954;
wire [53:0] u_ca_in_955;
wire [53:0] u_ca_in_956;
wire [53:0] u_ca_in_957;
wire [53:0] u_ca_in_958;
wire [53:0] u_ca_in_959;
wire [53:0] u_ca_in_960;
wire [53:0] u_ca_in_961;
wire [53:0] u_ca_in_962;
wire [53:0] u_ca_in_963;
wire [53:0] u_ca_in_964;
wire [53:0] u_ca_in_965;
wire [53:0] u_ca_in_966;
wire [53:0] u_ca_in_967;
wire [53:0] u_ca_in_968;
wire [53:0] u_ca_in_969;
wire [53:0] u_ca_in_970;
wire [53:0] u_ca_in_971;
wire [53:0] u_ca_in_972;
wire [53:0] u_ca_in_973;
wire [53:0] u_ca_in_974;
wire [53:0] u_ca_in_975;
wire [53:0] u_ca_in_976;
wire [53:0] u_ca_in_977;
wire [53:0] u_ca_in_978;
wire [53:0] u_ca_in_979;
wire [53:0] u_ca_in_980;
wire [53:0] u_ca_in_981;
wire [53:0] u_ca_in_982;
wire [53:0] u_ca_in_983;
wire [53:0] u_ca_in_984;
wire [53:0] u_ca_in_985;
wire [53:0] u_ca_in_986;
wire [53:0] u_ca_in_987;
wire [53:0] u_ca_in_988;
wire [53:0] u_ca_in_989;
wire [53:0] u_ca_in_990;
wire [53:0] u_ca_in_991;
wire [53:0] u_ca_in_992;
wire [53:0] u_ca_in_993;
wire [53:0] u_ca_in_994;
wire [53:0] u_ca_in_995;
wire [53:0] u_ca_in_996;
wire [53:0] u_ca_in_997;
wire [53:0] u_ca_in_998;
wire [53:0] u_ca_in_999;
wire [53:0] u_ca_in_1000;
wire [53:0] u_ca_in_1001;
wire [53:0] u_ca_in_1002;
wire [53:0] u_ca_in_1003;
wire [53:0] u_ca_in_1004;
wire [53:0] u_ca_in_1005;
wire [53:0] u_ca_in_1006;
wire [53:0] u_ca_in_1007;
wire [53:0] u_ca_in_1008;
wire [53:0] u_ca_in_1009;
wire [53:0] u_ca_in_1010;
wire [53:0] u_ca_in_1011;
wire [53:0] u_ca_in_1012;
wire [53:0] u_ca_in_1013;
wire [53:0] u_ca_in_1014;
wire [53:0] u_ca_in_1015;
wire [53:0] u_ca_in_1016;
wire [53:0] u_ca_in_1017;
wire [53:0] u_ca_in_1018;
wire [53:0] u_ca_in_1019;
wire [53:0] u_ca_in_1020;
wire [53:0] u_ca_in_1021;
wire [53:0] u_ca_in_1022;
wire [53:0] u_ca_in_1023;
wire [53:0] u_ca_in_1024;
wire [53:0] u_ca_in_1025;
wire [53:0] u_ca_in_1026;
wire [53:0] u_ca_in_1027;
wire [53:0] u_ca_in_1028;
wire [53:0] u_ca_in_1029;
wire [15:0] u_ca_out_0;
wire [15:0] u_ca_out_1;
wire [15:0] u_ca_out_2;
wire [15:0] u_ca_out_3;
wire [15:0] u_ca_out_4;
wire [15:0] u_ca_out_5;
wire [15:0] u_ca_out_6;
wire [15:0] u_ca_out_7;
wire [15:0] u_ca_out_8;
wire [15:0] u_ca_out_9;
wire [15:0] u_ca_out_10;
wire [15:0] u_ca_out_11;
wire [15:0] u_ca_out_12;
wire [15:0] u_ca_out_13;
wire [15:0] u_ca_out_14;
wire [15:0] u_ca_out_15;
wire [15:0] u_ca_out_16;
wire [15:0] u_ca_out_17;
wire [15:0] u_ca_out_18;
wire [15:0] u_ca_out_19;
wire [15:0] u_ca_out_20;
wire [15:0] u_ca_out_21;
wire [15:0] u_ca_out_22;
wire [15:0] u_ca_out_23;
wire [15:0] u_ca_out_24;
wire [15:0] u_ca_out_25;
wire [15:0] u_ca_out_26;
wire [15:0] u_ca_out_27;
wire [15:0] u_ca_out_28;
wire [15:0] u_ca_out_29;
wire [15:0] u_ca_out_30;
wire [15:0] u_ca_out_31;
wire [15:0] u_ca_out_32;
wire [15:0] u_ca_out_33;
wire [15:0] u_ca_out_34;
wire [15:0] u_ca_out_35;
wire [15:0] u_ca_out_36;
wire [15:0] u_ca_out_37;
wire [15:0] u_ca_out_38;
wire [15:0] u_ca_out_39;
wire [15:0] u_ca_out_40;
wire [15:0] u_ca_out_41;
wire [15:0] u_ca_out_42;
wire [15:0] u_ca_out_43;
wire [15:0] u_ca_out_44;
wire [15:0] u_ca_out_45;
wire [15:0] u_ca_out_46;
wire [15:0] u_ca_out_47;
wire [15:0] u_ca_out_48;
wire [15:0] u_ca_out_49;
wire [15:0] u_ca_out_50;
wire [15:0] u_ca_out_51;
wire [15:0] u_ca_out_52;
wire [15:0] u_ca_out_53;
wire [15:0] u_ca_out_54;
wire [15:0] u_ca_out_55;
wire [15:0] u_ca_out_56;
wire [15:0] u_ca_out_57;
wire [15:0] u_ca_out_58;
wire [15:0] u_ca_out_59;
wire [15:0] u_ca_out_60;
wire [15:0] u_ca_out_61;
wire [15:0] u_ca_out_62;
wire [15:0] u_ca_out_63;
wire [15:0] u_ca_out_64;
wire [15:0] u_ca_out_65;
wire [15:0] u_ca_out_66;
wire [15:0] u_ca_out_67;
wire [15:0] u_ca_out_68;
wire [15:0] u_ca_out_69;
wire [15:0] u_ca_out_70;
wire [15:0] u_ca_out_71;
wire [15:0] u_ca_out_72;
wire [15:0] u_ca_out_73;
wire [15:0] u_ca_out_74;
wire [15:0] u_ca_out_75;
wire [15:0] u_ca_out_76;
wire [15:0] u_ca_out_77;
wire [15:0] u_ca_out_78;
wire [15:0] u_ca_out_79;
wire [15:0] u_ca_out_80;
wire [15:0] u_ca_out_81;
wire [15:0] u_ca_out_82;
wire [15:0] u_ca_out_83;
wire [15:0] u_ca_out_84;
wire [15:0] u_ca_out_85;
wire [15:0] u_ca_out_86;
wire [15:0] u_ca_out_87;
wire [15:0] u_ca_out_88;
wire [15:0] u_ca_out_89;
wire [15:0] u_ca_out_90;
wire [15:0] u_ca_out_91;
wire [15:0] u_ca_out_92;
wire [15:0] u_ca_out_93;
wire [15:0] u_ca_out_94;
wire [15:0] u_ca_out_95;
wire [15:0] u_ca_out_96;
wire [15:0] u_ca_out_97;
wire [15:0] u_ca_out_98;
wire [15:0] u_ca_out_99;
wire [15:0] u_ca_out_100;
wire [15:0] u_ca_out_101;
wire [15:0] u_ca_out_102;
wire [15:0] u_ca_out_103;
wire [15:0] u_ca_out_104;
wire [15:0] u_ca_out_105;
wire [15:0] u_ca_out_106;
wire [15:0] u_ca_out_107;
wire [15:0] u_ca_out_108;
wire [15:0] u_ca_out_109;
wire [15:0] u_ca_out_110;
wire [15:0] u_ca_out_111;
wire [15:0] u_ca_out_112;
wire [15:0] u_ca_out_113;
wire [15:0] u_ca_out_114;
wire [15:0] u_ca_out_115;
wire [15:0] u_ca_out_116;
wire [15:0] u_ca_out_117;
wire [15:0] u_ca_out_118;
wire [15:0] u_ca_out_119;
wire [15:0] u_ca_out_120;
wire [15:0] u_ca_out_121;
wire [15:0] u_ca_out_122;
wire [15:0] u_ca_out_123;
wire [15:0] u_ca_out_124;
wire [15:0] u_ca_out_125;
wire [15:0] u_ca_out_126;
wire [15:0] u_ca_out_127;
wire [15:0] u_ca_out_128;
wire [15:0] u_ca_out_129;
wire [15:0] u_ca_out_130;
wire [15:0] u_ca_out_131;
wire [15:0] u_ca_out_132;
wire [15:0] u_ca_out_133;
wire [15:0] u_ca_out_134;
wire [15:0] u_ca_out_135;
wire [15:0] u_ca_out_136;
wire [15:0] u_ca_out_137;
wire [15:0] u_ca_out_138;
wire [15:0] u_ca_out_139;
wire [15:0] u_ca_out_140;
wire [15:0] u_ca_out_141;
wire [15:0] u_ca_out_142;
wire [15:0] u_ca_out_143;
wire [15:0] u_ca_out_144;
wire [15:0] u_ca_out_145;
wire [15:0] u_ca_out_146;
wire [15:0] u_ca_out_147;
wire [15:0] u_ca_out_148;
wire [15:0] u_ca_out_149;
wire [15:0] u_ca_out_150;
wire [15:0] u_ca_out_151;
wire [15:0] u_ca_out_152;
wire [15:0] u_ca_out_153;
wire [15:0] u_ca_out_154;
wire [15:0] u_ca_out_155;
wire [15:0] u_ca_out_156;
wire [15:0] u_ca_out_157;
wire [15:0] u_ca_out_158;
wire [15:0] u_ca_out_159;
wire [15:0] u_ca_out_160;
wire [15:0] u_ca_out_161;
wire [15:0] u_ca_out_162;
wire [15:0] u_ca_out_163;
wire [15:0] u_ca_out_164;
wire [15:0] u_ca_out_165;
wire [15:0] u_ca_out_166;
wire [15:0] u_ca_out_167;
wire [15:0] u_ca_out_168;
wire [15:0] u_ca_out_169;
wire [15:0] u_ca_out_170;
wire [15:0] u_ca_out_171;
wire [15:0] u_ca_out_172;
wire [15:0] u_ca_out_173;
wire [15:0] u_ca_out_174;
wire [15:0] u_ca_out_175;
wire [15:0] u_ca_out_176;
wire [15:0] u_ca_out_177;
wire [15:0] u_ca_out_178;
wire [15:0] u_ca_out_179;
wire [15:0] u_ca_out_180;
wire [15:0] u_ca_out_181;
wire [15:0] u_ca_out_182;
wire [15:0] u_ca_out_183;
wire [15:0] u_ca_out_184;
wire [15:0] u_ca_out_185;
wire [15:0] u_ca_out_186;
wire [15:0] u_ca_out_187;
wire [15:0] u_ca_out_188;
wire [15:0] u_ca_out_189;
wire [15:0] u_ca_out_190;
wire [15:0] u_ca_out_191;
wire [15:0] u_ca_out_192;
wire [15:0] u_ca_out_193;
wire [15:0] u_ca_out_194;
wire [15:0] u_ca_out_195;
wire [15:0] u_ca_out_196;
wire [15:0] u_ca_out_197;
wire [15:0] u_ca_out_198;
wire [15:0] u_ca_out_199;
wire [15:0] u_ca_out_200;
wire [15:0] u_ca_out_201;
wire [15:0] u_ca_out_202;
wire [15:0] u_ca_out_203;
wire [15:0] u_ca_out_204;
wire [15:0] u_ca_out_205;
wire [15:0] u_ca_out_206;
wire [15:0] u_ca_out_207;
wire [15:0] u_ca_out_208;
wire [15:0] u_ca_out_209;
wire [15:0] u_ca_out_210;
wire [15:0] u_ca_out_211;
wire [15:0] u_ca_out_212;
wire [15:0] u_ca_out_213;
wire [15:0] u_ca_out_214;
wire [15:0] u_ca_out_215;
wire [15:0] u_ca_out_216;
wire [15:0] u_ca_out_217;
wire [15:0] u_ca_out_218;
wire [15:0] u_ca_out_219;
wire [15:0] u_ca_out_220;
wire [15:0] u_ca_out_221;
wire [15:0] u_ca_out_222;
wire [15:0] u_ca_out_223;
wire [15:0] u_ca_out_224;
wire [15:0] u_ca_out_225;
wire [15:0] u_ca_out_226;
wire [15:0] u_ca_out_227;
wire [15:0] u_ca_out_228;
wire [15:0] u_ca_out_229;
wire [15:0] u_ca_out_230;
wire [15:0] u_ca_out_231;
wire [15:0] u_ca_out_232;
wire [15:0] u_ca_out_233;
wire [15:0] u_ca_out_234;
wire [15:0] u_ca_out_235;
wire [15:0] u_ca_out_236;
wire [15:0] u_ca_out_237;
wire [15:0] u_ca_out_238;
wire [15:0] u_ca_out_239;
wire [15:0] u_ca_out_240;
wire [15:0] u_ca_out_241;
wire [15:0] u_ca_out_242;
wire [15:0] u_ca_out_243;
wire [15:0] u_ca_out_244;
wire [15:0] u_ca_out_245;
wire [15:0] u_ca_out_246;
wire [15:0] u_ca_out_247;
wire [15:0] u_ca_out_248;
wire [15:0] u_ca_out_249;
wire [15:0] u_ca_out_250;
wire [15:0] u_ca_out_251;
wire [15:0] u_ca_out_252;
wire [15:0] u_ca_out_253;
wire [15:0] u_ca_out_254;
wire [15:0] u_ca_out_255;
wire [15:0] u_ca_out_256;
wire [15:0] u_ca_out_257;
wire [15:0] u_ca_out_258;
wire [15:0] u_ca_out_259;
wire [15:0] u_ca_out_260;
wire [15:0] u_ca_out_261;
wire [15:0] u_ca_out_262;
wire [15:0] u_ca_out_263;
wire [15:0] u_ca_out_264;
wire [15:0] u_ca_out_265;
wire [15:0] u_ca_out_266;
wire [15:0] u_ca_out_267;
wire [15:0] u_ca_out_268;
wire [15:0] u_ca_out_269;
wire [15:0] u_ca_out_270;
wire [15:0] u_ca_out_271;
wire [15:0] u_ca_out_272;
wire [15:0] u_ca_out_273;
wire [15:0] u_ca_out_274;
wire [15:0] u_ca_out_275;
wire [15:0] u_ca_out_276;
wire [15:0] u_ca_out_277;
wire [15:0] u_ca_out_278;
wire [15:0] u_ca_out_279;
wire [15:0] u_ca_out_280;
wire [15:0] u_ca_out_281;
wire [15:0] u_ca_out_282;
wire [15:0] u_ca_out_283;
wire [15:0] u_ca_out_284;
wire [15:0] u_ca_out_285;
wire [15:0] u_ca_out_286;
wire [15:0] u_ca_out_287;
wire [15:0] u_ca_out_288;
wire [15:0] u_ca_out_289;
wire [15:0] u_ca_out_290;
wire [15:0] u_ca_out_291;
wire [15:0] u_ca_out_292;
wire [15:0] u_ca_out_293;
wire [15:0] u_ca_out_294;
wire [15:0] u_ca_out_295;
wire [15:0] u_ca_out_296;
wire [15:0] u_ca_out_297;
wire [15:0] u_ca_out_298;
wire [15:0] u_ca_out_299;
wire [15:0] u_ca_out_300;
wire [15:0] u_ca_out_301;
wire [15:0] u_ca_out_302;
wire [15:0] u_ca_out_303;
wire [15:0] u_ca_out_304;
wire [15:0] u_ca_out_305;
wire [15:0] u_ca_out_306;
wire [15:0] u_ca_out_307;
wire [15:0] u_ca_out_308;
wire [15:0] u_ca_out_309;
wire [15:0] u_ca_out_310;
wire [15:0] u_ca_out_311;
wire [15:0] u_ca_out_312;
wire [15:0] u_ca_out_313;
wire [15:0] u_ca_out_314;
wire [15:0] u_ca_out_315;
wire [15:0] u_ca_out_316;
wire [15:0] u_ca_out_317;
wire [15:0] u_ca_out_318;
wire [15:0] u_ca_out_319;
wire [15:0] u_ca_out_320;
wire [15:0] u_ca_out_321;
wire [15:0] u_ca_out_322;
wire [15:0] u_ca_out_323;
wire [15:0] u_ca_out_324;
wire [15:0] u_ca_out_325;
wire [15:0] u_ca_out_326;
wire [15:0] u_ca_out_327;
wire [15:0] u_ca_out_328;
wire [15:0] u_ca_out_329;
wire [15:0] u_ca_out_330;
wire [15:0] u_ca_out_331;
wire [15:0] u_ca_out_332;
wire [15:0] u_ca_out_333;
wire [15:0] u_ca_out_334;
wire [15:0] u_ca_out_335;
wire [15:0] u_ca_out_336;
wire [15:0] u_ca_out_337;
wire [15:0] u_ca_out_338;
wire [15:0] u_ca_out_339;
wire [15:0] u_ca_out_340;
wire [15:0] u_ca_out_341;
wire [15:0] u_ca_out_342;
wire [15:0] u_ca_out_343;
wire [15:0] u_ca_out_344;
wire [15:0] u_ca_out_345;
wire [15:0] u_ca_out_346;
wire [15:0] u_ca_out_347;
wire [15:0] u_ca_out_348;
wire [15:0] u_ca_out_349;
wire [15:0] u_ca_out_350;
wire [15:0] u_ca_out_351;
wire [15:0] u_ca_out_352;
wire [15:0] u_ca_out_353;
wire [15:0] u_ca_out_354;
wire [15:0] u_ca_out_355;
wire [15:0] u_ca_out_356;
wire [15:0] u_ca_out_357;
wire [15:0] u_ca_out_358;
wire [15:0] u_ca_out_359;
wire [15:0] u_ca_out_360;
wire [15:0] u_ca_out_361;
wire [15:0] u_ca_out_362;
wire [15:0] u_ca_out_363;
wire [15:0] u_ca_out_364;
wire [15:0] u_ca_out_365;
wire [15:0] u_ca_out_366;
wire [15:0] u_ca_out_367;
wire [15:0] u_ca_out_368;
wire [15:0] u_ca_out_369;
wire [15:0] u_ca_out_370;
wire [15:0] u_ca_out_371;
wire [15:0] u_ca_out_372;
wire [15:0] u_ca_out_373;
wire [15:0] u_ca_out_374;
wire [15:0] u_ca_out_375;
wire [15:0] u_ca_out_376;
wire [15:0] u_ca_out_377;
wire [15:0] u_ca_out_378;
wire [15:0] u_ca_out_379;
wire [15:0] u_ca_out_380;
wire [15:0] u_ca_out_381;
wire [15:0] u_ca_out_382;
wire [15:0] u_ca_out_383;
wire [15:0] u_ca_out_384;
wire [15:0] u_ca_out_385;
wire [15:0] u_ca_out_386;
wire [15:0] u_ca_out_387;
wire [15:0] u_ca_out_388;
wire [15:0] u_ca_out_389;
wire [15:0] u_ca_out_390;
wire [15:0] u_ca_out_391;
wire [15:0] u_ca_out_392;
wire [15:0] u_ca_out_393;
wire [15:0] u_ca_out_394;
wire [15:0] u_ca_out_395;
wire [15:0] u_ca_out_396;
wire [15:0] u_ca_out_397;
wire [15:0] u_ca_out_398;
wire [15:0] u_ca_out_399;
wire [15:0] u_ca_out_400;
wire [15:0] u_ca_out_401;
wire [15:0] u_ca_out_402;
wire [15:0] u_ca_out_403;
wire [15:0] u_ca_out_404;
wire [15:0] u_ca_out_405;
wire [15:0] u_ca_out_406;
wire [15:0] u_ca_out_407;
wire [15:0] u_ca_out_408;
wire [15:0] u_ca_out_409;
wire [15:0] u_ca_out_410;
wire [15:0] u_ca_out_411;
wire [15:0] u_ca_out_412;
wire [15:0] u_ca_out_413;
wire [15:0] u_ca_out_414;
wire [15:0] u_ca_out_415;
wire [15:0] u_ca_out_416;
wire [15:0] u_ca_out_417;
wire [15:0] u_ca_out_418;
wire [15:0] u_ca_out_419;
wire [15:0] u_ca_out_420;
wire [15:0] u_ca_out_421;
wire [15:0] u_ca_out_422;
wire [15:0] u_ca_out_423;
wire [15:0] u_ca_out_424;
wire [15:0] u_ca_out_425;
wire [15:0] u_ca_out_426;
wire [15:0] u_ca_out_427;
wire [15:0] u_ca_out_428;
wire [15:0] u_ca_out_429;
wire [15:0] u_ca_out_430;
wire [15:0] u_ca_out_431;
wire [15:0] u_ca_out_432;
wire [15:0] u_ca_out_433;
wire [15:0] u_ca_out_434;
wire [15:0] u_ca_out_435;
wire [15:0] u_ca_out_436;
wire [15:0] u_ca_out_437;
wire [15:0] u_ca_out_438;
wire [15:0] u_ca_out_439;
wire [15:0] u_ca_out_440;
wire [15:0] u_ca_out_441;
wire [15:0] u_ca_out_442;
wire [15:0] u_ca_out_443;
wire [15:0] u_ca_out_444;
wire [15:0] u_ca_out_445;
wire [15:0] u_ca_out_446;
wire [15:0] u_ca_out_447;
wire [15:0] u_ca_out_448;
wire [15:0] u_ca_out_449;
wire [15:0] u_ca_out_450;
wire [15:0] u_ca_out_451;
wire [15:0] u_ca_out_452;
wire [15:0] u_ca_out_453;
wire [15:0] u_ca_out_454;
wire [15:0] u_ca_out_455;
wire [15:0] u_ca_out_456;
wire [15:0] u_ca_out_457;
wire [15:0] u_ca_out_458;
wire [15:0] u_ca_out_459;
wire [15:0] u_ca_out_460;
wire [15:0] u_ca_out_461;
wire [15:0] u_ca_out_462;
wire [15:0] u_ca_out_463;
wire [15:0] u_ca_out_464;
wire [15:0] u_ca_out_465;
wire [15:0] u_ca_out_466;
wire [15:0] u_ca_out_467;
wire [15:0] u_ca_out_468;
wire [15:0] u_ca_out_469;
wire [15:0] u_ca_out_470;
wire [15:0] u_ca_out_471;
wire [15:0] u_ca_out_472;
wire [15:0] u_ca_out_473;
wire [15:0] u_ca_out_474;
wire [15:0] u_ca_out_475;
wire [15:0] u_ca_out_476;
wire [15:0] u_ca_out_477;
wire [15:0] u_ca_out_478;
wire [15:0] u_ca_out_479;
wire [15:0] u_ca_out_480;
wire [15:0] u_ca_out_481;
wire [15:0] u_ca_out_482;
wire [15:0] u_ca_out_483;
wire [15:0] u_ca_out_484;
wire [15:0] u_ca_out_485;
wire [15:0] u_ca_out_486;
wire [15:0] u_ca_out_487;
wire [15:0] u_ca_out_488;
wire [15:0] u_ca_out_489;
wire [15:0] u_ca_out_490;
wire [15:0] u_ca_out_491;
wire [15:0] u_ca_out_492;
wire [15:0] u_ca_out_493;
wire [15:0] u_ca_out_494;
wire [15:0] u_ca_out_495;
wire [15:0] u_ca_out_496;
wire [15:0] u_ca_out_497;
wire [15:0] u_ca_out_498;
wire [15:0] u_ca_out_499;
wire [15:0] u_ca_out_500;
wire [15:0] u_ca_out_501;
wire [15:0] u_ca_out_502;
wire [15:0] u_ca_out_503;
wire [15:0] u_ca_out_504;
wire [15:0] u_ca_out_505;
wire [15:0] u_ca_out_506;
wire [15:0] u_ca_out_507;
wire [15:0] u_ca_out_508;
wire [15:0] u_ca_out_509;
wire [15:0] u_ca_out_510;
wire [15:0] u_ca_out_511;
wire [15:0] u_ca_out_512;
wire [15:0] u_ca_out_513;
wire [15:0] u_ca_out_514;
wire [15:0] u_ca_out_515;
wire [15:0] u_ca_out_516;
wire [15:0] u_ca_out_517;
wire [15:0] u_ca_out_518;
wire [15:0] u_ca_out_519;
wire [15:0] u_ca_out_520;
wire [15:0] u_ca_out_521;
wire [15:0] u_ca_out_522;
wire [15:0] u_ca_out_523;
wire [15:0] u_ca_out_524;
wire [15:0] u_ca_out_525;
wire [15:0] u_ca_out_526;
wire [15:0] u_ca_out_527;
wire [15:0] u_ca_out_528;
wire [15:0] u_ca_out_529;
wire [15:0] u_ca_out_530;
wire [15:0] u_ca_out_531;
wire [15:0] u_ca_out_532;
wire [15:0] u_ca_out_533;
wire [15:0] u_ca_out_534;
wire [15:0] u_ca_out_535;
wire [15:0] u_ca_out_536;
wire [15:0] u_ca_out_537;
wire [15:0] u_ca_out_538;
wire [15:0] u_ca_out_539;
wire [15:0] u_ca_out_540;
wire [15:0] u_ca_out_541;
wire [15:0] u_ca_out_542;
wire [15:0] u_ca_out_543;
wire [15:0] u_ca_out_544;
wire [15:0] u_ca_out_545;
wire [15:0] u_ca_out_546;
wire [15:0] u_ca_out_547;
wire [15:0] u_ca_out_548;
wire [15:0] u_ca_out_549;
wire [15:0] u_ca_out_550;
wire [15:0] u_ca_out_551;
wire [15:0] u_ca_out_552;
wire [15:0] u_ca_out_553;
wire [15:0] u_ca_out_554;
wire [15:0] u_ca_out_555;
wire [15:0] u_ca_out_556;
wire [15:0] u_ca_out_557;
wire [15:0] u_ca_out_558;
wire [15:0] u_ca_out_559;
wire [15:0] u_ca_out_560;
wire [15:0] u_ca_out_561;
wire [15:0] u_ca_out_562;
wire [15:0] u_ca_out_563;
wire [15:0] u_ca_out_564;
wire [15:0] u_ca_out_565;
wire [15:0] u_ca_out_566;
wire [15:0] u_ca_out_567;
wire [15:0] u_ca_out_568;
wire [15:0] u_ca_out_569;
wire [15:0] u_ca_out_570;
wire [15:0] u_ca_out_571;
wire [15:0] u_ca_out_572;
wire [15:0] u_ca_out_573;
wire [15:0] u_ca_out_574;
wire [15:0] u_ca_out_575;
wire [15:0] u_ca_out_576;
wire [15:0] u_ca_out_577;
wire [15:0] u_ca_out_578;
wire [15:0] u_ca_out_579;
wire [15:0] u_ca_out_580;
wire [15:0] u_ca_out_581;
wire [15:0] u_ca_out_582;
wire [15:0] u_ca_out_583;
wire [15:0] u_ca_out_584;
wire [15:0] u_ca_out_585;
wire [15:0] u_ca_out_586;
wire [15:0] u_ca_out_587;
wire [15:0] u_ca_out_588;
wire [15:0] u_ca_out_589;
wire [15:0] u_ca_out_590;
wire [15:0] u_ca_out_591;
wire [15:0] u_ca_out_592;
wire [15:0] u_ca_out_593;
wire [15:0] u_ca_out_594;
wire [15:0] u_ca_out_595;
wire [15:0] u_ca_out_596;
wire [15:0] u_ca_out_597;
wire [15:0] u_ca_out_598;
wire [15:0] u_ca_out_599;
wire [15:0] u_ca_out_600;
wire [15:0] u_ca_out_601;
wire [15:0] u_ca_out_602;
wire [15:0] u_ca_out_603;
wire [15:0] u_ca_out_604;
wire [15:0] u_ca_out_605;
wire [15:0] u_ca_out_606;
wire [15:0] u_ca_out_607;
wire [15:0] u_ca_out_608;
wire [15:0] u_ca_out_609;
wire [15:0] u_ca_out_610;
wire [15:0] u_ca_out_611;
wire [15:0] u_ca_out_612;
wire [15:0] u_ca_out_613;
wire [15:0] u_ca_out_614;
wire [15:0] u_ca_out_615;
wire [15:0] u_ca_out_616;
wire [15:0] u_ca_out_617;
wire [15:0] u_ca_out_618;
wire [15:0] u_ca_out_619;
wire [15:0] u_ca_out_620;
wire [15:0] u_ca_out_621;
wire [15:0] u_ca_out_622;
wire [15:0] u_ca_out_623;
wire [15:0] u_ca_out_624;
wire [15:0] u_ca_out_625;
wire [15:0] u_ca_out_626;
wire [15:0] u_ca_out_627;
wire [15:0] u_ca_out_628;
wire [15:0] u_ca_out_629;
wire [15:0] u_ca_out_630;
wire [15:0] u_ca_out_631;
wire [15:0] u_ca_out_632;
wire [15:0] u_ca_out_633;
wire [15:0] u_ca_out_634;
wire [15:0] u_ca_out_635;
wire [15:0] u_ca_out_636;
wire [15:0] u_ca_out_637;
wire [15:0] u_ca_out_638;
wire [15:0] u_ca_out_639;
wire [15:0] u_ca_out_640;
wire [15:0] u_ca_out_641;
wire [15:0] u_ca_out_642;
wire [15:0] u_ca_out_643;
wire [15:0] u_ca_out_644;
wire [15:0] u_ca_out_645;
wire [15:0] u_ca_out_646;
wire [15:0] u_ca_out_647;
wire [15:0] u_ca_out_648;
wire [15:0] u_ca_out_649;
wire [15:0] u_ca_out_650;
wire [15:0] u_ca_out_651;
wire [15:0] u_ca_out_652;
wire [15:0] u_ca_out_653;
wire [15:0] u_ca_out_654;
wire [15:0] u_ca_out_655;
wire [15:0] u_ca_out_656;
wire [15:0] u_ca_out_657;
wire [15:0] u_ca_out_658;
wire [15:0] u_ca_out_659;
wire [15:0] u_ca_out_660;
wire [15:0] u_ca_out_661;
wire [15:0] u_ca_out_662;
wire [15:0] u_ca_out_663;
wire [15:0] u_ca_out_664;
wire [15:0] u_ca_out_665;
wire [15:0] u_ca_out_666;
wire [15:0] u_ca_out_667;
wire [15:0] u_ca_out_668;
wire [15:0] u_ca_out_669;
wire [15:0] u_ca_out_670;
wire [15:0] u_ca_out_671;
wire [15:0] u_ca_out_672;
wire [15:0] u_ca_out_673;
wire [15:0] u_ca_out_674;
wire [15:0] u_ca_out_675;
wire [15:0] u_ca_out_676;
wire [15:0] u_ca_out_677;
wire [15:0] u_ca_out_678;
wire [15:0] u_ca_out_679;
wire [15:0] u_ca_out_680;
wire [15:0] u_ca_out_681;
wire [15:0] u_ca_out_682;
wire [15:0] u_ca_out_683;
wire [15:0] u_ca_out_684;
wire [15:0] u_ca_out_685;
wire [15:0] u_ca_out_686;
wire [15:0] u_ca_out_687;
wire [15:0] u_ca_out_688;
wire [15:0] u_ca_out_689;
wire [15:0] u_ca_out_690;
wire [15:0] u_ca_out_691;
wire [15:0] u_ca_out_692;
wire [15:0] u_ca_out_693;
wire [15:0] u_ca_out_694;
wire [15:0] u_ca_out_695;
wire [15:0] u_ca_out_696;
wire [15:0] u_ca_out_697;
wire [15:0] u_ca_out_698;
wire [15:0] u_ca_out_699;
wire [15:0] u_ca_out_700;
wire [15:0] u_ca_out_701;
wire [15:0] u_ca_out_702;
wire [15:0] u_ca_out_703;
wire [15:0] u_ca_out_704;
wire [15:0] u_ca_out_705;
wire [15:0] u_ca_out_706;
wire [15:0] u_ca_out_707;
wire [15:0] u_ca_out_708;
wire [15:0] u_ca_out_709;
wire [15:0] u_ca_out_710;
wire [15:0] u_ca_out_711;
wire [15:0] u_ca_out_712;
wire [15:0] u_ca_out_713;
wire [15:0] u_ca_out_714;
wire [15:0] u_ca_out_715;
wire [15:0] u_ca_out_716;
wire [15:0] u_ca_out_717;
wire [15:0] u_ca_out_718;
wire [15:0] u_ca_out_719;
wire [15:0] u_ca_out_720;
wire [15:0] u_ca_out_721;
wire [15:0] u_ca_out_722;
wire [15:0] u_ca_out_723;
wire [15:0] u_ca_out_724;
wire [15:0] u_ca_out_725;
wire [15:0] u_ca_out_726;
wire [15:0] u_ca_out_727;
wire [15:0] u_ca_out_728;
wire [15:0] u_ca_out_729;
wire [15:0] u_ca_out_730;
wire [15:0] u_ca_out_731;
wire [15:0] u_ca_out_732;
wire [15:0] u_ca_out_733;
wire [15:0] u_ca_out_734;
wire [15:0] u_ca_out_735;
wire [15:0] u_ca_out_736;
wire [15:0] u_ca_out_737;
wire [15:0] u_ca_out_738;
wire [15:0] u_ca_out_739;
wire [15:0] u_ca_out_740;
wire [15:0] u_ca_out_741;
wire [15:0] u_ca_out_742;
wire [15:0] u_ca_out_743;
wire [15:0] u_ca_out_744;
wire [15:0] u_ca_out_745;
wire [15:0] u_ca_out_746;
wire [15:0] u_ca_out_747;
wire [15:0] u_ca_out_748;
wire [15:0] u_ca_out_749;
wire [15:0] u_ca_out_750;
wire [15:0] u_ca_out_751;
wire [15:0] u_ca_out_752;
wire [15:0] u_ca_out_753;
wire [15:0] u_ca_out_754;
wire [15:0] u_ca_out_755;
wire [15:0] u_ca_out_756;
wire [15:0] u_ca_out_757;
wire [15:0] u_ca_out_758;
wire [15:0] u_ca_out_759;
wire [15:0] u_ca_out_760;
wire [15:0] u_ca_out_761;
wire [15:0] u_ca_out_762;
wire [15:0] u_ca_out_763;
wire [15:0] u_ca_out_764;
wire [15:0] u_ca_out_765;
wire [15:0] u_ca_out_766;
wire [15:0] u_ca_out_767;
wire [15:0] u_ca_out_768;
wire [15:0] u_ca_out_769;
wire [15:0] u_ca_out_770;
wire [15:0] u_ca_out_771;
wire [15:0] u_ca_out_772;
wire [15:0] u_ca_out_773;
wire [15:0] u_ca_out_774;
wire [15:0] u_ca_out_775;
wire [15:0] u_ca_out_776;
wire [15:0] u_ca_out_777;
wire [15:0] u_ca_out_778;
wire [15:0] u_ca_out_779;
wire [15:0] u_ca_out_780;
wire [15:0] u_ca_out_781;
wire [15:0] u_ca_out_782;
wire [15:0] u_ca_out_783;
wire [15:0] u_ca_out_784;
wire [15:0] u_ca_out_785;
wire [15:0] u_ca_out_786;
wire [15:0] u_ca_out_787;
wire [15:0] u_ca_out_788;
wire [15:0] u_ca_out_789;
wire [15:0] u_ca_out_790;
wire [15:0] u_ca_out_791;
wire [15:0] u_ca_out_792;
wire [15:0] u_ca_out_793;
wire [15:0] u_ca_out_794;
wire [15:0] u_ca_out_795;
wire [15:0] u_ca_out_796;
wire [15:0] u_ca_out_797;
wire [15:0] u_ca_out_798;
wire [15:0] u_ca_out_799;
wire [15:0] u_ca_out_800;
wire [15:0] u_ca_out_801;
wire [15:0] u_ca_out_802;
wire [15:0] u_ca_out_803;
wire [15:0] u_ca_out_804;
wire [15:0] u_ca_out_805;
wire [15:0] u_ca_out_806;
wire [15:0] u_ca_out_807;
wire [15:0] u_ca_out_808;
wire [15:0] u_ca_out_809;
wire [15:0] u_ca_out_810;
wire [15:0] u_ca_out_811;
wire [15:0] u_ca_out_812;
wire [15:0] u_ca_out_813;
wire [15:0] u_ca_out_814;
wire [15:0] u_ca_out_815;
wire [15:0] u_ca_out_816;
wire [15:0] u_ca_out_817;
wire [15:0] u_ca_out_818;
wire [15:0] u_ca_out_819;
wire [15:0] u_ca_out_820;
wire [15:0] u_ca_out_821;
wire [15:0] u_ca_out_822;
wire [15:0] u_ca_out_823;
wire [15:0] u_ca_out_824;
wire [15:0] u_ca_out_825;
wire [15:0] u_ca_out_826;
wire [15:0] u_ca_out_827;
wire [15:0] u_ca_out_828;
wire [15:0] u_ca_out_829;
wire [15:0] u_ca_out_830;
wire [15:0] u_ca_out_831;
wire [15:0] u_ca_out_832;
wire [15:0] u_ca_out_833;
wire [15:0] u_ca_out_834;
wire [15:0] u_ca_out_835;
wire [15:0] u_ca_out_836;
wire [15:0] u_ca_out_837;
wire [15:0] u_ca_out_838;
wire [15:0] u_ca_out_839;
wire [15:0] u_ca_out_840;
wire [15:0] u_ca_out_841;
wire [15:0] u_ca_out_842;
wire [15:0] u_ca_out_843;
wire [15:0] u_ca_out_844;
wire [15:0] u_ca_out_845;
wire [15:0] u_ca_out_846;
wire [15:0] u_ca_out_847;
wire [15:0] u_ca_out_848;
wire [15:0] u_ca_out_849;
wire [15:0] u_ca_out_850;
wire [15:0] u_ca_out_851;
wire [15:0] u_ca_out_852;
wire [15:0] u_ca_out_853;
wire [15:0] u_ca_out_854;
wire [15:0] u_ca_out_855;
wire [15:0] u_ca_out_856;
wire [15:0] u_ca_out_857;
wire [15:0] u_ca_out_858;
wire [15:0] u_ca_out_859;
wire [15:0] u_ca_out_860;
wire [15:0] u_ca_out_861;
wire [15:0] u_ca_out_862;
wire [15:0] u_ca_out_863;
wire [15:0] u_ca_out_864;
wire [15:0] u_ca_out_865;
wire [15:0] u_ca_out_866;
wire [15:0] u_ca_out_867;
wire [15:0] u_ca_out_868;
wire [15:0] u_ca_out_869;
wire [15:0] u_ca_out_870;
wire [15:0] u_ca_out_871;
wire [15:0] u_ca_out_872;
wire [15:0] u_ca_out_873;
wire [15:0] u_ca_out_874;
wire [15:0] u_ca_out_875;
wire [15:0] u_ca_out_876;
wire [15:0] u_ca_out_877;
wire [15:0] u_ca_out_878;
wire [15:0] u_ca_out_879;
wire [15:0] u_ca_out_880;
wire [15:0] u_ca_out_881;
wire [15:0] u_ca_out_882;
wire [15:0] u_ca_out_883;
wire [15:0] u_ca_out_884;
wire [15:0] u_ca_out_885;
wire [15:0] u_ca_out_886;
wire [15:0] u_ca_out_887;
wire [15:0] u_ca_out_888;
wire [15:0] u_ca_out_889;
wire [15:0] u_ca_out_890;
wire [15:0] u_ca_out_891;
wire [15:0] u_ca_out_892;
wire [15:0] u_ca_out_893;
wire [15:0] u_ca_out_894;
wire [15:0] u_ca_out_895;
wire [15:0] u_ca_out_896;
wire [15:0] u_ca_out_897;
wire [15:0] u_ca_out_898;
wire [15:0] u_ca_out_899;
wire [15:0] u_ca_out_900;
wire [15:0] u_ca_out_901;
wire [15:0] u_ca_out_902;
wire [15:0] u_ca_out_903;
wire [15:0] u_ca_out_904;
wire [15:0] u_ca_out_905;
wire [15:0] u_ca_out_906;
wire [15:0] u_ca_out_907;
wire [15:0] u_ca_out_908;
wire [15:0] u_ca_out_909;
wire [15:0] u_ca_out_910;
wire [15:0] u_ca_out_911;
wire [15:0] u_ca_out_912;
wire [15:0] u_ca_out_913;
wire [15:0] u_ca_out_914;
wire [15:0] u_ca_out_915;
wire [15:0] u_ca_out_916;
wire [15:0] u_ca_out_917;
wire [15:0] u_ca_out_918;
wire [15:0] u_ca_out_919;
wire [15:0] u_ca_out_920;
wire [15:0] u_ca_out_921;
wire [15:0] u_ca_out_922;
wire [15:0] u_ca_out_923;
wire [15:0] u_ca_out_924;
wire [15:0] u_ca_out_925;
wire [15:0] u_ca_out_926;
wire [15:0] u_ca_out_927;
wire [15:0] u_ca_out_928;
wire [15:0] u_ca_out_929;
wire [15:0] u_ca_out_930;
wire [15:0] u_ca_out_931;
wire [15:0] u_ca_out_932;
wire [15:0] u_ca_out_933;
wire [15:0] u_ca_out_934;
wire [15:0] u_ca_out_935;
wire [15:0] u_ca_out_936;
wire [15:0] u_ca_out_937;
wire [15:0] u_ca_out_938;
wire [15:0] u_ca_out_939;
wire [15:0] u_ca_out_940;
wire [15:0] u_ca_out_941;
wire [15:0] u_ca_out_942;
wire [15:0] u_ca_out_943;
wire [15:0] u_ca_out_944;
wire [15:0] u_ca_out_945;
wire [15:0] u_ca_out_946;
wire [15:0] u_ca_out_947;
wire [15:0] u_ca_out_948;
wire [15:0] u_ca_out_949;
wire [15:0] u_ca_out_950;
wire [15:0] u_ca_out_951;
wire [15:0] u_ca_out_952;
wire [15:0] u_ca_out_953;
wire [15:0] u_ca_out_954;
wire [15:0] u_ca_out_955;
wire [15:0] u_ca_out_956;
wire [15:0] u_ca_out_957;
wire [15:0] u_ca_out_958;
wire [15:0] u_ca_out_959;
wire [15:0] u_ca_out_960;
wire [15:0] u_ca_out_961;
wire [15:0] u_ca_out_962;
wire [15:0] u_ca_out_963;
wire [15:0] u_ca_out_964;
wire [15:0] u_ca_out_965;
wire [15:0] u_ca_out_966;
wire [15:0] u_ca_out_967;
wire [15:0] u_ca_out_968;
wire [15:0] u_ca_out_969;
wire [15:0] u_ca_out_970;
wire [15:0] u_ca_out_971;
wire [15:0] u_ca_out_972;
wire [15:0] u_ca_out_973;
wire [15:0] u_ca_out_974;
wire [15:0] u_ca_out_975;
wire [15:0] u_ca_out_976;
wire [15:0] u_ca_out_977;
wire [15:0] u_ca_out_978;
wire [15:0] u_ca_out_979;
wire [15:0] u_ca_out_980;
wire [15:0] u_ca_out_981;
wire [15:0] u_ca_out_982;
wire [15:0] u_ca_out_983;
wire [15:0] u_ca_out_984;
wire [15:0] u_ca_out_985;
wire [15:0] u_ca_out_986;
wire [15:0] u_ca_out_987;
wire [15:0] u_ca_out_988;
wire [15:0] u_ca_out_989;
wire [15:0] u_ca_out_990;
wire [15:0] u_ca_out_991;
wire [15:0] u_ca_out_992;
wire [15:0] u_ca_out_993;
wire [15:0] u_ca_out_994;
wire [15:0] u_ca_out_995;
wire [15:0] u_ca_out_996;
wire [15:0] u_ca_out_997;
wire [15:0] u_ca_out_998;
wire [15:0] u_ca_out_999;
wire [15:0] u_ca_out_1000;
wire [15:0] u_ca_out_1001;
wire [15:0] u_ca_out_1002;
wire [15:0] u_ca_out_1003;
wire [15:0] u_ca_out_1004;
wire [15:0] u_ca_out_1005;
wire [15:0] u_ca_out_1006;
wire [15:0] u_ca_out_1007;
wire [15:0] u_ca_out_1008;
wire [15:0] u_ca_out_1009;
wire [15:0] u_ca_out_1010;
wire [15:0] u_ca_out_1011;
wire [15:0] u_ca_out_1012;
wire [15:0] u_ca_out_1013;
wire [15:0] u_ca_out_1014;
wire [15:0] u_ca_out_1015;
wire [15:0] u_ca_out_1016;
wire [15:0] u_ca_out_1017;
wire [15:0] u_ca_out_1018;
wire [15:0] u_ca_out_1019;
wire [15:0] u_ca_out_1020;
wire [15:0] u_ca_out_1021;
wire [15:0] u_ca_out_1022;
wire [15:0] u_ca_out_1023;
wire [15:0] u_ca_out_1024;
wire [15:0] u_ca_out_1025;
wire [15:0] u_ca_out_1026;
wire [15:0] u_ca_out_1027;
wire [15:0] u_ca_out_1028;
wire [15:0] u_ca_out_1029;

assign u_ca_in_0 = {{6{1'b0}}, col_in_0};
assign u_ca_in_1 = {{6{1'b0}}, col_in_1};
assign u_ca_in_2 = {{6{1'b0}}, col_in_2};
assign u_ca_in_3 = {{6{1'b0}}, col_in_3};
assign u_ca_in_4 = {{6{1'b0}}, col_in_4};
assign u_ca_in_5 = {{6{1'b0}}, col_in_5};
assign u_ca_in_6 = {{6{1'b0}}, col_in_6};
assign u_ca_in_7 = {{6{1'b0}}, col_in_7};
assign u_ca_in_8 = {{6{1'b0}}, col_in_8};
assign u_ca_in_9 = {{6{1'b0}}, col_in_9};
assign u_ca_in_10 = {{6{1'b0}}, col_in_10};
assign u_ca_in_11 = {{6{1'b0}}, col_in_11};
assign u_ca_in_12 = {{6{1'b0}}, col_in_12};
assign u_ca_in_13 = {{6{1'b0}}, col_in_13};
assign u_ca_in_14 = {{6{1'b0}}, col_in_14};
assign u_ca_in_15 = {{6{1'b0}}, col_in_15};
assign u_ca_in_16 = {{6{1'b0}}, col_in_16};
assign u_ca_in_17 = {{6{1'b0}}, col_in_17};
assign u_ca_in_18 = {{6{1'b0}}, col_in_18};
assign u_ca_in_19 = {{6{1'b0}}, col_in_19};
assign u_ca_in_20 = {{6{1'b0}}, col_in_20};
assign u_ca_in_21 = {{6{1'b0}}, col_in_21};
assign u_ca_in_22 = {{6{1'b0}}, col_in_22};
assign u_ca_in_23 = {{6{1'b0}}, col_in_23};
assign u_ca_in_24 = {{6{1'b0}}, col_in_24};
assign u_ca_in_25 = {{6{1'b0}}, col_in_25};
assign u_ca_in_26 = {{6{1'b0}}, col_in_26};
assign u_ca_in_27 = {{6{1'b0}}, col_in_27};
assign u_ca_in_28 = {{6{1'b0}}, col_in_28};
assign u_ca_in_29 = {{6{1'b0}}, col_in_29};
assign u_ca_in_30 = {{6{1'b0}}, col_in_30};
assign u_ca_in_31 = {{6{1'b0}}, col_in_31};
assign u_ca_in_32 = {{6{1'b0}}, col_in_32};
assign u_ca_in_33 = {{6{1'b0}}, col_in_33};
assign u_ca_in_34 = {{6{1'b0}}, col_in_34};
assign u_ca_in_35 = {{6{1'b0}}, col_in_35};
assign u_ca_in_36 = {{6{1'b0}}, col_in_36};
assign u_ca_in_37 = {{6{1'b0}}, col_in_37};
assign u_ca_in_38 = {{6{1'b0}}, col_in_38};
assign u_ca_in_39 = {{6{1'b0}}, col_in_39};
assign u_ca_in_40 = {{6{1'b0}}, col_in_40};
assign u_ca_in_41 = {{6{1'b0}}, col_in_41};
assign u_ca_in_42 = {{6{1'b0}}, col_in_42};
assign u_ca_in_43 = {{6{1'b0}}, col_in_43};
assign u_ca_in_44 = {{6{1'b0}}, col_in_44};
assign u_ca_in_45 = {{6{1'b0}}, col_in_45};
assign u_ca_in_46 = {{6{1'b0}}, col_in_46};
assign u_ca_in_47 = {{6{1'b0}}, col_in_47};
assign u_ca_in_48 = {{6{1'b0}}, col_in_48};
assign u_ca_in_49 = {{6{1'b0}}, col_in_49};
assign u_ca_in_50 = {{6{1'b0}}, col_in_50};
assign u_ca_in_51 = {{6{1'b0}}, col_in_51};
assign u_ca_in_52 = {{6{1'b0}}, col_in_52};
assign u_ca_in_53 = {{6{1'b0}}, col_in_53};
assign u_ca_in_54 = {{6{1'b0}}, col_in_54};
assign u_ca_in_55 = {{6{1'b0}}, col_in_55};
assign u_ca_in_56 = {{6{1'b0}}, col_in_56};
assign u_ca_in_57 = {{6{1'b0}}, col_in_57};
assign u_ca_in_58 = {{6{1'b0}}, col_in_58};
assign u_ca_in_59 = {{6{1'b0}}, col_in_59};
assign u_ca_in_60 = {{6{1'b0}}, col_in_60};
assign u_ca_in_61 = {{6{1'b0}}, col_in_61};
assign u_ca_in_62 = {{6{1'b0}}, col_in_62};
assign u_ca_in_63 = {{6{1'b0}}, col_in_63};
assign u_ca_in_64 = {{6{1'b0}}, col_in_64};
assign u_ca_in_65 = {{6{1'b0}}, col_in_65};
assign u_ca_in_66 = {{6{1'b0}}, col_in_66};
assign u_ca_in_67 = {{6{1'b0}}, col_in_67};
assign u_ca_in_68 = {{6{1'b0}}, col_in_68};
assign u_ca_in_69 = {{6{1'b0}}, col_in_69};
assign u_ca_in_70 = {{6{1'b0}}, col_in_70};
assign u_ca_in_71 = {{6{1'b0}}, col_in_71};
assign u_ca_in_72 = {{6{1'b0}}, col_in_72};
assign u_ca_in_73 = {{6{1'b0}}, col_in_73};
assign u_ca_in_74 = {{6{1'b0}}, col_in_74};
assign u_ca_in_75 = {{6{1'b0}}, col_in_75};
assign u_ca_in_76 = {{6{1'b0}}, col_in_76};
assign u_ca_in_77 = {{6{1'b0}}, col_in_77};
assign u_ca_in_78 = {{6{1'b0}}, col_in_78};
assign u_ca_in_79 = {{6{1'b0}}, col_in_79};
assign u_ca_in_80 = {{6{1'b0}}, col_in_80};
assign u_ca_in_81 = {{6{1'b0}}, col_in_81};
assign u_ca_in_82 = {{6{1'b0}}, col_in_82};
assign u_ca_in_83 = {{6{1'b0}}, col_in_83};
assign u_ca_in_84 = {{6{1'b0}}, col_in_84};
assign u_ca_in_85 = {{6{1'b0}}, col_in_85};
assign u_ca_in_86 = {{6{1'b0}}, col_in_86};
assign u_ca_in_87 = {{6{1'b0}}, col_in_87};
assign u_ca_in_88 = {{6{1'b0}}, col_in_88};
assign u_ca_in_89 = {{6{1'b0}}, col_in_89};
assign u_ca_in_90 = {{6{1'b0}}, col_in_90};
assign u_ca_in_91 = {{6{1'b0}}, col_in_91};
assign u_ca_in_92 = {{6{1'b0}}, col_in_92};
assign u_ca_in_93 = {{6{1'b0}}, col_in_93};
assign u_ca_in_94 = {{6{1'b0}}, col_in_94};
assign u_ca_in_95 = {{6{1'b0}}, col_in_95};
assign u_ca_in_96 = {{6{1'b0}}, col_in_96};
assign u_ca_in_97 = {{6{1'b0}}, col_in_97};
assign u_ca_in_98 = {{6{1'b0}}, col_in_98};
assign u_ca_in_99 = {{6{1'b0}}, col_in_99};
assign u_ca_in_100 = {{6{1'b0}}, col_in_100};
assign u_ca_in_101 = {{6{1'b0}}, col_in_101};
assign u_ca_in_102 = {{6{1'b0}}, col_in_102};
assign u_ca_in_103 = {{6{1'b0}}, col_in_103};
assign u_ca_in_104 = {{6{1'b0}}, col_in_104};
assign u_ca_in_105 = {{6{1'b0}}, col_in_105};
assign u_ca_in_106 = {{6{1'b0}}, col_in_106};
assign u_ca_in_107 = {{6{1'b0}}, col_in_107};
assign u_ca_in_108 = {{6{1'b0}}, col_in_108};
assign u_ca_in_109 = {{6{1'b0}}, col_in_109};
assign u_ca_in_110 = {{6{1'b0}}, col_in_110};
assign u_ca_in_111 = {{6{1'b0}}, col_in_111};
assign u_ca_in_112 = {{6{1'b0}}, col_in_112};
assign u_ca_in_113 = {{6{1'b0}}, col_in_113};
assign u_ca_in_114 = {{6{1'b0}}, col_in_114};
assign u_ca_in_115 = {{6{1'b0}}, col_in_115};
assign u_ca_in_116 = {{6{1'b0}}, col_in_116};
assign u_ca_in_117 = {{6{1'b0}}, col_in_117};
assign u_ca_in_118 = {{6{1'b0}}, col_in_118};
assign u_ca_in_119 = {{6{1'b0}}, col_in_119};
assign u_ca_in_120 = {{6{1'b0}}, col_in_120};
assign u_ca_in_121 = {{6{1'b0}}, col_in_121};
assign u_ca_in_122 = {{6{1'b0}}, col_in_122};
assign u_ca_in_123 = {{6{1'b0}}, col_in_123};
assign u_ca_in_124 = {{6{1'b0}}, col_in_124};
assign u_ca_in_125 = {{6{1'b0}}, col_in_125};
assign u_ca_in_126 = {{6{1'b0}}, col_in_126};
assign u_ca_in_127 = {{6{1'b0}}, col_in_127};
assign u_ca_in_128 = {{6{1'b0}}, col_in_128};
assign u_ca_in_129 = {{6{1'b0}}, col_in_129};
assign u_ca_in_130 = {{6{1'b0}}, col_in_130};
assign u_ca_in_131 = {{6{1'b0}}, col_in_131};
assign u_ca_in_132 = {{6{1'b0}}, col_in_132};
assign u_ca_in_133 = {{6{1'b0}}, col_in_133};
assign u_ca_in_134 = {{6{1'b0}}, col_in_134};
assign u_ca_in_135 = {{6{1'b0}}, col_in_135};
assign u_ca_in_136 = {{6{1'b0}}, col_in_136};
assign u_ca_in_137 = {{6{1'b0}}, col_in_137};
assign u_ca_in_138 = {{6{1'b0}}, col_in_138};
assign u_ca_in_139 = {{6{1'b0}}, col_in_139};
assign u_ca_in_140 = {{6{1'b0}}, col_in_140};
assign u_ca_in_141 = {{6{1'b0}}, col_in_141};
assign u_ca_in_142 = {{6{1'b0}}, col_in_142};
assign u_ca_in_143 = {{6{1'b0}}, col_in_143};
assign u_ca_in_144 = {{6{1'b0}}, col_in_144};
assign u_ca_in_145 = {{6{1'b0}}, col_in_145};
assign u_ca_in_146 = {{6{1'b0}}, col_in_146};
assign u_ca_in_147 = {{6{1'b0}}, col_in_147};
assign u_ca_in_148 = {{6{1'b0}}, col_in_148};
assign u_ca_in_149 = {{6{1'b0}}, col_in_149};
assign u_ca_in_150 = {{6{1'b0}}, col_in_150};
assign u_ca_in_151 = {{6{1'b0}}, col_in_151};
assign u_ca_in_152 = {{6{1'b0}}, col_in_152};
assign u_ca_in_153 = {{6{1'b0}}, col_in_153};
assign u_ca_in_154 = {{6{1'b0}}, col_in_154};
assign u_ca_in_155 = {{6{1'b0}}, col_in_155};
assign u_ca_in_156 = {{6{1'b0}}, col_in_156};
assign u_ca_in_157 = {{6{1'b0}}, col_in_157};
assign u_ca_in_158 = {{6{1'b0}}, col_in_158};
assign u_ca_in_159 = {{6{1'b0}}, col_in_159};
assign u_ca_in_160 = {{6{1'b0}}, col_in_160};
assign u_ca_in_161 = {{6{1'b0}}, col_in_161};
assign u_ca_in_162 = {{6{1'b0}}, col_in_162};
assign u_ca_in_163 = {{6{1'b0}}, col_in_163};
assign u_ca_in_164 = {{6{1'b0}}, col_in_164};
assign u_ca_in_165 = {{6{1'b0}}, col_in_165};
assign u_ca_in_166 = {{6{1'b0}}, col_in_166};
assign u_ca_in_167 = {{6{1'b0}}, col_in_167};
assign u_ca_in_168 = {{6{1'b0}}, col_in_168};
assign u_ca_in_169 = {{6{1'b0}}, col_in_169};
assign u_ca_in_170 = {{6{1'b0}}, col_in_170};
assign u_ca_in_171 = {{6{1'b0}}, col_in_171};
assign u_ca_in_172 = {{6{1'b0}}, col_in_172};
assign u_ca_in_173 = {{6{1'b0}}, col_in_173};
assign u_ca_in_174 = {{6{1'b0}}, col_in_174};
assign u_ca_in_175 = {{6{1'b0}}, col_in_175};
assign u_ca_in_176 = {{6{1'b0}}, col_in_176};
assign u_ca_in_177 = {{6{1'b0}}, col_in_177};
assign u_ca_in_178 = {{6{1'b0}}, col_in_178};
assign u_ca_in_179 = {{6{1'b0}}, col_in_179};
assign u_ca_in_180 = {{6{1'b0}}, col_in_180};
assign u_ca_in_181 = {{6{1'b0}}, col_in_181};
assign u_ca_in_182 = {{6{1'b0}}, col_in_182};
assign u_ca_in_183 = {{6{1'b0}}, col_in_183};
assign u_ca_in_184 = {{6{1'b0}}, col_in_184};
assign u_ca_in_185 = {{6{1'b0}}, col_in_185};
assign u_ca_in_186 = {{6{1'b0}}, col_in_186};
assign u_ca_in_187 = {{6{1'b0}}, col_in_187};
assign u_ca_in_188 = {{6{1'b0}}, col_in_188};
assign u_ca_in_189 = {{6{1'b0}}, col_in_189};
assign u_ca_in_190 = {{6{1'b0}}, col_in_190};
assign u_ca_in_191 = {{6{1'b0}}, col_in_191};
assign u_ca_in_192 = {{6{1'b0}}, col_in_192};
assign u_ca_in_193 = {{6{1'b0}}, col_in_193};
assign u_ca_in_194 = {{6{1'b0}}, col_in_194};
assign u_ca_in_195 = {{6{1'b0}}, col_in_195};
assign u_ca_in_196 = {{6{1'b0}}, col_in_196};
assign u_ca_in_197 = {{6{1'b0}}, col_in_197};
assign u_ca_in_198 = {{6{1'b0}}, col_in_198};
assign u_ca_in_199 = {{6{1'b0}}, col_in_199};
assign u_ca_in_200 = {{6{1'b0}}, col_in_200};
assign u_ca_in_201 = {{6{1'b0}}, col_in_201};
assign u_ca_in_202 = {{6{1'b0}}, col_in_202};
assign u_ca_in_203 = {{6{1'b0}}, col_in_203};
assign u_ca_in_204 = {{6{1'b0}}, col_in_204};
assign u_ca_in_205 = {{6{1'b0}}, col_in_205};
assign u_ca_in_206 = {{6{1'b0}}, col_in_206};
assign u_ca_in_207 = {{6{1'b0}}, col_in_207};
assign u_ca_in_208 = {{6{1'b0}}, col_in_208};
assign u_ca_in_209 = {{6{1'b0}}, col_in_209};
assign u_ca_in_210 = {{6{1'b0}}, col_in_210};
assign u_ca_in_211 = {{6{1'b0}}, col_in_211};
assign u_ca_in_212 = {{6{1'b0}}, col_in_212};
assign u_ca_in_213 = {{6{1'b0}}, col_in_213};
assign u_ca_in_214 = {{6{1'b0}}, col_in_214};
assign u_ca_in_215 = {{6{1'b0}}, col_in_215};
assign u_ca_in_216 = {{6{1'b0}}, col_in_216};
assign u_ca_in_217 = {{6{1'b0}}, col_in_217};
assign u_ca_in_218 = {{6{1'b0}}, col_in_218};
assign u_ca_in_219 = {{6{1'b0}}, col_in_219};
assign u_ca_in_220 = {{6{1'b0}}, col_in_220};
assign u_ca_in_221 = {{6{1'b0}}, col_in_221};
assign u_ca_in_222 = {{6{1'b0}}, col_in_222};
assign u_ca_in_223 = {{6{1'b0}}, col_in_223};
assign u_ca_in_224 = {{6{1'b0}}, col_in_224};
assign u_ca_in_225 = {{6{1'b0}}, col_in_225};
assign u_ca_in_226 = {{6{1'b0}}, col_in_226};
assign u_ca_in_227 = {{6{1'b0}}, col_in_227};
assign u_ca_in_228 = {{6{1'b0}}, col_in_228};
assign u_ca_in_229 = {{6{1'b0}}, col_in_229};
assign u_ca_in_230 = {{6{1'b0}}, col_in_230};
assign u_ca_in_231 = {{6{1'b0}}, col_in_231};
assign u_ca_in_232 = {{6{1'b0}}, col_in_232};
assign u_ca_in_233 = {{6{1'b0}}, col_in_233};
assign u_ca_in_234 = {{6{1'b0}}, col_in_234};
assign u_ca_in_235 = {{6{1'b0}}, col_in_235};
assign u_ca_in_236 = {{6{1'b0}}, col_in_236};
assign u_ca_in_237 = {{6{1'b0}}, col_in_237};
assign u_ca_in_238 = {{6{1'b0}}, col_in_238};
assign u_ca_in_239 = {{6{1'b0}}, col_in_239};
assign u_ca_in_240 = {{6{1'b0}}, col_in_240};
assign u_ca_in_241 = {{6{1'b0}}, col_in_241};
assign u_ca_in_242 = {{6{1'b0}}, col_in_242};
assign u_ca_in_243 = {{6{1'b0}}, col_in_243};
assign u_ca_in_244 = {{6{1'b0}}, col_in_244};
assign u_ca_in_245 = {{6{1'b0}}, col_in_245};
assign u_ca_in_246 = {{6{1'b0}}, col_in_246};
assign u_ca_in_247 = {{6{1'b0}}, col_in_247};
assign u_ca_in_248 = {{6{1'b0}}, col_in_248};
assign u_ca_in_249 = {{6{1'b0}}, col_in_249};
assign u_ca_in_250 = {{6{1'b0}}, col_in_250};
assign u_ca_in_251 = {{6{1'b0}}, col_in_251};
assign u_ca_in_252 = {{6{1'b0}}, col_in_252};
assign u_ca_in_253 = {{6{1'b0}}, col_in_253};
assign u_ca_in_254 = {{6{1'b0}}, col_in_254};
assign u_ca_in_255 = {{6{1'b0}}, col_in_255};
assign u_ca_in_256 = {{6{1'b0}}, col_in_256};
assign u_ca_in_257 = {{6{1'b0}}, col_in_257};
assign u_ca_in_258 = {{6{1'b0}}, col_in_258};
assign u_ca_in_259 = {{6{1'b0}}, col_in_259};
assign u_ca_in_260 = {{6{1'b0}}, col_in_260};
assign u_ca_in_261 = {{6{1'b0}}, col_in_261};
assign u_ca_in_262 = {{6{1'b0}}, col_in_262};
assign u_ca_in_263 = {{6{1'b0}}, col_in_263};
assign u_ca_in_264 = {{6{1'b0}}, col_in_264};
assign u_ca_in_265 = {{6{1'b0}}, col_in_265};
assign u_ca_in_266 = {{6{1'b0}}, col_in_266};
assign u_ca_in_267 = {{6{1'b0}}, col_in_267};
assign u_ca_in_268 = {{6{1'b0}}, col_in_268};
assign u_ca_in_269 = {{6{1'b0}}, col_in_269};
assign u_ca_in_270 = {{6{1'b0}}, col_in_270};
assign u_ca_in_271 = {{6{1'b0}}, col_in_271};
assign u_ca_in_272 = {{6{1'b0}}, col_in_272};
assign u_ca_in_273 = {{6{1'b0}}, col_in_273};
assign u_ca_in_274 = {{6{1'b0}}, col_in_274};
assign u_ca_in_275 = {{6{1'b0}}, col_in_275};
assign u_ca_in_276 = {{6{1'b0}}, col_in_276};
assign u_ca_in_277 = {{6{1'b0}}, col_in_277};
assign u_ca_in_278 = {{6{1'b0}}, col_in_278};
assign u_ca_in_279 = {{6{1'b0}}, col_in_279};
assign u_ca_in_280 = {{6{1'b0}}, col_in_280};
assign u_ca_in_281 = {{6{1'b0}}, col_in_281};
assign u_ca_in_282 = {{6{1'b0}}, col_in_282};
assign u_ca_in_283 = {{6{1'b0}}, col_in_283};
assign u_ca_in_284 = {{6{1'b0}}, col_in_284};
assign u_ca_in_285 = {{6{1'b0}}, col_in_285};
assign u_ca_in_286 = {{6{1'b0}}, col_in_286};
assign u_ca_in_287 = {{6{1'b0}}, col_in_287};
assign u_ca_in_288 = {{6{1'b0}}, col_in_288};
assign u_ca_in_289 = {{6{1'b0}}, col_in_289};
assign u_ca_in_290 = {{6{1'b0}}, col_in_290};
assign u_ca_in_291 = {{6{1'b0}}, col_in_291};
assign u_ca_in_292 = {{6{1'b0}}, col_in_292};
assign u_ca_in_293 = {{6{1'b0}}, col_in_293};
assign u_ca_in_294 = {{6{1'b0}}, col_in_294};
assign u_ca_in_295 = {{6{1'b0}}, col_in_295};
assign u_ca_in_296 = {{6{1'b0}}, col_in_296};
assign u_ca_in_297 = {{6{1'b0}}, col_in_297};
assign u_ca_in_298 = {{6{1'b0}}, col_in_298};
assign u_ca_in_299 = {{6{1'b0}}, col_in_299};
assign u_ca_in_300 = {{6{1'b0}}, col_in_300};
assign u_ca_in_301 = {{6{1'b0}}, col_in_301};
assign u_ca_in_302 = {{6{1'b0}}, col_in_302};
assign u_ca_in_303 = {{6{1'b0}}, col_in_303};
assign u_ca_in_304 = {{6{1'b0}}, col_in_304};
assign u_ca_in_305 = {{6{1'b0}}, col_in_305};
assign u_ca_in_306 = {{6{1'b0}}, col_in_306};
assign u_ca_in_307 = {{6{1'b0}}, col_in_307};
assign u_ca_in_308 = {{6{1'b0}}, col_in_308};
assign u_ca_in_309 = {{6{1'b0}}, col_in_309};
assign u_ca_in_310 = {{6{1'b0}}, col_in_310};
assign u_ca_in_311 = {{6{1'b0}}, col_in_311};
assign u_ca_in_312 = {{6{1'b0}}, col_in_312};
assign u_ca_in_313 = {{6{1'b0}}, col_in_313};
assign u_ca_in_314 = {{6{1'b0}}, col_in_314};
assign u_ca_in_315 = {{6{1'b0}}, col_in_315};
assign u_ca_in_316 = {{6{1'b0}}, col_in_316};
assign u_ca_in_317 = {{6{1'b0}}, col_in_317};
assign u_ca_in_318 = {{6{1'b0}}, col_in_318};
assign u_ca_in_319 = {{6{1'b0}}, col_in_319};
assign u_ca_in_320 = {{6{1'b0}}, col_in_320};
assign u_ca_in_321 = {{6{1'b0}}, col_in_321};
assign u_ca_in_322 = {{6{1'b0}}, col_in_322};
assign u_ca_in_323 = {{6{1'b0}}, col_in_323};
assign u_ca_in_324 = {{6{1'b0}}, col_in_324};
assign u_ca_in_325 = {{6{1'b0}}, col_in_325};
assign u_ca_in_326 = {{6{1'b0}}, col_in_326};
assign u_ca_in_327 = {{6{1'b0}}, col_in_327};
assign u_ca_in_328 = {{6{1'b0}}, col_in_328};
assign u_ca_in_329 = {{6{1'b0}}, col_in_329};
assign u_ca_in_330 = {{6{1'b0}}, col_in_330};
assign u_ca_in_331 = {{6{1'b0}}, col_in_331};
assign u_ca_in_332 = {{6{1'b0}}, col_in_332};
assign u_ca_in_333 = {{6{1'b0}}, col_in_333};
assign u_ca_in_334 = {{6{1'b0}}, col_in_334};
assign u_ca_in_335 = {{6{1'b0}}, col_in_335};
assign u_ca_in_336 = {{6{1'b0}}, col_in_336};
assign u_ca_in_337 = {{6{1'b0}}, col_in_337};
assign u_ca_in_338 = {{6{1'b0}}, col_in_338};
assign u_ca_in_339 = {{6{1'b0}}, col_in_339};
assign u_ca_in_340 = {{6{1'b0}}, col_in_340};
assign u_ca_in_341 = {{6{1'b0}}, col_in_341};
assign u_ca_in_342 = {{6{1'b0}}, col_in_342};
assign u_ca_in_343 = {{6{1'b0}}, col_in_343};
assign u_ca_in_344 = {{6{1'b0}}, col_in_344};
assign u_ca_in_345 = {{6{1'b0}}, col_in_345};
assign u_ca_in_346 = {{6{1'b0}}, col_in_346};
assign u_ca_in_347 = {{6{1'b0}}, col_in_347};
assign u_ca_in_348 = {{6{1'b0}}, col_in_348};
assign u_ca_in_349 = {{6{1'b0}}, col_in_349};
assign u_ca_in_350 = {{6{1'b0}}, col_in_350};
assign u_ca_in_351 = {{6{1'b0}}, col_in_351};
assign u_ca_in_352 = {{6{1'b0}}, col_in_352};
assign u_ca_in_353 = {{6{1'b0}}, col_in_353};
assign u_ca_in_354 = {{6{1'b0}}, col_in_354};
assign u_ca_in_355 = {{6{1'b0}}, col_in_355};
assign u_ca_in_356 = {{6{1'b0}}, col_in_356};
assign u_ca_in_357 = {{6{1'b0}}, col_in_357};
assign u_ca_in_358 = {{6{1'b0}}, col_in_358};
assign u_ca_in_359 = {{6{1'b0}}, col_in_359};
assign u_ca_in_360 = {{6{1'b0}}, col_in_360};
assign u_ca_in_361 = {{6{1'b0}}, col_in_361};
assign u_ca_in_362 = {{6{1'b0}}, col_in_362};
assign u_ca_in_363 = {{6{1'b0}}, col_in_363};
assign u_ca_in_364 = {{6{1'b0}}, col_in_364};
assign u_ca_in_365 = {{6{1'b0}}, col_in_365};
assign u_ca_in_366 = {{6{1'b0}}, col_in_366};
assign u_ca_in_367 = {{6{1'b0}}, col_in_367};
assign u_ca_in_368 = {{6{1'b0}}, col_in_368};
assign u_ca_in_369 = {{6{1'b0}}, col_in_369};
assign u_ca_in_370 = {{6{1'b0}}, col_in_370};
assign u_ca_in_371 = {{6{1'b0}}, col_in_371};
assign u_ca_in_372 = {{6{1'b0}}, col_in_372};
assign u_ca_in_373 = {{6{1'b0}}, col_in_373};
assign u_ca_in_374 = {{6{1'b0}}, col_in_374};
assign u_ca_in_375 = {{6{1'b0}}, col_in_375};
assign u_ca_in_376 = {{6{1'b0}}, col_in_376};
assign u_ca_in_377 = {{6{1'b0}}, col_in_377};
assign u_ca_in_378 = {{6{1'b0}}, col_in_378};
assign u_ca_in_379 = {{6{1'b0}}, col_in_379};
assign u_ca_in_380 = {{6{1'b0}}, col_in_380};
assign u_ca_in_381 = {{6{1'b0}}, col_in_381};
assign u_ca_in_382 = {{6{1'b0}}, col_in_382};
assign u_ca_in_383 = {{6{1'b0}}, col_in_383};
assign u_ca_in_384 = {{6{1'b0}}, col_in_384};
assign u_ca_in_385 = {{6{1'b0}}, col_in_385};
assign u_ca_in_386 = {{6{1'b0}}, col_in_386};
assign u_ca_in_387 = {{6{1'b0}}, col_in_387};
assign u_ca_in_388 = {{6{1'b0}}, col_in_388};
assign u_ca_in_389 = {{6{1'b0}}, col_in_389};
assign u_ca_in_390 = {{6{1'b0}}, col_in_390};
assign u_ca_in_391 = {{6{1'b0}}, col_in_391};
assign u_ca_in_392 = {{6{1'b0}}, col_in_392};
assign u_ca_in_393 = {{6{1'b0}}, col_in_393};
assign u_ca_in_394 = {{6{1'b0}}, col_in_394};
assign u_ca_in_395 = {{6{1'b0}}, col_in_395};
assign u_ca_in_396 = {{6{1'b0}}, col_in_396};
assign u_ca_in_397 = {{6{1'b0}}, col_in_397};
assign u_ca_in_398 = {{6{1'b0}}, col_in_398};
assign u_ca_in_399 = {{6{1'b0}}, col_in_399};
assign u_ca_in_400 = {{6{1'b0}}, col_in_400};
assign u_ca_in_401 = {{6{1'b0}}, col_in_401};
assign u_ca_in_402 = {{6{1'b0}}, col_in_402};
assign u_ca_in_403 = {{6{1'b0}}, col_in_403};
assign u_ca_in_404 = {{6{1'b0}}, col_in_404};
assign u_ca_in_405 = {{6{1'b0}}, col_in_405};
assign u_ca_in_406 = {{6{1'b0}}, col_in_406};
assign u_ca_in_407 = {{6{1'b0}}, col_in_407};
assign u_ca_in_408 = {{6{1'b0}}, col_in_408};
assign u_ca_in_409 = {{6{1'b0}}, col_in_409};
assign u_ca_in_410 = {{6{1'b0}}, col_in_410};
assign u_ca_in_411 = {{6{1'b0}}, col_in_411};
assign u_ca_in_412 = {{6{1'b0}}, col_in_412};
assign u_ca_in_413 = {{6{1'b0}}, col_in_413};
assign u_ca_in_414 = {{6{1'b0}}, col_in_414};
assign u_ca_in_415 = {{6{1'b0}}, col_in_415};
assign u_ca_in_416 = {{6{1'b0}}, col_in_416};
assign u_ca_in_417 = {{6{1'b0}}, col_in_417};
assign u_ca_in_418 = {{6{1'b0}}, col_in_418};
assign u_ca_in_419 = {{6{1'b0}}, col_in_419};
assign u_ca_in_420 = {{6{1'b0}}, col_in_420};
assign u_ca_in_421 = {{6{1'b0}}, col_in_421};
assign u_ca_in_422 = {{6{1'b0}}, col_in_422};
assign u_ca_in_423 = {{6{1'b0}}, col_in_423};
assign u_ca_in_424 = {{6{1'b0}}, col_in_424};
assign u_ca_in_425 = {{6{1'b0}}, col_in_425};
assign u_ca_in_426 = {{6{1'b0}}, col_in_426};
assign u_ca_in_427 = {{6{1'b0}}, col_in_427};
assign u_ca_in_428 = {{6{1'b0}}, col_in_428};
assign u_ca_in_429 = {{6{1'b0}}, col_in_429};
assign u_ca_in_430 = {{6{1'b0}}, col_in_430};
assign u_ca_in_431 = {{6{1'b0}}, col_in_431};
assign u_ca_in_432 = {{6{1'b0}}, col_in_432};
assign u_ca_in_433 = {{6{1'b0}}, col_in_433};
assign u_ca_in_434 = {{6{1'b0}}, col_in_434};
assign u_ca_in_435 = {{6{1'b0}}, col_in_435};
assign u_ca_in_436 = {{6{1'b0}}, col_in_436};
assign u_ca_in_437 = {{6{1'b0}}, col_in_437};
assign u_ca_in_438 = {{6{1'b0}}, col_in_438};
assign u_ca_in_439 = {{6{1'b0}}, col_in_439};
assign u_ca_in_440 = {{6{1'b0}}, col_in_440};
assign u_ca_in_441 = {{6{1'b0}}, col_in_441};
assign u_ca_in_442 = {{6{1'b0}}, col_in_442};
assign u_ca_in_443 = {{6{1'b0}}, col_in_443};
assign u_ca_in_444 = {{6{1'b0}}, col_in_444};
assign u_ca_in_445 = {{6{1'b0}}, col_in_445};
assign u_ca_in_446 = {{6{1'b0}}, col_in_446};
assign u_ca_in_447 = {{6{1'b0}}, col_in_447};
assign u_ca_in_448 = {{6{1'b0}}, col_in_448};
assign u_ca_in_449 = {{6{1'b0}}, col_in_449};
assign u_ca_in_450 = {{6{1'b0}}, col_in_450};
assign u_ca_in_451 = {{6{1'b0}}, col_in_451};
assign u_ca_in_452 = {{6{1'b0}}, col_in_452};
assign u_ca_in_453 = {{6{1'b0}}, col_in_453};
assign u_ca_in_454 = {{6{1'b0}}, col_in_454};
assign u_ca_in_455 = {{6{1'b0}}, col_in_455};
assign u_ca_in_456 = {{6{1'b0}}, col_in_456};
assign u_ca_in_457 = {{6{1'b0}}, col_in_457};
assign u_ca_in_458 = {{6{1'b0}}, col_in_458};
assign u_ca_in_459 = {{6{1'b0}}, col_in_459};
assign u_ca_in_460 = {{6{1'b0}}, col_in_460};
assign u_ca_in_461 = {{6{1'b0}}, col_in_461};
assign u_ca_in_462 = {{6{1'b0}}, col_in_462};
assign u_ca_in_463 = {{6{1'b0}}, col_in_463};
assign u_ca_in_464 = {{6{1'b0}}, col_in_464};
assign u_ca_in_465 = {{6{1'b0}}, col_in_465};
assign u_ca_in_466 = {{6{1'b0}}, col_in_466};
assign u_ca_in_467 = {{6{1'b0}}, col_in_467};
assign u_ca_in_468 = {{6{1'b0}}, col_in_468};
assign u_ca_in_469 = {{6{1'b0}}, col_in_469};
assign u_ca_in_470 = {{6{1'b0}}, col_in_470};
assign u_ca_in_471 = {{6{1'b0}}, col_in_471};
assign u_ca_in_472 = {{6{1'b0}}, col_in_472};
assign u_ca_in_473 = {{6{1'b0}}, col_in_473};
assign u_ca_in_474 = {{6{1'b0}}, col_in_474};
assign u_ca_in_475 = {{6{1'b0}}, col_in_475};
assign u_ca_in_476 = {{6{1'b0}}, col_in_476};
assign u_ca_in_477 = {{6{1'b0}}, col_in_477};
assign u_ca_in_478 = {{6{1'b0}}, col_in_478};
assign u_ca_in_479 = {{6{1'b0}}, col_in_479};
assign u_ca_in_480 = {{6{1'b0}}, col_in_480};
assign u_ca_in_481 = {{6{1'b0}}, col_in_481};
assign u_ca_in_482 = {{6{1'b0}}, col_in_482};
assign u_ca_in_483 = {{6{1'b0}}, col_in_483};
assign u_ca_in_484 = {{6{1'b0}}, col_in_484};
assign u_ca_in_485 = {{6{1'b0}}, col_in_485};
assign u_ca_in_486 = {{6{1'b0}}, col_in_486};
assign u_ca_in_487 = {{6{1'b0}}, col_in_487};
assign u_ca_in_488 = {{6{1'b0}}, col_in_488};
assign u_ca_in_489 = {{6{1'b0}}, col_in_489};
assign u_ca_in_490 = {{6{1'b0}}, col_in_490};
assign u_ca_in_491 = {{6{1'b0}}, col_in_491};
assign u_ca_in_492 = {{6{1'b0}}, col_in_492};
assign u_ca_in_493 = {{6{1'b0}}, col_in_493};
assign u_ca_in_494 = {{6{1'b0}}, col_in_494};
assign u_ca_in_495 = {{6{1'b0}}, col_in_495};
assign u_ca_in_496 = {{6{1'b0}}, col_in_496};
assign u_ca_in_497 = {{6{1'b0}}, col_in_497};
assign u_ca_in_498 = {{6{1'b0}}, col_in_498};
assign u_ca_in_499 = {{6{1'b0}}, col_in_499};
assign u_ca_in_500 = {{6{1'b0}}, col_in_500};
assign u_ca_in_501 = {{6{1'b0}}, col_in_501};
assign u_ca_in_502 = {{6{1'b0}}, col_in_502};
assign u_ca_in_503 = {{6{1'b0}}, col_in_503};
assign u_ca_in_504 = {{6{1'b0}}, col_in_504};
assign u_ca_in_505 = {{6{1'b0}}, col_in_505};
assign u_ca_in_506 = {{6{1'b0}}, col_in_506};
assign u_ca_in_507 = {{6{1'b0}}, col_in_507};
assign u_ca_in_508 = {{6{1'b0}}, col_in_508};
assign u_ca_in_509 = {{6{1'b0}}, col_in_509};
assign u_ca_in_510 = {{6{1'b0}}, col_in_510};
assign u_ca_in_511 = {{6{1'b0}}, col_in_511};
assign u_ca_in_512 = {{6{1'b0}}, col_in_512};
assign u_ca_in_513 = {{6{1'b0}}, col_in_513};
assign u_ca_in_514 = {{6{1'b0}}, col_in_514};
assign u_ca_in_515 = {{6{1'b0}}, col_in_515};
assign u_ca_in_516 = {{6{1'b0}}, col_in_516};
assign u_ca_in_517 = {{6{1'b0}}, col_in_517};
assign u_ca_in_518 = {{6{1'b0}}, col_in_518};
assign u_ca_in_519 = {{6{1'b0}}, col_in_519};
assign u_ca_in_520 = {{6{1'b0}}, col_in_520};
assign u_ca_in_521 = {{6{1'b0}}, col_in_521};
assign u_ca_in_522 = {{6{1'b0}}, col_in_522};
assign u_ca_in_523 = {{6{1'b0}}, col_in_523};
assign u_ca_in_524 = {{6{1'b0}}, col_in_524};
assign u_ca_in_525 = {{6{1'b0}}, col_in_525};
assign u_ca_in_526 = {{6{1'b0}}, col_in_526};
assign u_ca_in_527 = {{6{1'b0}}, col_in_527};
assign u_ca_in_528 = {{6{1'b0}}, col_in_528};
assign u_ca_in_529 = {{6{1'b0}}, col_in_529};
assign u_ca_in_530 = {{6{1'b0}}, col_in_530};
assign u_ca_in_531 = {{6{1'b0}}, col_in_531};
assign u_ca_in_532 = {{6{1'b0}}, col_in_532};
assign u_ca_in_533 = {{6{1'b0}}, col_in_533};
assign u_ca_in_534 = {{6{1'b0}}, col_in_534};
assign u_ca_in_535 = {{6{1'b0}}, col_in_535};
assign u_ca_in_536 = {{6{1'b0}}, col_in_536};
assign u_ca_in_537 = {{6{1'b0}}, col_in_537};
assign u_ca_in_538 = {{6{1'b0}}, col_in_538};
assign u_ca_in_539 = {{6{1'b0}}, col_in_539};
assign u_ca_in_540 = {{6{1'b0}}, col_in_540};
assign u_ca_in_541 = {{6{1'b0}}, col_in_541};
assign u_ca_in_542 = {{6{1'b0}}, col_in_542};
assign u_ca_in_543 = {{6{1'b0}}, col_in_543};
assign u_ca_in_544 = {{6{1'b0}}, col_in_544};
assign u_ca_in_545 = {{6{1'b0}}, col_in_545};
assign u_ca_in_546 = {{6{1'b0}}, col_in_546};
assign u_ca_in_547 = {{6{1'b0}}, col_in_547};
assign u_ca_in_548 = {{6{1'b0}}, col_in_548};
assign u_ca_in_549 = {{6{1'b0}}, col_in_549};
assign u_ca_in_550 = {{6{1'b0}}, col_in_550};
assign u_ca_in_551 = {{6{1'b0}}, col_in_551};
assign u_ca_in_552 = {{6{1'b0}}, col_in_552};
assign u_ca_in_553 = {{6{1'b0}}, col_in_553};
assign u_ca_in_554 = {{6{1'b0}}, col_in_554};
assign u_ca_in_555 = {{6{1'b0}}, col_in_555};
assign u_ca_in_556 = {{6{1'b0}}, col_in_556};
assign u_ca_in_557 = {{6{1'b0}}, col_in_557};
assign u_ca_in_558 = {{6{1'b0}}, col_in_558};
assign u_ca_in_559 = {{6{1'b0}}, col_in_559};
assign u_ca_in_560 = {{6{1'b0}}, col_in_560};
assign u_ca_in_561 = {{6{1'b0}}, col_in_561};
assign u_ca_in_562 = {{6{1'b0}}, col_in_562};
assign u_ca_in_563 = {{6{1'b0}}, col_in_563};
assign u_ca_in_564 = {{6{1'b0}}, col_in_564};
assign u_ca_in_565 = {{6{1'b0}}, col_in_565};
assign u_ca_in_566 = {{6{1'b0}}, col_in_566};
assign u_ca_in_567 = {{6{1'b0}}, col_in_567};
assign u_ca_in_568 = {{6{1'b0}}, col_in_568};
assign u_ca_in_569 = {{6{1'b0}}, col_in_569};
assign u_ca_in_570 = {{6{1'b0}}, col_in_570};
assign u_ca_in_571 = {{6{1'b0}}, col_in_571};
assign u_ca_in_572 = {{6{1'b0}}, col_in_572};
assign u_ca_in_573 = {{6{1'b0}}, col_in_573};
assign u_ca_in_574 = {{6{1'b0}}, col_in_574};
assign u_ca_in_575 = {{6{1'b0}}, col_in_575};
assign u_ca_in_576 = {{6{1'b0}}, col_in_576};
assign u_ca_in_577 = {{6{1'b0}}, col_in_577};
assign u_ca_in_578 = {{6{1'b0}}, col_in_578};
assign u_ca_in_579 = {{6{1'b0}}, col_in_579};
assign u_ca_in_580 = {{6{1'b0}}, col_in_580};
assign u_ca_in_581 = {{6{1'b0}}, col_in_581};
assign u_ca_in_582 = {{6{1'b0}}, col_in_582};
assign u_ca_in_583 = {{6{1'b0}}, col_in_583};
assign u_ca_in_584 = {{6{1'b0}}, col_in_584};
assign u_ca_in_585 = {{6{1'b0}}, col_in_585};
assign u_ca_in_586 = {{6{1'b0}}, col_in_586};
assign u_ca_in_587 = {{6{1'b0}}, col_in_587};
assign u_ca_in_588 = {{6{1'b0}}, col_in_588};
assign u_ca_in_589 = {{6{1'b0}}, col_in_589};
assign u_ca_in_590 = {{6{1'b0}}, col_in_590};
assign u_ca_in_591 = {{6{1'b0}}, col_in_591};
assign u_ca_in_592 = {{6{1'b0}}, col_in_592};
assign u_ca_in_593 = {{6{1'b0}}, col_in_593};
assign u_ca_in_594 = {{6{1'b0}}, col_in_594};
assign u_ca_in_595 = {{6{1'b0}}, col_in_595};
assign u_ca_in_596 = {{6{1'b0}}, col_in_596};
assign u_ca_in_597 = {{6{1'b0}}, col_in_597};
assign u_ca_in_598 = {{6{1'b0}}, col_in_598};
assign u_ca_in_599 = {{6{1'b0}}, col_in_599};
assign u_ca_in_600 = {{6{1'b0}}, col_in_600};
assign u_ca_in_601 = {{6{1'b0}}, col_in_601};
assign u_ca_in_602 = {{6{1'b0}}, col_in_602};
assign u_ca_in_603 = {{6{1'b0}}, col_in_603};
assign u_ca_in_604 = {{6{1'b0}}, col_in_604};
assign u_ca_in_605 = {{6{1'b0}}, col_in_605};
assign u_ca_in_606 = {{6{1'b0}}, col_in_606};
assign u_ca_in_607 = {{6{1'b0}}, col_in_607};
assign u_ca_in_608 = {{6{1'b0}}, col_in_608};
assign u_ca_in_609 = {{6{1'b0}}, col_in_609};
assign u_ca_in_610 = {{6{1'b0}}, col_in_610};
assign u_ca_in_611 = {{6{1'b0}}, col_in_611};
assign u_ca_in_612 = {{6{1'b0}}, col_in_612};
assign u_ca_in_613 = {{6{1'b0}}, col_in_613};
assign u_ca_in_614 = {{6{1'b0}}, col_in_614};
assign u_ca_in_615 = {{6{1'b0}}, col_in_615};
assign u_ca_in_616 = {{6{1'b0}}, col_in_616};
assign u_ca_in_617 = {{6{1'b0}}, col_in_617};
assign u_ca_in_618 = {{6{1'b0}}, col_in_618};
assign u_ca_in_619 = {{6{1'b0}}, col_in_619};
assign u_ca_in_620 = {{6{1'b0}}, col_in_620};
assign u_ca_in_621 = {{6{1'b0}}, col_in_621};
assign u_ca_in_622 = {{6{1'b0}}, col_in_622};
assign u_ca_in_623 = {{6{1'b0}}, col_in_623};
assign u_ca_in_624 = {{6{1'b0}}, col_in_624};
assign u_ca_in_625 = {{6{1'b0}}, col_in_625};
assign u_ca_in_626 = {{6{1'b0}}, col_in_626};
assign u_ca_in_627 = {{6{1'b0}}, col_in_627};
assign u_ca_in_628 = {{6{1'b0}}, col_in_628};
assign u_ca_in_629 = {{6{1'b0}}, col_in_629};
assign u_ca_in_630 = {{6{1'b0}}, col_in_630};
assign u_ca_in_631 = {{6{1'b0}}, col_in_631};
assign u_ca_in_632 = {{6{1'b0}}, col_in_632};
assign u_ca_in_633 = {{6{1'b0}}, col_in_633};
assign u_ca_in_634 = {{6{1'b0}}, col_in_634};
assign u_ca_in_635 = {{6{1'b0}}, col_in_635};
assign u_ca_in_636 = {{6{1'b0}}, col_in_636};
assign u_ca_in_637 = {{6{1'b0}}, col_in_637};
assign u_ca_in_638 = {{6{1'b0}}, col_in_638};
assign u_ca_in_639 = {{6{1'b0}}, col_in_639};
assign u_ca_in_640 = {{6{1'b0}}, col_in_640};
assign u_ca_in_641 = {{6{1'b0}}, col_in_641};
assign u_ca_in_642 = {{6{1'b0}}, col_in_642};
assign u_ca_in_643 = {{6{1'b0}}, col_in_643};
assign u_ca_in_644 = {{6{1'b0}}, col_in_644};
assign u_ca_in_645 = {{6{1'b0}}, col_in_645};
assign u_ca_in_646 = {{6{1'b0}}, col_in_646};
assign u_ca_in_647 = {{6{1'b0}}, col_in_647};
assign u_ca_in_648 = {{6{1'b0}}, col_in_648};
assign u_ca_in_649 = {{6{1'b0}}, col_in_649};
assign u_ca_in_650 = {{6{1'b0}}, col_in_650};
assign u_ca_in_651 = {{6{1'b0}}, col_in_651};
assign u_ca_in_652 = {{6{1'b0}}, col_in_652};
assign u_ca_in_653 = {{6{1'b0}}, col_in_653};
assign u_ca_in_654 = {{6{1'b0}}, col_in_654};
assign u_ca_in_655 = {{6{1'b0}}, col_in_655};
assign u_ca_in_656 = {{6{1'b0}}, col_in_656};
assign u_ca_in_657 = {{6{1'b0}}, col_in_657};
assign u_ca_in_658 = {{6{1'b0}}, col_in_658};
assign u_ca_in_659 = {{6{1'b0}}, col_in_659};
assign u_ca_in_660 = {{6{1'b0}}, col_in_660};
assign u_ca_in_661 = {{6{1'b0}}, col_in_661};
assign u_ca_in_662 = {{6{1'b0}}, col_in_662};
assign u_ca_in_663 = {{6{1'b0}}, col_in_663};
assign u_ca_in_664 = {{6{1'b0}}, col_in_664};
assign u_ca_in_665 = {{6{1'b0}}, col_in_665};
assign u_ca_in_666 = {{6{1'b0}}, col_in_666};
assign u_ca_in_667 = {{6{1'b0}}, col_in_667};
assign u_ca_in_668 = {{6{1'b0}}, col_in_668};
assign u_ca_in_669 = {{6{1'b0}}, col_in_669};
assign u_ca_in_670 = {{6{1'b0}}, col_in_670};
assign u_ca_in_671 = {{6{1'b0}}, col_in_671};
assign u_ca_in_672 = {{6{1'b0}}, col_in_672};
assign u_ca_in_673 = {{6{1'b0}}, col_in_673};
assign u_ca_in_674 = {{6{1'b0}}, col_in_674};
assign u_ca_in_675 = {{6{1'b0}}, col_in_675};
assign u_ca_in_676 = {{6{1'b0}}, col_in_676};
assign u_ca_in_677 = {{6{1'b0}}, col_in_677};
assign u_ca_in_678 = {{6{1'b0}}, col_in_678};
assign u_ca_in_679 = {{6{1'b0}}, col_in_679};
assign u_ca_in_680 = {{6{1'b0}}, col_in_680};
assign u_ca_in_681 = {{6{1'b0}}, col_in_681};
assign u_ca_in_682 = {{6{1'b0}}, col_in_682};
assign u_ca_in_683 = {{6{1'b0}}, col_in_683};
assign u_ca_in_684 = {{6{1'b0}}, col_in_684};
assign u_ca_in_685 = {{6{1'b0}}, col_in_685};
assign u_ca_in_686 = {{6{1'b0}}, col_in_686};
assign u_ca_in_687 = {{6{1'b0}}, col_in_687};
assign u_ca_in_688 = {{6{1'b0}}, col_in_688};
assign u_ca_in_689 = {{6{1'b0}}, col_in_689};
assign u_ca_in_690 = {{6{1'b0}}, col_in_690};
assign u_ca_in_691 = {{6{1'b0}}, col_in_691};
assign u_ca_in_692 = {{6{1'b0}}, col_in_692};
assign u_ca_in_693 = {{6{1'b0}}, col_in_693};
assign u_ca_in_694 = {{6{1'b0}}, col_in_694};
assign u_ca_in_695 = {{6{1'b0}}, col_in_695};
assign u_ca_in_696 = {{6{1'b0}}, col_in_696};
assign u_ca_in_697 = {{6{1'b0}}, col_in_697};
assign u_ca_in_698 = {{6{1'b0}}, col_in_698};
assign u_ca_in_699 = {{6{1'b0}}, col_in_699};
assign u_ca_in_700 = {{6{1'b0}}, col_in_700};
assign u_ca_in_701 = {{6{1'b0}}, col_in_701};
assign u_ca_in_702 = {{6{1'b0}}, col_in_702};
assign u_ca_in_703 = {{6{1'b0}}, col_in_703};
assign u_ca_in_704 = {{6{1'b0}}, col_in_704};
assign u_ca_in_705 = {{6{1'b0}}, col_in_705};
assign u_ca_in_706 = {{6{1'b0}}, col_in_706};
assign u_ca_in_707 = {{6{1'b0}}, col_in_707};
assign u_ca_in_708 = {{6{1'b0}}, col_in_708};
assign u_ca_in_709 = {{6{1'b0}}, col_in_709};
assign u_ca_in_710 = {{6{1'b0}}, col_in_710};
assign u_ca_in_711 = {{6{1'b0}}, col_in_711};
assign u_ca_in_712 = {{6{1'b0}}, col_in_712};
assign u_ca_in_713 = {{6{1'b0}}, col_in_713};
assign u_ca_in_714 = {{6{1'b0}}, col_in_714};
assign u_ca_in_715 = {{6{1'b0}}, col_in_715};
assign u_ca_in_716 = {{6{1'b0}}, col_in_716};
assign u_ca_in_717 = {{6{1'b0}}, col_in_717};
assign u_ca_in_718 = {{6{1'b0}}, col_in_718};
assign u_ca_in_719 = {{6{1'b0}}, col_in_719};
assign u_ca_in_720 = {{6{1'b0}}, col_in_720};
assign u_ca_in_721 = {{6{1'b0}}, col_in_721};
assign u_ca_in_722 = {{6{1'b0}}, col_in_722};
assign u_ca_in_723 = {{6{1'b0}}, col_in_723};
assign u_ca_in_724 = {{6{1'b0}}, col_in_724};
assign u_ca_in_725 = {{6{1'b0}}, col_in_725};
assign u_ca_in_726 = {{6{1'b0}}, col_in_726};
assign u_ca_in_727 = {{6{1'b0}}, col_in_727};
assign u_ca_in_728 = {{6{1'b0}}, col_in_728};
assign u_ca_in_729 = {{6{1'b0}}, col_in_729};
assign u_ca_in_730 = {{6{1'b0}}, col_in_730};
assign u_ca_in_731 = {{6{1'b0}}, col_in_731};
assign u_ca_in_732 = {{6{1'b0}}, col_in_732};
assign u_ca_in_733 = {{6{1'b0}}, col_in_733};
assign u_ca_in_734 = {{6{1'b0}}, col_in_734};
assign u_ca_in_735 = {{6{1'b0}}, col_in_735};
assign u_ca_in_736 = {{6{1'b0}}, col_in_736};
assign u_ca_in_737 = {{6{1'b0}}, col_in_737};
assign u_ca_in_738 = {{6{1'b0}}, col_in_738};
assign u_ca_in_739 = {{6{1'b0}}, col_in_739};
assign u_ca_in_740 = {{6{1'b0}}, col_in_740};
assign u_ca_in_741 = {{6{1'b0}}, col_in_741};
assign u_ca_in_742 = {{6{1'b0}}, col_in_742};
assign u_ca_in_743 = {{6{1'b0}}, col_in_743};
assign u_ca_in_744 = {{6{1'b0}}, col_in_744};
assign u_ca_in_745 = {{6{1'b0}}, col_in_745};
assign u_ca_in_746 = {{6{1'b0}}, col_in_746};
assign u_ca_in_747 = {{6{1'b0}}, col_in_747};
assign u_ca_in_748 = {{6{1'b0}}, col_in_748};
assign u_ca_in_749 = {{6{1'b0}}, col_in_749};
assign u_ca_in_750 = {{6{1'b0}}, col_in_750};
assign u_ca_in_751 = {{6{1'b0}}, col_in_751};
assign u_ca_in_752 = {{6{1'b0}}, col_in_752};
assign u_ca_in_753 = {{6{1'b0}}, col_in_753};
assign u_ca_in_754 = {{6{1'b0}}, col_in_754};
assign u_ca_in_755 = {{6{1'b0}}, col_in_755};
assign u_ca_in_756 = {{6{1'b0}}, col_in_756};
assign u_ca_in_757 = {{6{1'b0}}, col_in_757};
assign u_ca_in_758 = {{6{1'b0}}, col_in_758};
assign u_ca_in_759 = {{6{1'b0}}, col_in_759};
assign u_ca_in_760 = {{6{1'b0}}, col_in_760};
assign u_ca_in_761 = {{6{1'b0}}, col_in_761};
assign u_ca_in_762 = {{6{1'b0}}, col_in_762};
assign u_ca_in_763 = {{6{1'b0}}, col_in_763};
assign u_ca_in_764 = {{6{1'b0}}, col_in_764};
assign u_ca_in_765 = {{6{1'b0}}, col_in_765};
assign u_ca_in_766 = {{6{1'b0}}, col_in_766};
assign u_ca_in_767 = {{6{1'b0}}, col_in_767};
assign u_ca_in_768 = {{6{1'b0}}, col_in_768};
assign u_ca_in_769 = {{6{1'b0}}, col_in_769};
assign u_ca_in_770 = {{6{1'b0}}, col_in_770};
assign u_ca_in_771 = {{6{1'b0}}, col_in_771};
assign u_ca_in_772 = {{6{1'b0}}, col_in_772};
assign u_ca_in_773 = {{6{1'b0}}, col_in_773};
assign u_ca_in_774 = {{6{1'b0}}, col_in_774};
assign u_ca_in_775 = {{6{1'b0}}, col_in_775};
assign u_ca_in_776 = {{6{1'b0}}, col_in_776};
assign u_ca_in_777 = {{6{1'b0}}, col_in_777};
assign u_ca_in_778 = {{6{1'b0}}, col_in_778};
assign u_ca_in_779 = {{6{1'b0}}, col_in_779};
assign u_ca_in_780 = {{6{1'b0}}, col_in_780};
assign u_ca_in_781 = {{6{1'b0}}, col_in_781};
assign u_ca_in_782 = {{6{1'b0}}, col_in_782};
assign u_ca_in_783 = {{6{1'b0}}, col_in_783};
assign u_ca_in_784 = {{6{1'b0}}, col_in_784};
assign u_ca_in_785 = {{6{1'b0}}, col_in_785};
assign u_ca_in_786 = {{6{1'b0}}, col_in_786};
assign u_ca_in_787 = {{6{1'b0}}, col_in_787};
assign u_ca_in_788 = {{6{1'b0}}, col_in_788};
assign u_ca_in_789 = {{6{1'b0}}, col_in_789};
assign u_ca_in_790 = {{6{1'b0}}, col_in_790};
assign u_ca_in_791 = {{6{1'b0}}, col_in_791};
assign u_ca_in_792 = {{6{1'b0}}, col_in_792};
assign u_ca_in_793 = {{6{1'b0}}, col_in_793};
assign u_ca_in_794 = {{6{1'b0}}, col_in_794};
assign u_ca_in_795 = {{6{1'b0}}, col_in_795};
assign u_ca_in_796 = {{6{1'b0}}, col_in_796};
assign u_ca_in_797 = {{6{1'b0}}, col_in_797};
assign u_ca_in_798 = {{6{1'b0}}, col_in_798};
assign u_ca_in_799 = {{6{1'b0}}, col_in_799};
assign u_ca_in_800 = {{6{1'b0}}, col_in_800};
assign u_ca_in_801 = {{6{1'b0}}, col_in_801};
assign u_ca_in_802 = {{6{1'b0}}, col_in_802};
assign u_ca_in_803 = {{6{1'b0}}, col_in_803};
assign u_ca_in_804 = {{6{1'b0}}, col_in_804};
assign u_ca_in_805 = {{6{1'b0}}, col_in_805};
assign u_ca_in_806 = {{6{1'b0}}, col_in_806};
assign u_ca_in_807 = {{6{1'b0}}, col_in_807};
assign u_ca_in_808 = {{6{1'b0}}, col_in_808};
assign u_ca_in_809 = {{6{1'b0}}, col_in_809};
assign u_ca_in_810 = {{6{1'b0}}, col_in_810};
assign u_ca_in_811 = {{6{1'b0}}, col_in_811};
assign u_ca_in_812 = {{6{1'b0}}, col_in_812};
assign u_ca_in_813 = {{6{1'b0}}, col_in_813};
assign u_ca_in_814 = {{6{1'b0}}, col_in_814};
assign u_ca_in_815 = {{6{1'b0}}, col_in_815};
assign u_ca_in_816 = {{6{1'b0}}, col_in_816};
assign u_ca_in_817 = {{6{1'b0}}, col_in_817};
assign u_ca_in_818 = {{6{1'b0}}, col_in_818};
assign u_ca_in_819 = {{6{1'b0}}, col_in_819};
assign u_ca_in_820 = {{6{1'b0}}, col_in_820};
assign u_ca_in_821 = {{6{1'b0}}, col_in_821};
assign u_ca_in_822 = {{6{1'b0}}, col_in_822};
assign u_ca_in_823 = {{6{1'b0}}, col_in_823};
assign u_ca_in_824 = {{6{1'b0}}, col_in_824};
assign u_ca_in_825 = {{6{1'b0}}, col_in_825};
assign u_ca_in_826 = {{6{1'b0}}, col_in_826};
assign u_ca_in_827 = {{6{1'b0}}, col_in_827};
assign u_ca_in_828 = {{6{1'b0}}, col_in_828};
assign u_ca_in_829 = {{6{1'b0}}, col_in_829};
assign u_ca_in_830 = {{6{1'b0}}, col_in_830};
assign u_ca_in_831 = {{6{1'b0}}, col_in_831};
assign u_ca_in_832 = {{6{1'b0}}, col_in_832};
assign u_ca_in_833 = {{6{1'b0}}, col_in_833};
assign u_ca_in_834 = {{6{1'b0}}, col_in_834};
assign u_ca_in_835 = {{6{1'b0}}, col_in_835};
assign u_ca_in_836 = {{6{1'b0}}, col_in_836};
assign u_ca_in_837 = {{6{1'b0}}, col_in_837};
assign u_ca_in_838 = {{6{1'b0}}, col_in_838};
assign u_ca_in_839 = {{6{1'b0}}, col_in_839};
assign u_ca_in_840 = {{6{1'b0}}, col_in_840};
assign u_ca_in_841 = {{6{1'b0}}, col_in_841};
assign u_ca_in_842 = {{6{1'b0}}, col_in_842};
assign u_ca_in_843 = {{6{1'b0}}, col_in_843};
assign u_ca_in_844 = {{6{1'b0}}, col_in_844};
assign u_ca_in_845 = {{6{1'b0}}, col_in_845};
assign u_ca_in_846 = {{6{1'b0}}, col_in_846};
assign u_ca_in_847 = {{6{1'b0}}, col_in_847};
assign u_ca_in_848 = {{6{1'b0}}, col_in_848};
assign u_ca_in_849 = {{6{1'b0}}, col_in_849};
assign u_ca_in_850 = {{6{1'b0}}, col_in_850};
assign u_ca_in_851 = {{6{1'b0}}, col_in_851};
assign u_ca_in_852 = {{6{1'b0}}, col_in_852};
assign u_ca_in_853 = {{6{1'b0}}, col_in_853};
assign u_ca_in_854 = {{6{1'b0}}, col_in_854};
assign u_ca_in_855 = {{6{1'b0}}, col_in_855};
assign u_ca_in_856 = {{6{1'b0}}, col_in_856};
assign u_ca_in_857 = {{6{1'b0}}, col_in_857};
assign u_ca_in_858 = {{6{1'b0}}, col_in_858};
assign u_ca_in_859 = {{6{1'b0}}, col_in_859};
assign u_ca_in_860 = {{6{1'b0}}, col_in_860};
assign u_ca_in_861 = {{6{1'b0}}, col_in_861};
assign u_ca_in_862 = {{6{1'b0}}, col_in_862};
assign u_ca_in_863 = {{6{1'b0}}, col_in_863};
assign u_ca_in_864 = {{6{1'b0}}, col_in_864};
assign u_ca_in_865 = {{6{1'b0}}, col_in_865};
assign u_ca_in_866 = {{6{1'b0}}, col_in_866};
assign u_ca_in_867 = {{6{1'b0}}, col_in_867};
assign u_ca_in_868 = {{6{1'b0}}, col_in_868};
assign u_ca_in_869 = {{6{1'b0}}, col_in_869};
assign u_ca_in_870 = {{6{1'b0}}, col_in_870};
assign u_ca_in_871 = {{6{1'b0}}, col_in_871};
assign u_ca_in_872 = {{6{1'b0}}, col_in_872};
assign u_ca_in_873 = {{6{1'b0}}, col_in_873};
assign u_ca_in_874 = {{6{1'b0}}, col_in_874};
assign u_ca_in_875 = {{6{1'b0}}, col_in_875};
assign u_ca_in_876 = {{6{1'b0}}, col_in_876};
assign u_ca_in_877 = {{6{1'b0}}, col_in_877};
assign u_ca_in_878 = {{6{1'b0}}, col_in_878};
assign u_ca_in_879 = {{6{1'b0}}, col_in_879};
assign u_ca_in_880 = {{6{1'b0}}, col_in_880};
assign u_ca_in_881 = {{6{1'b0}}, col_in_881};
assign u_ca_in_882 = {{6{1'b0}}, col_in_882};
assign u_ca_in_883 = {{6{1'b0}}, col_in_883};
assign u_ca_in_884 = {{6{1'b0}}, col_in_884};
assign u_ca_in_885 = {{6{1'b0}}, col_in_885};
assign u_ca_in_886 = {{6{1'b0}}, col_in_886};
assign u_ca_in_887 = {{6{1'b0}}, col_in_887};
assign u_ca_in_888 = {{6{1'b0}}, col_in_888};
assign u_ca_in_889 = {{6{1'b0}}, col_in_889};
assign u_ca_in_890 = {{6{1'b0}}, col_in_890};
assign u_ca_in_891 = {{6{1'b0}}, col_in_891};
assign u_ca_in_892 = {{6{1'b0}}, col_in_892};
assign u_ca_in_893 = {{6{1'b0}}, col_in_893};
assign u_ca_in_894 = {{6{1'b0}}, col_in_894};
assign u_ca_in_895 = {{6{1'b0}}, col_in_895};
assign u_ca_in_896 = {{6{1'b0}}, col_in_896};
assign u_ca_in_897 = {{6{1'b0}}, col_in_897};
assign u_ca_in_898 = {{6{1'b0}}, col_in_898};
assign u_ca_in_899 = {{6{1'b0}}, col_in_899};
assign u_ca_in_900 = {{6{1'b0}}, col_in_900};
assign u_ca_in_901 = {{6{1'b0}}, col_in_901};
assign u_ca_in_902 = {{6{1'b0}}, col_in_902};
assign u_ca_in_903 = {{6{1'b0}}, col_in_903};
assign u_ca_in_904 = {{6{1'b0}}, col_in_904};
assign u_ca_in_905 = {{6{1'b0}}, col_in_905};
assign u_ca_in_906 = {{6{1'b0}}, col_in_906};
assign u_ca_in_907 = {{6{1'b0}}, col_in_907};
assign u_ca_in_908 = {{6{1'b0}}, col_in_908};
assign u_ca_in_909 = {{6{1'b0}}, col_in_909};
assign u_ca_in_910 = {{6{1'b0}}, col_in_910};
assign u_ca_in_911 = {{6{1'b0}}, col_in_911};
assign u_ca_in_912 = {{6{1'b0}}, col_in_912};
assign u_ca_in_913 = {{6{1'b0}}, col_in_913};
assign u_ca_in_914 = {{6{1'b0}}, col_in_914};
assign u_ca_in_915 = {{6{1'b0}}, col_in_915};
assign u_ca_in_916 = {{6{1'b0}}, col_in_916};
assign u_ca_in_917 = {{6{1'b0}}, col_in_917};
assign u_ca_in_918 = {{6{1'b0}}, col_in_918};
assign u_ca_in_919 = {{6{1'b0}}, col_in_919};
assign u_ca_in_920 = {{6{1'b0}}, col_in_920};
assign u_ca_in_921 = {{6{1'b0}}, col_in_921};
assign u_ca_in_922 = {{6{1'b0}}, col_in_922};
assign u_ca_in_923 = {{6{1'b0}}, col_in_923};
assign u_ca_in_924 = {{6{1'b0}}, col_in_924};
assign u_ca_in_925 = {{6{1'b0}}, col_in_925};
assign u_ca_in_926 = {{6{1'b0}}, col_in_926};
assign u_ca_in_927 = {{6{1'b0}}, col_in_927};
assign u_ca_in_928 = {{6{1'b0}}, col_in_928};
assign u_ca_in_929 = {{6{1'b0}}, col_in_929};
assign u_ca_in_930 = {{6{1'b0}}, col_in_930};
assign u_ca_in_931 = {{6{1'b0}}, col_in_931};
assign u_ca_in_932 = {{6{1'b0}}, col_in_932};
assign u_ca_in_933 = {{6{1'b0}}, col_in_933};
assign u_ca_in_934 = {{6{1'b0}}, col_in_934};
assign u_ca_in_935 = {{6{1'b0}}, col_in_935};
assign u_ca_in_936 = {{6{1'b0}}, col_in_936};
assign u_ca_in_937 = {{6{1'b0}}, col_in_937};
assign u_ca_in_938 = {{6{1'b0}}, col_in_938};
assign u_ca_in_939 = {{6{1'b0}}, col_in_939};
assign u_ca_in_940 = {{6{1'b0}}, col_in_940};
assign u_ca_in_941 = {{6{1'b0}}, col_in_941};
assign u_ca_in_942 = {{6{1'b0}}, col_in_942};
assign u_ca_in_943 = {{6{1'b0}}, col_in_943};
assign u_ca_in_944 = {{6{1'b0}}, col_in_944};
assign u_ca_in_945 = {{6{1'b0}}, col_in_945};
assign u_ca_in_946 = {{6{1'b0}}, col_in_946};
assign u_ca_in_947 = {{6{1'b0}}, col_in_947};
assign u_ca_in_948 = {{6{1'b0}}, col_in_948};
assign u_ca_in_949 = {{6{1'b0}}, col_in_949};
assign u_ca_in_950 = {{6{1'b0}}, col_in_950};
assign u_ca_in_951 = {{6{1'b0}}, col_in_951};
assign u_ca_in_952 = {{6{1'b0}}, col_in_952};
assign u_ca_in_953 = {{6{1'b0}}, col_in_953};
assign u_ca_in_954 = {{6{1'b0}}, col_in_954};
assign u_ca_in_955 = {{6{1'b0}}, col_in_955};
assign u_ca_in_956 = {{6{1'b0}}, col_in_956};
assign u_ca_in_957 = {{6{1'b0}}, col_in_957};
assign u_ca_in_958 = {{6{1'b0}}, col_in_958};
assign u_ca_in_959 = {{6{1'b0}}, col_in_959};
assign u_ca_in_960 = {{6{1'b0}}, col_in_960};
assign u_ca_in_961 = {{6{1'b0}}, col_in_961};
assign u_ca_in_962 = {{6{1'b0}}, col_in_962};
assign u_ca_in_963 = {{6{1'b0}}, col_in_963};
assign u_ca_in_964 = {{6{1'b0}}, col_in_964};
assign u_ca_in_965 = {{6{1'b0}}, col_in_965};
assign u_ca_in_966 = {{6{1'b0}}, col_in_966};
assign u_ca_in_967 = {{6{1'b0}}, col_in_967};
assign u_ca_in_968 = {{6{1'b0}}, col_in_968};
assign u_ca_in_969 = {{6{1'b0}}, col_in_969};
assign u_ca_in_970 = {{6{1'b0}}, col_in_970};
assign u_ca_in_971 = {{6{1'b0}}, col_in_971};
assign u_ca_in_972 = {{6{1'b0}}, col_in_972};
assign u_ca_in_973 = {{6{1'b0}}, col_in_973};
assign u_ca_in_974 = {{6{1'b0}}, col_in_974};
assign u_ca_in_975 = {{6{1'b0}}, col_in_975};
assign u_ca_in_976 = {{6{1'b0}}, col_in_976};
assign u_ca_in_977 = {{6{1'b0}}, col_in_977};
assign u_ca_in_978 = {{6{1'b0}}, col_in_978};
assign u_ca_in_979 = {{6{1'b0}}, col_in_979};
assign u_ca_in_980 = {{6{1'b0}}, col_in_980};
assign u_ca_in_981 = {{6{1'b0}}, col_in_981};
assign u_ca_in_982 = {{6{1'b0}}, col_in_982};
assign u_ca_in_983 = {{6{1'b0}}, col_in_983};
assign u_ca_in_984 = {{6{1'b0}}, col_in_984};
assign u_ca_in_985 = {{6{1'b0}}, col_in_985};
assign u_ca_in_986 = {{6{1'b0}}, col_in_986};
assign u_ca_in_987 = {{6{1'b0}}, col_in_987};
assign u_ca_in_988 = {{6{1'b0}}, col_in_988};
assign u_ca_in_989 = {{6{1'b0}}, col_in_989};
assign u_ca_in_990 = {{6{1'b0}}, col_in_990};
assign u_ca_in_991 = {{6{1'b0}}, col_in_991};
assign u_ca_in_992 = {{6{1'b0}}, col_in_992};
assign u_ca_in_993 = {{6{1'b0}}, col_in_993};
assign u_ca_in_994 = {{6{1'b0}}, col_in_994};
assign u_ca_in_995 = {{6{1'b0}}, col_in_995};
assign u_ca_in_996 = {{6{1'b0}}, col_in_996};
assign u_ca_in_997 = {{6{1'b0}}, col_in_997};
assign u_ca_in_998 = {{6{1'b0}}, col_in_998};
assign u_ca_in_999 = {{6{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{6{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{6{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{6{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{6{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{6{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{6{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{6{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{6{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{6{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{6{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{6{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{6{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{6{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{6{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{6{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{6{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{6{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{6{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{6{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{6{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{6{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{6{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{6{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{6{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{6{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{6{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{6{1'b0}}, col_in_1026};
assign u_ca_in_1027 = {{6{1'b0}}, col_in_1027};
assign u_ca_in_1028 = {{6{1'b0}}, col_in_1028};
assign u_ca_in_1029 = {{6{1'b0}}, col_in_1029};

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_54_16 u_ca_54_16_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_54_16 u_ca_54_16_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_54_16 u_ca_54_16_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_54_16 u_ca_54_16_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_54_16 u_ca_54_16_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_54_16 u_ca_54_16_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_54_16 u_ca_54_16_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_54_16 u_ca_54_16_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_54_16 u_ca_54_16_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_54_16 u_ca_54_16_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_54_16 u_ca_54_16_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_54_16 u_ca_54_16_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_54_16 u_ca_54_16_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_54_16 u_ca_54_16_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_54_16 u_ca_54_16_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_54_16 u_ca_54_16_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_54_16 u_ca_54_16_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_54_16 u_ca_54_16_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_54_16 u_ca_54_16_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_54_16 u_ca_54_16_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_54_16 u_ca_54_16_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_54_16 u_ca_54_16_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_54_16 u_ca_54_16_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_54_16 u_ca_54_16_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_54_16 u_ca_54_16_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_54_16 u_ca_54_16_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_54_16 u_ca_54_16_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_54_16 u_ca_54_16_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_54_16 u_ca_54_16_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_54_16 u_ca_54_16_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_54_16 u_ca_54_16_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_54_16 u_ca_54_16_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_54_16 u_ca_54_16_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_54_16 u_ca_54_16_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_54_16 u_ca_54_16_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_54_16 u_ca_54_16_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_54_16 u_ca_54_16_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_54_16 u_ca_54_16_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_54_16 u_ca_54_16_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_54_16 u_ca_54_16_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_54_16 u_ca_54_16_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_54_16 u_ca_54_16_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_54_16 u_ca_54_16_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_54_16 u_ca_54_16_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_54_16 u_ca_54_16_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_54_16 u_ca_54_16_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_54_16 u_ca_54_16_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_54_16 u_ca_54_16_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_54_16 u_ca_54_16_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_54_16 u_ca_54_16_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_54_16 u_ca_54_16_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_54_16 u_ca_54_16_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_54_16 u_ca_54_16_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_54_16 u_ca_54_16_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_54_16 u_ca_54_16_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_54_16 u_ca_54_16_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_54_16 u_ca_54_16_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_54_16 u_ca_54_16_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_54_16 u_ca_54_16_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_54_16 u_ca_54_16_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_54_16 u_ca_54_16_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_54_16 u_ca_54_16_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_54_16 u_ca_54_16_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_54_16 u_ca_54_16_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_54_16 u_ca_54_16_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_54_16 u_ca_54_16_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_54_16 u_ca_54_16_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_54_16 u_ca_54_16_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_54_16 u_ca_54_16_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_54_16 u_ca_54_16_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_54_16 u_ca_54_16_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_54_16 u_ca_54_16_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_54_16 u_ca_54_16_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_54_16 u_ca_54_16_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_54_16 u_ca_54_16_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_54_16 u_ca_54_16_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_54_16 u_ca_54_16_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_54_16 u_ca_54_16_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_54_16 u_ca_54_16_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_54_16 u_ca_54_16_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_54_16 u_ca_54_16_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_54_16 u_ca_54_16_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_54_16 u_ca_54_16_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_54_16 u_ca_54_16_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_54_16 u_ca_54_16_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_54_16 u_ca_54_16_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_54_16 u_ca_54_16_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_54_16 u_ca_54_16_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_54_16 u_ca_54_16_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_54_16 u_ca_54_16_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_54_16 u_ca_54_16_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_54_16 u_ca_54_16_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_54_16 u_ca_54_16_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_54_16 u_ca_54_16_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_54_16 u_ca_54_16_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_54_16 u_ca_54_16_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_54_16 u_ca_54_16_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_54_16 u_ca_54_16_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_54_16 u_ca_54_16_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_54_16 u_ca_54_16_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_54_16 u_ca_54_16_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_54_16 u_ca_54_16_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_54_16 u_ca_54_16_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_54_16 u_ca_54_16_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_54_16 u_ca_54_16_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_54_16 u_ca_54_16_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_54_16 u_ca_54_16_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_54_16 u_ca_54_16_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_54_16 u_ca_54_16_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_54_16 u_ca_54_16_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_54_16 u_ca_54_16_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_54_16 u_ca_54_16_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_54_16 u_ca_54_16_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_54_16 u_ca_54_16_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_54_16 u_ca_54_16_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_54_16 u_ca_54_16_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_54_16 u_ca_54_16_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_54_16 u_ca_54_16_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_54_16 u_ca_54_16_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_54_16 u_ca_54_16_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_54_16 u_ca_54_16_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_54_16 u_ca_54_16_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_54_16 u_ca_54_16_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_54_16 u_ca_54_16_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_54_16 u_ca_54_16_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_54_16 u_ca_54_16_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_54_16 u_ca_54_16_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_54_16 u_ca_54_16_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_54_16 u_ca_54_16_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_54_16 u_ca_54_16_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_54_16 u_ca_54_16_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_54_16 u_ca_54_16_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_54_16 u_ca_54_16_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_54_16 u_ca_54_16_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_54_16 u_ca_54_16_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_54_16 u_ca_54_16_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_54_16 u_ca_54_16_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_54_16 u_ca_54_16_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_54_16 u_ca_54_16_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_54_16 u_ca_54_16_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_54_16 u_ca_54_16_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_54_16 u_ca_54_16_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_54_16 u_ca_54_16_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_54_16 u_ca_54_16_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_54_16 u_ca_54_16_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_54_16 u_ca_54_16_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_54_16 u_ca_54_16_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_54_16 u_ca_54_16_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_54_16 u_ca_54_16_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_54_16 u_ca_54_16_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_54_16 u_ca_54_16_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_54_16 u_ca_54_16_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_54_16 u_ca_54_16_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_54_16 u_ca_54_16_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_54_16 u_ca_54_16_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_54_16 u_ca_54_16_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_54_16 u_ca_54_16_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_54_16 u_ca_54_16_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_54_16 u_ca_54_16_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_54_16 u_ca_54_16_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_54_16 u_ca_54_16_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_54_16 u_ca_54_16_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_54_16 u_ca_54_16_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_54_16 u_ca_54_16_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_54_16 u_ca_54_16_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_54_16 u_ca_54_16_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_54_16 u_ca_54_16_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_54_16 u_ca_54_16_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_54_16 u_ca_54_16_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_54_16 u_ca_54_16_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_54_16 u_ca_54_16_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_54_16 u_ca_54_16_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_54_16 u_ca_54_16_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_54_16 u_ca_54_16_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_54_16 u_ca_54_16_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_54_16 u_ca_54_16_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_54_16 u_ca_54_16_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_54_16 u_ca_54_16_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_54_16 u_ca_54_16_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_54_16 u_ca_54_16_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_54_16 u_ca_54_16_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_54_16 u_ca_54_16_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_54_16 u_ca_54_16_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_54_16 u_ca_54_16_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_54_16 u_ca_54_16_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_54_16 u_ca_54_16_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_54_16 u_ca_54_16_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_54_16 u_ca_54_16_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_54_16 u_ca_54_16_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_54_16 u_ca_54_16_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_54_16 u_ca_54_16_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_54_16 u_ca_54_16_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_54_16 u_ca_54_16_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_54_16 u_ca_54_16_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_54_16 u_ca_54_16_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_54_16 u_ca_54_16_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_54_16 u_ca_54_16_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_54_16 u_ca_54_16_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_54_16 u_ca_54_16_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_54_16 u_ca_54_16_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_54_16 u_ca_54_16_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_54_16 u_ca_54_16_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_54_16 u_ca_54_16_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_54_16 u_ca_54_16_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_54_16 u_ca_54_16_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_54_16 u_ca_54_16_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_54_16 u_ca_54_16_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_54_16 u_ca_54_16_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_54_16 u_ca_54_16_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_54_16 u_ca_54_16_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_54_16 u_ca_54_16_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_54_16 u_ca_54_16_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_54_16 u_ca_54_16_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_54_16 u_ca_54_16_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_54_16 u_ca_54_16_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_54_16 u_ca_54_16_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_54_16 u_ca_54_16_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_54_16 u_ca_54_16_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_54_16 u_ca_54_16_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_54_16 u_ca_54_16_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_54_16 u_ca_54_16_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_54_16 u_ca_54_16_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_54_16 u_ca_54_16_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_54_16 u_ca_54_16_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_54_16 u_ca_54_16_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_54_16 u_ca_54_16_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_54_16 u_ca_54_16_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_54_16 u_ca_54_16_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_54_16 u_ca_54_16_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_54_16 u_ca_54_16_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_54_16 u_ca_54_16_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_54_16 u_ca_54_16_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_54_16 u_ca_54_16_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_54_16 u_ca_54_16_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_54_16 u_ca_54_16_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_54_16 u_ca_54_16_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_54_16 u_ca_54_16_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_54_16 u_ca_54_16_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_54_16 u_ca_54_16_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_54_16 u_ca_54_16_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_54_16 u_ca_54_16_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_54_16 u_ca_54_16_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_54_16 u_ca_54_16_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_54_16 u_ca_54_16_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_54_16 u_ca_54_16_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_54_16 u_ca_54_16_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_54_16 u_ca_54_16_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_54_16 u_ca_54_16_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_54_16 u_ca_54_16_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_54_16 u_ca_54_16_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_54_16 u_ca_54_16_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_54_16 u_ca_54_16_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_54_16 u_ca_54_16_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_54_16 u_ca_54_16_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_54_16 u_ca_54_16_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_54_16 u_ca_54_16_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_54_16 u_ca_54_16_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_54_16 u_ca_54_16_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_54_16 u_ca_54_16_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_54_16 u_ca_54_16_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_54_16 u_ca_54_16_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_54_16 u_ca_54_16_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_54_16 u_ca_54_16_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_54_16 u_ca_54_16_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_54_16 u_ca_54_16_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_54_16 u_ca_54_16_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_54_16 u_ca_54_16_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_54_16 u_ca_54_16_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_54_16 u_ca_54_16_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_54_16 u_ca_54_16_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_54_16 u_ca_54_16_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_54_16 u_ca_54_16_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_54_16 u_ca_54_16_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_54_16 u_ca_54_16_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_54_16 u_ca_54_16_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_54_16 u_ca_54_16_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_54_16 u_ca_54_16_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_54_16 u_ca_54_16_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_54_16 u_ca_54_16_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_54_16 u_ca_54_16_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_54_16 u_ca_54_16_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_54_16 u_ca_54_16_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_54_16 u_ca_54_16_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_54_16 u_ca_54_16_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_54_16 u_ca_54_16_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_54_16 u_ca_54_16_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_54_16 u_ca_54_16_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_54_16 u_ca_54_16_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_54_16 u_ca_54_16_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_54_16 u_ca_54_16_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_54_16 u_ca_54_16_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_54_16 u_ca_54_16_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_54_16 u_ca_54_16_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_54_16 u_ca_54_16_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_54_16 u_ca_54_16_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_54_16 u_ca_54_16_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_54_16 u_ca_54_16_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_54_16 u_ca_54_16_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_54_16 u_ca_54_16_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_54_16 u_ca_54_16_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_54_16 u_ca_54_16_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_54_16 u_ca_54_16_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_54_16 u_ca_54_16_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_54_16 u_ca_54_16_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_54_16 u_ca_54_16_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_54_16 u_ca_54_16_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_54_16 u_ca_54_16_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_54_16 u_ca_54_16_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_54_16 u_ca_54_16_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_54_16 u_ca_54_16_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_54_16 u_ca_54_16_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_54_16 u_ca_54_16_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_54_16 u_ca_54_16_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_54_16 u_ca_54_16_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_54_16 u_ca_54_16_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_54_16 u_ca_54_16_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_54_16 u_ca_54_16_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_54_16 u_ca_54_16_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_54_16 u_ca_54_16_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_54_16 u_ca_54_16_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_54_16 u_ca_54_16_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_54_16 u_ca_54_16_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_54_16 u_ca_54_16_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_54_16 u_ca_54_16_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_54_16 u_ca_54_16_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_54_16 u_ca_54_16_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_54_16 u_ca_54_16_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_54_16 u_ca_54_16_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_54_16 u_ca_54_16_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_54_16 u_ca_54_16_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_54_16 u_ca_54_16_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_54_16 u_ca_54_16_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_54_16 u_ca_54_16_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_54_16 u_ca_54_16_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_54_16 u_ca_54_16_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_54_16 u_ca_54_16_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_54_16 u_ca_54_16_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_54_16 u_ca_54_16_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_54_16 u_ca_54_16_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_54_16 u_ca_54_16_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_54_16 u_ca_54_16_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_54_16 u_ca_54_16_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_54_16 u_ca_54_16_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_54_16 u_ca_54_16_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_54_16 u_ca_54_16_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_54_16 u_ca_54_16_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_54_16 u_ca_54_16_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_54_16 u_ca_54_16_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_54_16 u_ca_54_16_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_54_16 u_ca_54_16_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_54_16 u_ca_54_16_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_54_16 u_ca_54_16_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_54_16 u_ca_54_16_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_54_16 u_ca_54_16_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_54_16 u_ca_54_16_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_54_16 u_ca_54_16_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_54_16 u_ca_54_16_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_54_16 u_ca_54_16_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_54_16 u_ca_54_16_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_54_16 u_ca_54_16_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_54_16 u_ca_54_16_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_54_16 u_ca_54_16_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_54_16 u_ca_54_16_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_54_16 u_ca_54_16_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_54_16 u_ca_54_16_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_54_16 u_ca_54_16_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_54_16 u_ca_54_16_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_54_16 u_ca_54_16_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_54_16 u_ca_54_16_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_54_16 u_ca_54_16_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_54_16 u_ca_54_16_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_54_16 u_ca_54_16_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_54_16 u_ca_54_16_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_54_16 u_ca_54_16_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_54_16 u_ca_54_16_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_54_16 u_ca_54_16_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_54_16 u_ca_54_16_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_54_16 u_ca_54_16_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_54_16 u_ca_54_16_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_54_16 u_ca_54_16_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_54_16 u_ca_54_16_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_54_16 u_ca_54_16_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_54_16 u_ca_54_16_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_54_16 u_ca_54_16_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_54_16 u_ca_54_16_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_54_16 u_ca_54_16_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_54_16 u_ca_54_16_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_54_16 u_ca_54_16_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_54_16 u_ca_54_16_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_54_16 u_ca_54_16_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_54_16 u_ca_54_16_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_54_16 u_ca_54_16_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_54_16 u_ca_54_16_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_54_16 u_ca_54_16_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_54_16 u_ca_54_16_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_54_16 u_ca_54_16_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_54_16 u_ca_54_16_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_54_16 u_ca_54_16_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_54_16 u_ca_54_16_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_54_16 u_ca_54_16_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_54_16 u_ca_54_16_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_54_16 u_ca_54_16_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_54_16 u_ca_54_16_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_54_16 u_ca_54_16_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_54_16 u_ca_54_16_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_54_16 u_ca_54_16_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_54_16 u_ca_54_16_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_54_16 u_ca_54_16_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_54_16 u_ca_54_16_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_54_16 u_ca_54_16_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_54_16 u_ca_54_16_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_54_16 u_ca_54_16_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_54_16 u_ca_54_16_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_54_16 u_ca_54_16_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_54_16 u_ca_54_16_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_54_16 u_ca_54_16_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_54_16 u_ca_54_16_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_54_16 u_ca_54_16_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_54_16 u_ca_54_16_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_54_16 u_ca_54_16_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_54_16 u_ca_54_16_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_54_16 u_ca_54_16_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_54_16 u_ca_54_16_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_54_16 u_ca_54_16_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_54_16 u_ca_54_16_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_54_16 u_ca_54_16_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_54_16 u_ca_54_16_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_54_16 u_ca_54_16_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_54_16 u_ca_54_16_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_54_16 u_ca_54_16_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_54_16 u_ca_54_16_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_54_16 u_ca_54_16_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_54_16 u_ca_54_16_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_54_16 u_ca_54_16_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_54_16 u_ca_54_16_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_54_16 u_ca_54_16_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_54_16 u_ca_54_16_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_54_16 u_ca_54_16_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_54_16 u_ca_54_16_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_54_16 u_ca_54_16_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_54_16 u_ca_54_16_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_54_16 u_ca_54_16_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_54_16 u_ca_54_16_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_54_16 u_ca_54_16_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_54_16 u_ca_54_16_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_54_16 u_ca_54_16_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_54_16 u_ca_54_16_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_54_16 u_ca_54_16_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_54_16 u_ca_54_16_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_54_16 u_ca_54_16_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_54_16 u_ca_54_16_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_54_16 u_ca_54_16_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_54_16 u_ca_54_16_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_54_16 u_ca_54_16_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_54_16 u_ca_54_16_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_54_16 u_ca_54_16_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_54_16 u_ca_54_16_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_54_16 u_ca_54_16_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_54_16 u_ca_54_16_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_54_16 u_ca_54_16_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_54_16 u_ca_54_16_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_54_16 u_ca_54_16_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_54_16 u_ca_54_16_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_54_16 u_ca_54_16_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_54_16 u_ca_54_16_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_54_16 u_ca_54_16_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_54_16 u_ca_54_16_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_54_16 u_ca_54_16_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_54_16 u_ca_54_16_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_54_16 u_ca_54_16_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_54_16 u_ca_54_16_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_54_16 u_ca_54_16_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_54_16 u_ca_54_16_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_54_16 u_ca_54_16_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_54_16 u_ca_54_16_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_54_16 u_ca_54_16_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_54_16 u_ca_54_16_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_54_16 u_ca_54_16_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_54_16 u_ca_54_16_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_54_16 u_ca_54_16_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_54_16 u_ca_54_16_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_54_16 u_ca_54_16_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_54_16 u_ca_54_16_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_54_16 u_ca_54_16_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_54_16 u_ca_54_16_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_54_16 u_ca_54_16_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_54_16 u_ca_54_16_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_54_16 u_ca_54_16_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_54_16 u_ca_54_16_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_54_16 u_ca_54_16_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_54_16 u_ca_54_16_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_54_16 u_ca_54_16_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_54_16 u_ca_54_16_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_54_16 u_ca_54_16_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_54_16 u_ca_54_16_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_54_16 u_ca_54_16_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_54_16 u_ca_54_16_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_54_16 u_ca_54_16_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_54_16 u_ca_54_16_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_54_16 u_ca_54_16_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_54_16 u_ca_54_16_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_54_16 u_ca_54_16_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_54_16 u_ca_54_16_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_54_16 u_ca_54_16_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_54_16 u_ca_54_16_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_54_16 u_ca_54_16_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_54_16 u_ca_54_16_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_54_16 u_ca_54_16_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_54_16 u_ca_54_16_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_54_16 u_ca_54_16_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_54_16 u_ca_54_16_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_54_16 u_ca_54_16_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_54_16 u_ca_54_16_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_54_16 u_ca_54_16_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_54_16 u_ca_54_16_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_54_16 u_ca_54_16_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_54_16 u_ca_54_16_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_54_16 u_ca_54_16_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_54_16 u_ca_54_16_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_54_16 u_ca_54_16_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_54_16 u_ca_54_16_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_54_16 u_ca_54_16_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_54_16 u_ca_54_16_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_54_16 u_ca_54_16_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_54_16 u_ca_54_16_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_54_16 u_ca_54_16_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_54_16 u_ca_54_16_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_54_16 u_ca_54_16_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_54_16 u_ca_54_16_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_54_16 u_ca_54_16_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_54_16 u_ca_54_16_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_54_16 u_ca_54_16_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_54_16 u_ca_54_16_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_54_16 u_ca_54_16_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_54_16 u_ca_54_16_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_54_16 u_ca_54_16_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_54_16 u_ca_54_16_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_54_16 u_ca_54_16_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_54_16 u_ca_54_16_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_54_16 u_ca_54_16_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_54_16 u_ca_54_16_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_54_16 u_ca_54_16_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_54_16 u_ca_54_16_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_54_16 u_ca_54_16_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_54_16 u_ca_54_16_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_54_16 u_ca_54_16_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_54_16 u_ca_54_16_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_54_16 u_ca_54_16_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_54_16 u_ca_54_16_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_54_16 u_ca_54_16_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_54_16 u_ca_54_16_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_54_16 u_ca_54_16_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_54_16 u_ca_54_16_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_54_16 u_ca_54_16_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_54_16 u_ca_54_16_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_54_16 u_ca_54_16_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_54_16 u_ca_54_16_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_54_16 u_ca_54_16_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_54_16 u_ca_54_16_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_54_16 u_ca_54_16_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_54_16 u_ca_54_16_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_54_16 u_ca_54_16_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_54_16 u_ca_54_16_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_54_16 u_ca_54_16_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_54_16 u_ca_54_16_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_54_16 u_ca_54_16_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_54_16 u_ca_54_16_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_54_16 u_ca_54_16_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_54_16 u_ca_54_16_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_54_16 u_ca_54_16_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_54_16 u_ca_54_16_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_54_16 u_ca_54_16_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_54_16 u_ca_54_16_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_54_16 u_ca_54_16_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_54_16 u_ca_54_16_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_54_16 u_ca_54_16_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_54_16 u_ca_54_16_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_54_16 u_ca_54_16_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_54_16 u_ca_54_16_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_54_16 u_ca_54_16_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_54_16 u_ca_54_16_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_54_16 u_ca_54_16_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_54_16 u_ca_54_16_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_54_16 u_ca_54_16_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_54_16 u_ca_54_16_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_54_16 u_ca_54_16_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_54_16 u_ca_54_16_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_54_16 u_ca_54_16_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_54_16 u_ca_54_16_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_54_16 u_ca_54_16_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_54_16 u_ca_54_16_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_54_16 u_ca_54_16_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_54_16 u_ca_54_16_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_54_16 u_ca_54_16_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_54_16 u_ca_54_16_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_54_16 u_ca_54_16_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_54_16 u_ca_54_16_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_54_16 u_ca_54_16_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_54_16 u_ca_54_16_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_54_16 u_ca_54_16_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_54_16 u_ca_54_16_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_54_16 u_ca_54_16_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_54_16 u_ca_54_16_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_54_16 u_ca_54_16_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_54_16 u_ca_54_16_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_54_16 u_ca_54_16_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_54_16 u_ca_54_16_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_54_16 u_ca_54_16_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_54_16 u_ca_54_16_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_54_16 u_ca_54_16_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_54_16 u_ca_54_16_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_54_16 u_ca_54_16_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_54_16 u_ca_54_16_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_54_16 u_ca_54_16_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_54_16 u_ca_54_16_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_54_16 u_ca_54_16_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_54_16 u_ca_54_16_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_54_16 u_ca_54_16_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_54_16 u_ca_54_16_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_54_16 u_ca_54_16_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_54_16 u_ca_54_16_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_54_16 u_ca_54_16_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_54_16 u_ca_54_16_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_54_16 u_ca_54_16_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_54_16 u_ca_54_16_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_54_16 u_ca_54_16_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_54_16 u_ca_54_16_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_54_16 u_ca_54_16_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_54_16 u_ca_54_16_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_54_16 u_ca_54_16_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_54_16 u_ca_54_16_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_54_16 u_ca_54_16_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_54_16 u_ca_54_16_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_54_16 u_ca_54_16_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_54_16 u_ca_54_16_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_54_16 u_ca_54_16_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_54_16 u_ca_54_16_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_54_16 u_ca_54_16_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_54_16 u_ca_54_16_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_54_16 u_ca_54_16_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_54_16 u_ca_54_16_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_54_16 u_ca_54_16_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_54_16 u_ca_54_16_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_54_16 u_ca_54_16_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_54_16 u_ca_54_16_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_54_16 u_ca_54_16_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_54_16 u_ca_54_16_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_54_16 u_ca_54_16_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_54_16 u_ca_54_16_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_54_16 u_ca_54_16_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_54_16 u_ca_54_16_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_54_16 u_ca_54_16_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_54_16 u_ca_54_16_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_54_16 u_ca_54_16_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_54_16 u_ca_54_16_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_54_16 u_ca_54_16_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_54_16 u_ca_54_16_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_54_16 u_ca_54_16_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_54_16 u_ca_54_16_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_54_16 u_ca_54_16_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_54_16 u_ca_54_16_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_54_16 u_ca_54_16_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_54_16 u_ca_54_16_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_54_16 u_ca_54_16_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_54_16 u_ca_54_16_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_54_16 u_ca_54_16_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_54_16 u_ca_54_16_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_54_16 u_ca_54_16_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_54_16 u_ca_54_16_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_54_16 u_ca_54_16_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_54_16 u_ca_54_16_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_54_16 u_ca_54_16_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_54_16 u_ca_54_16_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_54_16 u_ca_54_16_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_54_16 u_ca_54_16_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_54_16 u_ca_54_16_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_54_16 u_ca_54_16_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_54_16 u_ca_54_16_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_54_16 u_ca_54_16_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_54_16 u_ca_54_16_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_54_16 u_ca_54_16_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_54_16 u_ca_54_16_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_54_16 u_ca_54_16_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_54_16 u_ca_54_16_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_54_16 u_ca_54_16_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_54_16 u_ca_54_16_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_54_16 u_ca_54_16_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_54_16 u_ca_54_16_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_54_16 u_ca_54_16_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_54_16 u_ca_54_16_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_54_16 u_ca_54_16_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_54_16 u_ca_54_16_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_54_16 u_ca_54_16_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_54_16 u_ca_54_16_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_54_16 u_ca_54_16_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_54_16 u_ca_54_16_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_54_16 u_ca_54_16_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_54_16 u_ca_54_16_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_54_16 u_ca_54_16_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_54_16 u_ca_54_16_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_54_16 u_ca_54_16_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_54_16 u_ca_54_16_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_54_16 u_ca_54_16_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_54_16 u_ca_54_16_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_54_16 u_ca_54_16_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_54_16 u_ca_54_16_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_54_16 u_ca_54_16_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_54_16 u_ca_54_16_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_54_16 u_ca_54_16_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_54_16 u_ca_54_16_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_54_16 u_ca_54_16_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_54_16 u_ca_54_16_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_54_16 u_ca_54_16_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_54_16 u_ca_54_16_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_54_16 u_ca_54_16_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_54_16 u_ca_54_16_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_54_16 u_ca_54_16_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_54_16 u_ca_54_16_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_54_16 u_ca_54_16_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_54_16 u_ca_54_16_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_54_16 u_ca_54_16_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_54_16 u_ca_54_16_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_54_16 u_ca_54_16_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_54_16 u_ca_54_16_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_54_16 u_ca_54_16_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_54_16 u_ca_54_16_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_54_16 u_ca_54_16_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_54_16 u_ca_54_16_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_54_16 u_ca_54_16_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_54_16 u_ca_54_16_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_54_16 u_ca_54_16_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_54_16 u_ca_54_16_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_54_16 u_ca_54_16_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_54_16 u_ca_54_16_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_54_16 u_ca_54_16_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_54_16 u_ca_54_16_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_54_16 u_ca_54_16_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_54_16 u_ca_54_16_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_54_16 u_ca_54_16_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_54_16 u_ca_54_16_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_54_16 u_ca_54_16_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_54_16 u_ca_54_16_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_54_16 u_ca_54_16_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_54_16 u_ca_54_16_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_54_16 u_ca_54_16_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_54_16 u_ca_54_16_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_54_16 u_ca_54_16_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_54_16 u_ca_54_16_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_54_16 u_ca_54_16_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_54_16 u_ca_54_16_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_54_16 u_ca_54_16_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_54_16 u_ca_54_16_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_54_16 u_ca_54_16_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_54_16 u_ca_54_16_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_54_16 u_ca_54_16_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_54_16 u_ca_54_16_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_54_16 u_ca_54_16_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_54_16 u_ca_54_16_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_54_16 u_ca_54_16_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_54_16 u_ca_54_16_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_54_16 u_ca_54_16_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_54_16 u_ca_54_16_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_54_16 u_ca_54_16_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_54_16 u_ca_54_16_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_54_16 u_ca_54_16_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_54_16 u_ca_54_16_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_54_16 u_ca_54_16_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_54_16 u_ca_54_16_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_54_16 u_ca_54_16_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_54_16 u_ca_54_16_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_54_16 u_ca_54_16_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_54_16 u_ca_54_16_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_54_16 u_ca_54_16_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_54_16 u_ca_54_16_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_54_16 u_ca_54_16_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_54_16 u_ca_54_16_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_54_16 u_ca_54_16_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_54_16 u_ca_54_16_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_54_16 u_ca_54_16_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_54_16 u_ca_54_16_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_54_16 u_ca_54_16_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_54_16 u_ca_54_16_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_54_16 u_ca_54_16_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_54_16 u_ca_54_16_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_54_16 u_ca_54_16_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_54_16 u_ca_54_16_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_54_16 u_ca_54_16_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_54_16 u_ca_54_16_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_54_16 u_ca_54_16_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_54_16 u_ca_54_16_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_54_16 u_ca_54_16_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_54_16 u_ca_54_16_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_54_16 u_ca_54_16_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_54_16 u_ca_54_16_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_54_16 u_ca_54_16_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_54_16 u_ca_54_16_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_54_16 u_ca_54_16_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_54_16 u_ca_54_16_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_54_16 u_ca_54_16_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_54_16 u_ca_54_16_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_54_16 u_ca_54_16_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_54_16 u_ca_54_16_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_54_16 u_ca_54_16_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_54_16 u_ca_54_16_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_54_16 u_ca_54_16_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_54_16 u_ca_54_16_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_54_16 u_ca_54_16_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_54_16 u_ca_54_16_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_54_16 u_ca_54_16_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_54_16 u_ca_54_16_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_54_16 u_ca_54_16_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_54_16 u_ca_54_16_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_54_16 u_ca_54_16_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_54_16 u_ca_54_16_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_54_16 u_ca_54_16_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_54_16 u_ca_54_16_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_54_16 u_ca_54_16_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_54_16 u_ca_54_16_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_54_16 u_ca_54_16_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_54_16 u_ca_54_16_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_54_16 u_ca_54_16_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_54_16 u_ca_54_16_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_54_16 u_ca_54_16_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_54_16 u_ca_54_16_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_54_16 u_ca_54_16_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_54_16 u_ca_54_16_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_54_16 u_ca_54_16_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_54_16 u_ca_54_16_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_54_16 u_ca_54_16_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_54_16 u_ca_54_16_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_54_16 u_ca_54_16_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_54_16 u_ca_54_16_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_54_16 u_ca_54_16_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_54_16 u_ca_54_16_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_54_16 u_ca_54_16_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_54_16 u_ca_54_16_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_54_16 u_ca_54_16_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_54_16 u_ca_54_16_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_54_16 u_ca_54_16_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_54_16 u_ca_54_16_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_54_16 u_ca_54_16_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_54_16 u_ca_54_16_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_54_16 u_ca_54_16_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_54_16 u_ca_54_16_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_54_16 u_ca_54_16_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_54_16 u_ca_54_16_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_54_16 u_ca_54_16_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_54_16 u_ca_54_16_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_54_16 u_ca_54_16_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_54_16 u_ca_54_16_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_54_16 u_ca_54_16_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_54_16 u_ca_54_16_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_54_16 u_ca_54_16_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_54_16 u_ca_54_16_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_54_16 u_ca_54_16_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_54_16 u_ca_54_16_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_54_16 u_ca_54_16_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_54_16 u_ca_54_16_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_54_16 u_ca_54_16_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_54_16 u_ca_54_16_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_54_16 u_ca_54_16_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_54_16 u_ca_54_16_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_54_16 u_ca_54_16_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_54_16 u_ca_54_16_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_54_16 u_ca_54_16_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_54_16 u_ca_54_16_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_54_16 u_ca_54_16_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_54_16 u_ca_54_16_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_54_16 u_ca_54_16_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_54_16 u_ca_54_16_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_54_16 u_ca_54_16_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_54_16 u_ca_54_16_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_54_16 u_ca_54_16_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_54_16 u_ca_54_16_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_54_16 u_ca_54_16_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_54_16 u_ca_54_16_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_54_16 u_ca_54_16_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_54_16 u_ca_54_16_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_54_16 u_ca_54_16_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_54_16 u_ca_54_16_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_54_16 u_ca_54_16_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_54_16 u_ca_54_16_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_54_16 u_ca_54_16_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_54_16 u_ca_54_16_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_54_16 u_ca_54_16_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_54_16 u_ca_54_16_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_54_16 u_ca_54_16_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_54_16 u_ca_54_16_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_54_16 u_ca_54_16_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_54_16 u_ca_54_16_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_54_16 u_ca_54_16_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_54_16 u_ca_54_16_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_54_16 u_ca_54_16_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_54_16 u_ca_54_16_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_54_16 u_ca_54_16_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_54_16 u_ca_54_16_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_54_16 u_ca_54_16_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_54_16 u_ca_54_16_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_54_16 u_ca_54_16_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_54_16 u_ca_54_16_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_54_16 u_ca_54_16_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_54_16 u_ca_54_16_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_54_16 u_ca_54_16_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_54_16 u_ca_54_16_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_54_16 u_ca_54_16_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_54_16 u_ca_54_16_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_54_16 u_ca_54_16_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_54_16 u_ca_54_16_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_54_16 u_ca_54_16_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_54_16 u_ca_54_16_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_54_16 u_ca_54_16_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_54_16 u_ca_54_16_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_54_16 u_ca_54_16_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_54_16 u_ca_54_16_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_54_16 u_ca_54_16_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_54_16 u_ca_54_16_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_54_16 u_ca_54_16_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_54_16 u_ca_54_16_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_54_16 u_ca_54_16_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_54_16 u_ca_54_16_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_54_16 u_ca_54_16_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_54_16 u_ca_54_16_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_54_16 u_ca_54_16_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_54_16 u_ca_54_16_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_54_16 u_ca_54_16_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_54_16 u_ca_54_16_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_54_16 u_ca_54_16_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_54_16 u_ca_54_16_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_54_16 u_ca_54_16_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_54_16 u_ca_54_16_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_54_16 u_ca_54_16_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_54_16 u_ca_54_16_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_54_16 u_ca_54_16_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_54_16 u_ca_54_16_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_54_16 u_ca_54_16_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_54_16 u_ca_54_16_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_54_16 u_ca_54_16_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_54_16 u_ca_54_16_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_54_16 u_ca_54_16_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_54_16 u_ca_54_16_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_54_16 u_ca_54_16_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_54_16 u_ca_54_16_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_54_16 u_ca_54_16_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_54_16 u_ca_54_16_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_54_16 u_ca_54_16_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_54_16 u_ca_54_16_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_54_16 u_ca_54_16_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_54_16 u_ca_54_16_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_54_16 u_ca_54_16_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_54_16 u_ca_54_16_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_54_16 u_ca_54_16_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_54_16 u_ca_54_16_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_54_16 u_ca_54_16_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_54_16 u_ca_54_16_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_54_16 u_ca_54_16_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_54_16 u_ca_54_16_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_54_16 u_ca_54_16_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_54_16 u_ca_54_16_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_54_16 u_ca_54_16_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_54_16 u_ca_54_16_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_54_16 u_ca_54_16_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_54_16 u_ca_54_16_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_54_16 u_ca_54_16_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_54_16 u_ca_54_16_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_54_16 u_ca_54_16_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_54_16 u_ca_54_16_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_54_16 u_ca_54_16_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_54_16 u_ca_54_16_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_54_16 u_ca_54_16_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_54_16 u_ca_54_16_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_54_16 u_ca_54_16_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_54_16 u_ca_54_16_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_54_16 u_ca_54_16_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_54_16 u_ca_54_16_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_54_16 u_ca_54_16_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_54_16 u_ca_54_16_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_54_16 u_ca_54_16_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_54_16 u_ca_54_16_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_54_16 u_ca_54_16_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_54_16 u_ca_54_16_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_54_16 u_ca_54_16_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_54_16 u_ca_54_16_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_54_16 u_ca_54_16_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_54_16 u_ca_54_16_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_54_16 u_ca_54_16_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_54_16 u_ca_54_16_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_54_16 u_ca_54_16_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_54_16 u_ca_54_16_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_54_16 u_ca_54_16_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_54_16 u_ca_54_16_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_54_16 u_ca_54_16_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_54_16 u_ca_54_16_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_54_16 u_ca_54_16_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_54_16 u_ca_54_16_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_54_16 u_ca_54_16_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_54_16 u_ca_54_16_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_54_16 u_ca_54_16_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_54_16 u_ca_54_16_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_54_16 u_ca_54_16_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_54_16 u_ca_54_16_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_54_16 u_ca_54_16_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_54_16 u_ca_54_16_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_54_16 u_ca_54_16_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_54_16 u_ca_54_16_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_54_16 u_ca_54_16_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_54_16 u_ca_54_16_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_54_16 u_ca_54_16_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_54_16 u_ca_54_16_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_54_16 u_ca_54_16_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_54_16 u_ca_54_16_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_54_16 u_ca_54_16_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_54_16 u_ca_54_16_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_54_16 u_ca_54_16_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_54_16 u_ca_54_16_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_54_16 u_ca_54_16_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_54_16 u_ca_54_16_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_54_16 u_ca_54_16_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_54_16 u_ca_54_16_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_54_16 u_ca_54_16_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_54_16 u_ca_54_16_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_54_16 u_ca_54_16_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_54_16 u_ca_54_16_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_54_16 u_ca_54_16_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_54_16 u_ca_54_16_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_54_16 u_ca_54_16_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_54_16 u_ca_54_16_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_54_16 u_ca_54_16_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_54_16 u_ca_54_16_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_54_16 u_ca_54_16_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_54_16 u_ca_54_16_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{14{1'b0}}, u_ca_out_0[1:0]};
assign col_out_1 = {{8{1'b0}}, u_ca_out_1[1:0], u_ca_out_0[7:2]};
assign col_out_2 = {{2{1'b0}}, u_ca_out_2[1:0], u_ca_out_1[7:2], u_ca_out_0[13:8]};
assign col_out_3 = {u_ca_out_3[1:0],u_ca_out_2[7:2], u_ca_out_1[13:8], u_ca_out_0[15:14]};
assign col_out_4 = {u_ca_out_4[1:0],u_ca_out_3[7:2], u_ca_out_2[13:8], u_ca_out_1[15:14]};
assign col_out_5 = {u_ca_out_5[1:0],u_ca_out_4[7:2], u_ca_out_3[13:8], u_ca_out_2[15:14]};
assign col_out_6 = {u_ca_out_6[1:0],u_ca_out_5[7:2], u_ca_out_4[13:8], u_ca_out_3[15:14]};
assign col_out_7 = {u_ca_out_7[1:0],u_ca_out_6[7:2], u_ca_out_5[13:8], u_ca_out_4[15:14]};
assign col_out_8 = {u_ca_out_8[1:0],u_ca_out_7[7:2], u_ca_out_6[13:8], u_ca_out_5[15:14]};
assign col_out_9 = {u_ca_out_9[1:0],u_ca_out_8[7:2], u_ca_out_7[13:8], u_ca_out_6[15:14]};
assign col_out_10 = {u_ca_out_10[1:0],u_ca_out_9[7:2], u_ca_out_8[13:8], u_ca_out_7[15:14]};
assign col_out_11 = {u_ca_out_11[1:0],u_ca_out_10[7:2], u_ca_out_9[13:8], u_ca_out_8[15:14]};
assign col_out_12 = {u_ca_out_12[1:0],u_ca_out_11[7:2], u_ca_out_10[13:8], u_ca_out_9[15:14]};
assign col_out_13 = {u_ca_out_13[1:0],u_ca_out_12[7:2], u_ca_out_11[13:8], u_ca_out_10[15:14]};
assign col_out_14 = {u_ca_out_14[1:0],u_ca_out_13[7:2], u_ca_out_12[13:8], u_ca_out_11[15:14]};
assign col_out_15 = {u_ca_out_15[1:0],u_ca_out_14[7:2], u_ca_out_13[13:8], u_ca_out_12[15:14]};
assign col_out_16 = {u_ca_out_16[1:0],u_ca_out_15[7:2], u_ca_out_14[13:8], u_ca_out_13[15:14]};
assign col_out_17 = {u_ca_out_17[1:0],u_ca_out_16[7:2], u_ca_out_15[13:8], u_ca_out_14[15:14]};
assign col_out_18 = {u_ca_out_18[1:0],u_ca_out_17[7:2], u_ca_out_16[13:8], u_ca_out_15[15:14]};
assign col_out_19 = {u_ca_out_19[1:0],u_ca_out_18[7:2], u_ca_out_17[13:8], u_ca_out_16[15:14]};
assign col_out_20 = {u_ca_out_20[1:0],u_ca_out_19[7:2], u_ca_out_18[13:8], u_ca_out_17[15:14]};
assign col_out_21 = {u_ca_out_21[1:0],u_ca_out_20[7:2], u_ca_out_19[13:8], u_ca_out_18[15:14]};
assign col_out_22 = {u_ca_out_22[1:0],u_ca_out_21[7:2], u_ca_out_20[13:8], u_ca_out_19[15:14]};
assign col_out_23 = {u_ca_out_23[1:0],u_ca_out_22[7:2], u_ca_out_21[13:8], u_ca_out_20[15:14]};
assign col_out_24 = {u_ca_out_24[1:0],u_ca_out_23[7:2], u_ca_out_22[13:8], u_ca_out_21[15:14]};
assign col_out_25 = {u_ca_out_25[1:0],u_ca_out_24[7:2], u_ca_out_23[13:8], u_ca_out_22[15:14]};
assign col_out_26 = {u_ca_out_26[1:0],u_ca_out_25[7:2], u_ca_out_24[13:8], u_ca_out_23[15:14]};
assign col_out_27 = {u_ca_out_27[1:0],u_ca_out_26[7:2], u_ca_out_25[13:8], u_ca_out_24[15:14]};
assign col_out_28 = {u_ca_out_28[1:0],u_ca_out_27[7:2], u_ca_out_26[13:8], u_ca_out_25[15:14]};
assign col_out_29 = {u_ca_out_29[1:0],u_ca_out_28[7:2], u_ca_out_27[13:8], u_ca_out_26[15:14]};
assign col_out_30 = {u_ca_out_30[1:0],u_ca_out_29[7:2], u_ca_out_28[13:8], u_ca_out_27[15:14]};
assign col_out_31 = {u_ca_out_31[1:0],u_ca_out_30[7:2], u_ca_out_29[13:8], u_ca_out_28[15:14]};
assign col_out_32 = {u_ca_out_32[1:0],u_ca_out_31[7:2], u_ca_out_30[13:8], u_ca_out_29[15:14]};
assign col_out_33 = {u_ca_out_33[1:0],u_ca_out_32[7:2], u_ca_out_31[13:8], u_ca_out_30[15:14]};
assign col_out_34 = {u_ca_out_34[1:0],u_ca_out_33[7:2], u_ca_out_32[13:8], u_ca_out_31[15:14]};
assign col_out_35 = {u_ca_out_35[1:0],u_ca_out_34[7:2], u_ca_out_33[13:8], u_ca_out_32[15:14]};
assign col_out_36 = {u_ca_out_36[1:0],u_ca_out_35[7:2], u_ca_out_34[13:8], u_ca_out_33[15:14]};
assign col_out_37 = {u_ca_out_37[1:0],u_ca_out_36[7:2], u_ca_out_35[13:8], u_ca_out_34[15:14]};
assign col_out_38 = {u_ca_out_38[1:0],u_ca_out_37[7:2], u_ca_out_36[13:8], u_ca_out_35[15:14]};
assign col_out_39 = {u_ca_out_39[1:0],u_ca_out_38[7:2], u_ca_out_37[13:8], u_ca_out_36[15:14]};
assign col_out_40 = {u_ca_out_40[1:0],u_ca_out_39[7:2], u_ca_out_38[13:8], u_ca_out_37[15:14]};
assign col_out_41 = {u_ca_out_41[1:0],u_ca_out_40[7:2], u_ca_out_39[13:8], u_ca_out_38[15:14]};
assign col_out_42 = {u_ca_out_42[1:0],u_ca_out_41[7:2], u_ca_out_40[13:8], u_ca_out_39[15:14]};
assign col_out_43 = {u_ca_out_43[1:0],u_ca_out_42[7:2], u_ca_out_41[13:8], u_ca_out_40[15:14]};
assign col_out_44 = {u_ca_out_44[1:0],u_ca_out_43[7:2], u_ca_out_42[13:8], u_ca_out_41[15:14]};
assign col_out_45 = {u_ca_out_45[1:0],u_ca_out_44[7:2], u_ca_out_43[13:8], u_ca_out_42[15:14]};
assign col_out_46 = {u_ca_out_46[1:0],u_ca_out_45[7:2], u_ca_out_44[13:8], u_ca_out_43[15:14]};
assign col_out_47 = {u_ca_out_47[1:0],u_ca_out_46[7:2], u_ca_out_45[13:8], u_ca_out_44[15:14]};
assign col_out_48 = {u_ca_out_48[1:0],u_ca_out_47[7:2], u_ca_out_46[13:8], u_ca_out_45[15:14]};
assign col_out_49 = {u_ca_out_49[1:0],u_ca_out_48[7:2], u_ca_out_47[13:8], u_ca_out_46[15:14]};
assign col_out_50 = {u_ca_out_50[1:0],u_ca_out_49[7:2], u_ca_out_48[13:8], u_ca_out_47[15:14]};
assign col_out_51 = {u_ca_out_51[1:0],u_ca_out_50[7:2], u_ca_out_49[13:8], u_ca_out_48[15:14]};
assign col_out_52 = {u_ca_out_52[1:0],u_ca_out_51[7:2], u_ca_out_50[13:8], u_ca_out_49[15:14]};
assign col_out_53 = {u_ca_out_53[1:0],u_ca_out_52[7:2], u_ca_out_51[13:8], u_ca_out_50[15:14]};
assign col_out_54 = {u_ca_out_54[1:0],u_ca_out_53[7:2], u_ca_out_52[13:8], u_ca_out_51[15:14]};
assign col_out_55 = {u_ca_out_55[1:0],u_ca_out_54[7:2], u_ca_out_53[13:8], u_ca_out_52[15:14]};
assign col_out_56 = {u_ca_out_56[1:0],u_ca_out_55[7:2], u_ca_out_54[13:8], u_ca_out_53[15:14]};
assign col_out_57 = {u_ca_out_57[1:0],u_ca_out_56[7:2], u_ca_out_55[13:8], u_ca_out_54[15:14]};
assign col_out_58 = {u_ca_out_58[1:0],u_ca_out_57[7:2], u_ca_out_56[13:8], u_ca_out_55[15:14]};
assign col_out_59 = {u_ca_out_59[1:0],u_ca_out_58[7:2], u_ca_out_57[13:8], u_ca_out_56[15:14]};
assign col_out_60 = {u_ca_out_60[1:0],u_ca_out_59[7:2], u_ca_out_58[13:8], u_ca_out_57[15:14]};
assign col_out_61 = {u_ca_out_61[1:0],u_ca_out_60[7:2], u_ca_out_59[13:8], u_ca_out_58[15:14]};
assign col_out_62 = {u_ca_out_62[1:0],u_ca_out_61[7:2], u_ca_out_60[13:8], u_ca_out_59[15:14]};
assign col_out_63 = {u_ca_out_63[1:0],u_ca_out_62[7:2], u_ca_out_61[13:8], u_ca_out_60[15:14]};
assign col_out_64 = {u_ca_out_64[1:0],u_ca_out_63[7:2], u_ca_out_62[13:8], u_ca_out_61[15:14]};
assign col_out_65 = {u_ca_out_65[1:0],u_ca_out_64[7:2], u_ca_out_63[13:8], u_ca_out_62[15:14]};
assign col_out_66 = {u_ca_out_66[1:0],u_ca_out_65[7:2], u_ca_out_64[13:8], u_ca_out_63[15:14]};
assign col_out_67 = {u_ca_out_67[1:0],u_ca_out_66[7:2], u_ca_out_65[13:8], u_ca_out_64[15:14]};
assign col_out_68 = {u_ca_out_68[1:0],u_ca_out_67[7:2], u_ca_out_66[13:8], u_ca_out_65[15:14]};
assign col_out_69 = {u_ca_out_69[1:0],u_ca_out_68[7:2], u_ca_out_67[13:8], u_ca_out_66[15:14]};
assign col_out_70 = {u_ca_out_70[1:0],u_ca_out_69[7:2], u_ca_out_68[13:8], u_ca_out_67[15:14]};
assign col_out_71 = {u_ca_out_71[1:0],u_ca_out_70[7:2], u_ca_out_69[13:8], u_ca_out_68[15:14]};
assign col_out_72 = {u_ca_out_72[1:0],u_ca_out_71[7:2], u_ca_out_70[13:8], u_ca_out_69[15:14]};
assign col_out_73 = {u_ca_out_73[1:0],u_ca_out_72[7:2], u_ca_out_71[13:8], u_ca_out_70[15:14]};
assign col_out_74 = {u_ca_out_74[1:0],u_ca_out_73[7:2], u_ca_out_72[13:8], u_ca_out_71[15:14]};
assign col_out_75 = {u_ca_out_75[1:0],u_ca_out_74[7:2], u_ca_out_73[13:8], u_ca_out_72[15:14]};
assign col_out_76 = {u_ca_out_76[1:0],u_ca_out_75[7:2], u_ca_out_74[13:8], u_ca_out_73[15:14]};
assign col_out_77 = {u_ca_out_77[1:0],u_ca_out_76[7:2], u_ca_out_75[13:8], u_ca_out_74[15:14]};
assign col_out_78 = {u_ca_out_78[1:0],u_ca_out_77[7:2], u_ca_out_76[13:8], u_ca_out_75[15:14]};
assign col_out_79 = {u_ca_out_79[1:0],u_ca_out_78[7:2], u_ca_out_77[13:8], u_ca_out_76[15:14]};
assign col_out_80 = {u_ca_out_80[1:0],u_ca_out_79[7:2], u_ca_out_78[13:8], u_ca_out_77[15:14]};
assign col_out_81 = {u_ca_out_81[1:0],u_ca_out_80[7:2], u_ca_out_79[13:8], u_ca_out_78[15:14]};
assign col_out_82 = {u_ca_out_82[1:0],u_ca_out_81[7:2], u_ca_out_80[13:8], u_ca_out_79[15:14]};
assign col_out_83 = {u_ca_out_83[1:0],u_ca_out_82[7:2], u_ca_out_81[13:8], u_ca_out_80[15:14]};
assign col_out_84 = {u_ca_out_84[1:0],u_ca_out_83[7:2], u_ca_out_82[13:8], u_ca_out_81[15:14]};
assign col_out_85 = {u_ca_out_85[1:0],u_ca_out_84[7:2], u_ca_out_83[13:8], u_ca_out_82[15:14]};
assign col_out_86 = {u_ca_out_86[1:0],u_ca_out_85[7:2], u_ca_out_84[13:8], u_ca_out_83[15:14]};
assign col_out_87 = {u_ca_out_87[1:0],u_ca_out_86[7:2], u_ca_out_85[13:8], u_ca_out_84[15:14]};
assign col_out_88 = {u_ca_out_88[1:0],u_ca_out_87[7:2], u_ca_out_86[13:8], u_ca_out_85[15:14]};
assign col_out_89 = {u_ca_out_89[1:0],u_ca_out_88[7:2], u_ca_out_87[13:8], u_ca_out_86[15:14]};
assign col_out_90 = {u_ca_out_90[1:0],u_ca_out_89[7:2], u_ca_out_88[13:8], u_ca_out_87[15:14]};
assign col_out_91 = {u_ca_out_91[1:0],u_ca_out_90[7:2], u_ca_out_89[13:8], u_ca_out_88[15:14]};
assign col_out_92 = {u_ca_out_92[1:0],u_ca_out_91[7:2], u_ca_out_90[13:8], u_ca_out_89[15:14]};
assign col_out_93 = {u_ca_out_93[1:0],u_ca_out_92[7:2], u_ca_out_91[13:8], u_ca_out_90[15:14]};
assign col_out_94 = {u_ca_out_94[1:0],u_ca_out_93[7:2], u_ca_out_92[13:8], u_ca_out_91[15:14]};
assign col_out_95 = {u_ca_out_95[1:0],u_ca_out_94[7:2], u_ca_out_93[13:8], u_ca_out_92[15:14]};
assign col_out_96 = {u_ca_out_96[1:0],u_ca_out_95[7:2], u_ca_out_94[13:8], u_ca_out_93[15:14]};
assign col_out_97 = {u_ca_out_97[1:0],u_ca_out_96[7:2], u_ca_out_95[13:8], u_ca_out_94[15:14]};
assign col_out_98 = {u_ca_out_98[1:0],u_ca_out_97[7:2], u_ca_out_96[13:8], u_ca_out_95[15:14]};
assign col_out_99 = {u_ca_out_99[1:0],u_ca_out_98[7:2], u_ca_out_97[13:8], u_ca_out_96[15:14]};
assign col_out_100 = {u_ca_out_100[1:0],u_ca_out_99[7:2], u_ca_out_98[13:8], u_ca_out_97[15:14]};
assign col_out_101 = {u_ca_out_101[1:0],u_ca_out_100[7:2], u_ca_out_99[13:8], u_ca_out_98[15:14]};
assign col_out_102 = {u_ca_out_102[1:0],u_ca_out_101[7:2], u_ca_out_100[13:8], u_ca_out_99[15:14]};
assign col_out_103 = {u_ca_out_103[1:0],u_ca_out_102[7:2], u_ca_out_101[13:8], u_ca_out_100[15:14]};
assign col_out_104 = {u_ca_out_104[1:0],u_ca_out_103[7:2], u_ca_out_102[13:8], u_ca_out_101[15:14]};
assign col_out_105 = {u_ca_out_105[1:0],u_ca_out_104[7:2], u_ca_out_103[13:8], u_ca_out_102[15:14]};
assign col_out_106 = {u_ca_out_106[1:0],u_ca_out_105[7:2], u_ca_out_104[13:8], u_ca_out_103[15:14]};
assign col_out_107 = {u_ca_out_107[1:0],u_ca_out_106[7:2], u_ca_out_105[13:8], u_ca_out_104[15:14]};
assign col_out_108 = {u_ca_out_108[1:0],u_ca_out_107[7:2], u_ca_out_106[13:8], u_ca_out_105[15:14]};
assign col_out_109 = {u_ca_out_109[1:0],u_ca_out_108[7:2], u_ca_out_107[13:8], u_ca_out_106[15:14]};
assign col_out_110 = {u_ca_out_110[1:0],u_ca_out_109[7:2], u_ca_out_108[13:8], u_ca_out_107[15:14]};
assign col_out_111 = {u_ca_out_111[1:0],u_ca_out_110[7:2], u_ca_out_109[13:8], u_ca_out_108[15:14]};
assign col_out_112 = {u_ca_out_112[1:0],u_ca_out_111[7:2], u_ca_out_110[13:8], u_ca_out_109[15:14]};
assign col_out_113 = {u_ca_out_113[1:0],u_ca_out_112[7:2], u_ca_out_111[13:8], u_ca_out_110[15:14]};
assign col_out_114 = {u_ca_out_114[1:0],u_ca_out_113[7:2], u_ca_out_112[13:8], u_ca_out_111[15:14]};
assign col_out_115 = {u_ca_out_115[1:0],u_ca_out_114[7:2], u_ca_out_113[13:8], u_ca_out_112[15:14]};
assign col_out_116 = {u_ca_out_116[1:0],u_ca_out_115[7:2], u_ca_out_114[13:8], u_ca_out_113[15:14]};
assign col_out_117 = {u_ca_out_117[1:0],u_ca_out_116[7:2], u_ca_out_115[13:8], u_ca_out_114[15:14]};
assign col_out_118 = {u_ca_out_118[1:0],u_ca_out_117[7:2], u_ca_out_116[13:8], u_ca_out_115[15:14]};
assign col_out_119 = {u_ca_out_119[1:0],u_ca_out_118[7:2], u_ca_out_117[13:8], u_ca_out_116[15:14]};
assign col_out_120 = {u_ca_out_120[1:0],u_ca_out_119[7:2], u_ca_out_118[13:8], u_ca_out_117[15:14]};
assign col_out_121 = {u_ca_out_121[1:0],u_ca_out_120[7:2], u_ca_out_119[13:8], u_ca_out_118[15:14]};
assign col_out_122 = {u_ca_out_122[1:0],u_ca_out_121[7:2], u_ca_out_120[13:8], u_ca_out_119[15:14]};
assign col_out_123 = {u_ca_out_123[1:0],u_ca_out_122[7:2], u_ca_out_121[13:8], u_ca_out_120[15:14]};
assign col_out_124 = {u_ca_out_124[1:0],u_ca_out_123[7:2], u_ca_out_122[13:8], u_ca_out_121[15:14]};
assign col_out_125 = {u_ca_out_125[1:0],u_ca_out_124[7:2], u_ca_out_123[13:8], u_ca_out_122[15:14]};
assign col_out_126 = {u_ca_out_126[1:0],u_ca_out_125[7:2], u_ca_out_124[13:8], u_ca_out_123[15:14]};
assign col_out_127 = {u_ca_out_127[1:0],u_ca_out_126[7:2], u_ca_out_125[13:8], u_ca_out_124[15:14]};
assign col_out_128 = {u_ca_out_128[1:0],u_ca_out_127[7:2], u_ca_out_126[13:8], u_ca_out_125[15:14]};
assign col_out_129 = {u_ca_out_129[1:0],u_ca_out_128[7:2], u_ca_out_127[13:8], u_ca_out_126[15:14]};
assign col_out_130 = {u_ca_out_130[1:0],u_ca_out_129[7:2], u_ca_out_128[13:8], u_ca_out_127[15:14]};
assign col_out_131 = {u_ca_out_131[1:0],u_ca_out_130[7:2], u_ca_out_129[13:8], u_ca_out_128[15:14]};
assign col_out_132 = {u_ca_out_132[1:0],u_ca_out_131[7:2], u_ca_out_130[13:8], u_ca_out_129[15:14]};
assign col_out_133 = {u_ca_out_133[1:0],u_ca_out_132[7:2], u_ca_out_131[13:8], u_ca_out_130[15:14]};
assign col_out_134 = {u_ca_out_134[1:0],u_ca_out_133[7:2], u_ca_out_132[13:8], u_ca_out_131[15:14]};
assign col_out_135 = {u_ca_out_135[1:0],u_ca_out_134[7:2], u_ca_out_133[13:8], u_ca_out_132[15:14]};
assign col_out_136 = {u_ca_out_136[1:0],u_ca_out_135[7:2], u_ca_out_134[13:8], u_ca_out_133[15:14]};
assign col_out_137 = {u_ca_out_137[1:0],u_ca_out_136[7:2], u_ca_out_135[13:8], u_ca_out_134[15:14]};
assign col_out_138 = {u_ca_out_138[1:0],u_ca_out_137[7:2], u_ca_out_136[13:8], u_ca_out_135[15:14]};
assign col_out_139 = {u_ca_out_139[1:0],u_ca_out_138[7:2], u_ca_out_137[13:8], u_ca_out_136[15:14]};
assign col_out_140 = {u_ca_out_140[1:0],u_ca_out_139[7:2], u_ca_out_138[13:8], u_ca_out_137[15:14]};
assign col_out_141 = {u_ca_out_141[1:0],u_ca_out_140[7:2], u_ca_out_139[13:8], u_ca_out_138[15:14]};
assign col_out_142 = {u_ca_out_142[1:0],u_ca_out_141[7:2], u_ca_out_140[13:8], u_ca_out_139[15:14]};
assign col_out_143 = {u_ca_out_143[1:0],u_ca_out_142[7:2], u_ca_out_141[13:8], u_ca_out_140[15:14]};
assign col_out_144 = {u_ca_out_144[1:0],u_ca_out_143[7:2], u_ca_out_142[13:8], u_ca_out_141[15:14]};
assign col_out_145 = {u_ca_out_145[1:0],u_ca_out_144[7:2], u_ca_out_143[13:8], u_ca_out_142[15:14]};
assign col_out_146 = {u_ca_out_146[1:0],u_ca_out_145[7:2], u_ca_out_144[13:8], u_ca_out_143[15:14]};
assign col_out_147 = {u_ca_out_147[1:0],u_ca_out_146[7:2], u_ca_out_145[13:8], u_ca_out_144[15:14]};
assign col_out_148 = {u_ca_out_148[1:0],u_ca_out_147[7:2], u_ca_out_146[13:8], u_ca_out_145[15:14]};
assign col_out_149 = {u_ca_out_149[1:0],u_ca_out_148[7:2], u_ca_out_147[13:8], u_ca_out_146[15:14]};
assign col_out_150 = {u_ca_out_150[1:0],u_ca_out_149[7:2], u_ca_out_148[13:8], u_ca_out_147[15:14]};
assign col_out_151 = {u_ca_out_151[1:0],u_ca_out_150[7:2], u_ca_out_149[13:8], u_ca_out_148[15:14]};
assign col_out_152 = {u_ca_out_152[1:0],u_ca_out_151[7:2], u_ca_out_150[13:8], u_ca_out_149[15:14]};
assign col_out_153 = {u_ca_out_153[1:0],u_ca_out_152[7:2], u_ca_out_151[13:8], u_ca_out_150[15:14]};
assign col_out_154 = {u_ca_out_154[1:0],u_ca_out_153[7:2], u_ca_out_152[13:8], u_ca_out_151[15:14]};
assign col_out_155 = {u_ca_out_155[1:0],u_ca_out_154[7:2], u_ca_out_153[13:8], u_ca_out_152[15:14]};
assign col_out_156 = {u_ca_out_156[1:0],u_ca_out_155[7:2], u_ca_out_154[13:8], u_ca_out_153[15:14]};
assign col_out_157 = {u_ca_out_157[1:0],u_ca_out_156[7:2], u_ca_out_155[13:8], u_ca_out_154[15:14]};
assign col_out_158 = {u_ca_out_158[1:0],u_ca_out_157[7:2], u_ca_out_156[13:8], u_ca_out_155[15:14]};
assign col_out_159 = {u_ca_out_159[1:0],u_ca_out_158[7:2], u_ca_out_157[13:8], u_ca_out_156[15:14]};
assign col_out_160 = {u_ca_out_160[1:0],u_ca_out_159[7:2], u_ca_out_158[13:8], u_ca_out_157[15:14]};
assign col_out_161 = {u_ca_out_161[1:0],u_ca_out_160[7:2], u_ca_out_159[13:8], u_ca_out_158[15:14]};
assign col_out_162 = {u_ca_out_162[1:0],u_ca_out_161[7:2], u_ca_out_160[13:8], u_ca_out_159[15:14]};
assign col_out_163 = {u_ca_out_163[1:0],u_ca_out_162[7:2], u_ca_out_161[13:8], u_ca_out_160[15:14]};
assign col_out_164 = {u_ca_out_164[1:0],u_ca_out_163[7:2], u_ca_out_162[13:8], u_ca_out_161[15:14]};
assign col_out_165 = {u_ca_out_165[1:0],u_ca_out_164[7:2], u_ca_out_163[13:8], u_ca_out_162[15:14]};
assign col_out_166 = {u_ca_out_166[1:0],u_ca_out_165[7:2], u_ca_out_164[13:8], u_ca_out_163[15:14]};
assign col_out_167 = {u_ca_out_167[1:0],u_ca_out_166[7:2], u_ca_out_165[13:8], u_ca_out_164[15:14]};
assign col_out_168 = {u_ca_out_168[1:0],u_ca_out_167[7:2], u_ca_out_166[13:8], u_ca_out_165[15:14]};
assign col_out_169 = {u_ca_out_169[1:0],u_ca_out_168[7:2], u_ca_out_167[13:8], u_ca_out_166[15:14]};
assign col_out_170 = {u_ca_out_170[1:0],u_ca_out_169[7:2], u_ca_out_168[13:8], u_ca_out_167[15:14]};
assign col_out_171 = {u_ca_out_171[1:0],u_ca_out_170[7:2], u_ca_out_169[13:8], u_ca_out_168[15:14]};
assign col_out_172 = {u_ca_out_172[1:0],u_ca_out_171[7:2], u_ca_out_170[13:8], u_ca_out_169[15:14]};
assign col_out_173 = {u_ca_out_173[1:0],u_ca_out_172[7:2], u_ca_out_171[13:8], u_ca_out_170[15:14]};
assign col_out_174 = {u_ca_out_174[1:0],u_ca_out_173[7:2], u_ca_out_172[13:8], u_ca_out_171[15:14]};
assign col_out_175 = {u_ca_out_175[1:0],u_ca_out_174[7:2], u_ca_out_173[13:8], u_ca_out_172[15:14]};
assign col_out_176 = {u_ca_out_176[1:0],u_ca_out_175[7:2], u_ca_out_174[13:8], u_ca_out_173[15:14]};
assign col_out_177 = {u_ca_out_177[1:0],u_ca_out_176[7:2], u_ca_out_175[13:8], u_ca_out_174[15:14]};
assign col_out_178 = {u_ca_out_178[1:0],u_ca_out_177[7:2], u_ca_out_176[13:8], u_ca_out_175[15:14]};
assign col_out_179 = {u_ca_out_179[1:0],u_ca_out_178[7:2], u_ca_out_177[13:8], u_ca_out_176[15:14]};
assign col_out_180 = {u_ca_out_180[1:0],u_ca_out_179[7:2], u_ca_out_178[13:8], u_ca_out_177[15:14]};
assign col_out_181 = {u_ca_out_181[1:0],u_ca_out_180[7:2], u_ca_out_179[13:8], u_ca_out_178[15:14]};
assign col_out_182 = {u_ca_out_182[1:0],u_ca_out_181[7:2], u_ca_out_180[13:8], u_ca_out_179[15:14]};
assign col_out_183 = {u_ca_out_183[1:0],u_ca_out_182[7:2], u_ca_out_181[13:8], u_ca_out_180[15:14]};
assign col_out_184 = {u_ca_out_184[1:0],u_ca_out_183[7:2], u_ca_out_182[13:8], u_ca_out_181[15:14]};
assign col_out_185 = {u_ca_out_185[1:0],u_ca_out_184[7:2], u_ca_out_183[13:8], u_ca_out_182[15:14]};
assign col_out_186 = {u_ca_out_186[1:0],u_ca_out_185[7:2], u_ca_out_184[13:8], u_ca_out_183[15:14]};
assign col_out_187 = {u_ca_out_187[1:0],u_ca_out_186[7:2], u_ca_out_185[13:8], u_ca_out_184[15:14]};
assign col_out_188 = {u_ca_out_188[1:0],u_ca_out_187[7:2], u_ca_out_186[13:8], u_ca_out_185[15:14]};
assign col_out_189 = {u_ca_out_189[1:0],u_ca_out_188[7:2], u_ca_out_187[13:8], u_ca_out_186[15:14]};
assign col_out_190 = {u_ca_out_190[1:0],u_ca_out_189[7:2], u_ca_out_188[13:8], u_ca_out_187[15:14]};
assign col_out_191 = {u_ca_out_191[1:0],u_ca_out_190[7:2], u_ca_out_189[13:8], u_ca_out_188[15:14]};
assign col_out_192 = {u_ca_out_192[1:0],u_ca_out_191[7:2], u_ca_out_190[13:8], u_ca_out_189[15:14]};
assign col_out_193 = {u_ca_out_193[1:0],u_ca_out_192[7:2], u_ca_out_191[13:8], u_ca_out_190[15:14]};
assign col_out_194 = {u_ca_out_194[1:0],u_ca_out_193[7:2], u_ca_out_192[13:8], u_ca_out_191[15:14]};
assign col_out_195 = {u_ca_out_195[1:0],u_ca_out_194[7:2], u_ca_out_193[13:8], u_ca_out_192[15:14]};
assign col_out_196 = {u_ca_out_196[1:0],u_ca_out_195[7:2], u_ca_out_194[13:8], u_ca_out_193[15:14]};
assign col_out_197 = {u_ca_out_197[1:0],u_ca_out_196[7:2], u_ca_out_195[13:8], u_ca_out_194[15:14]};
assign col_out_198 = {u_ca_out_198[1:0],u_ca_out_197[7:2], u_ca_out_196[13:8], u_ca_out_195[15:14]};
assign col_out_199 = {u_ca_out_199[1:0],u_ca_out_198[7:2], u_ca_out_197[13:8], u_ca_out_196[15:14]};
assign col_out_200 = {u_ca_out_200[1:0],u_ca_out_199[7:2], u_ca_out_198[13:8], u_ca_out_197[15:14]};
assign col_out_201 = {u_ca_out_201[1:0],u_ca_out_200[7:2], u_ca_out_199[13:8], u_ca_out_198[15:14]};
assign col_out_202 = {u_ca_out_202[1:0],u_ca_out_201[7:2], u_ca_out_200[13:8], u_ca_out_199[15:14]};
assign col_out_203 = {u_ca_out_203[1:0],u_ca_out_202[7:2], u_ca_out_201[13:8], u_ca_out_200[15:14]};
assign col_out_204 = {u_ca_out_204[1:0],u_ca_out_203[7:2], u_ca_out_202[13:8], u_ca_out_201[15:14]};
assign col_out_205 = {u_ca_out_205[1:0],u_ca_out_204[7:2], u_ca_out_203[13:8], u_ca_out_202[15:14]};
assign col_out_206 = {u_ca_out_206[1:0],u_ca_out_205[7:2], u_ca_out_204[13:8], u_ca_out_203[15:14]};
assign col_out_207 = {u_ca_out_207[1:0],u_ca_out_206[7:2], u_ca_out_205[13:8], u_ca_out_204[15:14]};
assign col_out_208 = {u_ca_out_208[1:0],u_ca_out_207[7:2], u_ca_out_206[13:8], u_ca_out_205[15:14]};
assign col_out_209 = {u_ca_out_209[1:0],u_ca_out_208[7:2], u_ca_out_207[13:8], u_ca_out_206[15:14]};
assign col_out_210 = {u_ca_out_210[1:0],u_ca_out_209[7:2], u_ca_out_208[13:8], u_ca_out_207[15:14]};
assign col_out_211 = {u_ca_out_211[1:0],u_ca_out_210[7:2], u_ca_out_209[13:8], u_ca_out_208[15:14]};
assign col_out_212 = {u_ca_out_212[1:0],u_ca_out_211[7:2], u_ca_out_210[13:8], u_ca_out_209[15:14]};
assign col_out_213 = {u_ca_out_213[1:0],u_ca_out_212[7:2], u_ca_out_211[13:8], u_ca_out_210[15:14]};
assign col_out_214 = {u_ca_out_214[1:0],u_ca_out_213[7:2], u_ca_out_212[13:8], u_ca_out_211[15:14]};
assign col_out_215 = {u_ca_out_215[1:0],u_ca_out_214[7:2], u_ca_out_213[13:8], u_ca_out_212[15:14]};
assign col_out_216 = {u_ca_out_216[1:0],u_ca_out_215[7:2], u_ca_out_214[13:8], u_ca_out_213[15:14]};
assign col_out_217 = {u_ca_out_217[1:0],u_ca_out_216[7:2], u_ca_out_215[13:8], u_ca_out_214[15:14]};
assign col_out_218 = {u_ca_out_218[1:0],u_ca_out_217[7:2], u_ca_out_216[13:8], u_ca_out_215[15:14]};
assign col_out_219 = {u_ca_out_219[1:0],u_ca_out_218[7:2], u_ca_out_217[13:8], u_ca_out_216[15:14]};
assign col_out_220 = {u_ca_out_220[1:0],u_ca_out_219[7:2], u_ca_out_218[13:8], u_ca_out_217[15:14]};
assign col_out_221 = {u_ca_out_221[1:0],u_ca_out_220[7:2], u_ca_out_219[13:8], u_ca_out_218[15:14]};
assign col_out_222 = {u_ca_out_222[1:0],u_ca_out_221[7:2], u_ca_out_220[13:8], u_ca_out_219[15:14]};
assign col_out_223 = {u_ca_out_223[1:0],u_ca_out_222[7:2], u_ca_out_221[13:8], u_ca_out_220[15:14]};
assign col_out_224 = {u_ca_out_224[1:0],u_ca_out_223[7:2], u_ca_out_222[13:8], u_ca_out_221[15:14]};
assign col_out_225 = {u_ca_out_225[1:0],u_ca_out_224[7:2], u_ca_out_223[13:8], u_ca_out_222[15:14]};
assign col_out_226 = {u_ca_out_226[1:0],u_ca_out_225[7:2], u_ca_out_224[13:8], u_ca_out_223[15:14]};
assign col_out_227 = {u_ca_out_227[1:0],u_ca_out_226[7:2], u_ca_out_225[13:8], u_ca_out_224[15:14]};
assign col_out_228 = {u_ca_out_228[1:0],u_ca_out_227[7:2], u_ca_out_226[13:8], u_ca_out_225[15:14]};
assign col_out_229 = {u_ca_out_229[1:0],u_ca_out_228[7:2], u_ca_out_227[13:8], u_ca_out_226[15:14]};
assign col_out_230 = {u_ca_out_230[1:0],u_ca_out_229[7:2], u_ca_out_228[13:8], u_ca_out_227[15:14]};
assign col_out_231 = {u_ca_out_231[1:0],u_ca_out_230[7:2], u_ca_out_229[13:8], u_ca_out_228[15:14]};
assign col_out_232 = {u_ca_out_232[1:0],u_ca_out_231[7:2], u_ca_out_230[13:8], u_ca_out_229[15:14]};
assign col_out_233 = {u_ca_out_233[1:0],u_ca_out_232[7:2], u_ca_out_231[13:8], u_ca_out_230[15:14]};
assign col_out_234 = {u_ca_out_234[1:0],u_ca_out_233[7:2], u_ca_out_232[13:8], u_ca_out_231[15:14]};
assign col_out_235 = {u_ca_out_235[1:0],u_ca_out_234[7:2], u_ca_out_233[13:8], u_ca_out_232[15:14]};
assign col_out_236 = {u_ca_out_236[1:0],u_ca_out_235[7:2], u_ca_out_234[13:8], u_ca_out_233[15:14]};
assign col_out_237 = {u_ca_out_237[1:0],u_ca_out_236[7:2], u_ca_out_235[13:8], u_ca_out_234[15:14]};
assign col_out_238 = {u_ca_out_238[1:0],u_ca_out_237[7:2], u_ca_out_236[13:8], u_ca_out_235[15:14]};
assign col_out_239 = {u_ca_out_239[1:0],u_ca_out_238[7:2], u_ca_out_237[13:8], u_ca_out_236[15:14]};
assign col_out_240 = {u_ca_out_240[1:0],u_ca_out_239[7:2], u_ca_out_238[13:8], u_ca_out_237[15:14]};
assign col_out_241 = {u_ca_out_241[1:0],u_ca_out_240[7:2], u_ca_out_239[13:8], u_ca_out_238[15:14]};
assign col_out_242 = {u_ca_out_242[1:0],u_ca_out_241[7:2], u_ca_out_240[13:8], u_ca_out_239[15:14]};
assign col_out_243 = {u_ca_out_243[1:0],u_ca_out_242[7:2], u_ca_out_241[13:8], u_ca_out_240[15:14]};
assign col_out_244 = {u_ca_out_244[1:0],u_ca_out_243[7:2], u_ca_out_242[13:8], u_ca_out_241[15:14]};
assign col_out_245 = {u_ca_out_245[1:0],u_ca_out_244[7:2], u_ca_out_243[13:8], u_ca_out_242[15:14]};
assign col_out_246 = {u_ca_out_246[1:0],u_ca_out_245[7:2], u_ca_out_244[13:8], u_ca_out_243[15:14]};
assign col_out_247 = {u_ca_out_247[1:0],u_ca_out_246[7:2], u_ca_out_245[13:8], u_ca_out_244[15:14]};
assign col_out_248 = {u_ca_out_248[1:0],u_ca_out_247[7:2], u_ca_out_246[13:8], u_ca_out_245[15:14]};
assign col_out_249 = {u_ca_out_249[1:0],u_ca_out_248[7:2], u_ca_out_247[13:8], u_ca_out_246[15:14]};
assign col_out_250 = {u_ca_out_250[1:0],u_ca_out_249[7:2], u_ca_out_248[13:8], u_ca_out_247[15:14]};
assign col_out_251 = {u_ca_out_251[1:0],u_ca_out_250[7:2], u_ca_out_249[13:8], u_ca_out_248[15:14]};
assign col_out_252 = {u_ca_out_252[1:0],u_ca_out_251[7:2], u_ca_out_250[13:8], u_ca_out_249[15:14]};
assign col_out_253 = {u_ca_out_253[1:0],u_ca_out_252[7:2], u_ca_out_251[13:8], u_ca_out_250[15:14]};
assign col_out_254 = {u_ca_out_254[1:0],u_ca_out_253[7:2], u_ca_out_252[13:8], u_ca_out_251[15:14]};
assign col_out_255 = {u_ca_out_255[1:0],u_ca_out_254[7:2], u_ca_out_253[13:8], u_ca_out_252[15:14]};
assign col_out_256 = {u_ca_out_256[1:0],u_ca_out_255[7:2], u_ca_out_254[13:8], u_ca_out_253[15:14]};
assign col_out_257 = {u_ca_out_257[1:0],u_ca_out_256[7:2], u_ca_out_255[13:8], u_ca_out_254[15:14]};
assign col_out_258 = {u_ca_out_258[1:0],u_ca_out_257[7:2], u_ca_out_256[13:8], u_ca_out_255[15:14]};
assign col_out_259 = {u_ca_out_259[1:0],u_ca_out_258[7:2], u_ca_out_257[13:8], u_ca_out_256[15:14]};
assign col_out_260 = {u_ca_out_260[1:0],u_ca_out_259[7:2], u_ca_out_258[13:8], u_ca_out_257[15:14]};
assign col_out_261 = {u_ca_out_261[1:0],u_ca_out_260[7:2], u_ca_out_259[13:8], u_ca_out_258[15:14]};
assign col_out_262 = {u_ca_out_262[1:0],u_ca_out_261[7:2], u_ca_out_260[13:8], u_ca_out_259[15:14]};
assign col_out_263 = {u_ca_out_263[1:0],u_ca_out_262[7:2], u_ca_out_261[13:8], u_ca_out_260[15:14]};
assign col_out_264 = {u_ca_out_264[1:0],u_ca_out_263[7:2], u_ca_out_262[13:8], u_ca_out_261[15:14]};
assign col_out_265 = {u_ca_out_265[1:0],u_ca_out_264[7:2], u_ca_out_263[13:8], u_ca_out_262[15:14]};
assign col_out_266 = {u_ca_out_266[1:0],u_ca_out_265[7:2], u_ca_out_264[13:8], u_ca_out_263[15:14]};
assign col_out_267 = {u_ca_out_267[1:0],u_ca_out_266[7:2], u_ca_out_265[13:8], u_ca_out_264[15:14]};
assign col_out_268 = {u_ca_out_268[1:0],u_ca_out_267[7:2], u_ca_out_266[13:8], u_ca_out_265[15:14]};
assign col_out_269 = {u_ca_out_269[1:0],u_ca_out_268[7:2], u_ca_out_267[13:8], u_ca_out_266[15:14]};
assign col_out_270 = {u_ca_out_270[1:0],u_ca_out_269[7:2], u_ca_out_268[13:8], u_ca_out_267[15:14]};
assign col_out_271 = {u_ca_out_271[1:0],u_ca_out_270[7:2], u_ca_out_269[13:8], u_ca_out_268[15:14]};
assign col_out_272 = {u_ca_out_272[1:0],u_ca_out_271[7:2], u_ca_out_270[13:8], u_ca_out_269[15:14]};
assign col_out_273 = {u_ca_out_273[1:0],u_ca_out_272[7:2], u_ca_out_271[13:8], u_ca_out_270[15:14]};
assign col_out_274 = {u_ca_out_274[1:0],u_ca_out_273[7:2], u_ca_out_272[13:8], u_ca_out_271[15:14]};
assign col_out_275 = {u_ca_out_275[1:0],u_ca_out_274[7:2], u_ca_out_273[13:8], u_ca_out_272[15:14]};
assign col_out_276 = {u_ca_out_276[1:0],u_ca_out_275[7:2], u_ca_out_274[13:8], u_ca_out_273[15:14]};
assign col_out_277 = {u_ca_out_277[1:0],u_ca_out_276[7:2], u_ca_out_275[13:8], u_ca_out_274[15:14]};
assign col_out_278 = {u_ca_out_278[1:0],u_ca_out_277[7:2], u_ca_out_276[13:8], u_ca_out_275[15:14]};
assign col_out_279 = {u_ca_out_279[1:0],u_ca_out_278[7:2], u_ca_out_277[13:8], u_ca_out_276[15:14]};
assign col_out_280 = {u_ca_out_280[1:0],u_ca_out_279[7:2], u_ca_out_278[13:8], u_ca_out_277[15:14]};
assign col_out_281 = {u_ca_out_281[1:0],u_ca_out_280[7:2], u_ca_out_279[13:8], u_ca_out_278[15:14]};
assign col_out_282 = {u_ca_out_282[1:0],u_ca_out_281[7:2], u_ca_out_280[13:8], u_ca_out_279[15:14]};
assign col_out_283 = {u_ca_out_283[1:0],u_ca_out_282[7:2], u_ca_out_281[13:8], u_ca_out_280[15:14]};
assign col_out_284 = {u_ca_out_284[1:0],u_ca_out_283[7:2], u_ca_out_282[13:8], u_ca_out_281[15:14]};
assign col_out_285 = {u_ca_out_285[1:0],u_ca_out_284[7:2], u_ca_out_283[13:8], u_ca_out_282[15:14]};
assign col_out_286 = {u_ca_out_286[1:0],u_ca_out_285[7:2], u_ca_out_284[13:8], u_ca_out_283[15:14]};
assign col_out_287 = {u_ca_out_287[1:0],u_ca_out_286[7:2], u_ca_out_285[13:8], u_ca_out_284[15:14]};
assign col_out_288 = {u_ca_out_288[1:0],u_ca_out_287[7:2], u_ca_out_286[13:8], u_ca_out_285[15:14]};
assign col_out_289 = {u_ca_out_289[1:0],u_ca_out_288[7:2], u_ca_out_287[13:8], u_ca_out_286[15:14]};
assign col_out_290 = {u_ca_out_290[1:0],u_ca_out_289[7:2], u_ca_out_288[13:8], u_ca_out_287[15:14]};
assign col_out_291 = {u_ca_out_291[1:0],u_ca_out_290[7:2], u_ca_out_289[13:8], u_ca_out_288[15:14]};
assign col_out_292 = {u_ca_out_292[1:0],u_ca_out_291[7:2], u_ca_out_290[13:8], u_ca_out_289[15:14]};
assign col_out_293 = {u_ca_out_293[1:0],u_ca_out_292[7:2], u_ca_out_291[13:8], u_ca_out_290[15:14]};
assign col_out_294 = {u_ca_out_294[1:0],u_ca_out_293[7:2], u_ca_out_292[13:8], u_ca_out_291[15:14]};
assign col_out_295 = {u_ca_out_295[1:0],u_ca_out_294[7:2], u_ca_out_293[13:8], u_ca_out_292[15:14]};
assign col_out_296 = {u_ca_out_296[1:0],u_ca_out_295[7:2], u_ca_out_294[13:8], u_ca_out_293[15:14]};
assign col_out_297 = {u_ca_out_297[1:0],u_ca_out_296[7:2], u_ca_out_295[13:8], u_ca_out_294[15:14]};
assign col_out_298 = {u_ca_out_298[1:0],u_ca_out_297[7:2], u_ca_out_296[13:8], u_ca_out_295[15:14]};
assign col_out_299 = {u_ca_out_299[1:0],u_ca_out_298[7:2], u_ca_out_297[13:8], u_ca_out_296[15:14]};
assign col_out_300 = {u_ca_out_300[1:0],u_ca_out_299[7:2], u_ca_out_298[13:8], u_ca_out_297[15:14]};
assign col_out_301 = {u_ca_out_301[1:0],u_ca_out_300[7:2], u_ca_out_299[13:8], u_ca_out_298[15:14]};
assign col_out_302 = {u_ca_out_302[1:0],u_ca_out_301[7:2], u_ca_out_300[13:8], u_ca_out_299[15:14]};
assign col_out_303 = {u_ca_out_303[1:0],u_ca_out_302[7:2], u_ca_out_301[13:8], u_ca_out_300[15:14]};
assign col_out_304 = {u_ca_out_304[1:0],u_ca_out_303[7:2], u_ca_out_302[13:8], u_ca_out_301[15:14]};
assign col_out_305 = {u_ca_out_305[1:0],u_ca_out_304[7:2], u_ca_out_303[13:8], u_ca_out_302[15:14]};
assign col_out_306 = {u_ca_out_306[1:0],u_ca_out_305[7:2], u_ca_out_304[13:8], u_ca_out_303[15:14]};
assign col_out_307 = {u_ca_out_307[1:0],u_ca_out_306[7:2], u_ca_out_305[13:8], u_ca_out_304[15:14]};
assign col_out_308 = {u_ca_out_308[1:0],u_ca_out_307[7:2], u_ca_out_306[13:8], u_ca_out_305[15:14]};
assign col_out_309 = {u_ca_out_309[1:0],u_ca_out_308[7:2], u_ca_out_307[13:8], u_ca_out_306[15:14]};
assign col_out_310 = {u_ca_out_310[1:0],u_ca_out_309[7:2], u_ca_out_308[13:8], u_ca_out_307[15:14]};
assign col_out_311 = {u_ca_out_311[1:0],u_ca_out_310[7:2], u_ca_out_309[13:8], u_ca_out_308[15:14]};
assign col_out_312 = {u_ca_out_312[1:0],u_ca_out_311[7:2], u_ca_out_310[13:8], u_ca_out_309[15:14]};
assign col_out_313 = {u_ca_out_313[1:0],u_ca_out_312[7:2], u_ca_out_311[13:8], u_ca_out_310[15:14]};
assign col_out_314 = {u_ca_out_314[1:0],u_ca_out_313[7:2], u_ca_out_312[13:8], u_ca_out_311[15:14]};
assign col_out_315 = {u_ca_out_315[1:0],u_ca_out_314[7:2], u_ca_out_313[13:8], u_ca_out_312[15:14]};
assign col_out_316 = {u_ca_out_316[1:0],u_ca_out_315[7:2], u_ca_out_314[13:8], u_ca_out_313[15:14]};
assign col_out_317 = {u_ca_out_317[1:0],u_ca_out_316[7:2], u_ca_out_315[13:8], u_ca_out_314[15:14]};
assign col_out_318 = {u_ca_out_318[1:0],u_ca_out_317[7:2], u_ca_out_316[13:8], u_ca_out_315[15:14]};
assign col_out_319 = {u_ca_out_319[1:0],u_ca_out_318[7:2], u_ca_out_317[13:8], u_ca_out_316[15:14]};
assign col_out_320 = {u_ca_out_320[1:0],u_ca_out_319[7:2], u_ca_out_318[13:8], u_ca_out_317[15:14]};
assign col_out_321 = {u_ca_out_321[1:0],u_ca_out_320[7:2], u_ca_out_319[13:8], u_ca_out_318[15:14]};
assign col_out_322 = {u_ca_out_322[1:0],u_ca_out_321[7:2], u_ca_out_320[13:8], u_ca_out_319[15:14]};
assign col_out_323 = {u_ca_out_323[1:0],u_ca_out_322[7:2], u_ca_out_321[13:8], u_ca_out_320[15:14]};
assign col_out_324 = {u_ca_out_324[1:0],u_ca_out_323[7:2], u_ca_out_322[13:8], u_ca_out_321[15:14]};
assign col_out_325 = {u_ca_out_325[1:0],u_ca_out_324[7:2], u_ca_out_323[13:8], u_ca_out_322[15:14]};
assign col_out_326 = {u_ca_out_326[1:0],u_ca_out_325[7:2], u_ca_out_324[13:8], u_ca_out_323[15:14]};
assign col_out_327 = {u_ca_out_327[1:0],u_ca_out_326[7:2], u_ca_out_325[13:8], u_ca_out_324[15:14]};
assign col_out_328 = {u_ca_out_328[1:0],u_ca_out_327[7:2], u_ca_out_326[13:8], u_ca_out_325[15:14]};
assign col_out_329 = {u_ca_out_329[1:0],u_ca_out_328[7:2], u_ca_out_327[13:8], u_ca_out_326[15:14]};
assign col_out_330 = {u_ca_out_330[1:0],u_ca_out_329[7:2], u_ca_out_328[13:8], u_ca_out_327[15:14]};
assign col_out_331 = {u_ca_out_331[1:0],u_ca_out_330[7:2], u_ca_out_329[13:8], u_ca_out_328[15:14]};
assign col_out_332 = {u_ca_out_332[1:0],u_ca_out_331[7:2], u_ca_out_330[13:8], u_ca_out_329[15:14]};
assign col_out_333 = {u_ca_out_333[1:0],u_ca_out_332[7:2], u_ca_out_331[13:8], u_ca_out_330[15:14]};
assign col_out_334 = {u_ca_out_334[1:0],u_ca_out_333[7:2], u_ca_out_332[13:8], u_ca_out_331[15:14]};
assign col_out_335 = {u_ca_out_335[1:0],u_ca_out_334[7:2], u_ca_out_333[13:8], u_ca_out_332[15:14]};
assign col_out_336 = {u_ca_out_336[1:0],u_ca_out_335[7:2], u_ca_out_334[13:8], u_ca_out_333[15:14]};
assign col_out_337 = {u_ca_out_337[1:0],u_ca_out_336[7:2], u_ca_out_335[13:8], u_ca_out_334[15:14]};
assign col_out_338 = {u_ca_out_338[1:0],u_ca_out_337[7:2], u_ca_out_336[13:8], u_ca_out_335[15:14]};
assign col_out_339 = {u_ca_out_339[1:0],u_ca_out_338[7:2], u_ca_out_337[13:8], u_ca_out_336[15:14]};
assign col_out_340 = {u_ca_out_340[1:0],u_ca_out_339[7:2], u_ca_out_338[13:8], u_ca_out_337[15:14]};
assign col_out_341 = {u_ca_out_341[1:0],u_ca_out_340[7:2], u_ca_out_339[13:8], u_ca_out_338[15:14]};
assign col_out_342 = {u_ca_out_342[1:0],u_ca_out_341[7:2], u_ca_out_340[13:8], u_ca_out_339[15:14]};
assign col_out_343 = {u_ca_out_343[1:0],u_ca_out_342[7:2], u_ca_out_341[13:8], u_ca_out_340[15:14]};
assign col_out_344 = {u_ca_out_344[1:0],u_ca_out_343[7:2], u_ca_out_342[13:8], u_ca_out_341[15:14]};
assign col_out_345 = {u_ca_out_345[1:0],u_ca_out_344[7:2], u_ca_out_343[13:8], u_ca_out_342[15:14]};
assign col_out_346 = {u_ca_out_346[1:0],u_ca_out_345[7:2], u_ca_out_344[13:8], u_ca_out_343[15:14]};
assign col_out_347 = {u_ca_out_347[1:0],u_ca_out_346[7:2], u_ca_out_345[13:8], u_ca_out_344[15:14]};
assign col_out_348 = {u_ca_out_348[1:0],u_ca_out_347[7:2], u_ca_out_346[13:8], u_ca_out_345[15:14]};
assign col_out_349 = {u_ca_out_349[1:0],u_ca_out_348[7:2], u_ca_out_347[13:8], u_ca_out_346[15:14]};
assign col_out_350 = {u_ca_out_350[1:0],u_ca_out_349[7:2], u_ca_out_348[13:8], u_ca_out_347[15:14]};
assign col_out_351 = {u_ca_out_351[1:0],u_ca_out_350[7:2], u_ca_out_349[13:8], u_ca_out_348[15:14]};
assign col_out_352 = {u_ca_out_352[1:0],u_ca_out_351[7:2], u_ca_out_350[13:8], u_ca_out_349[15:14]};
assign col_out_353 = {u_ca_out_353[1:0],u_ca_out_352[7:2], u_ca_out_351[13:8], u_ca_out_350[15:14]};
assign col_out_354 = {u_ca_out_354[1:0],u_ca_out_353[7:2], u_ca_out_352[13:8], u_ca_out_351[15:14]};
assign col_out_355 = {u_ca_out_355[1:0],u_ca_out_354[7:2], u_ca_out_353[13:8], u_ca_out_352[15:14]};
assign col_out_356 = {u_ca_out_356[1:0],u_ca_out_355[7:2], u_ca_out_354[13:8], u_ca_out_353[15:14]};
assign col_out_357 = {u_ca_out_357[1:0],u_ca_out_356[7:2], u_ca_out_355[13:8], u_ca_out_354[15:14]};
assign col_out_358 = {u_ca_out_358[1:0],u_ca_out_357[7:2], u_ca_out_356[13:8], u_ca_out_355[15:14]};
assign col_out_359 = {u_ca_out_359[1:0],u_ca_out_358[7:2], u_ca_out_357[13:8], u_ca_out_356[15:14]};
assign col_out_360 = {u_ca_out_360[1:0],u_ca_out_359[7:2], u_ca_out_358[13:8], u_ca_out_357[15:14]};
assign col_out_361 = {u_ca_out_361[1:0],u_ca_out_360[7:2], u_ca_out_359[13:8], u_ca_out_358[15:14]};
assign col_out_362 = {u_ca_out_362[1:0],u_ca_out_361[7:2], u_ca_out_360[13:8], u_ca_out_359[15:14]};
assign col_out_363 = {u_ca_out_363[1:0],u_ca_out_362[7:2], u_ca_out_361[13:8], u_ca_out_360[15:14]};
assign col_out_364 = {u_ca_out_364[1:0],u_ca_out_363[7:2], u_ca_out_362[13:8], u_ca_out_361[15:14]};
assign col_out_365 = {u_ca_out_365[1:0],u_ca_out_364[7:2], u_ca_out_363[13:8], u_ca_out_362[15:14]};
assign col_out_366 = {u_ca_out_366[1:0],u_ca_out_365[7:2], u_ca_out_364[13:8], u_ca_out_363[15:14]};
assign col_out_367 = {u_ca_out_367[1:0],u_ca_out_366[7:2], u_ca_out_365[13:8], u_ca_out_364[15:14]};
assign col_out_368 = {u_ca_out_368[1:0],u_ca_out_367[7:2], u_ca_out_366[13:8], u_ca_out_365[15:14]};
assign col_out_369 = {u_ca_out_369[1:0],u_ca_out_368[7:2], u_ca_out_367[13:8], u_ca_out_366[15:14]};
assign col_out_370 = {u_ca_out_370[1:0],u_ca_out_369[7:2], u_ca_out_368[13:8], u_ca_out_367[15:14]};
assign col_out_371 = {u_ca_out_371[1:0],u_ca_out_370[7:2], u_ca_out_369[13:8], u_ca_out_368[15:14]};
assign col_out_372 = {u_ca_out_372[1:0],u_ca_out_371[7:2], u_ca_out_370[13:8], u_ca_out_369[15:14]};
assign col_out_373 = {u_ca_out_373[1:0],u_ca_out_372[7:2], u_ca_out_371[13:8], u_ca_out_370[15:14]};
assign col_out_374 = {u_ca_out_374[1:0],u_ca_out_373[7:2], u_ca_out_372[13:8], u_ca_out_371[15:14]};
assign col_out_375 = {u_ca_out_375[1:0],u_ca_out_374[7:2], u_ca_out_373[13:8], u_ca_out_372[15:14]};
assign col_out_376 = {u_ca_out_376[1:0],u_ca_out_375[7:2], u_ca_out_374[13:8], u_ca_out_373[15:14]};
assign col_out_377 = {u_ca_out_377[1:0],u_ca_out_376[7:2], u_ca_out_375[13:8], u_ca_out_374[15:14]};
assign col_out_378 = {u_ca_out_378[1:0],u_ca_out_377[7:2], u_ca_out_376[13:8], u_ca_out_375[15:14]};
assign col_out_379 = {u_ca_out_379[1:0],u_ca_out_378[7:2], u_ca_out_377[13:8], u_ca_out_376[15:14]};
assign col_out_380 = {u_ca_out_380[1:0],u_ca_out_379[7:2], u_ca_out_378[13:8], u_ca_out_377[15:14]};
assign col_out_381 = {u_ca_out_381[1:0],u_ca_out_380[7:2], u_ca_out_379[13:8], u_ca_out_378[15:14]};
assign col_out_382 = {u_ca_out_382[1:0],u_ca_out_381[7:2], u_ca_out_380[13:8], u_ca_out_379[15:14]};
assign col_out_383 = {u_ca_out_383[1:0],u_ca_out_382[7:2], u_ca_out_381[13:8], u_ca_out_380[15:14]};
assign col_out_384 = {u_ca_out_384[1:0],u_ca_out_383[7:2], u_ca_out_382[13:8], u_ca_out_381[15:14]};
assign col_out_385 = {u_ca_out_385[1:0],u_ca_out_384[7:2], u_ca_out_383[13:8], u_ca_out_382[15:14]};
assign col_out_386 = {u_ca_out_386[1:0],u_ca_out_385[7:2], u_ca_out_384[13:8], u_ca_out_383[15:14]};
assign col_out_387 = {u_ca_out_387[1:0],u_ca_out_386[7:2], u_ca_out_385[13:8], u_ca_out_384[15:14]};
assign col_out_388 = {u_ca_out_388[1:0],u_ca_out_387[7:2], u_ca_out_386[13:8], u_ca_out_385[15:14]};
assign col_out_389 = {u_ca_out_389[1:0],u_ca_out_388[7:2], u_ca_out_387[13:8], u_ca_out_386[15:14]};
assign col_out_390 = {u_ca_out_390[1:0],u_ca_out_389[7:2], u_ca_out_388[13:8], u_ca_out_387[15:14]};
assign col_out_391 = {u_ca_out_391[1:0],u_ca_out_390[7:2], u_ca_out_389[13:8], u_ca_out_388[15:14]};
assign col_out_392 = {u_ca_out_392[1:0],u_ca_out_391[7:2], u_ca_out_390[13:8], u_ca_out_389[15:14]};
assign col_out_393 = {u_ca_out_393[1:0],u_ca_out_392[7:2], u_ca_out_391[13:8], u_ca_out_390[15:14]};
assign col_out_394 = {u_ca_out_394[1:0],u_ca_out_393[7:2], u_ca_out_392[13:8], u_ca_out_391[15:14]};
assign col_out_395 = {u_ca_out_395[1:0],u_ca_out_394[7:2], u_ca_out_393[13:8], u_ca_out_392[15:14]};
assign col_out_396 = {u_ca_out_396[1:0],u_ca_out_395[7:2], u_ca_out_394[13:8], u_ca_out_393[15:14]};
assign col_out_397 = {u_ca_out_397[1:0],u_ca_out_396[7:2], u_ca_out_395[13:8], u_ca_out_394[15:14]};
assign col_out_398 = {u_ca_out_398[1:0],u_ca_out_397[7:2], u_ca_out_396[13:8], u_ca_out_395[15:14]};
assign col_out_399 = {u_ca_out_399[1:0],u_ca_out_398[7:2], u_ca_out_397[13:8], u_ca_out_396[15:14]};
assign col_out_400 = {u_ca_out_400[1:0],u_ca_out_399[7:2], u_ca_out_398[13:8], u_ca_out_397[15:14]};
assign col_out_401 = {u_ca_out_401[1:0],u_ca_out_400[7:2], u_ca_out_399[13:8], u_ca_out_398[15:14]};
assign col_out_402 = {u_ca_out_402[1:0],u_ca_out_401[7:2], u_ca_out_400[13:8], u_ca_out_399[15:14]};
assign col_out_403 = {u_ca_out_403[1:0],u_ca_out_402[7:2], u_ca_out_401[13:8], u_ca_out_400[15:14]};
assign col_out_404 = {u_ca_out_404[1:0],u_ca_out_403[7:2], u_ca_out_402[13:8], u_ca_out_401[15:14]};
assign col_out_405 = {u_ca_out_405[1:0],u_ca_out_404[7:2], u_ca_out_403[13:8], u_ca_out_402[15:14]};
assign col_out_406 = {u_ca_out_406[1:0],u_ca_out_405[7:2], u_ca_out_404[13:8], u_ca_out_403[15:14]};
assign col_out_407 = {u_ca_out_407[1:0],u_ca_out_406[7:2], u_ca_out_405[13:8], u_ca_out_404[15:14]};
assign col_out_408 = {u_ca_out_408[1:0],u_ca_out_407[7:2], u_ca_out_406[13:8], u_ca_out_405[15:14]};
assign col_out_409 = {u_ca_out_409[1:0],u_ca_out_408[7:2], u_ca_out_407[13:8], u_ca_out_406[15:14]};
assign col_out_410 = {u_ca_out_410[1:0],u_ca_out_409[7:2], u_ca_out_408[13:8], u_ca_out_407[15:14]};
assign col_out_411 = {u_ca_out_411[1:0],u_ca_out_410[7:2], u_ca_out_409[13:8], u_ca_out_408[15:14]};
assign col_out_412 = {u_ca_out_412[1:0],u_ca_out_411[7:2], u_ca_out_410[13:8], u_ca_out_409[15:14]};
assign col_out_413 = {u_ca_out_413[1:0],u_ca_out_412[7:2], u_ca_out_411[13:8], u_ca_out_410[15:14]};
assign col_out_414 = {u_ca_out_414[1:0],u_ca_out_413[7:2], u_ca_out_412[13:8], u_ca_out_411[15:14]};
assign col_out_415 = {u_ca_out_415[1:0],u_ca_out_414[7:2], u_ca_out_413[13:8], u_ca_out_412[15:14]};
assign col_out_416 = {u_ca_out_416[1:0],u_ca_out_415[7:2], u_ca_out_414[13:8], u_ca_out_413[15:14]};
assign col_out_417 = {u_ca_out_417[1:0],u_ca_out_416[7:2], u_ca_out_415[13:8], u_ca_out_414[15:14]};
assign col_out_418 = {u_ca_out_418[1:0],u_ca_out_417[7:2], u_ca_out_416[13:8], u_ca_out_415[15:14]};
assign col_out_419 = {u_ca_out_419[1:0],u_ca_out_418[7:2], u_ca_out_417[13:8], u_ca_out_416[15:14]};
assign col_out_420 = {u_ca_out_420[1:0],u_ca_out_419[7:2], u_ca_out_418[13:8], u_ca_out_417[15:14]};
assign col_out_421 = {u_ca_out_421[1:0],u_ca_out_420[7:2], u_ca_out_419[13:8], u_ca_out_418[15:14]};
assign col_out_422 = {u_ca_out_422[1:0],u_ca_out_421[7:2], u_ca_out_420[13:8], u_ca_out_419[15:14]};
assign col_out_423 = {u_ca_out_423[1:0],u_ca_out_422[7:2], u_ca_out_421[13:8], u_ca_out_420[15:14]};
assign col_out_424 = {u_ca_out_424[1:0],u_ca_out_423[7:2], u_ca_out_422[13:8], u_ca_out_421[15:14]};
assign col_out_425 = {u_ca_out_425[1:0],u_ca_out_424[7:2], u_ca_out_423[13:8], u_ca_out_422[15:14]};
assign col_out_426 = {u_ca_out_426[1:0],u_ca_out_425[7:2], u_ca_out_424[13:8], u_ca_out_423[15:14]};
assign col_out_427 = {u_ca_out_427[1:0],u_ca_out_426[7:2], u_ca_out_425[13:8], u_ca_out_424[15:14]};
assign col_out_428 = {u_ca_out_428[1:0],u_ca_out_427[7:2], u_ca_out_426[13:8], u_ca_out_425[15:14]};
assign col_out_429 = {u_ca_out_429[1:0],u_ca_out_428[7:2], u_ca_out_427[13:8], u_ca_out_426[15:14]};
assign col_out_430 = {u_ca_out_430[1:0],u_ca_out_429[7:2], u_ca_out_428[13:8], u_ca_out_427[15:14]};
assign col_out_431 = {u_ca_out_431[1:0],u_ca_out_430[7:2], u_ca_out_429[13:8], u_ca_out_428[15:14]};
assign col_out_432 = {u_ca_out_432[1:0],u_ca_out_431[7:2], u_ca_out_430[13:8], u_ca_out_429[15:14]};
assign col_out_433 = {u_ca_out_433[1:0],u_ca_out_432[7:2], u_ca_out_431[13:8], u_ca_out_430[15:14]};
assign col_out_434 = {u_ca_out_434[1:0],u_ca_out_433[7:2], u_ca_out_432[13:8], u_ca_out_431[15:14]};
assign col_out_435 = {u_ca_out_435[1:0],u_ca_out_434[7:2], u_ca_out_433[13:8], u_ca_out_432[15:14]};
assign col_out_436 = {u_ca_out_436[1:0],u_ca_out_435[7:2], u_ca_out_434[13:8], u_ca_out_433[15:14]};
assign col_out_437 = {u_ca_out_437[1:0],u_ca_out_436[7:2], u_ca_out_435[13:8], u_ca_out_434[15:14]};
assign col_out_438 = {u_ca_out_438[1:0],u_ca_out_437[7:2], u_ca_out_436[13:8], u_ca_out_435[15:14]};
assign col_out_439 = {u_ca_out_439[1:0],u_ca_out_438[7:2], u_ca_out_437[13:8], u_ca_out_436[15:14]};
assign col_out_440 = {u_ca_out_440[1:0],u_ca_out_439[7:2], u_ca_out_438[13:8], u_ca_out_437[15:14]};
assign col_out_441 = {u_ca_out_441[1:0],u_ca_out_440[7:2], u_ca_out_439[13:8], u_ca_out_438[15:14]};
assign col_out_442 = {u_ca_out_442[1:0],u_ca_out_441[7:2], u_ca_out_440[13:8], u_ca_out_439[15:14]};
assign col_out_443 = {u_ca_out_443[1:0],u_ca_out_442[7:2], u_ca_out_441[13:8], u_ca_out_440[15:14]};
assign col_out_444 = {u_ca_out_444[1:0],u_ca_out_443[7:2], u_ca_out_442[13:8], u_ca_out_441[15:14]};
assign col_out_445 = {u_ca_out_445[1:0],u_ca_out_444[7:2], u_ca_out_443[13:8], u_ca_out_442[15:14]};
assign col_out_446 = {u_ca_out_446[1:0],u_ca_out_445[7:2], u_ca_out_444[13:8], u_ca_out_443[15:14]};
assign col_out_447 = {u_ca_out_447[1:0],u_ca_out_446[7:2], u_ca_out_445[13:8], u_ca_out_444[15:14]};
assign col_out_448 = {u_ca_out_448[1:0],u_ca_out_447[7:2], u_ca_out_446[13:8], u_ca_out_445[15:14]};
assign col_out_449 = {u_ca_out_449[1:0],u_ca_out_448[7:2], u_ca_out_447[13:8], u_ca_out_446[15:14]};
assign col_out_450 = {u_ca_out_450[1:0],u_ca_out_449[7:2], u_ca_out_448[13:8], u_ca_out_447[15:14]};
assign col_out_451 = {u_ca_out_451[1:0],u_ca_out_450[7:2], u_ca_out_449[13:8], u_ca_out_448[15:14]};
assign col_out_452 = {u_ca_out_452[1:0],u_ca_out_451[7:2], u_ca_out_450[13:8], u_ca_out_449[15:14]};
assign col_out_453 = {u_ca_out_453[1:0],u_ca_out_452[7:2], u_ca_out_451[13:8], u_ca_out_450[15:14]};
assign col_out_454 = {u_ca_out_454[1:0],u_ca_out_453[7:2], u_ca_out_452[13:8], u_ca_out_451[15:14]};
assign col_out_455 = {u_ca_out_455[1:0],u_ca_out_454[7:2], u_ca_out_453[13:8], u_ca_out_452[15:14]};
assign col_out_456 = {u_ca_out_456[1:0],u_ca_out_455[7:2], u_ca_out_454[13:8], u_ca_out_453[15:14]};
assign col_out_457 = {u_ca_out_457[1:0],u_ca_out_456[7:2], u_ca_out_455[13:8], u_ca_out_454[15:14]};
assign col_out_458 = {u_ca_out_458[1:0],u_ca_out_457[7:2], u_ca_out_456[13:8], u_ca_out_455[15:14]};
assign col_out_459 = {u_ca_out_459[1:0],u_ca_out_458[7:2], u_ca_out_457[13:8], u_ca_out_456[15:14]};
assign col_out_460 = {u_ca_out_460[1:0],u_ca_out_459[7:2], u_ca_out_458[13:8], u_ca_out_457[15:14]};
assign col_out_461 = {u_ca_out_461[1:0],u_ca_out_460[7:2], u_ca_out_459[13:8], u_ca_out_458[15:14]};
assign col_out_462 = {u_ca_out_462[1:0],u_ca_out_461[7:2], u_ca_out_460[13:8], u_ca_out_459[15:14]};
assign col_out_463 = {u_ca_out_463[1:0],u_ca_out_462[7:2], u_ca_out_461[13:8], u_ca_out_460[15:14]};
assign col_out_464 = {u_ca_out_464[1:0],u_ca_out_463[7:2], u_ca_out_462[13:8], u_ca_out_461[15:14]};
assign col_out_465 = {u_ca_out_465[1:0],u_ca_out_464[7:2], u_ca_out_463[13:8], u_ca_out_462[15:14]};
assign col_out_466 = {u_ca_out_466[1:0],u_ca_out_465[7:2], u_ca_out_464[13:8], u_ca_out_463[15:14]};
assign col_out_467 = {u_ca_out_467[1:0],u_ca_out_466[7:2], u_ca_out_465[13:8], u_ca_out_464[15:14]};
assign col_out_468 = {u_ca_out_468[1:0],u_ca_out_467[7:2], u_ca_out_466[13:8], u_ca_out_465[15:14]};
assign col_out_469 = {u_ca_out_469[1:0],u_ca_out_468[7:2], u_ca_out_467[13:8], u_ca_out_466[15:14]};
assign col_out_470 = {u_ca_out_470[1:0],u_ca_out_469[7:2], u_ca_out_468[13:8], u_ca_out_467[15:14]};
assign col_out_471 = {u_ca_out_471[1:0],u_ca_out_470[7:2], u_ca_out_469[13:8], u_ca_out_468[15:14]};
assign col_out_472 = {u_ca_out_472[1:0],u_ca_out_471[7:2], u_ca_out_470[13:8], u_ca_out_469[15:14]};
assign col_out_473 = {u_ca_out_473[1:0],u_ca_out_472[7:2], u_ca_out_471[13:8], u_ca_out_470[15:14]};
assign col_out_474 = {u_ca_out_474[1:0],u_ca_out_473[7:2], u_ca_out_472[13:8], u_ca_out_471[15:14]};
assign col_out_475 = {u_ca_out_475[1:0],u_ca_out_474[7:2], u_ca_out_473[13:8], u_ca_out_472[15:14]};
assign col_out_476 = {u_ca_out_476[1:0],u_ca_out_475[7:2], u_ca_out_474[13:8], u_ca_out_473[15:14]};
assign col_out_477 = {u_ca_out_477[1:0],u_ca_out_476[7:2], u_ca_out_475[13:8], u_ca_out_474[15:14]};
assign col_out_478 = {u_ca_out_478[1:0],u_ca_out_477[7:2], u_ca_out_476[13:8], u_ca_out_475[15:14]};
assign col_out_479 = {u_ca_out_479[1:0],u_ca_out_478[7:2], u_ca_out_477[13:8], u_ca_out_476[15:14]};
assign col_out_480 = {u_ca_out_480[1:0],u_ca_out_479[7:2], u_ca_out_478[13:8], u_ca_out_477[15:14]};
assign col_out_481 = {u_ca_out_481[1:0],u_ca_out_480[7:2], u_ca_out_479[13:8], u_ca_out_478[15:14]};
assign col_out_482 = {u_ca_out_482[1:0],u_ca_out_481[7:2], u_ca_out_480[13:8], u_ca_out_479[15:14]};
assign col_out_483 = {u_ca_out_483[1:0],u_ca_out_482[7:2], u_ca_out_481[13:8], u_ca_out_480[15:14]};
assign col_out_484 = {u_ca_out_484[1:0],u_ca_out_483[7:2], u_ca_out_482[13:8], u_ca_out_481[15:14]};
assign col_out_485 = {u_ca_out_485[1:0],u_ca_out_484[7:2], u_ca_out_483[13:8], u_ca_out_482[15:14]};
assign col_out_486 = {u_ca_out_486[1:0],u_ca_out_485[7:2], u_ca_out_484[13:8], u_ca_out_483[15:14]};
assign col_out_487 = {u_ca_out_487[1:0],u_ca_out_486[7:2], u_ca_out_485[13:8], u_ca_out_484[15:14]};
assign col_out_488 = {u_ca_out_488[1:0],u_ca_out_487[7:2], u_ca_out_486[13:8], u_ca_out_485[15:14]};
assign col_out_489 = {u_ca_out_489[1:0],u_ca_out_488[7:2], u_ca_out_487[13:8], u_ca_out_486[15:14]};
assign col_out_490 = {u_ca_out_490[1:0],u_ca_out_489[7:2], u_ca_out_488[13:8], u_ca_out_487[15:14]};
assign col_out_491 = {u_ca_out_491[1:0],u_ca_out_490[7:2], u_ca_out_489[13:8], u_ca_out_488[15:14]};
assign col_out_492 = {u_ca_out_492[1:0],u_ca_out_491[7:2], u_ca_out_490[13:8], u_ca_out_489[15:14]};
assign col_out_493 = {u_ca_out_493[1:0],u_ca_out_492[7:2], u_ca_out_491[13:8], u_ca_out_490[15:14]};
assign col_out_494 = {u_ca_out_494[1:0],u_ca_out_493[7:2], u_ca_out_492[13:8], u_ca_out_491[15:14]};
assign col_out_495 = {u_ca_out_495[1:0],u_ca_out_494[7:2], u_ca_out_493[13:8], u_ca_out_492[15:14]};
assign col_out_496 = {u_ca_out_496[1:0],u_ca_out_495[7:2], u_ca_out_494[13:8], u_ca_out_493[15:14]};
assign col_out_497 = {u_ca_out_497[1:0],u_ca_out_496[7:2], u_ca_out_495[13:8], u_ca_out_494[15:14]};
assign col_out_498 = {u_ca_out_498[1:0],u_ca_out_497[7:2], u_ca_out_496[13:8], u_ca_out_495[15:14]};
assign col_out_499 = {u_ca_out_499[1:0],u_ca_out_498[7:2], u_ca_out_497[13:8], u_ca_out_496[15:14]};
assign col_out_500 = {u_ca_out_500[1:0],u_ca_out_499[7:2], u_ca_out_498[13:8], u_ca_out_497[15:14]};
assign col_out_501 = {u_ca_out_501[1:0],u_ca_out_500[7:2], u_ca_out_499[13:8], u_ca_out_498[15:14]};
assign col_out_502 = {u_ca_out_502[1:0],u_ca_out_501[7:2], u_ca_out_500[13:8], u_ca_out_499[15:14]};
assign col_out_503 = {u_ca_out_503[1:0],u_ca_out_502[7:2], u_ca_out_501[13:8], u_ca_out_500[15:14]};
assign col_out_504 = {u_ca_out_504[1:0],u_ca_out_503[7:2], u_ca_out_502[13:8], u_ca_out_501[15:14]};
assign col_out_505 = {u_ca_out_505[1:0],u_ca_out_504[7:2], u_ca_out_503[13:8], u_ca_out_502[15:14]};
assign col_out_506 = {u_ca_out_506[1:0],u_ca_out_505[7:2], u_ca_out_504[13:8], u_ca_out_503[15:14]};
assign col_out_507 = {u_ca_out_507[1:0],u_ca_out_506[7:2], u_ca_out_505[13:8], u_ca_out_504[15:14]};
assign col_out_508 = {u_ca_out_508[1:0],u_ca_out_507[7:2], u_ca_out_506[13:8], u_ca_out_505[15:14]};
assign col_out_509 = {u_ca_out_509[1:0],u_ca_out_508[7:2], u_ca_out_507[13:8], u_ca_out_506[15:14]};
assign col_out_510 = {u_ca_out_510[1:0],u_ca_out_509[7:2], u_ca_out_508[13:8], u_ca_out_507[15:14]};
assign col_out_511 = {u_ca_out_511[1:0],u_ca_out_510[7:2], u_ca_out_509[13:8], u_ca_out_508[15:14]};
assign col_out_512 = {u_ca_out_512[1:0],u_ca_out_511[7:2], u_ca_out_510[13:8], u_ca_out_509[15:14]};
assign col_out_513 = {u_ca_out_513[1:0],u_ca_out_512[7:2], u_ca_out_511[13:8], u_ca_out_510[15:14]};
assign col_out_514 = {u_ca_out_514[1:0],u_ca_out_513[7:2], u_ca_out_512[13:8], u_ca_out_511[15:14]};
assign col_out_515 = {u_ca_out_515[1:0],u_ca_out_514[7:2], u_ca_out_513[13:8], u_ca_out_512[15:14]};
assign col_out_516 = {u_ca_out_516[1:0],u_ca_out_515[7:2], u_ca_out_514[13:8], u_ca_out_513[15:14]};
assign col_out_517 = {u_ca_out_517[1:0],u_ca_out_516[7:2], u_ca_out_515[13:8], u_ca_out_514[15:14]};
assign col_out_518 = {u_ca_out_518[1:0],u_ca_out_517[7:2], u_ca_out_516[13:8], u_ca_out_515[15:14]};
assign col_out_519 = {u_ca_out_519[1:0],u_ca_out_518[7:2], u_ca_out_517[13:8], u_ca_out_516[15:14]};
assign col_out_520 = {u_ca_out_520[1:0],u_ca_out_519[7:2], u_ca_out_518[13:8], u_ca_out_517[15:14]};
assign col_out_521 = {u_ca_out_521[1:0],u_ca_out_520[7:2], u_ca_out_519[13:8], u_ca_out_518[15:14]};
assign col_out_522 = {u_ca_out_522[1:0],u_ca_out_521[7:2], u_ca_out_520[13:8], u_ca_out_519[15:14]};
assign col_out_523 = {u_ca_out_523[1:0],u_ca_out_522[7:2], u_ca_out_521[13:8], u_ca_out_520[15:14]};
assign col_out_524 = {u_ca_out_524[1:0],u_ca_out_523[7:2], u_ca_out_522[13:8], u_ca_out_521[15:14]};
assign col_out_525 = {u_ca_out_525[1:0],u_ca_out_524[7:2], u_ca_out_523[13:8], u_ca_out_522[15:14]};
assign col_out_526 = {u_ca_out_526[1:0],u_ca_out_525[7:2], u_ca_out_524[13:8], u_ca_out_523[15:14]};
assign col_out_527 = {u_ca_out_527[1:0],u_ca_out_526[7:2], u_ca_out_525[13:8], u_ca_out_524[15:14]};
assign col_out_528 = {u_ca_out_528[1:0],u_ca_out_527[7:2], u_ca_out_526[13:8], u_ca_out_525[15:14]};
assign col_out_529 = {u_ca_out_529[1:0],u_ca_out_528[7:2], u_ca_out_527[13:8], u_ca_out_526[15:14]};
assign col_out_530 = {u_ca_out_530[1:0],u_ca_out_529[7:2], u_ca_out_528[13:8], u_ca_out_527[15:14]};
assign col_out_531 = {u_ca_out_531[1:0],u_ca_out_530[7:2], u_ca_out_529[13:8], u_ca_out_528[15:14]};
assign col_out_532 = {u_ca_out_532[1:0],u_ca_out_531[7:2], u_ca_out_530[13:8], u_ca_out_529[15:14]};
assign col_out_533 = {u_ca_out_533[1:0],u_ca_out_532[7:2], u_ca_out_531[13:8], u_ca_out_530[15:14]};
assign col_out_534 = {u_ca_out_534[1:0],u_ca_out_533[7:2], u_ca_out_532[13:8], u_ca_out_531[15:14]};
assign col_out_535 = {u_ca_out_535[1:0],u_ca_out_534[7:2], u_ca_out_533[13:8], u_ca_out_532[15:14]};
assign col_out_536 = {u_ca_out_536[1:0],u_ca_out_535[7:2], u_ca_out_534[13:8], u_ca_out_533[15:14]};
assign col_out_537 = {u_ca_out_537[1:0],u_ca_out_536[7:2], u_ca_out_535[13:8], u_ca_out_534[15:14]};
assign col_out_538 = {u_ca_out_538[1:0],u_ca_out_537[7:2], u_ca_out_536[13:8], u_ca_out_535[15:14]};
assign col_out_539 = {u_ca_out_539[1:0],u_ca_out_538[7:2], u_ca_out_537[13:8], u_ca_out_536[15:14]};
assign col_out_540 = {u_ca_out_540[1:0],u_ca_out_539[7:2], u_ca_out_538[13:8], u_ca_out_537[15:14]};
assign col_out_541 = {u_ca_out_541[1:0],u_ca_out_540[7:2], u_ca_out_539[13:8], u_ca_out_538[15:14]};
assign col_out_542 = {u_ca_out_542[1:0],u_ca_out_541[7:2], u_ca_out_540[13:8], u_ca_out_539[15:14]};
assign col_out_543 = {u_ca_out_543[1:0],u_ca_out_542[7:2], u_ca_out_541[13:8], u_ca_out_540[15:14]};
assign col_out_544 = {u_ca_out_544[1:0],u_ca_out_543[7:2], u_ca_out_542[13:8], u_ca_out_541[15:14]};
assign col_out_545 = {u_ca_out_545[1:0],u_ca_out_544[7:2], u_ca_out_543[13:8], u_ca_out_542[15:14]};
assign col_out_546 = {u_ca_out_546[1:0],u_ca_out_545[7:2], u_ca_out_544[13:8], u_ca_out_543[15:14]};
assign col_out_547 = {u_ca_out_547[1:0],u_ca_out_546[7:2], u_ca_out_545[13:8], u_ca_out_544[15:14]};
assign col_out_548 = {u_ca_out_548[1:0],u_ca_out_547[7:2], u_ca_out_546[13:8], u_ca_out_545[15:14]};
assign col_out_549 = {u_ca_out_549[1:0],u_ca_out_548[7:2], u_ca_out_547[13:8], u_ca_out_546[15:14]};
assign col_out_550 = {u_ca_out_550[1:0],u_ca_out_549[7:2], u_ca_out_548[13:8], u_ca_out_547[15:14]};
assign col_out_551 = {u_ca_out_551[1:0],u_ca_out_550[7:2], u_ca_out_549[13:8], u_ca_out_548[15:14]};
assign col_out_552 = {u_ca_out_552[1:0],u_ca_out_551[7:2], u_ca_out_550[13:8], u_ca_out_549[15:14]};
assign col_out_553 = {u_ca_out_553[1:0],u_ca_out_552[7:2], u_ca_out_551[13:8], u_ca_out_550[15:14]};
assign col_out_554 = {u_ca_out_554[1:0],u_ca_out_553[7:2], u_ca_out_552[13:8], u_ca_out_551[15:14]};
assign col_out_555 = {u_ca_out_555[1:0],u_ca_out_554[7:2], u_ca_out_553[13:8], u_ca_out_552[15:14]};
assign col_out_556 = {u_ca_out_556[1:0],u_ca_out_555[7:2], u_ca_out_554[13:8], u_ca_out_553[15:14]};
assign col_out_557 = {u_ca_out_557[1:0],u_ca_out_556[7:2], u_ca_out_555[13:8], u_ca_out_554[15:14]};
assign col_out_558 = {u_ca_out_558[1:0],u_ca_out_557[7:2], u_ca_out_556[13:8], u_ca_out_555[15:14]};
assign col_out_559 = {u_ca_out_559[1:0],u_ca_out_558[7:2], u_ca_out_557[13:8], u_ca_out_556[15:14]};
assign col_out_560 = {u_ca_out_560[1:0],u_ca_out_559[7:2], u_ca_out_558[13:8], u_ca_out_557[15:14]};
assign col_out_561 = {u_ca_out_561[1:0],u_ca_out_560[7:2], u_ca_out_559[13:8], u_ca_out_558[15:14]};
assign col_out_562 = {u_ca_out_562[1:0],u_ca_out_561[7:2], u_ca_out_560[13:8], u_ca_out_559[15:14]};
assign col_out_563 = {u_ca_out_563[1:0],u_ca_out_562[7:2], u_ca_out_561[13:8], u_ca_out_560[15:14]};
assign col_out_564 = {u_ca_out_564[1:0],u_ca_out_563[7:2], u_ca_out_562[13:8], u_ca_out_561[15:14]};
assign col_out_565 = {u_ca_out_565[1:0],u_ca_out_564[7:2], u_ca_out_563[13:8], u_ca_out_562[15:14]};
assign col_out_566 = {u_ca_out_566[1:0],u_ca_out_565[7:2], u_ca_out_564[13:8], u_ca_out_563[15:14]};
assign col_out_567 = {u_ca_out_567[1:0],u_ca_out_566[7:2], u_ca_out_565[13:8], u_ca_out_564[15:14]};
assign col_out_568 = {u_ca_out_568[1:0],u_ca_out_567[7:2], u_ca_out_566[13:8], u_ca_out_565[15:14]};
assign col_out_569 = {u_ca_out_569[1:0],u_ca_out_568[7:2], u_ca_out_567[13:8], u_ca_out_566[15:14]};
assign col_out_570 = {u_ca_out_570[1:0],u_ca_out_569[7:2], u_ca_out_568[13:8], u_ca_out_567[15:14]};
assign col_out_571 = {u_ca_out_571[1:0],u_ca_out_570[7:2], u_ca_out_569[13:8], u_ca_out_568[15:14]};
assign col_out_572 = {u_ca_out_572[1:0],u_ca_out_571[7:2], u_ca_out_570[13:8], u_ca_out_569[15:14]};
assign col_out_573 = {u_ca_out_573[1:0],u_ca_out_572[7:2], u_ca_out_571[13:8], u_ca_out_570[15:14]};
assign col_out_574 = {u_ca_out_574[1:0],u_ca_out_573[7:2], u_ca_out_572[13:8], u_ca_out_571[15:14]};
assign col_out_575 = {u_ca_out_575[1:0],u_ca_out_574[7:2], u_ca_out_573[13:8], u_ca_out_572[15:14]};
assign col_out_576 = {u_ca_out_576[1:0],u_ca_out_575[7:2], u_ca_out_574[13:8], u_ca_out_573[15:14]};
assign col_out_577 = {u_ca_out_577[1:0],u_ca_out_576[7:2], u_ca_out_575[13:8], u_ca_out_574[15:14]};
assign col_out_578 = {u_ca_out_578[1:0],u_ca_out_577[7:2], u_ca_out_576[13:8], u_ca_out_575[15:14]};
assign col_out_579 = {u_ca_out_579[1:0],u_ca_out_578[7:2], u_ca_out_577[13:8], u_ca_out_576[15:14]};
assign col_out_580 = {u_ca_out_580[1:0],u_ca_out_579[7:2], u_ca_out_578[13:8], u_ca_out_577[15:14]};
assign col_out_581 = {u_ca_out_581[1:0],u_ca_out_580[7:2], u_ca_out_579[13:8], u_ca_out_578[15:14]};
assign col_out_582 = {u_ca_out_582[1:0],u_ca_out_581[7:2], u_ca_out_580[13:8], u_ca_out_579[15:14]};
assign col_out_583 = {u_ca_out_583[1:0],u_ca_out_582[7:2], u_ca_out_581[13:8], u_ca_out_580[15:14]};
assign col_out_584 = {u_ca_out_584[1:0],u_ca_out_583[7:2], u_ca_out_582[13:8], u_ca_out_581[15:14]};
assign col_out_585 = {u_ca_out_585[1:0],u_ca_out_584[7:2], u_ca_out_583[13:8], u_ca_out_582[15:14]};
assign col_out_586 = {u_ca_out_586[1:0],u_ca_out_585[7:2], u_ca_out_584[13:8], u_ca_out_583[15:14]};
assign col_out_587 = {u_ca_out_587[1:0],u_ca_out_586[7:2], u_ca_out_585[13:8], u_ca_out_584[15:14]};
assign col_out_588 = {u_ca_out_588[1:0],u_ca_out_587[7:2], u_ca_out_586[13:8], u_ca_out_585[15:14]};
assign col_out_589 = {u_ca_out_589[1:0],u_ca_out_588[7:2], u_ca_out_587[13:8], u_ca_out_586[15:14]};
assign col_out_590 = {u_ca_out_590[1:0],u_ca_out_589[7:2], u_ca_out_588[13:8], u_ca_out_587[15:14]};
assign col_out_591 = {u_ca_out_591[1:0],u_ca_out_590[7:2], u_ca_out_589[13:8], u_ca_out_588[15:14]};
assign col_out_592 = {u_ca_out_592[1:0],u_ca_out_591[7:2], u_ca_out_590[13:8], u_ca_out_589[15:14]};
assign col_out_593 = {u_ca_out_593[1:0],u_ca_out_592[7:2], u_ca_out_591[13:8], u_ca_out_590[15:14]};
assign col_out_594 = {u_ca_out_594[1:0],u_ca_out_593[7:2], u_ca_out_592[13:8], u_ca_out_591[15:14]};
assign col_out_595 = {u_ca_out_595[1:0],u_ca_out_594[7:2], u_ca_out_593[13:8], u_ca_out_592[15:14]};
assign col_out_596 = {u_ca_out_596[1:0],u_ca_out_595[7:2], u_ca_out_594[13:8], u_ca_out_593[15:14]};
assign col_out_597 = {u_ca_out_597[1:0],u_ca_out_596[7:2], u_ca_out_595[13:8], u_ca_out_594[15:14]};
assign col_out_598 = {u_ca_out_598[1:0],u_ca_out_597[7:2], u_ca_out_596[13:8], u_ca_out_595[15:14]};
assign col_out_599 = {u_ca_out_599[1:0],u_ca_out_598[7:2], u_ca_out_597[13:8], u_ca_out_596[15:14]};
assign col_out_600 = {u_ca_out_600[1:0],u_ca_out_599[7:2], u_ca_out_598[13:8], u_ca_out_597[15:14]};
assign col_out_601 = {u_ca_out_601[1:0],u_ca_out_600[7:2], u_ca_out_599[13:8], u_ca_out_598[15:14]};
assign col_out_602 = {u_ca_out_602[1:0],u_ca_out_601[7:2], u_ca_out_600[13:8], u_ca_out_599[15:14]};
assign col_out_603 = {u_ca_out_603[1:0],u_ca_out_602[7:2], u_ca_out_601[13:8], u_ca_out_600[15:14]};
assign col_out_604 = {u_ca_out_604[1:0],u_ca_out_603[7:2], u_ca_out_602[13:8], u_ca_out_601[15:14]};
assign col_out_605 = {u_ca_out_605[1:0],u_ca_out_604[7:2], u_ca_out_603[13:8], u_ca_out_602[15:14]};
assign col_out_606 = {u_ca_out_606[1:0],u_ca_out_605[7:2], u_ca_out_604[13:8], u_ca_out_603[15:14]};
assign col_out_607 = {u_ca_out_607[1:0],u_ca_out_606[7:2], u_ca_out_605[13:8], u_ca_out_604[15:14]};
assign col_out_608 = {u_ca_out_608[1:0],u_ca_out_607[7:2], u_ca_out_606[13:8], u_ca_out_605[15:14]};
assign col_out_609 = {u_ca_out_609[1:0],u_ca_out_608[7:2], u_ca_out_607[13:8], u_ca_out_606[15:14]};
assign col_out_610 = {u_ca_out_610[1:0],u_ca_out_609[7:2], u_ca_out_608[13:8], u_ca_out_607[15:14]};
assign col_out_611 = {u_ca_out_611[1:0],u_ca_out_610[7:2], u_ca_out_609[13:8], u_ca_out_608[15:14]};
assign col_out_612 = {u_ca_out_612[1:0],u_ca_out_611[7:2], u_ca_out_610[13:8], u_ca_out_609[15:14]};
assign col_out_613 = {u_ca_out_613[1:0],u_ca_out_612[7:2], u_ca_out_611[13:8], u_ca_out_610[15:14]};
assign col_out_614 = {u_ca_out_614[1:0],u_ca_out_613[7:2], u_ca_out_612[13:8], u_ca_out_611[15:14]};
assign col_out_615 = {u_ca_out_615[1:0],u_ca_out_614[7:2], u_ca_out_613[13:8], u_ca_out_612[15:14]};
assign col_out_616 = {u_ca_out_616[1:0],u_ca_out_615[7:2], u_ca_out_614[13:8], u_ca_out_613[15:14]};
assign col_out_617 = {u_ca_out_617[1:0],u_ca_out_616[7:2], u_ca_out_615[13:8], u_ca_out_614[15:14]};
assign col_out_618 = {u_ca_out_618[1:0],u_ca_out_617[7:2], u_ca_out_616[13:8], u_ca_out_615[15:14]};
assign col_out_619 = {u_ca_out_619[1:0],u_ca_out_618[7:2], u_ca_out_617[13:8], u_ca_out_616[15:14]};
assign col_out_620 = {u_ca_out_620[1:0],u_ca_out_619[7:2], u_ca_out_618[13:8], u_ca_out_617[15:14]};
assign col_out_621 = {u_ca_out_621[1:0],u_ca_out_620[7:2], u_ca_out_619[13:8], u_ca_out_618[15:14]};
assign col_out_622 = {u_ca_out_622[1:0],u_ca_out_621[7:2], u_ca_out_620[13:8], u_ca_out_619[15:14]};
assign col_out_623 = {u_ca_out_623[1:0],u_ca_out_622[7:2], u_ca_out_621[13:8], u_ca_out_620[15:14]};
assign col_out_624 = {u_ca_out_624[1:0],u_ca_out_623[7:2], u_ca_out_622[13:8], u_ca_out_621[15:14]};
assign col_out_625 = {u_ca_out_625[1:0],u_ca_out_624[7:2], u_ca_out_623[13:8], u_ca_out_622[15:14]};
assign col_out_626 = {u_ca_out_626[1:0],u_ca_out_625[7:2], u_ca_out_624[13:8], u_ca_out_623[15:14]};
assign col_out_627 = {u_ca_out_627[1:0],u_ca_out_626[7:2], u_ca_out_625[13:8], u_ca_out_624[15:14]};
assign col_out_628 = {u_ca_out_628[1:0],u_ca_out_627[7:2], u_ca_out_626[13:8], u_ca_out_625[15:14]};
assign col_out_629 = {u_ca_out_629[1:0],u_ca_out_628[7:2], u_ca_out_627[13:8], u_ca_out_626[15:14]};
assign col_out_630 = {u_ca_out_630[1:0],u_ca_out_629[7:2], u_ca_out_628[13:8], u_ca_out_627[15:14]};
assign col_out_631 = {u_ca_out_631[1:0],u_ca_out_630[7:2], u_ca_out_629[13:8], u_ca_out_628[15:14]};
assign col_out_632 = {u_ca_out_632[1:0],u_ca_out_631[7:2], u_ca_out_630[13:8], u_ca_out_629[15:14]};
assign col_out_633 = {u_ca_out_633[1:0],u_ca_out_632[7:2], u_ca_out_631[13:8], u_ca_out_630[15:14]};
assign col_out_634 = {u_ca_out_634[1:0],u_ca_out_633[7:2], u_ca_out_632[13:8], u_ca_out_631[15:14]};
assign col_out_635 = {u_ca_out_635[1:0],u_ca_out_634[7:2], u_ca_out_633[13:8], u_ca_out_632[15:14]};
assign col_out_636 = {u_ca_out_636[1:0],u_ca_out_635[7:2], u_ca_out_634[13:8], u_ca_out_633[15:14]};
assign col_out_637 = {u_ca_out_637[1:0],u_ca_out_636[7:2], u_ca_out_635[13:8], u_ca_out_634[15:14]};
assign col_out_638 = {u_ca_out_638[1:0],u_ca_out_637[7:2], u_ca_out_636[13:8], u_ca_out_635[15:14]};
assign col_out_639 = {u_ca_out_639[1:0],u_ca_out_638[7:2], u_ca_out_637[13:8], u_ca_out_636[15:14]};
assign col_out_640 = {u_ca_out_640[1:0],u_ca_out_639[7:2], u_ca_out_638[13:8], u_ca_out_637[15:14]};
assign col_out_641 = {u_ca_out_641[1:0],u_ca_out_640[7:2], u_ca_out_639[13:8], u_ca_out_638[15:14]};
assign col_out_642 = {u_ca_out_642[1:0],u_ca_out_641[7:2], u_ca_out_640[13:8], u_ca_out_639[15:14]};
assign col_out_643 = {u_ca_out_643[1:0],u_ca_out_642[7:2], u_ca_out_641[13:8], u_ca_out_640[15:14]};
assign col_out_644 = {u_ca_out_644[1:0],u_ca_out_643[7:2], u_ca_out_642[13:8], u_ca_out_641[15:14]};
assign col_out_645 = {u_ca_out_645[1:0],u_ca_out_644[7:2], u_ca_out_643[13:8], u_ca_out_642[15:14]};
assign col_out_646 = {u_ca_out_646[1:0],u_ca_out_645[7:2], u_ca_out_644[13:8], u_ca_out_643[15:14]};
assign col_out_647 = {u_ca_out_647[1:0],u_ca_out_646[7:2], u_ca_out_645[13:8], u_ca_out_644[15:14]};
assign col_out_648 = {u_ca_out_648[1:0],u_ca_out_647[7:2], u_ca_out_646[13:8], u_ca_out_645[15:14]};
assign col_out_649 = {u_ca_out_649[1:0],u_ca_out_648[7:2], u_ca_out_647[13:8], u_ca_out_646[15:14]};
assign col_out_650 = {u_ca_out_650[1:0],u_ca_out_649[7:2], u_ca_out_648[13:8], u_ca_out_647[15:14]};
assign col_out_651 = {u_ca_out_651[1:0],u_ca_out_650[7:2], u_ca_out_649[13:8], u_ca_out_648[15:14]};
assign col_out_652 = {u_ca_out_652[1:0],u_ca_out_651[7:2], u_ca_out_650[13:8], u_ca_out_649[15:14]};
assign col_out_653 = {u_ca_out_653[1:0],u_ca_out_652[7:2], u_ca_out_651[13:8], u_ca_out_650[15:14]};
assign col_out_654 = {u_ca_out_654[1:0],u_ca_out_653[7:2], u_ca_out_652[13:8], u_ca_out_651[15:14]};
assign col_out_655 = {u_ca_out_655[1:0],u_ca_out_654[7:2], u_ca_out_653[13:8], u_ca_out_652[15:14]};
assign col_out_656 = {u_ca_out_656[1:0],u_ca_out_655[7:2], u_ca_out_654[13:8], u_ca_out_653[15:14]};
assign col_out_657 = {u_ca_out_657[1:0],u_ca_out_656[7:2], u_ca_out_655[13:8], u_ca_out_654[15:14]};
assign col_out_658 = {u_ca_out_658[1:0],u_ca_out_657[7:2], u_ca_out_656[13:8], u_ca_out_655[15:14]};
assign col_out_659 = {u_ca_out_659[1:0],u_ca_out_658[7:2], u_ca_out_657[13:8], u_ca_out_656[15:14]};
assign col_out_660 = {u_ca_out_660[1:0],u_ca_out_659[7:2], u_ca_out_658[13:8], u_ca_out_657[15:14]};
assign col_out_661 = {u_ca_out_661[1:0],u_ca_out_660[7:2], u_ca_out_659[13:8], u_ca_out_658[15:14]};
assign col_out_662 = {u_ca_out_662[1:0],u_ca_out_661[7:2], u_ca_out_660[13:8], u_ca_out_659[15:14]};
assign col_out_663 = {u_ca_out_663[1:0],u_ca_out_662[7:2], u_ca_out_661[13:8], u_ca_out_660[15:14]};
assign col_out_664 = {u_ca_out_664[1:0],u_ca_out_663[7:2], u_ca_out_662[13:8], u_ca_out_661[15:14]};
assign col_out_665 = {u_ca_out_665[1:0],u_ca_out_664[7:2], u_ca_out_663[13:8], u_ca_out_662[15:14]};
assign col_out_666 = {u_ca_out_666[1:0],u_ca_out_665[7:2], u_ca_out_664[13:8], u_ca_out_663[15:14]};
assign col_out_667 = {u_ca_out_667[1:0],u_ca_out_666[7:2], u_ca_out_665[13:8], u_ca_out_664[15:14]};
assign col_out_668 = {u_ca_out_668[1:0],u_ca_out_667[7:2], u_ca_out_666[13:8], u_ca_out_665[15:14]};
assign col_out_669 = {u_ca_out_669[1:0],u_ca_out_668[7:2], u_ca_out_667[13:8], u_ca_out_666[15:14]};
assign col_out_670 = {u_ca_out_670[1:0],u_ca_out_669[7:2], u_ca_out_668[13:8], u_ca_out_667[15:14]};
assign col_out_671 = {u_ca_out_671[1:0],u_ca_out_670[7:2], u_ca_out_669[13:8], u_ca_out_668[15:14]};
assign col_out_672 = {u_ca_out_672[1:0],u_ca_out_671[7:2], u_ca_out_670[13:8], u_ca_out_669[15:14]};
assign col_out_673 = {u_ca_out_673[1:0],u_ca_out_672[7:2], u_ca_out_671[13:8], u_ca_out_670[15:14]};
assign col_out_674 = {u_ca_out_674[1:0],u_ca_out_673[7:2], u_ca_out_672[13:8], u_ca_out_671[15:14]};
assign col_out_675 = {u_ca_out_675[1:0],u_ca_out_674[7:2], u_ca_out_673[13:8], u_ca_out_672[15:14]};
assign col_out_676 = {u_ca_out_676[1:0],u_ca_out_675[7:2], u_ca_out_674[13:8], u_ca_out_673[15:14]};
assign col_out_677 = {u_ca_out_677[1:0],u_ca_out_676[7:2], u_ca_out_675[13:8], u_ca_out_674[15:14]};
assign col_out_678 = {u_ca_out_678[1:0],u_ca_out_677[7:2], u_ca_out_676[13:8], u_ca_out_675[15:14]};
assign col_out_679 = {u_ca_out_679[1:0],u_ca_out_678[7:2], u_ca_out_677[13:8], u_ca_out_676[15:14]};
assign col_out_680 = {u_ca_out_680[1:0],u_ca_out_679[7:2], u_ca_out_678[13:8], u_ca_out_677[15:14]};
assign col_out_681 = {u_ca_out_681[1:0],u_ca_out_680[7:2], u_ca_out_679[13:8], u_ca_out_678[15:14]};
assign col_out_682 = {u_ca_out_682[1:0],u_ca_out_681[7:2], u_ca_out_680[13:8], u_ca_out_679[15:14]};
assign col_out_683 = {u_ca_out_683[1:0],u_ca_out_682[7:2], u_ca_out_681[13:8], u_ca_out_680[15:14]};
assign col_out_684 = {u_ca_out_684[1:0],u_ca_out_683[7:2], u_ca_out_682[13:8], u_ca_out_681[15:14]};
assign col_out_685 = {u_ca_out_685[1:0],u_ca_out_684[7:2], u_ca_out_683[13:8], u_ca_out_682[15:14]};
assign col_out_686 = {u_ca_out_686[1:0],u_ca_out_685[7:2], u_ca_out_684[13:8], u_ca_out_683[15:14]};
assign col_out_687 = {u_ca_out_687[1:0],u_ca_out_686[7:2], u_ca_out_685[13:8], u_ca_out_684[15:14]};
assign col_out_688 = {u_ca_out_688[1:0],u_ca_out_687[7:2], u_ca_out_686[13:8], u_ca_out_685[15:14]};
assign col_out_689 = {u_ca_out_689[1:0],u_ca_out_688[7:2], u_ca_out_687[13:8], u_ca_out_686[15:14]};
assign col_out_690 = {u_ca_out_690[1:0],u_ca_out_689[7:2], u_ca_out_688[13:8], u_ca_out_687[15:14]};
assign col_out_691 = {u_ca_out_691[1:0],u_ca_out_690[7:2], u_ca_out_689[13:8], u_ca_out_688[15:14]};
assign col_out_692 = {u_ca_out_692[1:0],u_ca_out_691[7:2], u_ca_out_690[13:8], u_ca_out_689[15:14]};
assign col_out_693 = {u_ca_out_693[1:0],u_ca_out_692[7:2], u_ca_out_691[13:8], u_ca_out_690[15:14]};
assign col_out_694 = {u_ca_out_694[1:0],u_ca_out_693[7:2], u_ca_out_692[13:8], u_ca_out_691[15:14]};
assign col_out_695 = {u_ca_out_695[1:0],u_ca_out_694[7:2], u_ca_out_693[13:8], u_ca_out_692[15:14]};
assign col_out_696 = {u_ca_out_696[1:0],u_ca_out_695[7:2], u_ca_out_694[13:8], u_ca_out_693[15:14]};
assign col_out_697 = {u_ca_out_697[1:0],u_ca_out_696[7:2], u_ca_out_695[13:8], u_ca_out_694[15:14]};
assign col_out_698 = {u_ca_out_698[1:0],u_ca_out_697[7:2], u_ca_out_696[13:8], u_ca_out_695[15:14]};
assign col_out_699 = {u_ca_out_699[1:0],u_ca_out_698[7:2], u_ca_out_697[13:8], u_ca_out_696[15:14]};
assign col_out_700 = {u_ca_out_700[1:0],u_ca_out_699[7:2], u_ca_out_698[13:8], u_ca_out_697[15:14]};
assign col_out_701 = {u_ca_out_701[1:0],u_ca_out_700[7:2], u_ca_out_699[13:8], u_ca_out_698[15:14]};
assign col_out_702 = {u_ca_out_702[1:0],u_ca_out_701[7:2], u_ca_out_700[13:8], u_ca_out_699[15:14]};
assign col_out_703 = {u_ca_out_703[1:0],u_ca_out_702[7:2], u_ca_out_701[13:8], u_ca_out_700[15:14]};
assign col_out_704 = {u_ca_out_704[1:0],u_ca_out_703[7:2], u_ca_out_702[13:8], u_ca_out_701[15:14]};
assign col_out_705 = {u_ca_out_705[1:0],u_ca_out_704[7:2], u_ca_out_703[13:8], u_ca_out_702[15:14]};
assign col_out_706 = {u_ca_out_706[1:0],u_ca_out_705[7:2], u_ca_out_704[13:8], u_ca_out_703[15:14]};
assign col_out_707 = {u_ca_out_707[1:0],u_ca_out_706[7:2], u_ca_out_705[13:8], u_ca_out_704[15:14]};
assign col_out_708 = {u_ca_out_708[1:0],u_ca_out_707[7:2], u_ca_out_706[13:8], u_ca_out_705[15:14]};
assign col_out_709 = {u_ca_out_709[1:0],u_ca_out_708[7:2], u_ca_out_707[13:8], u_ca_out_706[15:14]};
assign col_out_710 = {u_ca_out_710[1:0],u_ca_out_709[7:2], u_ca_out_708[13:8], u_ca_out_707[15:14]};
assign col_out_711 = {u_ca_out_711[1:0],u_ca_out_710[7:2], u_ca_out_709[13:8], u_ca_out_708[15:14]};
assign col_out_712 = {u_ca_out_712[1:0],u_ca_out_711[7:2], u_ca_out_710[13:8], u_ca_out_709[15:14]};
assign col_out_713 = {u_ca_out_713[1:0],u_ca_out_712[7:2], u_ca_out_711[13:8], u_ca_out_710[15:14]};
assign col_out_714 = {u_ca_out_714[1:0],u_ca_out_713[7:2], u_ca_out_712[13:8], u_ca_out_711[15:14]};
assign col_out_715 = {u_ca_out_715[1:0],u_ca_out_714[7:2], u_ca_out_713[13:8], u_ca_out_712[15:14]};
assign col_out_716 = {u_ca_out_716[1:0],u_ca_out_715[7:2], u_ca_out_714[13:8], u_ca_out_713[15:14]};
assign col_out_717 = {u_ca_out_717[1:0],u_ca_out_716[7:2], u_ca_out_715[13:8], u_ca_out_714[15:14]};
assign col_out_718 = {u_ca_out_718[1:0],u_ca_out_717[7:2], u_ca_out_716[13:8], u_ca_out_715[15:14]};
assign col_out_719 = {u_ca_out_719[1:0],u_ca_out_718[7:2], u_ca_out_717[13:8], u_ca_out_716[15:14]};
assign col_out_720 = {u_ca_out_720[1:0],u_ca_out_719[7:2], u_ca_out_718[13:8], u_ca_out_717[15:14]};
assign col_out_721 = {u_ca_out_721[1:0],u_ca_out_720[7:2], u_ca_out_719[13:8], u_ca_out_718[15:14]};
assign col_out_722 = {u_ca_out_722[1:0],u_ca_out_721[7:2], u_ca_out_720[13:8], u_ca_out_719[15:14]};
assign col_out_723 = {u_ca_out_723[1:0],u_ca_out_722[7:2], u_ca_out_721[13:8], u_ca_out_720[15:14]};
assign col_out_724 = {u_ca_out_724[1:0],u_ca_out_723[7:2], u_ca_out_722[13:8], u_ca_out_721[15:14]};
assign col_out_725 = {u_ca_out_725[1:0],u_ca_out_724[7:2], u_ca_out_723[13:8], u_ca_out_722[15:14]};
assign col_out_726 = {u_ca_out_726[1:0],u_ca_out_725[7:2], u_ca_out_724[13:8], u_ca_out_723[15:14]};
assign col_out_727 = {u_ca_out_727[1:0],u_ca_out_726[7:2], u_ca_out_725[13:8], u_ca_out_724[15:14]};
assign col_out_728 = {u_ca_out_728[1:0],u_ca_out_727[7:2], u_ca_out_726[13:8], u_ca_out_725[15:14]};
assign col_out_729 = {u_ca_out_729[1:0],u_ca_out_728[7:2], u_ca_out_727[13:8], u_ca_out_726[15:14]};
assign col_out_730 = {u_ca_out_730[1:0],u_ca_out_729[7:2], u_ca_out_728[13:8], u_ca_out_727[15:14]};
assign col_out_731 = {u_ca_out_731[1:0],u_ca_out_730[7:2], u_ca_out_729[13:8], u_ca_out_728[15:14]};
assign col_out_732 = {u_ca_out_732[1:0],u_ca_out_731[7:2], u_ca_out_730[13:8], u_ca_out_729[15:14]};
assign col_out_733 = {u_ca_out_733[1:0],u_ca_out_732[7:2], u_ca_out_731[13:8], u_ca_out_730[15:14]};
assign col_out_734 = {u_ca_out_734[1:0],u_ca_out_733[7:2], u_ca_out_732[13:8], u_ca_out_731[15:14]};
assign col_out_735 = {u_ca_out_735[1:0],u_ca_out_734[7:2], u_ca_out_733[13:8], u_ca_out_732[15:14]};
assign col_out_736 = {u_ca_out_736[1:0],u_ca_out_735[7:2], u_ca_out_734[13:8], u_ca_out_733[15:14]};
assign col_out_737 = {u_ca_out_737[1:0],u_ca_out_736[7:2], u_ca_out_735[13:8], u_ca_out_734[15:14]};
assign col_out_738 = {u_ca_out_738[1:0],u_ca_out_737[7:2], u_ca_out_736[13:8], u_ca_out_735[15:14]};
assign col_out_739 = {u_ca_out_739[1:0],u_ca_out_738[7:2], u_ca_out_737[13:8], u_ca_out_736[15:14]};
assign col_out_740 = {u_ca_out_740[1:0],u_ca_out_739[7:2], u_ca_out_738[13:8], u_ca_out_737[15:14]};
assign col_out_741 = {u_ca_out_741[1:0],u_ca_out_740[7:2], u_ca_out_739[13:8], u_ca_out_738[15:14]};
assign col_out_742 = {u_ca_out_742[1:0],u_ca_out_741[7:2], u_ca_out_740[13:8], u_ca_out_739[15:14]};
assign col_out_743 = {u_ca_out_743[1:0],u_ca_out_742[7:2], u_ca_out_741[13:8], u_ca_out_740[15:14]};
assign col_out_744 = {u_ca_out_744[1:0],u_ca_out_743[7:2], u_ca_out_742[13:8], u_ca_out_741[15:14]};
assign col_out_745 = {u_ca_out_745[1:0],u_ca_out_744[7:2], u_ca_out_743[13:8], u_ca_out_742[15:14]};
assign col_out_746 = {u_ca_out_746[1:0],u_ca_out_745[7:2], u_ca_out_744[13:8], u_ca_out_743[15:14]};
assign col_out_747 = {u_ca_out_747[1:0],u_ca_out_746[7:2], u_ca_out_745[13:8], u_ca_out_744[15:14]};
assign col_out_748 = {u_ca_out_748[1:0],u_ca_out_747[7:2], u_ca_out_746[13:8], u_ca_out_745[15:14]};
assign col_out_749 = {u_ca_out_749[1:0],u_ca_out_748[7:2], u_ca_out_747[13:8], u_ca_out_746[15:14]};
assign col_out_750 = {u_ca_out_750[1:0],u_ca_out_749[7:2], u_ca_out_748[13:8], u_ca_out_747[15:14]};
assign col_out_751 = {u_ca_out_751[1:0],u_ca_out_750[7:2], u_ca_out_749[13:8], u_ca_out_748[15:14]};
assign col_out_752 = {u_ca_out_752[1:0],u_ca_out_751[7:2], u_ca_out_750[13:8], u_ca_out_749[15:14]};
assign col_out_753 = {u_ca_out_753[1:0],u_ca_out_752[7:2], u_ca_out_751[13:8], u_ca_out_750[15:14]};
assign col_out_754 = {u_ca_out_754[1:0],u_ca_out_753[7:2], u_ca_out_752[13:8], u_ca_out_751[15:14]};
assign col_out_755 = {u_ca_out_755[1:0],u_ca_out_754[7:2], u_ca_out_753[13:8], u_ca_out_752[15:14]};
assign col_out_756 = {u_ca_out_756[1:0],u_ca_out_755[7:2], u_ca_out_754[13:8], u_ca_out_753[15:14]};
assign col_out_757 = {u_ca_out_757[1:0],u_ca_out_756[7:2], u_ca_out_755[13:8], u_ca_out_754[15:14]};
assign col_out_758 = {u_ca_out_758[1:0],u_ca_out_757[7:2], u_ca_out_756[13:8], u_ca_out_755[15:14]};
assign col_out_759 = {u_ca_out_759[1:0],u_ca_out_758[7:2], u_ca_out_757[13:8], u_ca_out_756[15:14]};
assign col_out_760 = {u_ca_out_760[1:0],u_ca_out_759[7:2], u_ca_out_758[13:8], u_ca_out_757[15:14]};
assign col_out_761 = {u_ca_out_761[1:0],u_ca_out_760[7:2], u_ca_out_759[13:8], u_ca_out_758[15:14]};
assign col_out_762 = {u_ca_out_762[1:0],u_ca_out_761[7:2], u_ca_out_760[13:8], u_ca_out_759[15:14]};
assign col_out_763 = {u_ca_out_763[1:0],u_ca_out_762[7:2], u_ca_out_761[13:8], u_ca_out_760[15:14]};
assign col_out_764 = {u_ca_out_764[1:0],u_ca_out_763[7:2], u_ca_out_762[13:8], u_ca_out_761[15:14]};
assign col_out_765 = {u_ca_out_765[1:0],u_ca_out_764[7:2], u_ca_out_763[13:8], u_ca_out_762[15:14]};
assign col_out_766 = {u_ca_out_766[1:0],u_ca_out_765[7:2], u_ca_out_764[13:8], u_ca_out_763[15:14]};
assign col_out_767 = {u_ca_out_767[1:0],u_ca_out_766[7:2], u_ca_out_765[13:8], u_ca_out_764[15:14]};
assign col_out_768 = {u_ca_out_768[1:0],u_ca_out_767[7:2], u_ca_out_766[13:8], u_ca_out_765[15:14]};
assign col_out_769 = {u_ca_out_769[1:0],u_ca_out_768[7:2], u_ca_out_767[13:8], u_ca_out_766[15:14]};
assign col_out_770 = {u_ca_out_770[1:0],u_ca_out_769[7:2], u_ca_out_768[13:8], u_ca_out_767[15:14]};
assign col_out_771 = {u_ca_out_771[1:0],u_ca_out_770[7:2], u_ca_out_769[13:8], u_ca_out_768[15:14]};
assign col_out_772 = {u_ca_out_772[1:0],u_ca_out_771[7:2], u_ca_out_770[13:8], u_ca_out_769[15:14]};
assign col_out_773 = {u_ca_out_773[1:0],u_ca_out_772[7:2], u_ca_out_771[13:8], u_ca_out_770[15:14]};
assign col_out_774 = {u_ca_out_774[1:0],u_ca_out_773[7:2], u_ca_out_772[13:8], u_ca_out_771[15:14]};
assign col_out_775 = {u_ca_out_775[1:0],u_ca_out_774[7:2], u_ca_out_773[13:8], u_ca_out_772[15:14]};
assign col_out_776 = {u_ca_out_776[1:0],u_ca_out_775[7:2], u_ca_out_774[13:8], u_ca_out_773[15:14]};
assign col_out_777 = {u_ca_out_777[1:0],u_ca_out_776[7:2], u_ca_out_775[13:8], u_ca_out_774[15:14]};
assign col_out_778 = {u_ca_out_778[1:0],u_ca_out_777[7:2], u_ca_out_776[13:8], u_ca_out_775[15:14]};
assign col_out_779 = {u_ca_out_779[1:0],u_ca_out_778[7:2], u_ca_out_777[13:8], u_ca_out_776[15:14]};
assign col_out_780 = {u_ca_out_780[1:0],u_ca_out_779[7:2], u_ca_out_778[13:8], u_ca_out_777[15:14]};
assign col_out_781 = {u_ca_out_781[1:0],u_ca_out_780[7:2], u_ca_out_779[13:8], u_ca_out_778[15:14]};
assign col_out_782 = {u_ca_out_782[1:0],u_ca_out_781[7:2], u_ca_out_780[13:8], u_ca_out_779[15:14]};
assign col_out_783 = {u_ca_out_783[1:0],u_ca_out_782[7:2], u_ca_out_781[13:8], u_ca_out_780[15:14]};
assign col_out_784 = {u_ca_out_784[1:0],u_ca_out_783[7:2], u_ca_out_782[13:8], u_ca_out_781[15:14]};
assign col_out_785 = {u_ca_out_785[1:0],u_ca_out_784[7:2], u_ca_out_783[13:8], u_ca_out_782[15:14]};
assign col_out_786 = {u_ca_out_786[1:0],u_ca_out_785[7:2], u_ca_out_784[13:8], u_ca_out_783[15:14]};
assign col_out_787 = {u_ca_out_787[1:0],u_ca_out_786[7:2], u_ca_out_785[13:8], u_ca_out_784[15:14]};
assign col_out_788 = {u_ca_out_788[1:0],u_ca_out_787[7:2], u_ca_out_786[13:8], u_ca_out_785[15:14]};
assign col_out_789 = {u_ca_out_789[1:0],u_ca_out_788[7:2], u_ca_out_787[13:8], u_ca_out_786[15:14]};
assign col_out_790 = {u_ca_out_790[1:0],u_ca_out_789[7:2], u_ca_out_788[13:8], u_ca_out_787[15:14]};
assign col_out_791 = {u_ca_out_791[1:0],u_ca_out_790[7:2], u_ca_out_789[13:8], u_ca_out_788[15:14]};
assign col_out_792 = {u_ca_out_792[1:0],u_ca_out_791[7:2], u_ca_out_790[13:8], u_ca_out_789[15:14]};
assign col_out_793 = {u_ca_out_793[1:0],u_ca_out_792[7:2], u_ca_out_791[13:8], u_ca_out_790[15:14]};
assign col_out_794 = {u_ca_out_794[1:0],u_ca_out_793[7:2], u_ca_out_792[13:8], u_ca_out_791[15:14]};
assign col_out_795 = {u_ca_out_795[1:0],u_ca_out_794[7:2], u_ca_out_793[13:8], u_ca_out_792[15:14]};
assign col_out_796 = {u_ca_out_796[1:0],u_ca_out_795[7:2], u_ca_out_794[13:8], u_ca_out_793[15:14]};
assign col_out_797 = {u_ca_out_797[1:0],u_ca_out_796[7:2], u_ca_out_795[13:8], u_ca_out_794[15:14]};
assign col_out_798 = {u_ca_out_798[1:0],u_ca_out_797[7:2], u_ca_out_796[13:8], u_ca_out_795[15:14]};
assign col_out_799 = {u_ca_out_799[1:0],u_ca_out_798[7:2], u_ca_out_797[13:8], u_ca_out_796[15:14]};
assign col_out_800 = {u_ca_out_800[1:0],u_ca_out_799[7:2], u_ca_out_798[13:8], u_ca_out_797[15:14]};
assign col_out_801 = {u_ca_out_801[1:0],u_ca_out_800[7:2], u_ca_out_799[13:8], u_ca_out_798[15:14]};
assign col_out_802 = {u_ca_out_802[1:0],u_ca_out_801[7:2], u_ca_out_800[13:8], u_ca_out_799[15:14]};
assign col_out_803 = {u_ca_out_803[1:0],u_ca_out_802[7:2], u_ca_out_801[13:8], u_ca_out_800[15:14]};
assign col_out_804 = {u_ca_out_804[1:0],u_ca_out_803[7:2], u_ca_out_802[13:8], u_ca_out_801[15:14]};
assign col_out_805 = {u_ca_out_805[1:0],u_ca_out_804[7:2], u_ca_out_803[13:8], u_ca_out_802[15:14]};
assign col_out_806 = {u_ca_out_806[1:0],u_ca_out_805[7:2], u_ca_out_804[13:8], u_ca_out_803[15:14]};
assign col_out_807 = {u_ca_out_807[1:0],u_ca_out_806[7:2], u_ca_out_805[13:8], u_ca_out_804[15:14]};
assign col_out_808 = {u_ca_out_808[1:0],u_ca_out_807[7:2], u_ca_out_806[13:8], u_ca_out_805[15:14]};
assign col_out_809 = {u_ca_out_809[1:0],u_ca_out_808[7:2], u_ca_out_807[13:8], u_ca_out_806[15:14]};
assign col_out_810 = {u_ca_out_810[1:0],u_ca_out_809[7:2], u_ca_out_808[13:8], u_ca_out_807[15:14]};
assign col_out_811 = {u_ca_out_811[1:0],u_ca_out_810[7:2], u_ca_out_809[13:8], u_ca_out_808[15:14]};
assign col_out_812 = {u_ca_out_812[1:0],u_ca_out_811[7:2], u_ca_out_810[13:8], u_ca_out_809[15:14]};
assign col_out_813 = {u_ca_out_813[1:0],u_ca_out_812[7:2], u_ca_out_811[13:8], u_ca_out_810[15:14]};
assign col_out_814 = {u_ca_out_814[1:0],u_ca_out_813[7:2], u_ca_out_812[13:8], u_ca_out_811[15:14]};
assign col_out_815 = {u_ca_out_815[1:0],u_ca_out_814[7:2], u_ca_out_813[13:8], u_ca_out_812[15:14]};
assign col_out_816 = {u_ca_out_816[1:0],u_ca_out_815[7:2], u_ca_out_814[13:8], u_ca_out_813[15:14]};
assign col_out_817 = {u_ca_out_817[1:0],u_ca_out_816[7:2], u_ca_out_815[13:8], u_ca_out_814[15:14]};
assign col_out_818 = {u_ca_out_818[1:0],u_ca_out_817[7:2], u_ca_out_816[13:8], u_ca_out_815[15:14]};
assign col_out_819 = {u_ca_out_819[1:0],u_ca_out_818[7:2], u_ca_out_817[13:8], u_ca_out_816[15:14]};
assign col_out_820 = {u_ca_out_820[1:0],u_ca_out_819[7:2], u_ca_out_818[13:8], u_ca_out_817[15:14]};
assign col_out_821 = {u_ca_out_821[1:0],u_ca_out_820[7:2], u_ca_out_819[13:8], u_ca_out_818[15:14]};
assign col_out_822 = {u_ca_out_822[1:0],u_ca_out_821[7:2], u_ca_out_820[13:8], u_ca_out_819[15:14]};
assign col_out_823 = {u_ca_out_823[1:0],u_ca_out_822[7:2], u_ca_out_821[13:8], u_ca_out_820[15:14]};
assign col_out_824 = {u_ca_out_824[1:0],u_ca_out_823[7:2], u_ca_out_822[13:8], u_ca_out_821[15:14]};
assign col_out_825 = {u_ca_out_825[1:0],u_ca_out_824[7:2], u_ca_out_823[13:8], u_ca_out_822[15:14]};
assign col_out_826 = {u_ca_out_826[1:0],u_ca_out_825[7:2], u_ca_out_824[13:8], u_ca_out_823[15:14]};
assign col_out_827 = {u_ca_out_827[1:0],u_ca_out_826[7:2], u_ca_out_825[13:8], u_ca_out_824[15:14]};
assign col_out_828 = {u_ca_out_828[1:0],u_ca_out_827[7:2], u_ca_out_826[13:8], u_ca_out_825[15:14]};
assign col_out_829 = {u_ca_out_829[1:0],u_ca_out_828[7:2], u_ca_out_827[13:8], u_ca_out_826[15:14]};
assign col_out_830 = {u_ca_out_830[1:0],u_ca_out_829[7:2], u_ca_out_828[13:8], u_ca_out_827[15:14]};
assign col_out_831 = {u_ca_out_831[1:0],u_ca_out_830[7:2], u_ca_out_829[13:8], u_ca_out_828[15:14]};
assign col_out_832 = {u_ca_out_832[1:0],u_ca_out_831[7:2], u_ca_out_830[13:8], u_ca_out_829[15:14]};
assign col_out_833 = {u_ca_out_833[1:0],u_ca_out_832[7:2], u_ca_out_831[13:8], u_ca_out_830[15:14]};
assign col_out_834 = {u_ca_out_834[1:0],u_ca_out_833[7:2], u_ca_out_832[13:8], u_ca_out_831[15:14]};
assign col_out_835 = {u_ca_out_835[1:0],u_ca_out_834[7:2], u_ca_out_833[13:8], u_ca_out_832[15:14]};
assign col_out_836 = {u_ca_out_836[1:0],u_ca_out_835[7:2], u_ca_out_834[13:8], u_ca_out_833[15:14]};
assign col_out_837 = {u_ca_out_837[1:0],u_ca_out_836[7:2], u_ca_out_835[13:8], u_ca_out_834[15:14]};
assign col_out_838 = {u_ca_out_838[1:0],u_ca_out_837[7:2], u_ca_out_836[13:8], u_ca_out_835[15:14]};
assign col_out_839 = {u_ca_out_839[1:0],u_ca_out_838[7:2], u_ca_out_837[13:8], u_ca_out_836[15:14]};
assign col_out_840 = {u_ca_out_840[1:0],u_ca_out_839[7:2], u_ca_out_838[13:8], u_ca_out_837[15:14]};
assign col_out_841 = {u_ca_out_841[1:0],u_ca_out_840[7:2], u_ca_out_839[13:8], u_ca_out_838[15:14]};
assign col_out_842 = {u_ca_out_842[1:0],u_ca_out_841[7:2], u_ca_out_840[13:8], u_ca_out_839[15:14]};
assign col_out_843 = {u_ca_out_843[1:0],u_ca_out_842[7:2], u_ca_out_841[13:8], u_ca_out_840[15:14]};
assign col_out_844 = {u_ca_out_844[1:0],u_ca_out_843[7:2], u_ca_out_842[13:8], u_ca_out_841[15:14]};
assign col_out_845 = {u_ca_out_845[1:0],u_ca_out_844[7:2], u_ca_out_843[13:8], u_ca_out_842[15:14]};
assign col_out_846 = {u_ca_out_846[1:0],u_ca_out_845[7:2], u_ca_out_844[13:8], u_ca_out_843[15:14]};
assign col_out_847 = {u_ca_out_847[1:0],u_ca_out_846[7:2], u_ca_out_845[13:8], u_ca_out_844[15:14]};
assign col_out_848 = {u_ca_out_848[1:0],u_ca_out_847[7:2], u_ca_out_846[13:8], u_ca_out_845[15:14]};
assign col_out_849 = {u_ca_out_849[1:0],u_ca_out_848[7:2], u_ca_out_847[13:8], u_ca_out_846[15:14]};
assign col_out_850 = {u_ca_out_850[1:0],u_ca_out_849[7:2], u_ca_out_848[13:8], u_ca_out_847[15:14]};
assign col_out_851 = {u_ca_out_851[1:0],u_ca_out_850[7:2], u_ca_out_849[13:8], u_ca_out_848[15:14]};
assign col_out_852 = {u_ca_out_852[1:0],u_ca_out_851[7:2], u_ca_out_850[13:8], u_ca_out_849[15:14]};
assign col_out_853 = {u_ca_out_853[1:0],u_ca_out_852[7:2], u_ca_out_851[13:8], u_ca_out_850[15:14]};
assign col_out_854 = {u_ca_out_854[1:0],u_ca_out_853[7:2], u_ca_out_852[13:8], u_ca_out_851[15:14]};
assign col_out_855 = {u_ca_out_855[1:0],u_ca_out_854[7:2], u_ca_out_853[13:8], u_ca_out_852[15:14]};
assign col_out_856 = {u_ca_out_856[1:0],u_ca_out_855[7:2], u_ca_out_854[13:8], u_ca_out_853[15:14]};
assign col_out_857 = {u_ca_out_857[1:0],u_ca_out_856[7:2], u_ca_out_855[13:8], u_ca_out_854[15:14]};
assign col_out_858 = {u_ca_out_858[1:0],u_ca_out_857[7:2], u_ca_out_856[13:8], u_ca_out_855[15:14]};
assign col_out_859 = {u_ca_out_859[1:0],u_ca_out_858[7:2], u_ca_out_857[13:8], u_ca_out_856[15:14]};
assign col_out_860 = {u_ca_out_860[1:0],u_ca_out_859[7:2], u_ca_out_858[13:8], u_ca_out_857[15:14]};
assign col_out_861 = {u_ca_out_861[1:0],u_ca_out_860[7:2], u_ca_out_859[13:8], u_ca_out_858[15:14]};
assign col_out_862 = {u_ca_out_862[1:0],u_ca_out_861[7:2], u_ca_out_860[13:8], u_ca_out_859[15:14]};
assign col_out_863 = {u_ca_out_863[1:0],u_ca_out_862[7:2], u_ca_out_861[13:8], u_ca_out_860[15:14]};
assign col_out_864 = {u_ca_out_864[1:0],u_ca_out_863[7:2], u_ca_out_862[13:8], u_ca_out_861[15:14]};
assign col_out_865 = {u_ca_out_865[1:0],u_ca_out_864[7:2], u_ca_out_863[13:8], u_ca_out_862[15:14]};
assign col_out_866 = {u_ca_out_866[1:0],u_ca_out_865[7:2], u_ca_out_864[13:8], u_ca_out_863[15:14]};
assign col_out_867 = {u_ca_out_867[1:0],u_ca_out_866[7:2], u_ca_out_865[13:8], u_ca_out_864[15:14]};
assign col_out_868 = {u_ca_out_868[1:0],u_ca_out_867[7:2], u_ca_out_866[13:8], u_ca_out_865[15:14]};
assign col_out_869 = {u_ca_out_869[1:0],u_ca_out_868[7:2], u_ca_out_867[13:8], u_ca_out_866[15:14]};
assign col_out_870 = {u_ca_out_870[1:0],u_ca_out_869[7:2], u_ca_out_868[13:8], u_ca_out_867[15:14]};
assign col_out_871 = {u_ca_out_871[1:0],u_ca_out_870[7:2], u_ca_out_869[13:8], u_ca_out_868[15:14]};
assign col_out_872 = {u_ca_out_872[1:0],u_ca_out_871[7:2], u_ca_out_870[13:8], u_ca_out_869[15:14]};
assign col_out_873 = {u_ca_out_873[1:0],u_ca_out_872[7:2], u_ca_out_871[13:8], u_ca_out_870[15:14]};
assign col_out_874 = {u_ca_out_874[1:0],u_ca_out_873[7:2], u_ca_out_872[13:8], u_ca_out_871[15:14]};
assign col_out_875 = {u_ca_out_875[1:0],u_ca_out_874[7:2], u_ca_out_873[13:8], u_ca_out_872[15:14]};
assign col_out_876 = {u_ca_out_876[1:0],u_ca_out_875[7:2], u_ca_out_874[13:8], u_ca_out_873[15:14]};
assign col_out_877 = {u_ca_out_877[1:0],u_ca_out_876[7:2], u_ca_out_875[13:8], u_ca_out_874[15:14]};
assign col_out_878 = {u_ca_out_878[1:0],u_ca_out_877[7:2], u_ca_out_876[13:8], u_ca_out_875[15:14]};
assign col_out_879 = {u_ca_out_879[1:0],u_ca_out_878[7:2], u_ca_out_877[13:8], u_ca_out_876[15:14]};
assign col_out_880 = {u_ca_out_880[1:0],u_ca_out_879[7:2], u_ca_out_878[13:8], u_ca_out_877[15:14]};
assign col_out_881 = {u_ca_out_881[1:0],u_ca_out_880[7:2], u_ca_out_879[13:8], u_ca_out_878[15:14]};
assign col_out_882 = {u_ca_out_882[1:0],u_ca_out_881[7:2], u_ca_out_880[13:8], u_ca_out_879[15:14]};
assign col_out_883 = {u_ca_out_883[1:0],u_ca_out_882[7:2], u_ca_out_881[13:8], u_ca_out_880[15:14]};
assign col_out_884 = {u_ca_out_884[1:0],u_ca_out_883[7:2], u_ca_out_882[13:8], u_ca_out_881[15:14]};
assign col_out_885 = {u_ca_out_885[1:0],u_ca_out_884[7:2], u_ca_out_883[13:8], u_ca_out_882[15:14]};
assign col_out_886 = {u_ca_out_886[1:0],u_ca_out_885[7:2], u_ca_out_884[13:8], u_ca_out_883[15:14]};
assign col_out_887 = {u_ca_out_887[1:0],u_ca_out_886[7:2], u_ca_out_885[13:8], u_ca_out_884[15:14]};
assign col_out_888 = {u_ca_out_888[1:0],u_ca_out_887[7:2], u_ca_out_886[13:8], u_ca_out_885[15:14]};
assign col_out_889 = {u_ca_out_889[1:0],u_ca_out_888[7:2], u_ca_out_887[13:8], u_ca_out_886[15:14]};
assign col_out_890 = {u_ca_out_890[1:0],u_ca_out_889[7:2], u_ca_out_888[13:8], u_ca_out_887[15:14]};
assign col_out_891 = {u_ca_out_891[1:0],u_ca_out_890[7:2], u_ca_out_889[13:8], u_ca_out_888[15:14]};
assign col_out_892 = {u_ca_out_892[1:0],u_ca_out_891[7:2], u_ca_out_890[13:8], u_ca_out_889[15:14]};
assign col_out_893 = {u_ca_out_893[1:0],u_ca_out_892[7:2], u_ca_out_891[13:8], u_ca_out_890[15:14]};
assign col_out_894 = {u_ca_out_894[1:0],u_ca_out_893[7:2], u_ca_out_892[13:8], u_ca_out_891[15:14]};
assign col_out_895 = {u_ca_out_895[1:0],u_ca_out_894[7:2], u_ca_out_893[13:8], u_ca_out_892[15:14]};
assign col_out_896 = {u_ca_out_896[1:0],u_ca_out_895[7:2], u_ca_out_894[13:8], u_ca_out_893[15:14]};
assign col_out_897 = {u_ca_out_897[1:0],u_ca_out_896[7:2], u_ca_out_895[13:8], u_ca_out_894[15:14]};
assign col_out_898 = {u_ca_out_898[1:0],u_ca_out_897[7:2], u_ca_out_896[13:8], u_ca_out_895[15:14]};
assign col_out_899 = {u_ca_out_899[1:0],u_ca_out_898[7:2], u_ca_out_897[13:8], u_ca_out_896[15:14]};
assign col_out_900 = {u_ca_out_900[1:0],u_ca_out_899[7:2], u_ca_out_898[13:8], u_ca_out_897[15:14]};
assign col_out_901 = {u_ca_out_901[1:0],u_ca_out_900[7:2], u_ca_out_899[13:8], u_ca_out_898[15:14]};
assign col_out_902 = {u_ca_out_902[1:0],u_ca_out_901[7:2], u_ca_out_900[13:8], u_ca_out_899[15:14]};
assign col_out_903 = {u_ca_out_903[1:0],u_ca_out_902[7:2], u_ca_out_901[13:8], u_ca_out_900[15:14]};
assign col_out_904 = {u_ca_out_904[1:0],u_ca_out_903[7:2], u_ca_out_902[13:8], u_ca_out_901[15:14]};
assign col_out_905 = {u_ca_out_905[1:0],u_ca_out_904[7:2], u_ca_out_903[13:8], u_ca_out_902[15:14]};
assign col_out_906 = {u_ca_out_906[1:0],u_ca_out_905[7:2], u_ca_out_904[13:8], u_ca_out_903[15:14]};
assign col_out_907 = {u_ca_out_907[1:0],u_ca_out_906[7:2], u_ca_out_905[13:8], u_ca_out_904[15:14]};
assign col_out_908 = {u_ca_out_908[1:0],u_ca_out_907[7:2], u_ca_out_906[13:8], u_ca_out_905[15:14]};
assign col_out_909 = {u_ca_out_909[1:0],u_ca_out_908[7:2], u_ca_out_907[13:8], u_ca_out_906[15:14]};
assign col_out_910 = {u_ca_out_910[1:0],u_ca_out_909[7:2], u_ca_out_908[13:8], u_ca_out_907[15:14]};
assign col_out_911 = {u_ca_out_911[1:0],u_ca_out_910[7:2], u_ca_out_909[13:8], u_ca_out_908[15:14]};
assign col_out_912 = {u_ca_out_912[1:0],u_ca_out_911[7:2], u_ca_out_910[13:8], u_ca_out_909[15:14]};
assign col_out_913 = {u_ca_out_913[1:0],u_ca_out_912[7:2], u_ca_out_911[13:8], u_ca_out_910[15:14]};
assign col_out_914 = {u_ca_out_914[1:0],u_ca_out_913[7:2], u_ca_out_912[13:8], u_ca_out_911[15:14]};
assign col_out_915 = {u_ca_out_915[1:0],u_ca_out_914[7:2], u_ca_out_913[13:8], u_ca_out_912[15:14]};
assign col_out_916 = {u_ca_out_916[1:0],u_ca_out_915[7:2], u_ca_out_914[13:8], u_ca_out_913[15:14]};
assign col_out_917 = {u_ca_out_917[1:0],u_ca_out_916[7:2], u_ca_out_915[13:8], u_ca_out_914[15:14]};
assign col_out_918 = {u_ca_out_918[1:0],u_ca_out_917[7:2], u_ca_out_916[13:8], u_ca_out_915[15:14]};
assign col_out_919 = {u_ca_out_919[1:0],u_ca_out_918[7:2], u_ca_out_917[13:8], u_ca_out_916[15:14]};
assign col_out_920 = {u_ca_out_920[1:0],u_ca_out_919[7:2], u_ca_out_918[13:8], u_ca_out_917[15:14]};
assign col_out_921 = {u_ca_out_921[1:0],u_ca_out_920[7:2], u_ca_out_919[13:8], u_ca_out_918[15:14]};
assign col_out_922 = {u_ca_out_922[1:0],u_ca_out_921[7:2], u_ca_out_920[13:8], u_ca_out_919[15:14]};
assign col_out_923 = {u_ca_out_923[1:0],u_ca_out_922[7:2], u_ca_out_921[13:8], u_ca_out_920[15:14]};
assign col_out_924 = {u_ca_out_924[1:0],u_ca_out_923[7:2], u_ca_out_922[13:8], u_ca_out_921[15:14]};
assign col_out_925 = {u_ca_out_925[1:0],u_ca_out_924[7:2], u_ca_out_923[13:8], u_ca_out_922[15:14]};
assign col_out_926 = {u_ca_out_926[1:0],u_ca_out_925[7:2], u_ca_out_924[13:8], u_ca_out_923[15:14]};
assign col_out_927 = {u_ca_out_927[1:0],u_ca_out_926[7:2], u_ca_out_925[13:8], u_ca_out_924[15:14]};
assign col_out_928 = {u_ca_out_928[1:0],u_ca_out_927[7:2], u_ca_out_926[13:8], u_ca_out_925[15:14]};
assign col_out_929 = {u_ca_out_929[1:0],u_ca_out_928[7:2], u_ca_out_927[13:8], u_ca_out_926[15:14]};
assign col_out_930 = {u_ca_out_930[1:0],u_ca_out_929[7:2], u_ca_out_928[13:8], u_ca_out_927[15:14]};
assign col_out_931 = {u_ca_out_931[1:0],u_ca_out_930[7:2], u_ca_out_929[13:8], u_ca_out_928[15:14]};
assign col_out_932 = {u_ca_out_932[1:0],u_ca_out_931[7:2], u_ca_out_930[13:8], u_ca_out_929[15:14]};
assign col_out_933 = {u_ca_out_933[1:0],u_ca_out_932[7:2], u_ca_out_931[13:8], u_ca_out_930[15:14]};
assign col_out_934 = {u_ca_out_934[1:0],u_ca_out_933[7:2], u_ca_out_932[13:8], u_ca_out_931[15:14]};
assign col_out_935 = {u_ca_out_935[1:0],u_ca_out_934[7:2], u_ca_out_933[13:8], u_ca_out_932[15:14]};
assign col_out_936 = {u_ca_out_936[1:0],u_ca_out_935[7:2], u_ca_out_934[13:8], u_ca_out_933[15:14]};
assign col_out_937 = {u_ca_out_937[1:0],u_ca_out_936[7:2], u_ca_out_935[13:8], u_ca_out_934[15:14]};
assign col_out_938 = {u_ca_out_938[1:0],u_ca_out_937[7:2], u_ca_out_936[13:8], u_ca_out_935[15:14]};
assign col_out_939 = {u_ca_out_939[1:0],u_ca_out_938[7:2], u_ca_out_937[13:8], u_ca_out_936[15:14]};
assign col_out_940 = {u_ca_out_940[1:0],u_ca_out_939[7:2], u_ca_out_938[13:8], u_ca_out_937[15:14]};
assign col_out_941 = {u_ca_out_941[1:0],u_ca_out_940[7:2], u_ca_out_939[13:8], u_ca_out_938[15:14]};
assign col_out_942 = {u_ca_out_942[1:0],u_ca_out_941[7:2], u_ca_out_940[13:8], u_ca_out_939[15:14]};
assign col_out_943 = {u_ca_out_943[1:0],u_ca_out_942[7:2], u_ca_out_941[13:8], u_ca_out_940[15:14]};
assign col_out_944 = {u_ca_out_944[1:0],u_ca_out_943[7:2], u_ca_out_942[13:8], u_ca_out_941[15:14]};
assign col_out_945 = {u_ca_out_945[1:0],u_ca_out_944[7:2], u_ca_out_943[13:8], u_ca_out_942[15:14]};
assign col_out_946 = {u_ca_out_946[1:0],u_ca_out_945[7:2], u_ca_out_944[13:8], u_ca_out_943[15:14]};
assign col_out_947 = {u_ca_out_947[1:0],u_ca_out_946[7:2], u_ca_out_945[13:8], u_ca_out_944[15:14]};
assign col_out_948 = {u_ca_out_948[1:0],u_ca_out_947[7:2], u_ca_out_946[13:8], u_ca_out_945[15:14]};
assign col_out_949 = {u_ca_out_949[1:0],u_ca_out_948[7:2], u_ca_out_947[13:8], u_ca_out_946[15:14]};
assign col_out_950 = {u_ca_out_950[1:0],u_ca_out_949[7:2], u_ca_out_948[13:8], u_ca_out_947[15:14]};
assign col_out_951 = {u_ca_out_951[1:0],u_ca_out_950[7:2], u_ca_out_949[13:8], u_ca_out_948[15:14]};
assign col_out_952 = {u_ca_out_952[1:0],u_ca_out_951[7:2], u_ca_out_950[13:8], u_ca_out_949[15:14]};
assign col_out_953 = {u_ca_out_953[1:0],u_ca_out_952[7:2], u_ca_out_951[13:8], u_ca_out_950[15:14]};
assign col_out_954 = {u_ca_out_954[1:0],u_ca_out_953[7:2], u_ca_out_952[13:8], u_ca_out_951[15:14]};
assign col_out_955 = {u_ca_out_955[1:0],u_ca_out_954[7:2], u_ca_out_953[13:8], u_ca_out_952[15:14]};
assign col_out_956 = {u_ca_out_956[1:0],u_ca_out_955[7:2], u_ca_out_954[13:8], u_ca_out_953[15:14]};
assign col_out_957 = {u_ca_out_957[1:0],u_ca_out_956[7:2], u_ca_out_955[13:8], u_ca_out_954[15:14]};
assign col_out_958 = {u_ca_out_958[1:0],u_ca_out_957[7:2], u_ca_out_956[13:8], u_ca_out_955[15:14]};
assign col_out_959 = {u_ca_out_959[1:0],u_ca_out_958[7:2], u_ca_out_957[13:8], u_ca_out_956[15:14]};
assign col_out_960 = {u_ca_out_960[1:0],u_ca_out_959[7:2], u_ca_out_958[13:8], u_ca_out_957[15:14]};
assign col_out_961 = {u_ca_out_961[1:0],u_ca_out_960[7:2], u_ca_out_959[13:8], u_ca_out_958[15:14]};
assign col_out_962 = {u_ca_out_962[1:0],u_ca_out_961[7:2], u_ca_out_960[13:8], u_ca_out_959[15:14]};
assign col_out_963 = {u_ca_out_963[1:0],u_ca_out_962[7:2], u_ca_out_961[13:8], u_ca_out_960[15:14]};
assign col_out_964 = {u_ca_out_964[1:0],u_ca_out_963[7:2], u_ca_out_962[13:8], u_ca_out_961[15:14]};
assign col_out_965 = {u_ca_out_965[1:0],u_ca_out_964[7:2], u_ca_out_963[13:8], u_ca_out_962[15:14]};
assign col_out_966 = {u_ca_out_966[1:0],u_ca_out_965[7:2], u_ca_out_964[13:8], u_ca_out_963[15:14]};
assign col_out_967 = {u_ca_out_967[1:0],u_ca_out_966[7:2], u_ca_out_965[13:8], u_ca_out_964[15:14]};
assign col_out_968 = {u_ca_out_968[1:0],u_ca_out_967[7:2], u_ca_out_966[13:8], u_ca_out_965[15:14]};
assign col_out_969 = {u_ca_out_969[1:0],u_ca_out_968[7:2], u_ca_out_967[13:8], u_ca_out_966[15:14]};
assign col_out_970 = {u_ca_out_970[1:0],u_ca_out_969[7:2], u_ca_out_968[13:8], u_ca_out_967[15:14]};
assign col_out_971 = {u_ca_out_971[1:0],u_ca_out_970[7:2], u_ca_out_969[13:8], u_ca_out_968[15:14]};
assign col_out_972 = {u_ca_out_972[1:0],u_ca_out_971[7:2], u_ca_out_970[13:8], u_ca_out_969[15:14]};
assign col_out_973 = {u_ca_out_973[1:0],u_ca_out_972[7:2], u_ca_out_971[13:8], u_ca_out_970[15:14]};
assign col_out_974 = {u_ca_out_974[1:0],u_ca_out_973[7:2], u_ca_out_972[13:8], u_ca_out_971[15:14]};
assign col_out_975 = {u_ca_out_975[1:0],u_ca_out_974[7:2], u_ca_out_973[13:8], u_ca_out_972[15:14]};
assign col_out_976 = {u_ca_out_976[1:0],u_ca_out_975[7:2], u_ca_out_974[13:8], u_ca_out_973[15:14]};
assign col_out_977 = {u_ca_out_977[1:0],u_ca_out_976[7:2], u_ca_out_975[13:8], u_ca_out_974[15:14]};
assign col_out_978 = {u_ca_out_978[1:0],u_ca_out_977[7:2], u_ca_out_976[13:8], u_ca_out_975[15:14]};
assign col_out_979 = {u_ca_out_979[1:0],u_ca_out_978[7:2], u_ca_out_977[13:8], u_ca_out_976[15:14]};
assign col_out_980 = {u_ca_out_980[1:0],u_ca_out_979[7:2], u_ca_out_978[13:8], u_ca_out_977[15:14]};
assign col_out_981 = {u_ca_out_981[1:0],u_ca_out_980[7:2], u_ca_out_979[13:8], u_ca_out_978[15:14]};
assign col_out_982 = {u_ca_out_982[1:0],u_ca_out_981[7:2], u_ca_out_980[13:8], u_ca_out_979[15:14]};
assign col_out_983 = {u_ca_out_983[1:0],u_ca_out_982[7:2], u_ca_out_981[13:8], u_ca_out_980[15:14]};
assign col_out_984 = {u_ca_out_984[1:0],u_ca_out_983[7:2], u_ca_out_982[13:8], u_ca_out_981[15:14]};
assign col_out_985 = {u_ca_out_985[1:0],u_ca_out_984[7:2], u_ca_out_983[13:8], u_ca_out_982[15:14]};
assign col_out_986 = {u_ca_out_986[1:0],u_ca_out_985[7:2], u_ca_out_984[13:8], u_ca_out_983[15:14]};
assign col_out_987 = {u_ca_out_987[1:0],u_ca_out_986[7:2], u_ca_out_985[13:8], u_ca_out_984[15:14]};
assign col_out_988 = {u_ca_out_988[1:0],u_ca_out_987[7:2], u_ca_out_986[13:8], u_ca_out_985[15:14]};
assign col_out_989 = {u_ca_out_989[1:0],u_ca_out_988[7:2], u_ca_out_987[13:8], u_ca_out_986[15:14]};
assign col_out_990 = {u_ca_out_990[1:0],u_ca_out_989[7:2], u_ca_out_988[13:8], u_ca_out_987[15:14]};
assign col_out_991 = {u_ca_out_991[1:0],u_ca_out_990[7:2], u_ca_out_989[13:8], u_ca_out_988[15:14]};
assign col_out_992 = {u_ca_out_992[1:0],u_ca_out_991[7:2], u_ca_out_990[13:8], u_ca_out_989[15:14]};
assign col_out_993 = {u_ca_out_993[1:0],u_ca_out_992[7:2], u_ca_out_991[13:8], u_ca_out_990[15:14]};
assign col_out_994 = {u_ca_out_994[1:0],u_ca_out_993[7:2], u_ca_out_992[13:8], u_ca_out_991[15:14]};
assign col_out_995 = {u_ca_out_995[1:0],u_ca_out_994[7:2], u_ca_out_993[13:8], u_ca_out_992[15:14]};
assign col_out_996 = {u_ca_out_996[1:0],u_ca_out_995[7:2], u_ca_out_994[13:8], u_ca_out_993[15:14]};
assign col_out_997 = {u_ca_out_997[1:0],u_ca_out_996[7:2], u_ca_out_995[13:8], u_ca_out_994[15:14]};
assign col_out_998 = {u_ca_out_998[1:0],u_ca_out_997[7:2], u_ca_out_996[13:8], u_ca_out_995[15:14]};
assign col_out_999 = {u_ca_out_999[1:0],u_ca_out_998[7:2], u_ca_out_997[13:8], u_ca_out_996[15:14]};
assign col_out_1000 = {u_ca_out_1000[1:0],u_ca_out_999[7:2], u_ca_out_998[13:8], u_ca_out_997[15:14]};
assign col_out_1001 = {u_ca_out_1001[1:0],u_ca_out_1000[7:2], u_ca_out_999[13:8], u_ca_out_998[15:14]};
assign col_out_1002 = {u_ca_out_1002[1:0],u_ca_out_1001[7:2], u_ca_out_1000[13:8], u_ca_out_999[15:14]};
assign col_out_1003 = {u_ca_out_1003[1:0],u_ca_out_1002[7:2], u_ca_out_1001[13:8], u_ca_out_1000[15:14]};
assign col_out_1004 = {u_ca_out_1004[1:0],u_ca_out_1003[7:2], u_ca_out_1002[13:8], u_ca_out_1001[15:14]};
assign col_out_1005 = {u_ca_out_1005[1:0],u_ca_out_1004[7:2], u_ca_out_1003[13:8], u_ca_out_1002[15:14]};
assign col_out_1006 = {u_ca_out_1006[1:0],u_ca_out_1005[7:2], u_ca_out_1004[13:8], u_ca_out_1003[15:14]};
assign col_out_1007 = {u_ca_out_1007[1:0],u_ca_out_1006[7:2], u_ca_out_1005[13:8], u_ca_out_1004[15:14]};
assign col_out_1008 = {u_ca_out_1008[1:0],u_ca_out_1007[7:2], u_ca_out_1006[13:8], u_ca_out_1005[15:14]};
assign col_out_1009 = {u_ca_out_1009[1:0],u_ca_out_1008[7:2], u_ca_out_1007[13:8], u_ca_out_1006[15:14]};
assign col_out_1010 = {u_ca_out_1010[1:0],u_ca_out_1009[7:2], u_ca_out_1008[13:8], u_ca_out_1007[15:14]};
assign col_out_1011 = {u_ca_out_1011[1:0],u_ca_out_1010[7:2], u_ca_out_1009[13:8], u_ca_out_1008[15:14]};
assign col_out_1012 = {u_ca_out_1012[1:0],u_ca_out_1011[7:2], u_ca_out_1010[13:8], u_ca_out_1009[15:14]};
assign col_out_1013 = {u_ca_out_1013[1:0],u_ca_out_1012[7:2], u_ca_out_1011[13:8], u_ca_out_1010[15:14]};
assign col_out_1014 = {u_ca_out_1014[1:0],u_ca_out_1013[7:2], u_ca_out_1012[13:8], u_ca_out_1011[15:14]};
assign col_out_1015 = {u_ca_out_1015[1:0],u_ca_out_1014[7:2], u_ca_out_1013[13:8], u_ca_out_1012[15:14]};
assign col_out_1016 = {u_ca_out_1016[1:0],u_ca_out_1015[7:2], u_ca_out_1014[13:8], u_ca_out_1013[15:14]};
assign col_out_1017 = {u_ca_out_1017[1:0],u_ca_out_1016[7:2], u_ca_out_1015[13:8], u_ca_out_1014[15:14]};
assign col_out_1018 = {u_ca_out_1018[1:0],u_ca_out_1017[7:2], u_ca_out_1016[13:8], u_ca_out_1015[15:14]};
assign col_out_1019 = {u_ca_out_1019[1:0],u_ca_out_1018[7:2], u_ca_out_1017[13:8], u_ca_out_1016[15:14]};
assign col_out_1020 = {u_ca_out_1020[1:0],u_ca_out_1019[7:2], u_ca_out_1018[13:8], u_ca_out_1017[15:14]};
assign col_out_1021 = {u_ca_out_1021[1:0],u_ca_out_1020[7:2], u_ca_out_1019[13:8], u_ca_out_1018[15:14]};
assign col_out_1022 = {u_ca_out_1022[1:0],u_ca_out_1021[7:2], u_ca_out_1020[13:8], u_ca_out_1019[15:14]};
assign col_out_1023 = {u_ca_out_1023[1:0],u_ca_out_1022[7:2], u_ca_out_1021[13:8], u_ca_out_1020[15:14]};
assign col_out_1024 = {u_ca_out_1024[1:0],u_ca_out_1023[7:2], u_ca_out_1022[13:8], u_ca_out_1021[15:14]};
assign col_out_1025 = {u_ca_out_1025[1:0],u_ca_out_1024[7:2], u_ca_out_1023[13:8], u_ca_out_1022[15:14]};
assign col_out_1026 = {u_ca_out_1026[1:0],u_ca_out_1025[7:2], u_ca_out_1024[13:8], u_ca_out_1023[15:14]};
assign col_out_1027 = {u_ca_out_1027[1:0],u_ca_out_1026[7:2], u_ca_out_1025[13:8], u_ca_out_1024[15:14]};
assign col_out_1028 = {u_ca_out_1028[1:0],u_ca_out_1027[7:2], u_ca_out_1026[13:8], u_ca_out_1025[15:14]};
assign col_out_1029 = {u_ca_out_1029[1:0],u_ca_out_1028[7:2], u_ca_out_1027[13:8], u_ca_out_1026[15:14]};
assign col_out_1030 = {{2{1'b0}}, u_ca_out_1029[7:2], u_ca_out_1028[13:8], u_ca_out_1027[15:14]};
assign col_out_1031 = {{8{1'b0}}, u_ca_out_1029[13:8], u_ca_out_1028[15:14]};
assign col_out_1032 = {{14{1'b0}}, u_ca_out_1029[15:14]};

//---------------------------------------------------------


endmodule
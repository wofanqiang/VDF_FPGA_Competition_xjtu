module xpb_5_840
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h94d69e055f6d4eaa4e81729c53c2aa5c16637515c725ebc27f3c9a9a7fd1ce9c1c1a2a16d29bcc068b475cb0dba6ef70f954e3e9189a7c40bab967cc97cb9ae659070361afeda489ad543e5b734c755f5c28bc024f0c1f2a44896ac01ec539f5d434397d5da303a8e1ab18f99121ecf028c6bbeb55f7062658381a4be01c05e3;
    5'b00010 : xpb = 1024'h78fff6b4fcec688bd1fd6d61972b0d66bb50e6fab8d4370d809c7bdf4ca0f03034ebd6b4db11197e77307a1ad3efce178e8f9fec0e822835c4d3903af4c4c11b3dbed214b04a4bce480e7a144dbd268dc44c7e6c11921143d3864385835fd1597960e0d10a7d0ec43c964b142a73b3b702b398f45ba2af1c6a00b9933755a55b;
    5'b00011 : xpb = 1024'h5d294f649a6b826d55796826da937071603e58dfaa82825881fc5d24197011c44dbd8352e38666f663199784cc38acbe23ca5bef0469d42aceedb8a951bde7502276a0c7b0a6f312e2c8b5cd282dd7bc2c7040d5d418035d62831c4ae7fa68bd1e8d8824b75719df97817d2ec3c57a7ddca075fd614e58127bc958da8e8f44d3;
    5'b00100 : xpb = 1024'h4152a81437ea9c4ed8f562ec1dfbd37c052bcac49c30cda3835c3e68e63f3358668f2ff0ebfbb46e4f02b4eec4818b64b90517f1fa51801fd907e117aeb70d85072e6f7ab1039a577d82f186029e88ea9494033f969df576f17ff5104c950020c3ba2f78643124faf26caf495d174144b68d530666fa01088d91f821e5c8e44b;
    5'b00101 : xpb = 1024'h257c00c3d569b6305c715db161643686aa193ca98ddf18ee84bc1fadb30e54ec7f60dc8ef47101e63aebd258bcca6a0b4e3fd3f4f0392c14e32209860bb033b9ebe63e2db160419c183d2d3edd0f3a18fcb7c5a95923e790807ccdd5b12f978468e6d6cc110b30164d57e163f669080b907a300f6ca5a9fe9f5a97693d0283c3;
    5'b00110 : xpb = 1024'h9a5597372e8d011dfed5876a4cc99914f06ae8e7f8d6439861c00f27fdd76809832892cfce64f5e26d4efc2b51348b1e37a8ff7e620d809ed3c31f468a959eed09e0ce0b1bce8e0b2f768f7b77feb4764db88131ba9d9aa0f79a69b15ca2ee80e137e1fbde53b31a843137e8fbaced26a670d18725152f4b12336b0943c233b;
    5'b00111 : xpb = 1024'h9e7bf778d2561ebc2e6ecb12f88f43ed656a23a446b34ffc05589b8cffaf451cb44cb343cf821b64b21c4c7390ba3822dccf73e0febb544aa7f599c10074f4d529a5104261aa8d6a604ba7532acc60a6c10444156ab5f8d45403115b348f68dde247b79d1b883eda89ee2c7820dcbbc2932dc903c848591b095b50fc7458291e;
    5'b01000 : xpb = 1024'h82a550286fd5389db1eac5d83bf7a6f80a57958938619b4706b87cd1cc7e66b0cd1e5fe1d7f768dc9e0569dd890316c9720a2fe3f4a3003fb20fc22f5d6e1b0a0e5cdef5620734aefb05e30c053d11d52928067f2d3beaede2ffea20992a004187745ef0c86249f5e4d95e92ba2e82896d1aa60ccdf402111b23f043cb91c896;
    5'b01001 : xpb = 1024'h66cea8d80d54527f3566c09d7f600a02af45076e2a0fe69208185e16994d8844e5f00c7fe06cb65489ee8747814bf5700744ebe6ea8aac34bc29ea9dba67413ef314ada86263dbf395c01ec4dfadc303914bc8e8efc1dd0771fcc2e5fdc497a52ca10644753c55113fc490ad5380495047078315d39fab072cec8f8b22cb680e;
    5'b01010 : xpb = 1024'h4af80187aad36c60b8e2bb62c2c86d0d543279531bbe31dd09783f5b661ca9d8fec1b91de8e203cc75d7a4b17994d4169c7fa7e9e0725829c644130c17606773d7cc7c5b62c08338307a5a7dba1e7431f96f8b52b247cf2100f99bab625f2f08d1cdad982216602c9aafc2c7ecd2101720f4601ed94b53fd3eb52ed27a050786;
    5'b01011 : xpb = 1024'h2f215a37485286423c5eb6280630d017f91feb380d6c7d280ad820a032ebcb6d179365bbf157514461c0c21b71ddb2bd31ba63ecd65a041ed05e3b7a74598da8bc844b0e631d2a7ccb349636948f256061934dbc74cdc13a8ff67470c6f9c66c76fa54ebcef06b47f59af4e28623d6ddfae13d27def6fcf3507dce19d13ea6fe;
    5'b01100 : xpb = 1024'h134ab2e6e5d1a023bfdab0ed499933229e0d5d1cff1ac8730c3801e4ffbaed0130651259f9cc9ebc4da9df856a269163c6f51fefcc41b013da7863e8d152b3dda13c19c16379d1c165eed1ef6effd68ec9b710263753b3541ef34d362b945dd01c26fc3f7bca7663508626fd1f759da4d4ce1a30e4a2a5e962466d6128784676;
    5'b01101 : xpb = 1024'ha82150ec453eeece0e5c23899d5bdd7eb470d232c640b4358b749c7f7f8cbb9d4c7f3c70cc686ac2d8f13c3645cd80d4c04a03d8e4dc2c549531cbb5691e4ec3fa431d231367764b1343104ae24c4bee25dfcc28865fd27e637cb7f64a5997c5f05b35bcd96d7a0c32313ff6b0978a94fd94d61c3a99ac0fba7e87ad08944c59;
    5'b01110 : xpb = 1024'h8c4aa99be2be08af91d81e4ee0c44089595e4417b7eeff808cd47dc44c5bdd316550e90ed4ddb83ac4da59a03e165f7b5584bfdbdac3d8499f4bf423c61774f8defaebd613c41d8fadfd4c03bcbcfd1c8e038e9248e5c497f27990bbaef42f299587dd10864785278d1c721149e9515bd781b32540455505cc4726f45fcdebd1;
    5'b01111 : xpb = 1024'h7074024b803d229115541914242ca393fe4bb5fca99d4acb8e345f09192afec57e2295acdd5305b2b0c3770a365f3e21eabf7bded0ab843ea9661c9223109b2dc3b2ba891420c4d448b787bc972dae4af62750fc0b6bb6b181766981138ec68d3ab4846433219042e807a42be33b1822b16e902e45f0fdfbde0fc63bb7078b49;
    5'b10000 : xpb = 1024'h549d5afb1dbc3c7298d013d96795069ea33927e19b4b96168f94404de5fa205996f4424ae5c8532a9cac94742ea81cc87ffa37e1c6933033b38045008009c162a86a893c147d6c18e371c375719e5f795e4b1365cdf1a8cb1073424678295df0dfe12bb7dffb9b5e42f2d6467c8cdee98b5b6d374b9ca6f1efd865830e412ac1;
    5'b10001 : xpb = 1024'h38c6b3aabb3b56541c4c0e9eaafd69a9482699c68cf9e16190f42192b2c941edafc5eee8ee3da0a28895b1de26f0fb6f1534f3e4bc7adc28bd9a6d6edd02e7978d2257ef14da135d7e2bff2e4c0f10a7c66ed5cf90779ae49f701b0bdcc3f554850dd30b8cd5a6799dde086115dea5b065484a4051484fe801a104ca657aca39;
    5'b10010 : xpb = 1024'h1cf00c5a58ba70359fc80963ee65ccb3ed140bab7ea82cac925402d77f986381c8979b86f6b2ee1a747ecf481f39da15aa6fafe7b262881dc7b495dd39fc0dcc71da26a21536baa218e63ae7267fc1d62e92983952fd8cfe2e6cf3d1415e8cb82a3a7a5f39afb194f8c93a7baf306c773f35274956f3f8de1369a411bcb469b1;
    5'b10011 : xpb = 1024'h1196509f6398a172344042931ce2fbe92017d90705677f793b3e41c4c678515e1694824ff283b926067ecb21782b8bc3faa6beaa84a3412d1cebe4b96f534015691f555159361e6b3a076a000f0730496b65aa315837f17bd69cc96a5f9241bcf6721b2e689bcb053b46c964882333e192204525c9fa1d42532435913ee0929;
    5'b10100 : xpb = 1024'h95f0030f55a6d8c171c576c58590da1aa864f2a6377c63ba12f07eb6cc3953b1fd83723bd1c40798ebaf4962f329a82d38ff4fd3c0e4b0538c8826182ec0cee7af98f8b6c581067060f4b4fb743ce863f2df16a5648f9e4201f33756c4be5e11a39b5b30442cc059355f858fd9a4202e41e8c03db296a7fa7d6a5da4f40a0f0c;
    5'b10101 : xpb = 1024'h7a195bbef325f2a2f541718ac8f93d254d52648b292aaf0514505ffb9908754616551ed9da395510d79866cceb7286d3ce3a0bd6b6cc5c4896a24e868bb9f51c9450c769c5ddadb4fbaef0b44ead99925b02d90f2715905b90f0101c2958f57548c80283f106cb74904ab7aa72f5e6f51bd59d46b84250f08f32fcec4b43ae84;
    5'b10110 : xpb = 1024'h5e42b46e90a50c8478bd6c500c61a02ff23fd6701ad8fa5015b0414065d796da2f26cb77e2aea288c3818436e3bb657a6374c7d9acb4083da0bc76f4e8b31b517908961cc63a54f996692c6d291e4ac0c3269b78e99b82751fece8e18df38cd8edf4a9d79de0d68feb35e9c50c47adbbf5c27a4fbdedf9e6a0fb9c33a27d4dfc;
    5'b10111 : xpb = 1024'h426c0d1e2e242665fc3967154fca033a972d48550c87459b1710228532a6b86e47f87815eb23f000af6aa1a0dc044420f8af83dca29bb432aad69f6345ac41865dc064cfc696fc3e31236826038efbef2b4a5de2ac21748eaee9c1a6f28e243c9321512b4abae1ab46211bdfa5997482cfaf5758c399a2dcb2c43b7af9b6ed74;
    5'b11000 : xpb = 1024'h269565cdcba340477fb561da933266453c1aba39fe3590e6187003c9ff75da0260ca24b3f3993d789b53bf0ad44d22c78dea3fdf98836027b4f0c7d1a2a567bb42783382c6f3a382cbdda3deddffad1d936e204c6ea766a83de69a6c5728bba0384df87ef794ecc6a10c4dfa3eeb3b49a99c3461c9454bd2c48cdac250f08cec;
    5'b11001 : xpb = 1024'habebe7d69225a2903315c9fd69ac94fe1082c1eefe3dc3119cfe50ecc44fb96799bd151fc0e8af0873cdc74cc96016e2324fbe28e6b0c1cbf0af03fff9e8df027300235c7504ac76697df97b8705e4bfb91e2b6312d58c1cce37331bbc35303dd7a9fd2a46ef7e1fbf78014d83d02108389116acef0f4c8d6557a09a82a2c64;
    5'b11010 : xpb = 1024'h9f955c82c88fa8d351b2cf3c2a5d73abf76ba134b709c7f3990c7fa94c16ca3295b5fb68ceaa56f712843925a83cf0df1c79dfcba705885d79c4580c976a28d680370597773def5113ec1df32bbcd3ab57ba9eb8803977ec116cddf1da888cf9b1aed9500211fb8adda2990e695eef00ac4fcd5624e7faef2e8d945588463247;
    5'b11011 : xpb = 1024'h83beb532660ec2b4d52eca016dc5d6b69c591319a8b8133e9a6c60ee18e5ebc6ae87a806d71fa46efe6d568fa085cf85b1b49bce9ced345283de807af4634f0b64eed44a779a9695aea659ac062d84d9bfde612242bf6a05a069b6b73f23245d56db80a3aeec06a6388dcb2902b0b5c7863caa5f2a93a3e54056339cdf7fd1bf;
    5'b11100 : xpb = 1024'h67e80de2038ddc9658aac4c6b12e39c1414684fe9a665e899bcc4232e5b50d5ac75954a4df94f1e6ea5673f998ceae2c46ef57d192d4e0478df8a8e9515c754049a6a2fd77f73dda49609564e09e36082802238c05455c1f2f668f7ca3bdbbc0fc0827f75bc611c19378fd439c027c8e60298768303f4cdb521ed2e436b97137;
    5'b11101 : xpb = 1024'h4c116691a10cf677dc26bf8bf4969ccbe633f6e38c14a9d49d2c2377b2842eeee02b0142e80a3f5ed63f916391178cd2dc2a13d488bc8c3c9812d157ae559b752e5e71b07853e51ee41ad11dbb0ee7369025e5f5c7cb4e38be63684208585324a134cf4b08a01cdcee642f5e355443553a16647135eaf5d163e7722b8df310af;
    5'b11110 : xpb = 1024'h303abf413e8c10595fa2ba5137feffd68b2168c87dc2f51f9e8c04bc7f535082f8fcade0f07f8cd6c228aecd89606b797164cfd77ea43831a22cf9c60b4ec1aa1316406378b08c637ed50cd6957f9864f849a85f8a5140524d6041076cf2ea884661769eb57a27f8494f6178cea60a1c1403417a3b969ec775b01172e52cb027;
    5'b11111 : xpb = 1024'h146417f0dc0b2a3ae31eb5167b6762e1300edaad6f71406a9febe6014c22721711ce5a7ef8f4da4eae11cc3781a94a20069f8bda748be426ac4722346847e7def7ce0f16790d33a8198f488f6ff04993606d6ac94cd7326bdc5d19ccd18d81ebeb8e1df262543313a43a939367f7d0e2edf01e83414247bd8778b0ba3c664f9f;
    endcase
end

endmodule

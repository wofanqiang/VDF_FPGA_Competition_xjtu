module xpb_5_40
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h344995ed4933391b103e5f2852b9a4d8adfae8a1d9ba1c2af9d169d320ef76325cfbc69e4026a91dd21e92ab2fef94c70b172d30d20a47692c8243dda0c98787d1f9a535f65dbb58d9016f1c9e99da79244d90cd3060d3a63de502d6cf4c64a44ec774d3d1360b497f023b558cd67358c09eb94b3cba0cbea869a5be923d6422;
    5'b00010 : xpb = 1024'h68932bda92667236207cbe50a57349b15bf5d143b3743855f3a2d3a641deec64b9f78d3c804d523ba43d25565fdf298e162e5a61a4148ed2590487bb41930f0fa3f34a6becbb76b1b202de393d33b4f2489b219a60c1a74c7bca05ad9e98c9489d8ee9a7a26c1692fe0476ab19ace6b1813d72967974197d50d34b7d247ac844;
    5'b00011 : xpb = 1024'h9cdcc1c7db99ab5130bb1d78f82cee8a09f0b9e58d2e5480ed743d7962ce629716f353dac073fb59765bb8018fcebe5521458792761ed63b8586cb98e25c969775ecefa1e319320a8b044d55dbcd8f6b6ce8b26791227af2b9af08846de52decec565e7b73a221dc7d06b200a6835a0a41dc2be1b62e263bf93cf13bb6b82c66;
    5'b00100 : xpb = 1024'h2079125f62deafa375f404ca3a8c4c1146759f569170d0346968edf6d0bb2bc170a69d00367425e8a91c0b65dc604251c8428cdd25764d590169d0184853a96dd397602929e5f01e516bb9cfe18ba5b39d31499c34fd2188420779608306efff0c164125940f3498754906773b89a739b3a1064aa29cd5ca5b371bf5c0132a1d;
    5'b00101 : xpb = 1024'h54c2a84cac11e8be863263f28d45f0e9f47087f86b2aec5f633a57c9f1aaa1f3cda2639e769acf067b3a9e110c4fd718d359ba0df78094c22dec13f5e91d30f5a591055f2043ab772a6d28ec8025802cc17eda69655df52e7fec7c37525354a35addb5f965453fe1f44b41ccc8601a92743fbf95df56e28903a0c1b452508e3f;
    5'b00110 : xpb = 1024'h890c3e39f54521d99670c31adfff95c2a26b709a44e5088a5d0bc19d129a18262a9e2a3cb6c178244d5930bc3c3f6bdfde70e73ec98adc2b5a6e57d389e6b87d778aaa9516a166d0036e98091ebf5aa5e5cc6b3695bec8d4bdd17f0e219fb947a9a52acd367b4b2b734d7d2255368deb34de78e11c10ef47ac0a6772e48df261;
    5'b00111 : xpb = 1024'hca88ed17c8a262bdba9aa6c225ef349def0560b4927843dd900721a8086e150845173622cc1a2b38019842088d0efdc856dec8978e25348d6515c52efddcb53d5351b1c5d6e24e3c9d60483247d70ee1615026b39996f6a4629efea36c17b59c9650d7756e85de76b8fd198ea3cdb1aa6a3534a087f9ed60e04922cede8f018;
    5'b01000 : xpb = 1024'h40f224bec5bd5f46ebe80994751898228ceb3ead22e1a068d2d1dbeda1765782e14d3a006ce84bd1523816cbb8c084a3908519ba4aec9ab202d3a03090a752dba72ec05253cbe03ca2d7739fc3174b673a62933869fa4310840ef2c1060ddffe182c824b281e6930ea920cee77134e7367420c954539ab94b66e37eb8026543a;
    5'b01001 : xpb = 1024'h753bbaac0ef09861fc2668bcc7d23cfb3ae6274efc9bbc93cca345c0c265cdb53e49009ead0ef4ef2456a976e8b0196a9b9c46eb1cf6e21b2f55e40e3170da63792865884a299b957bd8e2bc61b125e05eb024059a5b16b6c1f3f597d55a44a266f3f71ef954747a6994484403e9c1cc27e0c5e081f3b8535ed7ddaa1263b85c;
    5'b01010 : xpb = 1024'ha98550995823d17d0c64c7e51a8be1d3e8e10ff0d655d8bec674af93e35543e79b44c73ced359e0cf6753c22189fae31a6b3741bef0129845bd827ebd23a61eb4b220abe408756ee54da51d9004b005982fdb4d2cabbea5cffd8f86ea4a6a946b5bb6bf2ca8a7fc3e896839990c03524e87f7f2bbeadc51207418368a4a11c7e;
    5'b01011 : xpb = 1024'h2d21a130df68d5cf519daf365ceb3f5b2565f561da9854724269601151420d11f4f810626335c89c29358f866531322e4db079669e58a0a1d7bb2c6b383174c1a8cc7b45875415021b41be53060916a1b3464c076e9690f28831694ab9c86b58d57b4e9ceaf7927fe0d8d81025c682545a445994ab1c74a0693bae22adfc1a35;
    5'b01100 : xpb = 1024'h616b371e289c0eea61dc0e5eafa4e433d360de03b452709d3c3ac9e47231834451f3d700a35c71b9fb5422319520c6f558c7a6977062e80b043d7048d8fafc497ac6207b7db1d05af4432d6fa4a2f11ad793dcd49ef76498c6166c218914cffd2442c370bc2d9dc95fdb1365b29cf5ad1ae312dfe7d6815f11a553e140397e57;
    5'b01101 : xpb = 1024'h95b4cd0b71cf4805721a6d87025e890c815bc6a58e0c8cc8360c33b79320f976aeef9d9ee3831ad7cd72b4dcc5105bbc63ded3c8426d2f7430bfb42679c483d14cbfc5b1740f8bb3cd449c8c433ccb93fbe16da1cf58383f03fb6ef8586134a1730a38448d63a912dedd4ebb3f736905db81cc2b24908e1dba0ef99fd276e279;
    5'b01110 : xpb = 1024'h19511da2f9144c57b75354d844bde693bde0ac16924f087bb200e435010dc2a108a2e6c4598345670033084111a1dfb90adbd912f1c4a691aca2b8a5dfbb96a7aa6a3638badc49c793ac090648fae1dc2c2a04d67332ded48c53dfd46d82f6b392ca1aeeadd0bbced71fa331d479b6354d46a69410ff3dac1c092459dbd1e030;
    5'b01111 : xpb = 1024'h4d9ab39042478572c791b40097778b6c6bdb94b86c0924a6abd24e0821fd38d3659ead6299a9ee84d2519aec4191748015f30643c3ceedfad924fc8380851e2f7c63db6eb13a05206cad7822e794bc55507795a3a393b27aca38e2ab3ccf5b57e1918fc27f06c7185621de876150298e0de55fdf4db94a6ac472ca186e0f4452;
    5'b10000 : xpb = 1024'h81e4497d8b7abe8dd7d01328ea31304519d67d5a45c340d1a5a3b7db42ecaf05c29a7400d9d097a2a4702d9771810947210a337495d9356405a74061214ea5b74e5d80a4a797c07945aee73f862e96ce74c52670d3f48621081de5820c1bbffc30590496503cd261d52419dcee269ce6ce84192a8a7357296cdc6fd7004ca874;
    5'b10001 : xpb = 1024'h5809a1512bfc2e01d08fa7a2c908dcc565b62cb4a05bc8521986858b0d978301c4dbd264fd0c231d73080fbbe128d43c80738bf4530ac81818a44e08745b88dac07f12bee647e8d0c1653b98becad16a50dbda577cf2cb69076565e213d820e5018e74070a9e51dcd666e53832cea164048f39376e206b7ced69a9109a7a62b;
    5'b10010 : xpb = 1024'h39ca30025bf2fbfb2d4759a27f4a32a504564b6d23bfd8b01b69d22bd1c8ee62794983c48ff76b4fa94f13a6ee02220ad31e65f0173af3eaae0c88be280f40157e019661e4c239e5e517c2d62a86878fc95b4e72a830005cce5b5934f089e6b29ee05c1441dff0674c68a9a910035d6f00e7acdeb39c13767740404f9be50a4d;
    5'b10011 : xpb = 1024'h6e13c5efa52635163d85b8cad203d77db251340efd79f4db153b3bfef2b86494d6454a62d01e146d7b6da6521df1b6d1de359320e9453b53da8ecc9bc8d8c79d4ffb3b97db1ff53ebe1931f2c9206208eda8df3fd890d4030c405c0bbfd64b56eda7d0e81315fbb0cb6ae4fe9cd9d0c7c1866629f05620351fa9e60e2e226e6f;
    5'b10100 : xpb = 1024'ha25d5bdcee596e314dc417f324bd7c56604c1cb0d73411060f0ca5d213a7dac7334111011044bd8b4d8c38fd4de14b98e94cc051bb4f82bd0711107969a24f2521f4e0cdd17db097971aa10f67ba3c8211f6700d08f1a7a94a255ee28f22affb3c6f45bbe44c06fa4a6d205429b0442082251f752d102cf3c8138bccc05fd291;
    5'b10101 : xpb = 1024'h25f9ac74759e728392fcff44671cd9dd9cd10221db768cb98b01564f8194a3f18cf45a268644e81a804c8c619a72cf959049c59c6aa6f9da82f414f8cf9961fb7f9f5155184a6eab5d820d896d7852ca423f0741accc4e3ed27dcfbea444720d5c2f286604b919b642af74cabeb6914ff3e9f9de197edc822a0db686c9bad048;
    5'b10110 : xpb = 1024'h5a434261bed1ab9ea33b5e6cb9d67eb64acbeac3b530a8e484d2c022a2841a23e9f020c4c66b9138526b1f0cca62645c9b60f2cd3cb14143af7658d67062e9835198f68b0ea82a0436837ca60c122d43668c980edd2d21e51062d2957390d6b1aaf69d39d5ef24ffc1b1b0204b8d04a8b488b3295638e940d2775c455bf8346a;
    5'b10111 : xpb = 1024'h8e8cd84f0804e4b9b379bd950c90238ef8c6d3658eeac50f7ea429f5c373905646ebe76306923a562489b1b7fa51f923a6781ffe0ebb88acdbf89cb4112c710b23929bc10505e55d0f84ebc2aaac07bc8ada28dc0d8df58b4e47d56c42dd3b55f9be120da725304940b3eb75d863780175276c7492f2f5ff7ae10203ee35988c;
    5'b11000 : xpb = 1024'h122928e68f49e90bf8b2a4e64eef8116354bb8d6932d40c2fa98da7331605980a09f30887c9264e5574a051c46e37d204d752548be12ffca57dba133772383e1813d0c484bd2a370d5ec583cb06a1e04bb22c010b1689c20d6a0464857fefd68197df4b7c792430538f63fec6d69c530e6ec46dd7f61a58ddcdb2cbdf7909643;
    5'b11001 : xpb = 1024'h4672bed3d87d222708f1040ea1a925eee346a1786ce75cedf46a4446524fcfb2fd9af726bcb90e03296897c776d311e7588c5279901d4733845de51117ed0b695336b17e42305ec9aeedc7594f03f87ddf7050dde1c96fc71485491f274b620c6845698b98c84e4eb7f87b41fa403889a78b0028bc1bb24c8544d27c89cdfa65;
    5'b11010 : xpb = 1024'h7abc54c121b05b42192f6336f462cac791418a1a46a17918ee3bae19733f45e55a96bdc4fcdfb720fb872a72a6c2a6ae63a37faa62278e9cb0e028eeb8b692f1253056b4388e1a2287ef3675ed9dd2f703bde1ab122a436d526a4bf5f697c6b0b70cde5f69fe599836fab6978716abe26829b973f8d5bf0b2dae783b1c0b5e87;
    5'b11011 : xpb = 1024'haf05eaae6ae3945d296dc25f471c6fa03f3c72bc205b9543e80d17ec942ebc17b79284633d06603ecda5bd1dd6b23b756ebaacdb3431d605dd626ccc59801a78f729fbea2eebd57b60f0a5928c37ad70280b7278428b1713904f4eccc5e42b5505d453333b3464e1b5fcf1ed13ed1f3b28c872bf358fcbc9d6181df9ae48c2a9;
    5'b11100 : xpb = 1024'h32a23b45f22898af6ea6a9b0897bcd277bc1582d249e10f76401c86a021b85421145cd88b3068ace006610822343bf7215b7b225e3894d235945714bbf772d4f54d46c7175b8938f2758120c91f5c3b8585409ace665bda918a7bfa8db05ed67259435dd5ba1779dae3f4663a8f36c6a9a8d4d2821fe7b58381248b3b7a3c060;
    5'b11101 : xpb = 1024'h66ebd1333b5bd1ca7ee508d8dc35720029bc40cefe582d225dd3323d230afb746e419426f32d33ebd284a32d5333543920cedf56b593948c85c7b5296040b4d726ce11a76c164ee800598129308f9e317ca19a7a16c6914f568cc27faa52520b745baab12cd782e72d4181b935c9dfc35b2c06735eb88816e07bee7249e12482;
    5'b11110 : xpb = 1024'h9b356720848f0ae58f2368012eef16d8d7b72970d812494d57a49c1043fa71a6cb3d5ac53353dd09a4a335d88322e9002be60c87879ddbf5b249f907010a3c5ef8c7b6dd62740a40d95af045cf2978aaa0ef2b47472764f59471c556799eb6afc3231f84fe0d8e30ac43bd0ec2a0531c1bcabfbe9b7294d588e59430dc1e88a4;
    5'b11111 : xpb = 1024'h1ed1b7b80bd40f37d45c4f52714e7460143c0ee1dc54c500d3994c8db1e73ad124f0a3eaa9540798d763893ccfb46cfcd2e311d236f553132e2cfd8667014f3556722764a940c8549fc25cbfd4e78ef2d137c27beb020b8b1cca36328ec078c1e2e3022f1e7aa0eca486118557a6a04b8d8f9a2787e14463eadfbeeae579865b;
    endcase
end

endmodule

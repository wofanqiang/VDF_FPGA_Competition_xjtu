module xpb_5_225
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h789c737ca21fede86da3b5bd8613acdeb7fa3cc71d7ebf4b33d5eab3ca1fde310c16bf0091b8acf75f6da197ebd1f26b513021c38c0c7effdca19415eb72b20ad18cbc41efe9a940dbc4a1be80a9486cd516bafe3c0ff643cc8f8829f4301e0ef286bf94c861290ecbe683c0d54a70319ee943d7a60da770ad77ffbf74e16367;
    5'b00010 : xpb = 1024'h408ba1a38251a7081041f3a3fbcd126bfe7e765d6585de1ee9cf1c11e13d0f5a14e50088594adb601f7d03e8f445d40c3e461ba0f5662db408a3e8cd9c12ef642eca43d53042553ca4ef40da6876cca8b6287c63eb99bf76e3927e592e35998bb605ecffdff95990110d20a2b2c4ba39eef8a8ccfbcff1b11480847a60e06063;
    5'b00011 : xpb = 1024'h87acfca62836027b2e0318a718677f94502aff3ad8cfcf29fc84d6ff85a40831db3421020dd09c8df8c6639fcb9b5ad2b5c157e5ebfdc6834a63d854cb32cbd8c07cb68709b01386e19dff6504450e4973a3dc99b2388a9fa957488683b150879851a6af7918a115633bd84903f04423f080dc251923bf17b8909354cdf5d5f;
    5'b00100 : xpb = 1024'h8117434704a34e102083e747f79a24d7fcfcecbacb0bbc3dd39e3823c27a1eb429ca0110b295b6c03efa07d1e88ba8187c8c3741eacc5b681147d19b3825dec85d9487aa6084aa7949de81b4d0ed99516c50f8c7d7337eedc724fcb25c6b33176c0bd9ffbff2b320221a414565897473ddf15199f79fe362290108f4c1c0c0c6;
    5'b00101 : xpb = 1024'h4906716de4d5072fc322252e6d538a65438126511312db1189976981d9974fdd329842987a27e528ff096a22f0ff89b969a2311f54260a1c3d4a2652e8c61c21bad20f3da0dd5675130920d0b8bb1d8d4d62ba2d86bd4820de27f2e19670ae942f8b076ad78ae3a16740de274303be7c2e00b68f4d622da290098dafadbfbdc2;
    5'b00110 : xpb = 1024'h10f59f94c506c04f65c06314e30ceff28a055fe75b19f9e53f909adff0b481063b66842041ba1391bf18cc73f9736b5a56b82afcbd7fb8d0694c7b0a9966597b180f96d0e1360270dc33bfeca088a1c92e747b9336471153f52ae910d0762a10f30a34d5ef231422ac677b09207e08847e101b84a32477e2f712126a99bebabe;
    5'b00111 : xpb = 1024'h899213116726ae37d36418d269209cd141ff9cae7898b93073668593bad45f37477d4320d372c0891e866e0be5455dc5a7e84cc0498c37d045ee0f2084d90b85e99c5312d11fabb1b7f861ab2131ea36038b369172570797c1ba713ac4a6481fe590f46ab7843d31784dfec9f5c878b61cf95f5c49321f53a48a122a0ea01e25;
    5'b01000 : xpb = 1024'h5181413847586757760256b8deda025e8883d644c09fd804295fb6f1d1f19060504b84a89b04eef1de95d05cedb93f6694fe469db2e5e68471f063d8357948df46d9daa6117857ad812300c708ff6e71e49cf7f721e0d0cad8bd6769feabc39ca91021d5cf1c6db2bd749babd342c2be6d08c4519ef469940b9296e4fa9f1b21;
    5'b01001 : xpb = 1024'h19706f5f278a207718a0949f549367ebcf080fdb08a6f6d7df58e84fe90ec1895919c63062971d5a9ea532adf62d21078214407b1c3f95389df2b88fe6198638a417623951d103a94a4d9fe2f0ccf2adc5aeb95cd16a99fdefc05d9938b13f196c8f4f40e6b49e34029b388db0bd0cc6bd182946f4b6b3d4729b1b9fe69e181d;
    5'b01010 : xpb = 1024'h920ce2dbc9aa0e5f86444a5cdaa714ca87024ca22625b623132ed303b32e9fba65308530f44fca51fe12d445e1ff1372d344623ea84c14387a944ca5d18c384375a41e7b41baacea261241a171763b1a9ac5745b0d7a9041bc4fe5c32ce15d285f160ed5af15c742ce81bc4e86077cf85c016d1e9ac45b4520131b5f5b7f7b84;
    5'b01011 : xpb = 1024'h59fc1102a9dbc77f28e2884350607a57cd8686386e2cd4f6c9280461ca4bd0e36dfec6b8bbe1f8babe223696ea72f513c05a5c1c11a5c2eca696a15d822c759cd2e1a60e821358e5ef3ce0bd5943bf567bd735c0bd045974d352dbf266e6d8a522953c40c6adf7c413a859306381c700ac10d213f086a585871ba01a477e7880;
    5'b01100 : xpb = 1024'h21eb3f298a0d809ecb80c629c619dfe5140abfceb633f3ca7f2135bfe169020c76cd0840837427237e3198e7f2e6d6b4ad7055f97aff71a0d298f61532ccb2f6301f2da1c26c04e1b8677fd9411143925ce8f7266c8e22a7ea55d221a0ec5421e61469abde46284558cef61240fc1108fc2037094648efc5ee2424d5337d757c;
    5'b01101 : xpb = 1024'h9a87b2a62c2d6e8739247be74c2d8cc3cc04fc95d3b2b315b2f72073ab88e03d82e3c741152cd41add9f3a7fdeb8c91ffea077bd070bf0a0af3a8a2b1e3f650101abe9e3b255ae22942c2197c1ba8bff31ffb224a89e18ebb6e55a4b951c7230d89b2940a6a7515424b579d31646813a9b097ae0ec5697369b9c2494a85ed8e3;
    5'b01110 : xpb = 1024'h6276e0cd0c5f27a6dbc2b9cdc1e6f2511289362c1bb9d1e968f051d1c2a611668bb208c8dcbf02839dae9cd0e72caac0ebb6719a70659f54db3cdee2cedfa25a5ee97176f2ae5a1e5d56c0b3a988103b1311738a5827e21ecde8507acf21edad9c1a56abbe3f81d569dc16b4f3c0cb42eb18dfd64218e17702a4a94f945dd5df;
    5'b01111 : xpb = 1024'h2a660ef3ec90e0c67e60f7b437a057de590d6fc263c0f0bd1ee9832fd9c3428f94804a50a45130ec5dbdff21efa08c61d8cc6b77d9bf4e09073f339a7f7fdfb3bc26f90a3307061a26815fcf91559476f42334f007b1ab51e4eb46aa0927692a5f998416d5d7b256af02b396d13b154b3b2844cb97db2bb769ad2e0a805cd2db;
    5'b10000 : xpb = 1024'ha30282708eb0ceaeec04ad71bdb404bd1107ac89813fb00852bf6de3a3e320c0a09709513609dde3bd2ba0b9db727ecd29fc8d3b65cbcd08e3e0c7b06af291be8db3b54c22f0af5b0246018e11fedce3c939efee43c1a195b17aced3fd578739522043ab9e38db657ae93757a685857cda1188a33de8d32817252dc9f53e3642;
    5'b10001 : xpb = 1024'h6af1b0976ee287ce8ea2eb58336d6a4a578be61fc946cedc08b89f41bb0051e9a9654ad8fd9c0c4c7d3b030ae3e6606e17128718cf257bbd0fe31c681b92cf17eaf13cdf63495b56cb70a0a9f9cc611faa4bb153f34b6ac8c87dc503375d02b6159f7116b5d10be6c00fd43983ffcf852a20ed9893ab1d687e2db284e13d333e;
    5'b10010 : xpb = 1024'h32e0debe4f1440ee3141293ea926cfd79e101fb6114dedafbeb1d09fd21d8312b2338c60c52e3ab53d4a655bec5a420f042880f6387f2a713be5711fcc330c71482ec472a3a20752949b3fc5e199e55b8b5d72b9a2d533fbdf80bb3271627e32d91e9e81cd693c680536711b617a198d7a30528de96d67a8e536373fcd3c303a;
    5'b10011 : xpb = 1024'hab7d523af1342ed69ee4defc2f3a7cb6560a5c7d2eccacfaf287bb539c3d6143be4a4b6156e6e7ac9cb806f3d82c347a5558a2b9c48ba97118870535b7a5be7c19bb80b4938bb093705fe18462432dc860742db7dee52a3fac10435c65929c41cba55e1695ca6576d11cf4dc36c489bf191996658f7b0f1992ae36ff421d93a1;
    5'b10100 : xpb = 1024'h736c8061d165e7f641831ce2a4f3e2439c8e961376d3cbcea880ecb1b35a926cc7188ce91e7916155cc76944e0a0161b426e9c972de55825448959ed6845fbd576f90847d3e45c8f398a80a04a10b2044185ef1d8e6ef372c313398b9f9817be8f248b81ad6295f8164391be143ed3c76928fb5ae53d5959f9b6bbba2e1c909d;
    5'b10101 : xpb = 1024'h3b5bae88b197a115e4215ac91aad47d0e312cfa9bedaeaa25e7a1e0fca77c395cfe6ce70e60b447e1cd6cb95e913f7bc2f849674973f06d9708baea518e6392ed4368fdb143d088b02b51fbc31de36402297b0833df8bca5da162fbad99d933b52a3b8ecc4fac6795b6a2e9ff1b91dcfb93860503affa39a60bf40751a1b8d99;
    5'b10110 : xpb = 1024'h34adcaf91c95a3586bf98af9066ad5e2997094006e2097614734f6de194f4bed8b50ff8ad9d72e6dce62de6f187d95d1c9a90520098b58d9c8e035cc98676883174176e5495b486cbdfbed819abba7c03a971e8ed8285d8f11925ea13a30eb81622e657dc92f6faa090cb81cf3367d80947c54590c1eddac7c7c530061a8a95;
    5'b10111 : xpb = 1024'h7be7502c33e9481df4634e6d167a5a3ce19146072460c8c148493a21abb4d2efe4cbcef93f561fde3c53cf7edd59cbc86dcab2158ca5348d792f9772b4f928930300d3b0447f5dc7a7a460969a5502e8d8c02ce729927c1cbda8ae1407d32cc708a9a5eca4f420096c774f42a47dd809a831091d36cf954b753fc4ef7afbedfc;
    5'b11000 : xpb = 1024'h43d67e53141b013d97018c538c33bfca28157f9d6c67e794fe426b7fc2d20418ed9a108106e84e46fc6331cfe5cdad695ae0abf2f5fee341a531ec2a659965ec603e5b4384d809c370ceffb282228724b9d1ee4cd91c454fd4aba44341d8a843cc28d357bc8c508ab19dec2481f82211f8406e128c91df8bdc4849aa66faeaf8;
    5'b11001 : xpb = 1024'hbc5ac79f44cba5d399fca3a01ed25576e99b933b46f0668b43b9cddd9ef3541f6685208ce7a7cafbc729420ee418f0a47f6a5d05f5891f5d13440e21639a345bd7be2d6c530b5bf39f99ece69f00b609ae3afb288a60e82ebae9a727bde23c08fa800c2d424810bf6c489065f726c1a484fd307e25429cc4350ce6552f9e7f4;
    5'b11010 : xpb = 1024'h84621ff6966ca845a7437ff78800d2362693f5fad1edc5b3e8118791a40f1373027f1109603329a71be035b8da1381759926c793eb6510f5add5d4f801ac55508f089f18b51a5f0015be408cea9953cd6ffa6ab0c4b604c6b83e229c700e41cf822ec0579c85aa1ac2ab0cc734bcdc4be73916df8861d13cf0c8ce24c7db4b5b;
    5'b11011 : xpb = 1024'h4c514e1d769e616549e1bdddfdba37c36d182f9119f4e4879e0ab8efbb2c449c0b4d529127c5580fdbef9809e2876316863cc17154bebfa9d9d829afb24c92a9ec4626abf5730afbdee8dfa8d266d809510c2c16743fcdf9cf4118cbaa13bd4c45adedc2b41dda9c07d1a9a91237265437487bd4de241b7d57d152dfb3da4857;
    5'b11100 : xpb = 1024'h14407c4456d01a84ec7ffbc473739d50b39c692761fc035b5403ea4dd24975c5141b9418ef5786789bfefa5aeafb44b77352bb4ebe186e5e05da7e6762ecd0034983ae3f35cbb6f7a8137ec4ba345c45321ded7c23c9972ce6440efae41938c9092d1b2dcbb60b1d4cf8468aefb1705c8757e0ca33e665bdbed9d79a9fd94553;
    5'b11101 : xpb = 1024'h8cdcefc0f8f0086d5a23b181f9874a2f6b96a5ee7f7ac2a687d9d5019c6953f6203253198110336ffb6c9bf2d6cd3722c482dd124a24ed5de27c127d4e5f820e1b106a8125b5603883d820833adda4b20734a87a5fd98d70b2d39724d84956d7fbb3dac29417342c18deca4bc4fbe08e264124a1d9f40d2e6c51d75a14baa8ba;
    5'b11110 : xpb = 1024'h54cc1de7d921c18cfcc1ef686f40afbcb21adf84c781e17a3dd3065fb386851f290094a148a261d8bb7bfe43df4118c3b198d6efb37e9c120e7e6734feffbf67784df214660e0c344d02bf9f22ab28ede84669e00f6356a3c9d68d54124ed254bf33082dabaf64ad5e05672da2762a96765089972fb6576ed35a5c1500b9a5b6;
    5'b11111 : xpb = 1024'h1cbb4c0eb9537aac9f602d4ee4fa1549f89f191b0f89004df3cc37bdcaa3b64831ced629103490417b8b6094e7b4fa649eaed0cd1cd84ac63a80bbecaf9ffcc0d58b79a7a666b830162d5ebb0a78ad29c9582b45beed1fd6e0d983834c544dd182b23598c347952ea32c040f7ff0749ec65fee8c8578a1af3a62e0cfecb8a2b2;
    endcase
end

endmodule

module compressor_array_512_152_1024
(
    input  [511:0] col_in_0,
    input  [511:0] col_in_1,
    input  [511:0] col_in_2,
    input  [511:0] col_in_3,
    input  [511:0] col_in_4,
    input  [511:0] col_in_5,
    input  [511:0] col_in_6,
    input  [511:0] col_in_7,
    input  [511:0] col_in_8,
    input  [511:0] col_in_9,
    input  [511:0] col_in_10,
    input  [511:0] col_in_11,
    input  [511:0] col_in_12,
    input  [511:0] col_in_13,
    input  [511:0] col_in_14,
    input  [511:0] col_in_15,
    input  [511:0] col_in_16,
    input  [511:0] col_in_17,
    input  [511:0] col_in_18,
    input  [511:0] col_in_19,
    input  [511:0] col_in_20,
    input  [511:0] col_in_21,
    input  [511:0] col_in_22,
    input  [511:0] col_in_23,
    input  [511:0] col_in_24,
    input  [511:0] col_in_25,
    input  [511:0] col_in_26,
    input  [511:0] col_in_27,
    input  [511:0] col_in_28,
    input  [511:0] col_in_29,
    input  [511:0] col_in_30,
    input  [511:0] col_in_31,
    input  [511:0] col_in_32,
    input  [511:0] col_in_33,
    input  [511:0] col_in_34,
    input  [511:0] col_in_35,
    input  [511:0] col_in_36,
    input  [511:0] col_in_37,
    input  [511:0] col_in_38,
    input  [511:0] col_in_39,
    input  [511:0] col_in_40,
    input  [511:0] col_in_41,
    input  [511:0] col_in_42,
    input  [511:0] col_in_43,
    input  [511:0] col_in_44,
    input  [511:0] col_in_45,
    input  [511:0] col_in_46,
    input  [511:0] col_in_47,
    input  [511:0] col_in_48,
    input  [511:0] col_in_49,
    input  [511:0] col_in_50,
    input  [511:0] col_in_51,
    input  [511:0] col_in_52,
    input  [511:0] col_in_53,
    input  [511:0] col_in_54,
    input  [511:0] col_in_55,
    input  [511:0] col_in_56,
    input  [511:0] col_in_57,
    input  [511:0] col_in_58,
    input  [511:0] col_in_59,
    input  [511:0] col_in_60,
    input  [511:0] col_in_61,
    input  [511:0] col_in_62,
    input  [511:0] col_in_63,
    input  [511:0] col_in_64,
    input  [511:0] col_in_65,
    input  [511:0] col_in_66,
    input  [511:0] col_in_67,
    input  [511:0] col_in_68,
    input  [511:0] col_in_69,
    input  [511:0] col_in_70,
    input  [511:0] col_in_71,
    input  [511:0] col_in_72,
    input  [511:0] col_in_73,
    input  [511:0] col_in_74,
    input  [511:0] col_in_75,
    input  [511:0] col_in_76,
    input  [511:0] col_in_77,
    input  [511:0] col_in_78,
    input  [511:0] col_in_79,
    input  [511:0] col_in_80,
    input  [511:0] col_in_81,
    input  [511:0] col_in_82,
    input  [511:0] col_in_83,
    input  [511:0] col_in_84,
    input  [511:0] col_in_85,
    input  [511:0] col_in_86,
    input  [511:0] col_in_87,
    input  [511:0] col_in_88,
    input  [511:0] col_in_89,
    input  [511:0] col_in_90,
    input  [511:0] col_in_91,
    input  [511:0] col_in_92,
    input  [511:0] col_in_93,
    input  [511:0] col_in_94,
    input  [511:0] col_in_95,
    input  [511:0] col_in_96,
    input  [511:0] col_in_97,
    input  [511:0] col_in_98,
    input  [511:0] col_in_99,
    input  [511:0] col_in_100,
    input  [511:0] col_in_101,
    input  [511:0] col_in_102,
    input  [511:0] col_in_103,
    input  [511:0] col_in_104,
    input  [511:0] col_in_105,
    input  [511:0] col_in_106,
    input  [511:0] col_in_107,
    input  [511:0] col_in_108,
    input  [511:0] col_in_109,
    input  [511:0] col_in_110,
    input  [511:0] col_in_111,
    input  [511:0] col_in_112,
    input  [511:0] col_in_113,
    input  [511:0] col_in_114,
    input  [511:0] col_in_115,
    input  [511:0] col_in_116,
    input  [511:0] col_in_117,
    input  [511:0] col_in_118,
    input  [511:0] col_in_119,
    input  [511:0] col_in_120,
    input  [511:0] col_in_121,
    input  [511:0] col_in_122,
    input  [511:0] col_in_123,
    input  [511:0] col_in_124,
    input  [511:0] col_in_125,
    input  [511:0] col_in_126,
    input  [511:0] col_in_127,
    input  [511:0] col_in_128,
    input  [511:0] col_in_129,
    input  [511:0] col_in_130,
    input  [511:0] col_in_131,
    input  [511:0] col_in_132,
    input  [511:0] col_in_133,
    input  [511:0] col_in_134,
    input  [511:0] col_in_135,
    input  [511:0] col_in_136,
    input  [511:0] col_in_137,
    input  [511:0] col_in_138,
    input  [511:0] col_in_139,
    input  [511:0] col_in_140,
    input  [511:0] col_in_141,
    input  [511:0] col_in_142,
    input  [511:0] col_in_143,
    input  [511:0] col_in_144,
    input  [511:0] col_in_145,
    input  [511:0] col_in_146,
    input  [511:0] col_in_147,
    input  [511:0] col_in_148,
    input  [511:0] col_in_149,
    input  [511:0] col_in_150,
    input  [511:0] col_in_151,
    input  [511:0] col_in_152,
    input  [511:0] col_in_153,
    input  [511:0] col_in_154,
    input  [511:0] col_in_155,
    input  [511:0] col_in_156,
    input  [511:0] col_in_157,
    input  [511:0] col_in_158,
    input  [511:0] col_in_159,
    input  [511:0] col_in_160,
    input  [511:0] col_in_161,
    input  [511:0] col_in_162,
    input  [511:0] col_in_163,
    input  [511:0] col_in_164,
    input  [511:0] col_in_165,
    input  [511:0] col_in_166,
    input  [511:0] col_in_167,
    input  [511:0] col_in_168,
    input  [511:0] col_in_169,
    input  [511:0] col_in_170,
    input  [511:0] col_in_171,
    input  [511:0] col_in_172,
    input  [511:0] col_in_173,
    input  [511:0] col_in_174,
    input  [511:0] col_in_175,
    input  [511:0] col_in_176,
    input  [511:0] col_in_177,
    input  [511:0] col_in_178,
    input  [511:0] col_in_179,
    input  [511:0] col_in_180,
    input  [511:0] col_in_181,
    input  [511:0] col_in_182,
    input  [511:0] col_in_183,
    input  [511:0] col_in_184,
    input  [511:0] col_in_185,
    input  [511:0] col_in_186,
    input  [511:0] col_in_187,
    input  [511:0] col_in_188,
    input  [511:0] col_in_189,
    input  [511:0] col_in_190,
    input  [511:0] col_in_191,
    input  [511:0] col_in_192,
    input  [511:0] col_in_193,
    input  [511:0] col_in_194,
    input  [511:0] col_in_195,
    input  [511:0] col_in_196,
    input  [511:0] col_in_197,
    input  [511:0] col_in_198,
    input  [511:0] col_in_199,
    input  [511:0] col_in_200,
    input  [511:0] col_in_201,
    input  [511:0] col_in_202,
    input  [511:0] col_in_203,
    input  [511:0] col_in_204,
    input  [511:0] col_in_205,
    input  [511:0] col_in_206,
    input  [511:0] col_in_207,
    input  [511:0] col_in_208,
    input  [511:0] col_in_209,
    input  [511:0] col_in_210,
    input  [511:0] col_in_211,
    input  [511:0] col_in_212,
    input  [511:0] col_in_213,
    input  [511:0] col_in_214,
    input  [511:0] col_in_215,
    input  [511:0] col_in_216,
    input  [511:0] col_in_217,
    input  [511:0] col_in_218,
    input  [511:0] col_in_219,
    input  [511:0] col_in_220,
    input  [511:0] col_in_221,
    input  [511:0] col_in_222,
    input  [511:0] col_in_223,
    input  [511:0] col_in_224,
    input  [511:0] col_in_225,
    input  [511:0] col_in_226,
    input  [511:0] col_in_227,
    input  [511:0] col_in_228,
    input  [511:0] col_in_229,
    input  [511:0] col_in_230,
    input  [511:0] col_in_231,
    input  [511:0] col_in_232,
    input  [511:0] col_in_233,
    input  [511:0] col_in_234,
    input  [511:0] col_in_235,
    input  [511:0] col_in_236,
    input  [511:0] col_in_237,
    input  [511:0] col_in_238,
    input  [511:0] col_in_239,
    input  [511:0] col_in_240,
    input  [511:0] col_in_241,
    input  [511:0] col_in_242,
    input  [511:0] col_in_243,
    input  [511:0] col_in_244,
    input  [511:0] col_in_245,
    input  [511:0] col_in_246,
    input  [511:0] col_in_247,
    input  [511:0] col_in_248,
    input  [511:0] col_in_249,
    input  [511:0] col_in_250,
    input  [511:0] col_in_251,
    input  [511:0] col_in_252,
    input  [511:0] col_in_253,
    input  [511:0] col_in_254,
    input  [511:0] col_in_255,
    input  [511:0] col_in_256,
    input  [511:0] col_in_257,
    input  [511:0] col_in_258,
    input  [511:0] col_in_259,
    input  [511:0] col_in_260,
    input  [511:0] col_in_261,
    input  [511:0] col_in_262,
    input  [511:0] col_in_263,
    input  [511:0] col_in_264,
    input  [511:0] col_in_265,
    input  [511:0] col_in_266,
    input  [511:0] col_in_267,
    input  [511:0] col_in_268,
    input  [511:0] col_in_269,
    input  [511:0] col_in_270,
    input  [511:0] col_in_271,
    input  [511:0] col_in_272,
    input  [511:0] col_in_273,
    input  [511:0] col_in_274,
    input  [511:0] col_in_275,
    input  [511:0] col_in_276,
    input  [511:0] col_in_277,
    input  [511:0] col_in_278,
    input  [511:0] col_in_279,
    input  [511:0] col_in_280,
    input  [511:0] col_in_281,
    input  [511:0] col_in_282,
    input  [511:0] col_in_283,
    input  [511:0] col_in_284,
    input  [511:0] col_in_285,
    input  [511:0] col_in_286,
    input  [511:0] col_in_287,
    input  [511:0] col_in_288,
    input  [511:0] col_in_289,
    input  [511:0] col_in_290,
    input  [511:0] col_in_291,
    input  [511:0] col_in_292,
    input  [511:0] col_in_293,
    input  [511:0] col_in_294,
    input  [511:0] col_in_295,
    input  [511:0] col_in_296,
    input  [511:0] col_in_297,
    input  [511:0] col_in_298,
    input  [511:0] col_in_299,
    input  [511:0] col_in_300,
    input  [511:0] col_in_301,
    input  [511:0] col_in_302,
    input  [511:0] col_in_303,
    input  [511:0] col_in_304,
    input  [511:0] col_in_305,
    input  [511:0] col_in_306,
    input  [511:0] col_in_307,
    input  [511:0] col_in_308,
    input  [511:0] col_in_309,
    input  [511:0] col_in_310,
    input  [511:0] col_in_311,
    input  [511:0] col_in_312,
    input  [511:0] col_in_313,
    input  [511:0] col_in_314,
    input  [511:0] col_in_315,
    input  [511:0] col_in_316,
    input  [511:0] col_in_317,
    input  [511:0] col_in_318,
    input  [511:0] col_in_319,
    input  [511:0] col_in_320,
    input  [511:0] col_in_321,
    input  [511:0] col_in_322,
    input  [511:0] col_in_323,
    input  [511:0] col_in_324,
    input  [511:0] col_in_325,
    input  [511:0] col_in_326,
    input  [511:0] col_in_327,
    input  [511:0] col_in_328,
    input  [511:0] col_in_329,
    input  [511:0] col_in_330,
    input  [511:0] col_in_331,
    input  [511:0] col_in_332,
    input  [511:0] col_in_333,
    input  [511:0] col_in_334,
    input  [511:0] col_in_335,
    input  [511:0] col_in_336,
    input  [511:0] col_in_337,
    input  [511:0] col_in_338,
    input  [511:0] col_in_339,
    input  [511:0] col_in_340,
    input  [511:0] col_in_341,
    input  [511:0] col_in_342,
    input  [511:0] col_in_343,
    input  [511:0] col_in_344,
    input  [511:0] col_in_345,
    input  [511:0] col_in_346,
    input  [511:0] col_in_347,
    input  [511:0] col_in_348,
    input  [511:0] col_in_349,
    input  [511:0] col_in_350,
    input  [511:0] col_in_351,
    input  [511:0] col_in_352,
    input  [511:0] col_in_353,
    input  [511:0] col_in_354,
    input  [511:0] col_in_355,
    input  [511:0] col_in_356,
    input  [511:0] col_in_357,
    input  [511:0] col_in_358,
    input  [511:0] col_in_359,
    input  [511:0] col_in_360,
    input  [511:0] col_in_361,
    input  [511:0] col_in_362,
    input  [511:0] col_in_363,
    input  [511:0] col_in_364,
    input  [511:0] col_in_365,
    input  [511:0] col_in_366,
    input  [511:0] col_in_367,
    input  [511:0] col_in_368,
    input  [511:0] col_in_369,
    input  [511:0] col_in_370,
    input  [511:0] col_in_371,
    input  [511:0] col_in_372,
    input  [511:0] col_in_373,
    input  [511:0] col_in_374,
    input  [511:0] col_in_375,
    input  [511:0] col_in_376,
    input  [511:0] col_in_377,
    input  [511:0] col_in_378,
    input  [511:0] col_in_379,
    input  [511:0] col_in_380,
    input  [511:0] col_in_381,
    input  [511:0] col_in_382,
    input  [511:0] col_in_383,
    input  [511:0] col_in_384,
    input  [511:0] col_in_385,
    input  [511:0] col_in_386,
    input  [511:0] col_in_387,
    input  [511:0] col_in_388,
    input  [511:0] col_in_389,
    input  [511:0] col_in_390,
    input  [511:0] col_in_391,
    input  [511:0] col_in_392,
    input  [511:0] col_in_393,
    input  [511:0] col_in_394,
    input  [511:0] col_in_395,
    input  [511:0] col_in_396,
    input  [511:0] col_in_397,
    input  [511:0] col_in_398,
    input  [511:0] col_in_399,
    input  [511:0] col_in_400,
    input  [511:0] col_in_401,
    input  [511:0] col_in_402,
    input  [511:0] col_in_403,
    input  [511:0] col_in_404,
    input  [511:0] col_in_405,
    input  [511:0] col_in_406,
    input  [511:0] col_in_407,
    input  [511:0] col_in_408,
    input  [511:0] col_in_409,
    input  [511:0] col_in_410,
    input  [511:0] col_in_411,
    input  [511:0] col_in_412,
    input  [511:0] col_in_413,
    input  [511:0] col_in_414,
    input  [511:0] col_in_415,
    input  [511:0] col_in_416,
    input  [511:0] col_in_417,
    input  [511:0] col_in_418,
    input  [511:0] col_in_419,
    input  [511:0] col_in_420,
    input  [511:0] col_in_421,
    input  [511:0] col_in_422,
    input  [511:0] col_in_423,
    input  [511:0] col_in_424,
    input  [511:0] col_in_425,
    input  [511:0] col_in_426,
    input  [511:0] col_in_427,
    input  [511:0] col_in_428,
    input  [511:0] col_in_429,
    input  [511:0] col_in_430,
    input  [511:0] col_in_431,
    input  [511:0] col_in_432,
    input  [511:0] col_in_433,
    input  [511:0] col_in_434,
    input  [511:0] col_in_435,
    input  [511:0] col_in_436,
    input  [511:0] col_in_437,
    input  [511:0] col_in_438,
    input  [511:0] col_in_439,
    input  [511:0] col_in_440,
    input  [511:0] col_in_441,
    input  [511:0] col_in_442,
    input  [511:0] col_in_443,
    input  [511:0] col_in_444,
    input  [511:0] col_in_445,
    input  [511:0] col_in_446,
    input  [511:0] col_in_447,
    input  [511:0] col_in_448,
    input  [511:0] col_in_449,
    input  [511:0] col_in_450,
    input  [511:0] col_in_451,
    input  [511:0] col_in_452,
    input  [511:0] col_in_453,
    input  [511:0] col_in_454,
    input  [511:0] col_in_455,
    input  [511:0] col_in_456,
    input  [511:0] col_in_457,
    input  [511:0] col_in_458,
    input  [511:0] col_in_459,
    input  [511:0] col_in_460,
    input  [511:0] col_in_461,
    input  [511:0] col_in_462,
    input  [511:0] col_in_463,
    input  [511:0] col_in_464,
    input  [511:0] col_in_465,
    input  [511:0] col_in_466,
    input  [511:0] col_in_467,
    input  [511:0] col_in_468,
    input  [511:0] col_in_469,
    input  [511:0] col_in_470,
    input  [511:0] col_in_471,
    input  [511:0] col_in_472,
    input  [511:0] col_in_473,
    input  [511:0] col_in_474,
    input  [511:0] col_in_475,
    input  [511:0] col_in_476,
    input  [511:0] col_in_477,
    input  [511:0] col_in_478,
    input  [511:0] col_in_479,
    input  [511:0] col_in_480,
    input  [511:0] col_in_481,
    input  [511:0] col_in_482,
    input  [511:0] col_in_483,
    input  [511:0] col_in_484,
    input  [511:0] col_in_485,
    input  [511:0] col_in_486,
    input  [511:0] col_in_487,
    input  [511:0] col_in_488,
    input  [511:0] col_in_489,
    input  [511:0] col_in_490,
    input  [511:0] col_in_491,
    input  [511:0] col_in_492,
    input  [511:0] col_in_493,
    input  [511:0] col_in_494,
    input  [511:0] col_in_495,
    input  [511:0] col_in_496,
    input  [511:0] col_in_497,
    input  [511:0] col_in_498,
    input  [511:0] col_in_499,
    input  [511:0] col_in_500,
    input  [511:0] col_in_501,
    input  [511:0] col_in_502,
    input  [511:0] col_in_503,
    input  [511:0] col_in_504,
    input  [511:0] col_in_505,
    input  [511:0] col_in_506,
    input  [511:0] col_in_507,
    input  [511:0] col_in_508,
    input  [511:0] col_in_509,
    input  [511:0] col_in_510,
    input  [511:0] col_in_511,
    input  [511:0] col_in_512,
    input  [511:0] col_in_513,
    input  [511:0] col_in_514,
    input  [511:0] col_in_515,
    input  [511:0] col_in_516,
    input  [511:0] col_in_517,
    input  [511:0] col_in_518,
    input  [511:0] col_in_519,
    input  [511:0] col_in_520,
    input  [511:0] col_in_521,
    input  [511:0] col_in_522,
    input  [511:0] col_in_523,
    input  [511:0] col_in_524,
    input  [511:0] col_in_525,
    input  [511:0] col_in_526,
    input  [511:0] col_in_527,
    input  [511:0] col_in_528,
    input  [511:0] col_in_529,
    input  [511:0] col_in_530,
    input  [511:0] col_in_531,
    input  [511:0] col_in_532,
    input  [511:0] col_in_533,
    input  [511:0] col_in_534,
    input  [511:0] col_in_535,
    input  [511:0] col_in_536,
    input  [511:0] col_in_537,
    input  [511:0] col_in_538,
    input  [511:0] col_in_539,
    input  [511:0] col_in_540,
    input  [511:0] col_in_541,
    input  [511:0] col_in_542,
    input  [511:0] col_in_543,
    input  [511:0] col_in_544,
    input  [511:0] col_in_545,
    input  [511:0] col_in_546,
    input  [511:0] col_in_547,
    input  [511:0] col_in_548,
    input  [511:0] col_in_549,
    input  [511:0] col_in_550,
    input  [511:0] col_in_551,
    input  [511:0] col_in_552,
    input  [511:0] col_in_553,
    input  [511:0] col_in_554,
    input  [511:0] col_in_555,
    input  [511:0] col_in_556,
    input  [511:0] col_in_557,
    input  [511:0] col_in_558,
    input  [511:0] col_in_559,
    input  [511:0] col_in_560,
    input  [511:0] col_in_561,
    input  [511:0] col_in_562,
    input  [511:0] col_in_563,
    input  [511:0] col_in_564,
    input  [511:0] col_in_565,
    input  [511:0] col_in_566,
    input  [511:0] col_in_567,
    input  [511:0] col_in_568,
    input  [511:0] col_in_569,
    input  [511:0] col_in_570,
    input  [511:0] col_in_571,
    input  [511:0] col_in_572,
    input  [511:0] col_in_573,
    input  [511:0] col_in_574,
    input  [511:0] col_in_575,
    input  [511:0] col_in_576,
    input  [511:0] col_in_577,
    input  [511:0] col_in_578,
    input  [511:0] col_in_579,
    input  [511:0] col_in_580,
    input  [511:0] col_in_581,
    input  [511:0] col_in_582,
    input  [511:0] col_in_583,
    input  [511:0] col_in_584,
    input  [511:0] col_in_585,
    input  [511:0] col_in_586,
    input  [511:0] col_in_587,
    input  [511:0] col_in_588,
    input  [511:0] col_in_589,
    input  [511:0] col_in_590,
    input  [511:0] col_in_591,
    input  [511:0] col_in_592,
    input  [511:0] col_in_593,
    input  [511:0] col_in_594,
    input  [511:0] col_in_595,
    input  [511:0] col_in_596,
    input  [511:0] col_in_597,
    input  [511:0] col_in_598,
    input  [511:0] col_in_599,
    input  [511:0] col_in_600,
    input  [511:0] col_in_601,
    input  [511:0] col_in_602,
    input  [511:0] col_in_603,
    input  [511:0] col_in_604,
    input  [511:0] col_in_605,
    input  [511:0] col_in_606,
    input  [511:0] col_in_607,
    input  [511:0] col_in_608,
    input  [511:0] col_in_609,
    input  [511:0] col_in_610,
    input  [511:0] col_in_611,
    input  [511:0] col_in_612,
    input  [511:0] col_in_613,
    input  [511:0] col_in_614,
    input  [511:0] col_in_615,
    input  [511:0] col_in_616,
    input  [511:0] col_in_617,
    input  [511:0] col_in_618,
    input  [511:0] col_in_619,
    input  [511:0] col_in_620,
    input  [511:0] col_in_621,
    input  [511:0] col_in_622,
    input  [511:0] col_in_623,
    input  [511:0] col_in_624,
    input  [511:0] col_in_625,
    input  [511:0] col_in_626,
    input  [511:0] col_in_627,
    input  [511:0] col_in_628,
    input  [511:0] col_in_629,
    input  [511:0] col_in_630,
    input  [511:0] col_in_631,
    input  [511:0] col_in_632,
    input  [511:0] col_in_633,
    input  [511:0] col_in_634,
    input  [511:0] col_in_635,
    input  [511:0] col_in_636,
    input  [511:0] col_in_637,
    input  [511:0] col_in_638,
    input  [511:0] col_in_639,
    input  [511:0] col_in_640,
    input  [511:0] col_in_641,
    input  [511:0] col_in_642,
    input  [511:0] col_in_643,
    input  [511:0] col_in_644,
    input  [511:0] col_in_645,
    input  [511:0] col_in_646,
    input  [511:0] col_in_647,
    input  [511:0] col_in_648,
    input  [511:0] col_in_649,
    input  [511:0] col_in_650,
    input  [511:0] col_in_651,
    input  [511:0] col_in_652,
    input  [511:0] col_in_653,
    input  [511:0] col_in_654,
    input  [511:0] col_in_655,
    input  [511:0] col_in_656,
    input  [511:0] col_in_657,
    input  [511:0] col_in_658,
    input  [511:0] col_in_659,
    input  [511:0] col_in_660,
    input  [511:0] col_in_661,
    input  [511:0] col_in_662,
    input  [511:0] col_in_663,
    input  [511:0] col_in_664,
    input  [511:0] col_in_665,
    input  [511:0] col_in_666,
    input  [511:0] col_in_667,
    input  [511:0] col_in_668,
    input  [511:0] col_in_669,
    input  [511:0] col_in_670,
    input  [511:0] col_in_671,
    input  [511:0] col_in_672,
    input  [511:0] col_in_673,
    input  [511:0] col_in_674,
    input  [511:0] col_in_675,
    input  [511:0] col_in_676,
    input  [511:0] col_in_677,
    input  [511:0] col_in_678,
    input  [511:0] col_in_679,
    input  [511:0] col_in_680,
    input  [511:0] col_in_681,
    input  [511:0] col_in_682,
    input  [511:0] col_in_683,
    input  [511:0] col_in_684,
    input  [511:0] col_in_685,
    input  [511:0] col_in_686,
    input  [511:0] col_in_687,
    input  [511:0] col_in_688,
    input  [511:0] col_in_689,
    input  [511:0] col_in_690,
    input  [511:0] col_in_691,
    input  [511:0] col_in_692,
    input  [511:0] col_in_693,
    input  [511:0] col_in_694,
    input  [511:0] col_in_695,
    input  [511:0] col_in_696,
    input  [511:0] col_in_697,
    input  [511:0] col_in_698,
    input  [511:0] col_in_699,
    input  [511:0] col_in_700,
    input  [511:0] col_in_701,
    input  [511:0] col_in_702,
    input  [511:0] col_in_703,
    input  [511:0] col_in_704,
    input  [511:0] col_in_705,
    input  [511:0] col_in_706,
    input  [511:0] col_in_707,
    input  [511:0] col_in_708,
    input  [511:0] col_in_709,
    input  [511:0] col_in_710,
    input  [511:0] col_in_711,
    input  [511:0] col_in_712,
    input  [511:0] col_in_713,
    input  [511:0] col_in_714,
    input  [511:0] col_in_715,
    input  [511:0] col_in_716,
    input  [511:0] col_in_717,
    input  [511:0] col_in_718,
    input  [511:0] col_in_719,
    input  [511:0] col_in_720,
    input  [511:0] col_in_721,
    input  [511:0] col_in_722,
    input  [511:0] col_in_723,
    input  [511:0] col_in_724,
    input  [511:0] col_in_725,
    input  [511:0] col_in_726,
    input  [511:0] col_in_727,
    input  [511:0] col_in_728,
    input  [511:0] col_in_729,
    input  [511:0] col_in_730,
    input  [511:0] col_in_731,
    input  [511:0] col_in_732,
    input  [511:0] col_in_733,
    input  [511:0] col_in_734,
    input  [511:0] col_in_735,
    input  [511:0] col_in_736,
    input  [511:0] col_in_737,
    input  [511:0] col_in_738,
    input  [511:0] col_in_739,
    input  [511:0] col_in_740,
    input  [511:0] col_in_741,
    input  [511:0] col_in_742,
    input  [511:0] col_in_743,
    input  [511:0] col_in_744,
    input  [511:0] col_in_745,
    input  [511:0] col_in_746,
    input  [511:0] col_in_747,
    input  [511:0] col_in_748,
    input  [511:0] col_in_749,
    input  [511:0] col_in_750,
    input  [511:0] col_in_751,
    input  [511:0] col_in_752,
    input  [511:0] col_in_753,
    input  [511:0] col_in_754,
    input  [511:0] col_in_755,
    input  [511:0] col_in_756,
    input  [511:0] col_in_757,
    input  [511:0] col_in_758,
    input  [511:0] col_in_759,
    input  [511:0] col_in_760,
    input  [511:0] col_in_761,
    input  [511:0] col_in_762,
    input  [511:0] col_in_763,
    input  [511:0] col_in_764,
    input  [511:0] col_in_765,
    input  [511:0] col_in_766,
    input  [511:0] col_in_767,
    input  [511:0] col_in_768,
    input  [511:0] col_in_769,
    input  [511:0] col_in_770,
    input  [511:0] col_in_771,
    input  [511:0] col_in_772,
    input  [511:0] col_in_773,
    input  [511:0] col_in_774,
    input  [511:0] col_in_775,
    input  [511:0] col_in_776,
    input  [511:0] col_in_777,
    input  [511:0] col_in_778,
    input  [511:0] col_in_779,
    input  [511:0] col_in_780,
    input  [511:0] col_in_781,
    input  [511:0] col_in_782,
    input  [511:0] col_in_783,
    input  [511:0] col_in_784,
    input  [511:0] col_in_785,
    input  [511:0] col_in_786,
    input  [511:0] col_in_787,
    input  [511:0] col_in_788,
    input  [511:0] col_in_789,
    input  [511:0] col_in_790,
    input  [511:0] col_in_791,
    input  [511:0] col_in_792,
    input  [511:0] col_in_793,
    input  [511:0] col_in_794,
    input  [511:0] col_in_795,
    input  [511:0] col_in_796,
    input  [511:0] col_in_797,
    input  [511:0] col_in_798,
    input  [511:0] col_in_799,
    input  [511:0] col_in_800,
    input  [511:0] col_in_801,
    input  [511:0] col_in_802,
    input  [511:0] col_in_803,
    input  [511:0] col_in_804,
    input  [511:0] col_in_805,
    input  [511:0] col_in_806,
    input  [511:0] col_in_807,
    input  [511:0] col_in_808,
    input  [511:0] col_in_809,
    input  [511:0] col_in_810,
    input  [511:0] col_in_811,
    input  [511:0] col_in_812,
    input  [511:0] col_in_813,
    input  [511:0] col_in_814,
    input  [511:0] col_in_815,
    input  [511:0] col_in_816,
    input  [511:0] col_in_817,
    input  [511:0] col_in_818,
    input  [511:0] col_in_819,
    input  [511:0] col_in_820,
    input  [511:0] col_in_821,
    input  [511:0] col_in_822,
    input  [511:0] col_in_823,
    input  [511:0] col_in_824,
    input  [511:0] col_in_825,
    input  [511:0] col_in_826,
    input  [511:0] col_in_827,
    input  [511:0] col_in_828,
    input  [511:0] col_in_829,
    input  [511:0] col_in_830,
    input  [511:0] col_in_831,
    input  [511:0] col_in_832,
    input  [511:0] col_in_833,
    input  [511:0] col_in_834,
    input  [511:0] col_in_835,
    input  [511:0] col_in_836,
    input  [511:0] col_in_837,
    input  [511:0] col_in_838,
    input  [511:0] col_in_839,
    input  [511:0] col_in_840,
    input  [511:0] col_in_841,
    input  [511:0] col_in_842,
    input  [511:0] col_in_843,
    input  [511:0] col_in_844,
    input  [511:0] col_in_845,
    input  [511:0] col_in_846,
    input  [511:0] col_in_847,
    input  [511:0] col_in_848,
    input  [511:0] col_in_849,
    input  [511:0] col_in_850,
    input  [511:0] col_in_851,
    input  [511:0] col_in_852,
    input  [511:0] col_in_853,
    input  [511:0] col_in_854,
    input  [511:0] col_in_855,
    input  [511:0] col_in_856,
    input  [511:0] col_in_857,
    input  [511:0] col_in_858,
    input  [511:0] col_in_859,
    input  [511:0] col_in_860,
    input  [511:0] col_in_861,
    input  [511:0] col_in_862,
    input  [511:0] col_in_863,
    input  [511:0] col_in_864,
    input  [511:0] col_in_865,
    input  [511:0] col_in_866,
    input  [511:0] col_in_867,
    input  [511:0] col_in_868,
    input  [511:0] col_in_869,
    input  [511:0] col_in_870,
    input  [511:0] col_in_871,
    input  [511:0] col_in_872,
    input  [511:0] col_in_873,
    input  [511:0] col_in_874,
    input  [511:0] col_in_875,
    input  [511:0] col_in_876,
    input  [511:0] col_in_877,
    input  [511:0] col_in_878,
    input  [511:0] col_in_879,
    input  [511:0] col_in_880,
    input  [511:0] col_in_881,
    input  [511:0] col_in_882,
    input  [511:0] col_in_883,
    input  [511:0] col_in_884,
    input  [511:0] col_in_885,
    input  [511:0] col_in_886,
    input  [511:0] col_in_887,
    input  [511:0] col_in_888,
    input  [511:0] col_in_889,
    input  [511:0] col_in_890,
    input  [511:0] col_in_891,
    input  [511:0] col_in_892,
    input  [511:0] col_in_893,
    input  [511:0] col_in_894,
    input  [511:0] col_in_895,
    input  [511:0] col_in_896,
    input  [511:0] col_in_897,
    input  [511:0] col_in_898,
    input  [511:0] col_in_899,
    input  [511:0] col_in_900,
    input  [511:0] col_in_901,
    input  [511:0] col_in_902,
    input  [511:0] col_in_903,
    input  [511:0] col_in_904,
    input  [511:0] col_in_905,
    input  [511:0] col_in_906,
    input  [511:0] col_in_907,
    input  [511:0] col_in_908,
    input  [511:0] col_in_909,
    input  [511:0] col_in_910,
    input  [511:0] col_in_911,
    input  [511:0] col_in_912,
    input  [511:0] col_in_913,
    input  [511:0] col_in_914,
    input  [511:0] col_in_915,
    input  [511:0] col_in_916,
    input  [511:0] col_in_917,
    input  [511:0] col_in_918,
    input  [511:0] col_in_919,
    input  [511:0] col_in_920,
    input  [511:0] col_in_921,
    input  [511:0] col_in_922,
    input  [511:0] col_in_923,
    input  [511:0] col_in_924,
    input  [511:0] col_in_925,
    input  [511:0] col_in_926,
    input  [511:0] col_in_927,
    input  [511:0] col_in_928,
    input  [511:0] col_in_929,
    input  [511:0] col_in_930,
    input  [511:0] col_in_931,
    input  [511:0] col_in_932,
    input  [511:0] col_in_933,
    input  [511:0] col_in_934,
    input  [511:0] col_in_935,
    input  [511:0] col_in_936,
    input  [511:0] col_in_937,
    input  [511:0] col_in_938,
    input  [511:0] col_in_939,
    input  [511:0] col_in_940,
    input  [511:0] col_in_941,
    input  [511:0] col_in_942,
    input  [511:0] col_in_943,
    input  [511:0] col_in_944,
    input  [511:0] col_in_945,
    input  [511:0] col_in_946,
    input  [511:0] col_in_947,
    input  [511:0] col_in_948,
    input  [511:0] col_in_949,
    input  [511:0] col_in_950,
    input  [511:0] col_in_951,
    input  [511:0] col_in_952,
    input  [511:0] col_in_953,
    input  [511:0] col_in_954,
    input  [511:0] col_in_955,
    input  [511:0] col_in_956,
    input  [511:0] col_in_957,
    input  [511:0] col_in_958,
    input  [511:0] col_in_959,
    input  [511:0] col_in_960,
    input  [511:0] col_in_961,
    input  [511:0] col_in_962,
    input  [511:0] col_in_963,
    input  [511:0] col_in_964,
    input  [511:0] col_in_965,
    input  [511:0] col_in_966,
    input  [511:0] col_in_967,
    input  [511:0] col_in_968,
    input  [511:0] col_in_969,
    input  [511:0] col_in_970,
    input  [511:0] col_in_971,
    input  [511:0] col_in_972,
    input  [511:0] col_in_973,
    input  [511:0] col_in_974,
    input  [511:0] col_in_975,
    input  [511:0] col_in_976,
    input  [511:0] col_in_977,
    input  [511:0] col_in_978,
    input  [511:0] col_in_979,
    input  [511:0] col_in_980,
    input  [511:0] col_in_981,
    input  [511:0] col_in_982,
    input  [511:0] col_in_983,
    input  [511:0] col_in_984,
    input  [511:0] col_in_985,
    input  [511:0] col_in_986,
    input  [511:0] col_in_987,
    input  [511:0] col_in_988,
    input  [511:0] col_in_989,
    input  [511:0] col_in_990,
    input  [511:0] col_in_991,
    input  [511:0] col_in_992,
    input  [511:0] col_in_993,
    input  [511:0] col_in_994,
    input  [511:0] col_in_995,
    input  [511:0] col_in_996,
    input  [511:0] col_in_997,
    input  [511:0] col_in_998,
    input  [511:0] col_in_999,
    input  [511:0] col_in_1000,
    input  [511:0] col_in_1001,
    input  [511:0] col_in_1002,
    input  [511:0] col_in_1003,
    input  [511:0] col_in_1004,
    input  [511:0] col_in_1005,
    input  [511:0] col_in_1006,
    input  [511:0] col_in_1007,
    input  [511:0] col_in_1008,
    input  [511:0] col_in_1009,
    input  [511:0] col_in_1010,
    input  [511:0] col_in_1011,
    input  [511:0] col_in_1012,
    input  [511:0] col_in_1013,
    input  [511:0] col_in_1014,
    input  [511:0] col_in_1015,
    input  [511:0] col_in_1016,
    input  [511:0] col_in_1017,
    input  [511:0] col_in_1018,
    input  [511:0] col_in_1019,
    input  [511:0] col_in_1020,
    input  [511:0] col_in_1021,
    input  [511:0] col_in_1022,
    input  [511:0] col_in_1023,

    output [151:0] col_out_0,
    output [151:0] col_out_1,
    output [151:0] col_out_2,
    output [151:0] col_out_3,
    output [151:0] col_out_4,
    output [151:0] col_out_5,
    output [151:0] col_out_6,
    output [151:0] col_out_7,
    output [151:0] col_out_8,
    output [151:0] col_out_9,
    output [151:0] col_out_10,
    output [151:0] col_out_11,
    output [151:0] col_out_12,
    output [151:0] col_out_13,
    output [151:0] col_out_14,
    output [151:0] col_out_15,
    output [151:0] col_out_16,
    output [151:0] col_out_17,
    output [151:0] col_out_18,
    output [151:0] col_out_19,
    output [151:0] col_out_20,
    output [151:0] col_out_21,
    output [151:0] col_out_22,
    output [151:0] col_out_23,
    output [151:0] col_out_24,
    output [151:0] col_out_25,
    output [151:0] col_out_26,
    output [151:0] col_out_27,
    output [151:0] col_out_28,
    output [151:0] col_out_29,
    output [151:0] col_out_30,
    output [151:0] col_out_31,
    output [151:0] col_out_32,
    output [151:0] col_out_33,
    output [151:0] col_out_34,
    output [151:0] col_out_35,
    output [151:0] col_out_36,
    output [151:0] col_out_37,
    output [151:0] col_out_38,
    output [151:0] col_out_39,
    output [151:0] col_out_40,
    output [151:0] col_out_41,
    output [151:0] col_out_42,
    output [151:0] col_out_43,
    output [151:0] col_out_44,
    output [151:0] col_out_45,
    output [151:0] col_out_46,
    output [151:0] col_out_47,
    output [151:0] col_out_48,
    output [151:0] col_out_49,
    output [151:0] col_out_50,
    output [151:0] col_out_51,
    output [151:0] col_out_52,
    output [151:0] col_out_53,
    output [151:0] col_out_54,
    output [151:0] col_out_55,
    output [151:0] col_out_56,
    output [151:0] col_out_57,
    output [151:0] col_out_58,
    output [151:0] col_out_59,
    output [151:0] col_out_60,
    output [151:0] col_out_61,
    output [151:0] col_out_62,
    output [151:0] col_out_63,
    output [151:0] col_out_64,
    output [151:0] col_out_65,
    output [151:0] col_out_66,
    output [151:0] col_out_67,
    output [151:0] col_out_68,
    output [151:0] col_out_69,
    output [151:0] col_out_70,
    output [151:0] col_out_71,
    output [151:0] col_out_72,
    output [151:0] col_out_73,
    output [151:0] col_out_74,
    output [151:0] col_out_75,
    output [151:0] col_out_76,
    output [151:0] col_out_77,
    output [151:0] col_out_78,
    output [151:0] col_out_79,
    output [151:0] col_out_80,
    output [151:0] col_out_81,
    output [151:0] col_out_82,
    output [151:0] col_out_83,
    output [151:0] col_out_84,
    output [151:0] col_out_85,
    output [151:0] col_out_86,
    output [151:0] col_out_87,
    output [151:0] col_out_88,
    output [151:0] col_out_89,
    output [151:0] col_out_90,
    output [151:0] col_out_91,
    output [151:0] col_out_92,
    output [151:0] col_out_93,
    output [151:0] col_out_94,
    output [151:0] col_out_95,
    output [151:0] col_out_96,
    output [151:0] col_out_97,
    output [151:0] col_out_98,
    output [151:0] col_out_99,
    output [151:0] col_out_100,
    output [151:0] col_out_101,
    output [151:0] col_out_102,
    output [151:0] col_out_103,
    output [151:0] col_out_104,
    output [151:0] col_out_105,
    output [151:0] col_out_106,
    output [151:0] col_out_107,
    output [151:0] col_out_108,
    output [151:0] col_out_109,
    output [151:0] col_out_110,
    output [151:0] col_out_111,
    output [151:0] col_out_112,
    output [151:0] col_out_113,
    output [151:0] col_out_114,
    output [151:0] col_out_115,
    output [151:0] col_out_116,
    output [151:0] col_out_117,
    output [151:0] col_out_118,
    output [151:0] col_out_119,
    output [151:0] col_out_120,
    output [151:0] col_out_121,
    output [151:0] col_out_122,
    output [151:0] col_out_123,
    output [151:0] col_out_124,
    output [151:0] col_out_125,
    output [151:0] col_out_126,
    output [151:0] col_out_127,
    output [151:0] col_out_128,
    output [151:0] col_out_129,
    output [151:0] col_out_130,
    output [151:0] col_out_131,
    output [151:0] col_out_132,
    output [151:0] col_out_133,
    output [151:0] col_out_134,
    output [151:0] col_out_135,
    output [151:0] col_out_136,
    output [151:0] col_out_137,
    output [151:0] col_out_138,
    output [151:0] col_out_139,
    output [151:0] col_out_140,
    output [151:0] col_out_141,
    output [151:0] col_out_142,
    output [151:0] col_out_143,
    output [151:0] col_out_144,
    output [151:0] col_out_145,
    output [151:0] col_out_146,
    output [151:0] col_out_147,
    output [151:0] col_out_148,
    output [151:0] col_out_149,
    output [151:0] col_out_150,
    output [151:0] col_out_151,
    output [151:0] col_out_152,
    output [151:0] col_out_153,
    output [151:0] col_out_154,
    output [151:0] col_out_155,
    output [151:0] col_out_156,
    output [151:0] col_out_157,
    output [151:0] col_out_158,
    output [151:0] col_out_159,
    output [151:0] col_out_160,
    output [151:0] col_out_161,
    output [151:0] col_out_162,
    output [151:0] col_out_163,
    output [151:0] col_out_164,
    output [151:0] col_out_165,
    output [151:0] col_out_166,
    output [151:0] col_out_167,
    output [151:0] col_out_168,
    output [151:0] col_out_169,
    output [151:0] col_out_170,
    output [151:0] col_out_171,
    output [151:0] col_out_172,
    output [151:0] col_out_173,
    output [151:0] col_out_174,
    output [151:0] col_out_175,
    output [151:0] col_out_176,
    output [151:0] col_out_177,
    output [151:0] col_out_178,
    output [151:0] col_out_179,
    output [151:0] col_out_180,
    output [151:0] col_out_181,
    output [151:0] col_out_182,
    output [151:0] col_out_183,
    output [151:0] col_out_184,
    output [151:0] col_out_185,
    output [151:0] col_out_186,
    output [151:0] col_out_187,
    output [151:0] col_out_188,
    output [151:0] col_out_189,
    output [151:0] col_out_190,
    output [151:0] col_out_191,
    output [151:0] col_out_192,
    output [151:0] col_out_193,
    output [151:0] col_out_194,
    output [151:0] col_out_195,
    output [151:0] col_out_196,
    output [151:0] col_out_197,
    output [151:0] col_out_198,
    output [151:0] col_out_199,
    output [151:0] col_out_200,
    output [151:0] col_out_201,
    output [151:0] col_out_202,
    output [151:0] col_out_203,
    output [151:0] col_out_204,
    output [151:0] col_out_205,
    output [151:0] col_out_206,
    output [151:0] col_out_207,
    output [151:0] col_out_208,
    output [151:0] col_out_209,
    output [151:0] col_out_210,
    output [151:0] col_out_211,
    output [151:0] col_out_212,
    output [151:0] col_out_213,
    output [151:0] col_out_214,
    output [151:0] col_out_215,
    output [151:0] col_out_216,
    output [151:0] col_out_217,
    output [151:0] col_out_218,
    output [151:0] col_out_219,
    output [151:0] col_out_220,
    output [151:0] col_out_221,
    output [151:0] col_out_222,
    output [151:0] col_out_223,
    output [151:0] col_out_224,
    output [151:0] col_out_225,
    output [151:0] col_out_226,
    output [151:0] col_out_227,
    output [151:0] col_out_228,
    output [151:0] col_out_229,
    output [151:0] col_out_230,
    output [151:0] col_out_231,
    output [151:0] col_out_232,
    output [151:0] col_out_233,
    output [151:0] col_out_234,
    output [151:0] col_out_235,
    output [151:0] col_out_236,
    output [151:0] col_out_237,
    output [151:0] col_out_238,
    output [151:0] col_out_239,
    output [151:0] col_out_240,
    output [151:0] col_out_241,
    output [151:0] col_out_242,
    output [151:0] col_out_243,
    output [151:0] col_out_244,
    output [151:0] col_out_245,
    output [151:0] col_out_246,
    output [151:0] col_out_247,
    output [151:0] col_out_248,
    output [151:0] col_out_249,
    output [151:0] col_out_250,
    output [151:0] col_out_251,
    output [151:0] col_out_252,
    output [151:0] col_out_253,
    output [151:0] col_out_254,
    output [151:0] col_out_255,
    output [151:0] col_out_256,
    output [151:0] col_out_257,
    output [151:0] col_out_258,
    output [151:0] col_out_259,
    output [151:0] col_out_260,
    output [151:0] col_out_261,
    output [151:0] col_out_262,
    output [151:0] col_out_263,
    output [151:0] col_out_264,
    output [151:0] col_out_265,
    output [151:0] col_out_266,
    output [151:0] col_out_267,
    output [151:0] col_out_268,
    output [151:0] col_out_269,
    output [151:0] col_out_270,
    output [151:0] col_out_271,
    output [151:0] col_out_272,
    output [151:0] col_out_273,
    output [151:0] col_out_274,
    output [151:0] col_out_275,
    output [151:0] col_out_276,
    output [151:0] col_out_277,
    output [151:0] col_out_278,
    output [151:0] col_out_279,
    output [151:0] col_out_280,
    output [151:0] col_out_281,
    output [151:0] col_out_282,
    output [151:0] col_out_283,
    output [151:0] col_out_284,
    output [151:0] col_out_285,
    output [151:0] col_out_286,
    output [151:0] col_out_287,
    output [151:0] col_out_288,
    output [151:0] col_out_289,
    output [151:0] col_out_290,
    output [151:0] col_out_291,
    output [151:0] col_out_292,
    output [151:0] col_out_293,
    output [151:0] col_out_294,
    output [151:0] col_out_295,
    output [151:0] col_out_296,
    output [151:0] col_out_297,
    output [151:0] col_out_298,
    output [151:0] col_out_299,
    output [151:0] col_out_300,
    output [151:0] col_out_301,
    output [151:0] col_out_302,
    output [151:0] col_out_303,
    output [151:0] col_out_304,
    output [151:0] col_out_305,
    output [151:0] col_out_306,
    output [151:0] col_out_307,
    output [151:0] col_out_308,
    output [151:0] col_out_309,
    output [151:0] col_out_310,
    output [151:0] col_out_311,
    output [151:0] col_out_312,
    output [151:0] col_out_313,
    output [151:0] col_out_314,
    output [151:0] col_out_315,
    output [151:0] col_out_316,
    output [151:0] col_out_317,
    output [151:0] col_out_318,
    output [151:0] col_out_319,
    output [151:0] col_out_320,
    output [151:0] col_out_321,
    output [151:0] col_out_322,
    output [151:0] col_out_323,
    output [151:0] col_out_324,
    output [151:0] col_out_325,
    output [151:0] col_out_326,
    output [151:0] col_out_327,
    output [151:0] col_out_328,
    output [151:0] col_out_329,
    output [151:0] col_out_330,
    output [151:0] col_out_331,
    output [151:0] col_out_332,
    output [151:0] col_out_333,
    output [151:0] col_out_334,
    output [151:0] col_out_335,
    output [151:0] col_out_336,
    output [151:0] col_out_337,
    output [151:0] col_out_338,
    output [151:0] col_out_339,
    output [151:0] col_out_340,
    output [151:0] col_out_341,
    output [151:0] col_out_342,
    output [151:0] col_out_343,
    output [151:0] col_out_344,
    output [151:0] col_out_345,
    output [151:0] col_out_346,
    output [151:0] col_out_347,
    output [151:0] col_out_348,
    output [151:0] col_out_349,
    output [151:0] col_out_350,
    output [151:0] col_out_351,
    output [151:0] col_out_352,
    output [151:0] col_out_353,
    output [151:0] col_out_354,
    output [151:0] col_out_355,
    output [151:0] col_out_356,
    output [151:0] col_out_357,
    output [151:0] col_out_358,
    output [151:0] col_out_359,
    output [151:0] col_out_360,
    output [151:0] col_out_361,
    output [151:0] col_out_362,
    output [151:0] col_out_363,
    output [151:0] col_out_364,
    output [151:0] col_out_365,
    output [151:0] col_out_366,
    output [151:0] col_out_367,
    output [151:0] col_out_368,
    output [151:0] col_out_369,
    output [151:0] col_out_370,
    output [151:0] col_out_371,
    output [151:0] col_out_372,
    output [151:0] col_out_373,
    output [151:0] col_out_374,
    output [151:0] col_out_375,
    output [151:0] col_out_376,
    output [151:0] col_out_377,
    output [151:0] col_out_378,
    output [151:0] col_out_379,
    output [151:0] col_out_380,
    output [151:0] col_out_381,
    output [151:0] col_out_382,
    output [151:0] col_out_383,
    output [151:0] col_out_384,
    output [151:0] col_out_385,
    output [151:0] col_out_386,
    output [151:0] col_out_387,
    output [151:0] col_out_388,
    output [151:0] col_out_389,
    output [151:0] col_out_390,
    output [151:0] col_out_391,
    output [151:0] col_out_392,
    output [151:0] col_out_393,
    output [151:0] col_out_394,
    output [151:0] col_out_395,
    output [151:0] col_out_396,
    output [151:0] col_out_397,
    output [151:0] col_out_398,
    output [151:0] col_out_399,
    output [151:0] col_out_400,
    output [151:0] col_out_401,
    output [151:0] col_out_402,
    output [151:0] col_out_403,
    output [151:0] col_out_404,
    output [151:0] col_out_405,
    output [151:0] col_out_406,
    output [151:0] col_out_407,
    output [151:0] col_out_408,
    output [151:0] col_out_409,
    output [151:0] col_out_410,
    output [151:0] col_out_411,
    output [151:0] col_out_412,
    output [151:0] col_out_413,
    output [151:0] col_out_414,
    output [151:0] col_out_415,
    output [151:0] col_out_416,
    output [151:0] col_out_417,
    output [151:0] col_out_418,
    output [151:0] col_out_419,
    output [151:0] col_out_420,
    output [151:0] col_out_421,
    output [151:0] col_out_422,
    output [151:0] col_out_423,
    output [151:0] col_out_424,
    output [151:0] col_out_425,
    output [151:0] col_out_426,
    output [151:0] col_out_427,
    output [151:0] col_out_428,
    output [151:0] col_out_429,
    output [151:0] col_out_430,
    output [151:0] col_out_431,
    output [151:0] col_out_432,
    output [151:0] col_out_433,
    output [151:0] col_out_434,
    output [151:0] col_out_435,
    output [151:0] col_out_436,
    output [151:0] col_out_437,
    output [151:0] col_out_438,
    output [151:0] col_out_439,
    output [151:0] col_out_440,
    output [151:0] col_out_441,
    output [151:0] col_out_442,
    output [151:0] col_out_443,
    output [151:0] col_out_444,
    output [151:0] col_out_445,
    output [151:0] col_out_446,
    output [151:0] col_out_447,
    output [151:0] col_out_448,
    output [151:0] col_out_449,
    output [151:0] col_out_450,
    output [151:0] col_out_451,
    output [151:0] col_out_452,
    output [151:0] col_out_453,
    output [151:0] col_out_454,
    output [151:0] col_out_455,
    output [151:0] col_out_456,
    output [151:0] col_out_457,
    output [151:0] col_out_458,
    output [151:0] col_out_459,
    output [151:0] col_out_460,
    output [151:0] col_out_461,
    output [151:0] col_out_462,
    output [151:0] col_out_463,
    output [151:0] col_out_464,
    output [151:0] col_out_465,
    output [151:0] col_out_466,
    output [151:0] col_out_467,
    output [151:0] col_out_468,
    output [151:0] col_out_469,
    output [151:0] col_out_470,
    output [151:0] col_out_471,
    output [151:0] col_out_472,
    output [151:0] col_out_473,
    output [151:0] col_out_474,
    output [151:0] col_out_475,
    output [151:0] col_out_476,
    output [151:0] col_out_477,
    output [151:0] col_out_478,
    output [151:0] col_out_479,
    output [151:0] col_out_480,
    output [151:0] col_out_481,
    output [151:0] col_out_482,
    output [151:0] col_out_483,
    output [151:0] col_out_484,
    output [151:0] col_out_485,
    output [151:0] col_out_486,
    output [151:0] col_out_487,
    output [151:0] col_out_488,
    output [151:0] col_out_489,
    output [151:0] col_out_490,
    output [151:0] col_out_491,
    output [151:0] col_out_492,
    output [151:0] col_out_493,
    output [151:0] col_out_494,
    output [151:0] col_out_495,
    output [151:0] col_out_496,
    output [151:0] col_out_497,
    output [151:0] col_out_498,
    output [151:0] col_out_499,
    output [151:0] col_out_500,
    output [151:0] col_out_501,
    output [151:0] col_out_502,
    output [151:0] col_out_503,
    output [151:0] col_out_504,
    output [151:0] col_out_505,
    output [151:0] col_out_506,
    output [151:0] col_out_507,
    output [151:0] col_out_508,
    output [151:0] col_out_509,
    output [151:0] col_out_510,
    output [151:0] col_out_511,
    output [151:0] col_out_512,
    output [151:0] col_out_513,
    output [151:0] col_out_514,
    output [151:0] col_out_515,
    output [151:0] col_out_516,
    output [151:0] col_out_517,
    output [151:0] col_out_518,
    output [151:0] col_out_519,
    output [151:0] col_out_520,
    output [151:0] col_out_521,
    output [151:0] col_out_522,
    output [151:0] col_out_523,
    output [151:0] col_out_524,
    output [151:0] col_out_525,
    output [151:0] col_out_526,
    output [151:0] col_out_527,
    output [151:0] col_out_528,
    output [151:0] col_out_529,
    output [151:0] col_out_530,
    output [151:0] col_out_531,
    output [151:0] col_out_532,
    output [151:0] col_out_533,
    output [151:0] col_out_534,
    output [151:0] col_out_535,
    output [151:0] col_out_536,
    output [151:0] col_out_537,
    output [151:0] col_out_538,
    output [151:0] col_out_539,
    output [151:0] col_out_540,
    output [151:0] col_out_541,
    output [151:0] col_out_542,
    output [151:0] col_out_543,
    output [151:0] col_out_544,
    output [151:0] col_out_545,
    output [151:0] col_out_546,
    output [151:0] col_out_547,
    output [151:0] col_out_548,
    output [151:0] col_out_549,
    output [151:0] col_out_550,
    output [151:0] col_out_551,
    output [151:0] col_out_552,
    output [151:0] col_out_553,
    output [151:0] col_out_554,
    output [151:0] col_out_555,
    output [151:0] col_out_556,
    output [151:0] col_out_557,
    output [151:0] col_out_558,
    output [151:0] col_out_559,
    output [151:0] col_out_560,
    output [151:0] col_out_561,
    output [151:0] col_out_562,
    output [151:0] col_out_563,
    output [151:0] col_out_564,
    output [151:0] col_out_565,
    output [151:0] col_out_566,
    output [151:0] col_out_567,
    output [151:0] col_out_568,
    output [151:0] col_out_569,
    output [151:0] col_out_570,
    output [151:0] col_out_571,
    output [151:0] col_out_572,
    output [151:0] col_out_573,
    output [151:0] col_out_574,
    output [151:0] col_out_575,
    output [151:0] col_out_576,
    output [151:0] col_out_577,
    output [151:0] col_out_578,
    output [151:0] col_out_579,
    output [151:0] col_out_580,
    output [151:0] col_out_581,
    output [151:0] col_out_582,
    output [151:0] col_out_583,
    output [151:0] col_out_584,
    output [151:0] col_out_585,
    output [151:0] col_out_586,
    output [151:0] col_out_587,
    output [151:0] col_out_588,
    output [151:0] col_out_589,
    output [151:0] col_out_590,
    output [151:0] col_out_591,
    output [151:0] col_out_592,
    output [151:0] col_out_593,
    output [151:0] col_out_594,
    output [151:0] col_out_595,
    output [151:0] col_out_596,
    output [151:0] col_out_597,
    output [151:0] col_out_598,
    output [151:0] col_out_599,
    output [151:0] col_out_600,
    output [151:0] col_out_601,
    output [151:0] col_out_602,
    output [151:0] col_out_603,
    output [151:0] col_out_604,
    output [151:0] col_out_605,
    output [151:0] col_out_606,
    output [151:0] col_out_607,
    output [151:0] col_out_608,
    output [151:0] col_out_609,
    output [151:0] col_out_610,
    output [151:0] col_out_611,
    output [151:0] col_out_612,
    output [151:0] col_out_613,
    output [151:0] col_out_614,
    output [151:0] col_out_615,
    output [151:0] col_out_616,
    output [151:0] col_out_617,
    output [151:0] col_out_618,
    output [151:0] col_out_619,
    output [151:0] col_out_620,
    output [151:0] col_out_621,
    output [151:0] col_out_622,
    output [151:0] col_out_623,
    output [151:0] col_out_624,
    output [151:0] col_out_625,
    output [151:0] col_out_626,
    output [151:0] col_out_627,
    output [151:0] col_out_628,
    output [151:0] col_out_629,
    output [151:0] col_out_630,
    output [151:0] col_out_631,
    output [151:0] col_out_632,
    output [151:0] col_out_633,
    output [151:0] col_out_634,
    output [151:0] col_out_635,
    output [151:0] col_out_636,
    output [151:0] col_out_637,
    output [151:0] col_out_638,
    output [151:0] col_out_639,
    output [151:0] col_out_640,
    output [151:0] col_out_641,
    output [151:0] col_out_642,
    output [151:0] col_out_643,
    output [151:0] col_out_644,
    output [151:0] col_out_645,
    output [151:0] col_out_646,
    output [151:0] col_out_647,
    output [151:0] col_out_648,
    output [151:0] col_out_649,
    output [151:0] col_out_650,
    output [151:0] col_out_651,
    output [151:0] col_out_652,
    output [151:0] col_out_653,
    output [151:0] col_out_654,
    output [151:0] col_out_655,
    output [151:0] col_out_656,
    output [151:0] col_out_657,
    output [151:0] col_out_658,
    output [151:0] col_out_659,
    output [151:0] col_out_660,
    output [151:0] col_out_661,
    output [151:0] col_out_662,
    output [151:0] col_out_663,
    output [151:0] col_out_664,
    output [151:0] col_out_665,
    output [151:0] col_out_666,
    output [151:0] col_out_667,
    output [151:0] col_out_668,
    output [151:0] col_out_669,
    output [151:0] col_out_670,
    output [151:0] col_out_671,
    output [151:0] col_out_672,
    output [151:0] col_out_673,
    output [151:0] col_out_674,
    output [151:0] col_out_675,
    output [151:0] col_out_676,
    output [151:0] col_out_677,
    output [151:0] col_out_678,
    output [151:0] col_out_679,
    output [151:0] col_out_680,
    output [151:0] col_out_681,
    output [151:0] col_out_682,
    output [151:0] col_out_683,
    output [151:0] col_out_684,
    output [151:0] col_out_685,
    output [151:0] col_out_686,
    output [151:0] col_out_687,
    output [151:0] col_out_688,
    output [151:0] col_out_689,
    output [151:0] col_out_690,
    output [151:0] col_out_691,
    output [151:0] col_out_692,
    output [151:0] col_out_693,
    output [151:0] col_out_694,
    output [151:0] col_out_695,
    output [151:0] col_out_696,
    output [151:0] col_out_697,
    output [151:0] col_out_698,
    output [151:0] col_out_699,
    output [151:0] col_out_700,
    output [151:0] col_out_701,
    output [151:0] col_out_702,
    output [151:0] col_out_703,
    output [151:0] col_out_704,
    output [151:0] col_out_705,
    output [151:0] col_out_706,
    output [151:0] col_out_707,
    output [151:0] col_out_708,
    output [151:0] col_out_709,
    output [151:0] col_out_710,
    output [151:0] col_out_711,
    output [151:0] col_out_712,
    output [151:0] col_out_713,
    output [151:0] col_out_714,
    output [151:0] col_out_715,
    output [151:0] col_out_716,
    output [151:0] col_out_717,
    output [151:0] col_out_718,
    output [151:0] col_out_719,
    output [151:0] col_out_720,
    output [151:0] col_out_721,
    output [151:0] col_out_722,
    output [151:0] col_out_723,
    output [151:0] col_out_724,
    output [151:0] col_out_725,
    output [151:0] col_out_726,
    output [151:0] col_out_727,
    output [151:0] col_out_728,
    output [151:0] col_out_729,
    output [151:0] col_out_730,
    output [151:0] col_out_731,
    output [151:0] col_out_732,
    output [151:0] col_out_733,
    output [151:0] col_out_734,
    output [151:0] col_out_735,
    output [151:0] col_out_736,
    output [151:0] col_out_737,
    output [151:0] col_out_738,
    output [151:0] col_out_739,
    output [151:0] col_out_740,
    output [151:0] col_out_741,
    output [151:0] col_out_742,
    output [151:0] col_out_743,
    output [151:0] col_out_744,
    output [151:0] col_out_745,
    output [151:0] col_out_746,
    output [151:0] col_out_747,
    output [151:0] col_out_748,
    output [151:0] col_out_749,
    output [151:0] col_out_750,
    output [151:0] col_out_751,
    output [151:0] col_out_752,
    output [151:0] col_out_753,
    output [151:0] col_out_754,
    output [151:0] col_out_755,
    output [151:0] col_out_756,
    output [151:0] col_out_757,
    output [151:0] col_out_758,
    output [151:0] col_out_759,
    output [151:0] col_out_760,
    output [151:0] col_out_761,
    output [151:0] col_out_762,
    output [151:0] col_out_763,
    output [151:0] col_out_764,
    output [151:0] col_out_765,
    output [151:0] col_out_766,
    output [151:0] col_out_767,
    output [151:0] col_out_768,
    output [151:0] col_out_769,
    output [151:0] col_out_770,
    output [151:0] col_out_771,
    output [151:0] col_out_772,
    output [151:0] col_out_773,
    output [151:0] col_out_774,
    output [151:0] col_out_775,
    output [151:0] col_out_776,
    output [151:0] col_out_777,
    output [151:0] col_out_778,
    output [151:0] col_out_779,
    output [151:0] col_out_780,
    output [151:0] col_out_781,
    output [151:0] col_out_782,
    output [151:0] col_out_783,
    output [151:0] col_out_784,
    output [151:0] col_out_785,
    output [151:0] col_out_786,
    output [151:0] col_out_787,
    output [151:0] col_out_788,
    output [151:0] col_out_789,
    output [151:0] col_out_790,
    output [151:0] col_out_791,
    output [151:0] col_out_792,
    output [151:0] col_out_793,
    output [151:0] col_out_794,
    output [151:0] col_out_795,
    output [151:0] col_out_796,
    output [151:0] col_out_797,
    output [151:0] col_out_798,
    output [151:0] col_out_799,
    output [151:0] col_out_800,
    output [151:0] col_out_801,
    output [151:0] col_out_802,
    output [151:0] col_out_803,
    output [151:0] col_out_804,
    output [151:0] col_out_805,
    output [151:0] col_out_806,
    output [151:0] col_out_807,
    output [151:0] col_out_808,
    output [151:0] col_out_809,
    output [151:0] col_out_810,
    output [151:0] col_out_811,
    output [151:0] col_out_812,
    output [151:0] col_out_813,
    output [151:0] col_out_814,
    output [151:0] col_out_815,
    output [151:0] col_out_816,
    output [151:0] col_out_817,
    output [151:0] col_out_818,
    output [151:0] col_out_819,
    output [151:0] col_out_820,
    output [151:0] col_out_821,
    output [151:0] col_out_822,
    output [151:0] col_out_823,
    output [151:0] col_out_824,
    output [151:0] col_out_825,
    output [151:0] col_out_826,
    output [151:0] col_out_827,
    output [151:0] col_out_828,
    output [151:0] col_out_829,
    output [151:0] col_out_830,
    output [151:0] col_out_831,
    output [151:0] col_out_832,
    output [151:0] col_out_833,
    output [151:0] col_out_834,
    output [151:0] col_out_835,
    output [151:0] col_out_836,
    output [151:0] col_out_837,
    output [151:0] col_out_838,
    output [151:0] col_out_839,
    output [151:0] col_out_840,
    output [151:0] col_out_841,
    output [151:0] col_out_842,
    output [151:0] col_out_843,
    output [151:0] col_out_844,
    output [151:0] col_out_845,
    output [151:0] col_out_846,
    output [151:0] col_out_847,
    output [151:0] col_out_848,
    output [151:0] col_out_849,
    output [151:0] col_out_850,
    output [151:0] col_out_851,
    output [151:0] col_out_852,
    output [151:0] col_out_853,
    output [151:0] col_out_854,
    output [151:0] col_out_855,
    output [151:0] col_out_856,
    output [151:0] col_out_857,
    output [151:0] col_out_858,
    output [151:0] col_out_859,
    output [151:0] col_out_860,
    output [151:0] col_out_861,
    output [151:0] col_out_862,
    output [151:0] col_out_863,
    output [151:0] col_out_864,
    output [151:0] col_out_865,
    output [151:0] col_out_866,
    output [151:0] col_out_867,
    output [151:0] col_out_868,
    output [151:0] col_out_869,
    output [151:0] col_out_870,
    output [151:0] col_out_871,
    output [151:0] col_out_872,
    output [151:0] col_out_873,
    output [151:0] col_out_874,
    output [151:0] col_out_875,
    output [151:0] col_out_876,
    output [151:0] col_out_877,
    output [151:0] col_out_878,
    output [151:0] col_out_879,
    output [151:0] col_out_880,
    output [151:0] col_out_881,
    output [151:0] col_out_882,
    output [151:0] col_out_883,
    output [151:0] col_out_884,
    output [151:0] col_out_885,
    output [151:0] col_out_886,
    output [151:0] col_out_887,
    output [151:0] col_out_888,
    output [151:0] col_out_889,
    output [151:0] col_out_890,
    output [151:0] col_out_891,
    output [151:0] col_out_892,
    output [151:0] col_out_893,
    output [151:0] col_out_894,
    output [151:0] col_out_895,
    output [151:0] col_out_896,
    output [151:0] col_out_897,
    output [151:0] col_out_898,
    output [151:0] col_out_899,
    output [151:0] col_out_900,
    output [151:0] col_out_901,
    output [151:0] col_out_902,
    output [151:0] col_out_903,
    output [151:0] col_out_904,
    output [151:0] col_out_905,
    output [151:0] col_out_906,
    output [151:0] col_out_907,
    output [151:0] col_out_908,
    output [151:0] col_out_909,
    output [151:0] col_out_910,
    output [151:0] col_out_911,
    output [151:0] col_out_912,
    output [151:0] col_out_913,
    output [151:0] col_out_914,
    output [151:0] col_out_915,
    output [151:0] col_out_916,
    output [151:0] col_out_917,
    output [151:0] col_out_918,
    output [151:0] col_out_919,
    output [151:0] col_out_920,
    output [151:0] col_out_921,
    output [151:0] col_out_922,
    output [151:0] col_out_923,
    output [151:0] col_out_924,
    output [151:0] col_out_925,
    output [151:0] col_out_926,
    output [151:0] col_out_927,
    output [151:0] col_out_928,
    output [151:0] col_out_929,
    output [151:0] col_out_930,
    output [151:0] col_out_931,
    output [151:0] col_out_932,
    output [151:0] col_out_933,
    output [151:0] col_out_934,
    output [151:0] col_out_935,
    output [151:0] col_out_936,
    output [151:0] col_out_937,
    output [151:0] col_out_938,
    output [151:0] col_out_939,
    output [151:0] col_out_940,
    output [151:0] col_out_941,
    output [151:0] col_out_942,
    output [151:0] col_out_943,
    output [151:0] col_out_944,
    output [151:0] col_out_945,
    output [151:0] col_out_946,
    output [151:0] col_out_947,
    output [151:0] col_out_948,
    output [151:0] col_out_949,
    output [151:0] col_out_950,
    output [151:0] col_out_951,
    output [151:0] col_out_952,
    output [151:0] col_out_953,
    output [151:0] col_out_954,
    output [151:0] col_out_955,
    output [151:0] col_out_956,
    output [151:0] col_out_957,
    output [151:0] col_out_958,
    output [151:0] col_out_959,
    output [151:0] col_out_960,
    output [151:0] col_out_961,
    output [151:0] col_out_962,
    output [151:0] col_out_963,
    output [151:0] col_out_964,
    output [151:0] col_out_965,
    output [151:0] col_out_966,
    output [151:0] col_out_967,
    output [151:0] col_out_968,
    output [151:0] col_out_969,
    output [151:0] col_out_970,
    output [151:0] col_out_971,
    output [151:0] col_out_972,
    output [151:0] col_out_973,
    output [151:0] col_out_974,
    output [151:0] col_out_975,
    output [151:0] col_out_976,
    output [151:0] col_out_977,
    output [151:0] col_out_978,
    output [151:0] col_out_979,
    output [151:0] col_out_980,
    output [151:0] col_out_981,
    output [151:0] col_out_982,
    output [151:0] col_out_983,
    output [151:0] col_out_984,
    output [151:0] col_out_985,
    output [151:0] col_out_986,
    output [151:0] col_out_987,
    output [151:0] col_out_988,
    output [151:0] col_out_989,
    output [151:0] col_out_990,
    output [151:0] col_out_991,
    output [151:0] col_out_992,
    output [151:0] col_out_993,
    output [151:0] col_out_994,
    output [151:0] col_out_995,
    output [151:0] col_out_996,
    output [151:0] col_out_997,
    output [151:0] col_out_998,
    output [151:0] col_out_999,
    output [151:0] col_out_1000,
    output [151:0] col_out_1001,
    output [151:0] col_out_1002,
    output [151:0] col_out_1003,
    output [151:0] col_out_1004,
    output [151:0] col_out_1005,
    output [151:0] col_out_1006,
    output [151:0] col_out_1007,
    output [151:0] col_out_1008,
    output [151:0] col_out_1009,
    output [151:0] col_out_1010,
    output [151:0] col_out_1011,
    output [151:0] col_out_1012,
    output [151:0] col_out_1013,
    output [151:0] col_out_1014,
    output [151:0] col_out_1015,
    output [151:0] col_out_1016,
    output [151:0] col_out_1017,
    output [151:0] col_out_1018,
    output [151:0] col_out_1019,
    output [151:0] col_out_1020,
    output [151:0] col_out_1021,
    output [151:0] col_out_1022,
    output [151:0] col_out_1023,
    output [151:0] col_out_1024,
    output [151:0] col_out_1025,
    output [151:0] col_out_1026
);



//--compressor_array input and output----------------------

wire [512:0] u_ca_in_0;
wire [512:0] u_ca_in_1;
wire [512:0] u_ca_in_2;
wire [512:0] u_ca_in_3;
wire [512:0] u_ca_in_4;
wire [512:0] u_ca_in_5;
wire [512:0] u_ca_in_6;
wire [512:0] u_ca_in_7;
wire [512:0] u_ca_in_8;
wire [512:0] u_ca_in_9;
wire [512:0] u_ca_in_10;
wire [512:0] u_ca_in_11;
wire [512:0] u_ca_in_12;
wire [512:0] u_ca_in_13;
wire [512:0] u_ca_in_14;
wire [512:0] u_ca_in_15;
wire [512:0] u_ca_in_16;
wire [512:0] u_ca_in_17;
wire [512:0] u_ca_in_18;
wire [512:0] u_ca_in_19;
wire [512:0] u_ca_in_20;
wire [512:0] u_ca_in_21;
wire [512:0] u_ca_in_22;
wire [512:0] u_ca_in_23;
wire [512:0] u_ca_in_24;
wire [512:0] u_ca_in_25;
wire [512:0] u_ca_in_26;
wire [512:0] u_ca_in_27;
wire [512:0] u_ca_in_28;
wire [512:0] u_ca_in_29;
wire [512:0] u_ca_in_30;
wire [512:0] u_ca_in_31;
wire [512:0] u_ca_in_32;
wire [512:0] u_ca_in_33;
wire [512:0] u_ca_in_34;
wire [512:0] u_ca_in_35;
wire [512:0] u_ca_in_36;
wire [512:0] u_ca_in_37;
wire [512:0] u_ca_in_38;
wire [512:0] u_ca_in_39;
wire [512:0] u_ca_in_40;
wire [512:0] u_ca_in_41;
wire [512:0] u_ca_in_42;
wire [512:0] u_ca_in_43;
wire [512:0] u_ca_in_44;
wire [512:0] u_ca_in_45;
wire [512:0] u_ca_in_46;
wire [512:0] u_ca_in_47;
wire [512:0] u_ca_in_48;
wire [512:0] u_ca_in_49;
wire [512:0] u_ca_in_50;
wire [512:0] u_ca_in_51;
wire [512:0] u_ca_in_52;
wire [512:0] u_ca_in_53;
wire [512:0] u_ca_in_54;
wire [512:0] u_ca_in_55;
wire [512:0] u_ca_in_56;
wire [512:0] u_ca_in_57;
wire [512:0] u_ca_in_58;
wire [512:0] u_ca_in_59;
wire [512:0] u_ca_in_60;
wire [512:0] u_ca_in_61;
wire [512:0] u_ca_in_62;
wire [512:0] u_ca_in_63;
wire [512:0] u_ca_in_64;
wire [512:0] u_ca_in_65;
wire [512:0] u_ca_in_66;
wire [512:0] u_ca_in_67;
wire [512:0] u_ca_in_68;
wire [512:0] u_ca_in_69;
wire [512:0] u_ca_in_70;
wire [512:0] u_ca_in_71;
wire [512:0] u_ca_in_72;
wire [512:0] u_ca_in_73;
wire [512:0] u_ca_in_74;
wire [512:0] u_ca_in_75;
wire [512:0] u_ca_in_76;
wire [512:0] u_ca_in_77;
wire [512:0] u_ca_in_78;
wire [512:0] u_ca_in_79;
wire [512:0] u_ca_in_80;
wire [512:0] u_ca_in_81;
wire [512:0] u_ca_in_82;
wire [512:0] u_ca_in_83;
wire [512:0] u_ca_in_84;
wire [512:0] u_ca_in_85;
wire [512:0] u_ca_in_86;
wire [512:0] u_ca_in_87;
wire [512:0] u_ca_in_88;
wire [512:0] u_ca_in_89;
wire [512:0] u_ca_in_90;
wire [512:0] u_ca_in_91;
wire [512:0] u_ca_in_92;
wire [512:0] u_ca_in_93;
wire [512:0] u_ca_in_94;
wire [512:0] u_ca_in_95;
wire [512:0] u_ca_in_96;
wire [512:0] u_ca_in_97;
wire [512:0] u_ca_in_98;
wire [512:0] u_ca_in_99;
wire [512:0] u_ca_in_100;
wire [512:0] u_ca_in_101;
wire [512:0] u_ca_in_102;
wire [512:0] u_ca_in_103;
wire [512:0] u_ca_in_104;
wire [512:0] u_ca_in_105;
wire [512:0] u_ca_in_106;
wire [512:0] u_ca_in_107;
wire [512:0] u_ca_in_108;
wire [512:0] u_ca_in_109;
wire [512:0] u_ca_in_110;
wire [512:0] u_ca_in_111;
wire [512:0] u_ca_in_112;
wire [512:0] u_ca_in_113;
wire [512:0] u_ca_in_114;
wire [512:0] u_ca_in_115;
wire [512:0] u_ca_in_116;
wire [512:0] u_ca_in_117;
wire [512:0] u_ca_in_118;
wire [512:0] u_ca_in_119;
wire [512:0] u_ca_in_120;
wire [512:0] u_ca_in_121;
wire [512:0] u_ca_in_122;
wire [512:0] u_ca_in_123;
wire [512:0] u_ca_in_124;
wire [512:0] u_ca_in_125;
wire [512:0] u_ca_in_126;
wire [512:0] u_ca_in_127;
wire [512:0] u_ca_in_128;
wire [512:0] u_ca_in_129;
wire [512:0] u_ca_in_130;
wire [512:0] u_ca_in_131;
wire [512:0] u_ca_in_132;
wire [512:0] u_ca_in_133;
wire [512:0] u_ca_in_134;
wire [512:0] u_ca_in_135;
wire [512:0] u_ca_in_136;
wire [512:0] u_ca_in_137;
wire [512:0] u_ca_in_138;
wire [512:0] u_ca_in_139;
wire [512:0] u_ca_in_140;
wire [512:0] u_ca_in_141;
wire [512:0] u_ca_in_142;
wire [512:0] u_ca_in_143;
wire [512:0] u_ca_in_144;
wire [512:0] u_ca_in_145;
wire [512:0] u_ca_in_146;
wire [512:0] u_ca_in_147;
wire [512:0] u_ca_in_148;
wire [512:0] u_ca_in_149;
wire [512:0] u_ca_in_150;
wire [512:0] u_ca_in_151;
wire [512:0] u_ca_in_152;
wire [512:0] u_ca_in_153;
wire [512:0] u_ca_in_154;
wire [512:0] u_ca_in_155;
wire [512:0] u_ca_in_156;
wire [512:0] u_ca_in_157;
wire [512:0] u_ca_in_158;
wire [512:0] u_ca_in_159;
wire [512:0] u_ca_in_160;
wire [512:0] u_ca_in_161;
wire [512:0] u_ca_in_162;
wire [512:0] u_ca_in_163;
wire [512:0] u_ca_in_164;
wire [512:0] u_ca_in_165;
wire [512:0] u_ca_in_166;
wire [512:0] u_ca_in_167;
wire [512:0] u_ca_in_168;
wire [512:0] u_ca_in_169;
wire [512:0] u_ca_in_170;
wire [512:0] u_ca_in_171;
wire [512:0] u_ca_in_172;
wire [512:0] u_ca_in_173;
wire [512:0] u_ca_in_174;
wire [512:0] u_ca_in_175;
wire [512:0] u_ca_in_176;
wire [512:0] u_ca_in_177;
wire [512:0] u_ca_in_178;
wire [512:0] u_ca_in_179;
wire [512:0] u_ca_in_180;
wire [512:0] u_ca_in_181;
wire [512:0] u_ca_in_182;
wire [512:0] u_ca_in_183;
wire [512:0] u_ca_in_184;
wire [512:0] u_ca_in_185;
wire [512:0] u_ca_in_186;
wire [512:0] u_ca_in_187;
wire [512:0] u_ca_in_188;
wire [512:0] u_ca_in_189;
wire [512:0] u_ca_in_190;
wire [512:0] u_ca_in_191;
wire [512:0] u_ca_in_192;
wire [512:0] u_ca_in_193;
wire [512:0] u_ca_in_194;
wire [512:0] u_ca_in_195;
wire [512:0] u_ca_in_196;
wire [512:0] u_ca_in_197;
wire [512:0] u_ca_in_198;
wire [512:0] u_ca_in_199;
wire [512:0] u_ca_in_200;
wire [512:0] u_ca_in_201;
wire [512:0] u_ca_in_202;
wire [512:0] u_ca_in_203;
wire [512:0] u_ca_in_204;
wire [512:0] u_ca_in_205;
wire [512:0] u_ca_in_206;
wire [512:0] u_ca_in_207;
wire [512:0] u_ca_in_208;
wire [512:0] u_ca_in_209;
wire [512:0] u_ca_in_210;
wire [512:0] u_ca_in_211;
wire [512:0] u_ca_in_212;
wire [512:0] u_ca_in_213;
wire [512:0] u_ca_in_214;
wire [512:0] u_ca_in_215;
wire [512:0] u_ca_in_216;
wire [512:0] u_ca_in_217;
wire [512:0] u_ca_in_218;
wire [512:0] u_ca_in_219;
wire [512:0] u_ca_in_220;
wire [512:0] u_ca_in_221;
wire [512:0] u_ca_in_222;
wire [512:0] u_ca_in_223;
wire [512:0] u_ca_in_224;
wire [512:0] u_ca_in_225;
wire [512:0] u_ca_in_226;
wire [512:0] u_ca_in_227;
wire [512:0] u_ca_in_228;
wire [512:0] u_ca_in_229;
wire [512:0] u_ca_in_230;
wire [512:0] u_ca_in_231;
wire [512:0] u_ca_in_232;
wire [512:0] u_ca_in_233;
wire [512:0] u_ca_in_234;
wire [512:0] u_ca_in_235;
wire [512:0] u_ca_in_236;
wire [512:0] u_ca_in_237;
wire [512:0] u_ca_in_238;
wire [512:0] u_ca_in_239;
wire [512:0] u_ca_in_240;
wire [512:0] u_ca_in_241;
wire [512:0] u_ca_in_242;
wire [512:0] u_ca_in_243;
wire [512:0] u_ca_in_244;
wire [512:0] u_ca_in_245;
wire [512:0] u_ca_in_246;
wire [512:0] u_ca_in_247;
wire [512:0] u_ca_in_248;
wire [512:0] u_ca_in_249;
wire [512:0] u_ca_in_250;
wire [512:0] u_ca_in_251;
wire [512:0] u_ca_in_252;
wire [512:0] u_ca_in_253;
wire [512:0] u_ca_in_254;
wire [512:0] u_ca_in_255;
wire [512:0] u_ca_in_256;
wire [512:0] u_ca_in_257;
wire [512:0] u_ca_in_258;
wire [512:0] u_ca_in_259;
wire [512:0] u_ca_in_260;
wire [512:0] u_ca_in_261;
wire [512:0] u_ca_in_262;
wire [512:0] u_ca_in_263;
wire [512:0] u_ca_in_264;
wire [512:0] u_ca_in_265;
wire [512:0] u_ca_in_266;
wire [512:0] u_ca_in_267;
wire [512:0] u_ca_in_268;
wire [512:0] u_ca_in_269;
wire [512:0] u_ca_in_270;
wire [512:0] u_ca_in_271;
wire [512:0] u_ca_in_272;
wire [512:0] u_ca_in_273;
wire [512:0] u_ca_in_274;
wire [512:0] u_ca_in_275;
wire [512:0] u_ca_in_276;
wire [512:0] u_ca_in_277;
wire [512:0] u_ca_in_278;
wire [512:0] u_ca_in_279;
wire [512:0] u_ca_in_280;
wire [512:0] u_ca_in_281;
wire [512:0] u_ca_in_282;
wire [512:0] u_ca_in_283;
wire [512:0] u_ca_in_284;
wire [512:0] u_ca_in_285;
wire [512:0] u_ca_in_286;
wire [512:0] u_ca_in_287;
wire [512:0] u_ca_in_288;
wire [512:0] u_ca_in_289;
wire [512:0] u_ca_in_290;
wire [512:0] u_ca_in_291;
wire [512:0] u_ca_in_292;
wire [512:0] u_ca_in_293;
wire [512:0] u_ca_in_294;
wire [512:0] u_ca_in_295;
wire [512:0] u_ca_in_296;
wire [512:0] u_ca_in_297;
wire [512:0] u_ca_in_298;
wire [512:0] u_ca_in_299;
wire [512:0] u_ca_in_300;
wire [512:0] u_ca_in_301;
wire [512:0] u_ca_in_302;
wire [512:0] u_ca_in_303;
wire [512:0] u_ca_in_304;
wire [512:0] u_ca_in_305;
wire [512:0] u_ca_in_306;
wire [512:0] u_ca_in_307;
wire [512:0] u_ca_in_308;
wire [512:0] u_ca_in_309;
wire [512:0] u_ca_in_310;
wire [512:0] u_ca_in_311;
wire [512:0] u_ca_in_312;
wire [512:0] u_ca_in_313;
wire [512:0] u_ca_in_314;
wire [512:0] u_ca_in_315;
wire [512:0] u_ca_in_316;
wire [512:0] u_ca_in_317;
wire [512:0] u_ca_in_318;
wire [512:0] u_ca_in_319;
wire [512:0] u_ca_in_320;
wire [512:0] u_ca_in_321;
wire [512:0] u_ca_in_322;
wire [512:0] u_ca_in_323;
wire [512:0] u_ca_in_324;
wire [512:0] u_ca_in_325;
wire [512:0] u_ca_in_326;
wire [512:0] u_ca_in_327;
wire [512:0] u_ca_in_328;
wire [512:0] u_ca_in_329;
wire [512:0] u_ca_in_330;
wire [512:0] u_ca_in_331;
wire [512:0] u_ca_in_332;
wire [512:0] u_ca_in_333;
wire [512:0] u_ca_in_334;
wire [512:0] u_ca_in_335;
wire [512:0] u_ca_in_336;
wire [512:0] u_ca_in_337;
wire [512:0] u_ca_in_338;
wire [512:0] u_ca_in_339;
wire [512:0] u_ca_in_340;
wire [512:0] u_ca_in_341;
wire [512:0] u_ca_in_342;
wire [512:0] u_ca_in_343;
wire [512:0] u_ca_in_344;
wire [512:0] u_ca_in_345;
wire [512:0] u_ca_in_346;
wire [512:0] u_ca_in_347;
wire [512:0] u_ca_in_348;
wire [512:0] u_ca_in_349;
wire [512:0] u_ca_in_350;
wire [512:0] u_ca_in_351;
wire [512:0] u_ca_in_352;
wire [512:0] u_ca_in_353;
wire [512:0] u_ca_in_354;
wire [512:0] u_ca_in_355;
wire [512:0] u_ca_in_356;
wire [512:0] u_ca_in_357;
wire [512:0] u_ca_in_358;
wire [512:0] u_ca_in_359;
wire [512:0] u_ca_in_360;
wire [512:0] u_ca_in_361;
wire [512:0] u_ca_in_362;
wire [512:0] u_ca_in_363;
wire [512:0] u_ca_in_364;
wire [512:0] u_ca_in_365;
wire [512:0] u_ca_in_366;
wire [512:0] u_ca_in_367;
wire [512:0] u_ca_in_368;
wire [512:0] u_ca_in_369;
wire [512:0] u_ca_in_370;
wire [512:0] u_ca_in_371;
wire [512:0] u_ca_in_372;
wire [512:0] u_ca_in_373;
wire [512:0] u_ca_in_374;
wire [512:0] u_ca_in_375;
wire [512:0] u_ca_in_376;
wire [512:0] u_ca_in_377;
wire [512:0] u_ca_in_378;
wire [512:0] u_ca_in_379;
wire [512:0] u_ca_in_380;
wire [512:0] u_ca_in_381;
wire [512:0] u_ca_in_382;
wire [512:0] u_ca_in_383;
wire [512:0] u_ca_in_384;
wire [512:0] u_ca_in_385;
wire [512:0] u_ca_in_386;
wire [512:0] u_ca_in_387;
wire [512:0] u_ca_in_388;
wire [512:0] u_ca_in_389;
wire [512:0] u_ca_in_390;
wire [512:0] u_ca_in_391;
wire [512:0] u_ca_in_392;
wire [512:0] u_ca_in_393;
wire [512:0] u_ca_in_394;
wire [512:0] u_ca_in_395;
wire [512:0] u_ca_in_396;
wire [512:0] u_ca_in_397;
wire [512:0] u_ca_in_398;
wire [512:0] u_ca_in_399;
wire [512:0] u_ca_in_400;
wire [512:0] u_ca_in_401;
wire [512:0] u_ca_in_402;
wire [512:0] u_ca_in_403;
wire [512:0] u_ca_in_404;
wire [512:0] u_ca_in_405;
wire [512:0] u_ca_in_406;
wire [512:0] u_ca_in_407;
wire [512:0] u_ca_in_408;
wire [512:0] u_ca_in_409;
wire [512:0] u_ca_in_410;
wire [512:0] u_ca_in_411;
wire [512:0] u_ca_in_412;
wire [512:0] u_ca_in_413;
wire [512:0] u_ca_in_414;
wire [512:0] u_ca_in_415;
wire [512:0] u_ca_in_416;
wire [512:0] u_ca_in_417;
wire [512:0] u_ca_in_418;
wire [512:0] u_ca_in_419;
wire [512:0] u_ca_in_420;
wire [512:0] u_ca_in_421;
wire [512:0] u_ca_in_422;
wire [512:0] u_ca_in_423;
wire [512:0] u_ca_in_424;
wire [512:0] u_ca_in_425;
wire [512:0] u_ca_in_426;
wire [512:0] u_ca_in_427;
wire [512:0] u_ca_in_428;
wire [512:0] u_ca_in_429;
wire [512:0] u_ca_in_430;
wire [512:0] u_ca_in_431;
wire [512:0] u_ca_in_432;
wire [512:0] u_ca_in_433;
wire [512:0] u_ca_in_434;
wire [512:0] u_ca_in_435;
wire [512:0] u_ca_in_436;
wire [512:0] u_ca_in_437;
wire [512:0] u_ca_in_438;
wire [512:0] u_ca_in_439;
wire [512:0] u_ca_in_440;
wire [512:0] u_ca_in_441;
wire [512:0] u_ca_in_442;
wire [512:0] u_ca_in_443;
wire [512:0] u_ca_in_444;
wire [512:0] u_ca_in_445;
wire [512:0] u_ca_in_446;
wire [512:0] u_ca_in_447;
wire [512:0] u_ca_in_448;
wire [512:0] u_ca_in_449;
wire [512:0] u_ca_in_450;
wire [512:0] u_ca_in_451;
wire [512:0] u_ca_in_452;
wire [512:0] u_ca_in_453;
wire [512:0] u_ca_in_454;
wire [512:0] u_ca_in_455;
wire [512:0] u_ca_in_456;
wire [512:0] u_ca_in_457;
wire [512:0] u_ca_in_458;
wire [512:0] u_ca_in_459;
wire [512:0] u_ca_in_460;
wire [512:0] u_ca_in_461;
wire [512:0] u_ca_in_462;
wire [512:0] u_ca_in_463;
wire [512:0] u_ca_in_464;
wire [512:0] u_ca_in_465;
wire [512:0] u_ca_in_466;
wire [512:0] u_ca_in_467;
wire [512:0] u_ca_in_468;
wire [512:0] u_ca_in_469;
wire [512:0] u_ca_in_470;
wire [512:0] u_ca_in_471;
wire [512:0] u_ca_in_472;
wire [512:0] u_ca_in_473;
wire [512:0] u_ca_in_474;
wire [512:0] u_ca_in_475;
wire [512:0] u_ca_in_476;
wire [512:0] u_ca_in_477;
wire [512:0] u_ca_in_478;
wire [512:0] u_ca_in_479;
wire [512:0] u_ca_in_480;
wire [512:0] u_ca_in_481;
wire [512:0] u_ca_in_482;
wire [512:0] u_ca_in_483;
wire [512:0] u_ca_in_484;
wire [512:0] u_ca_in_485;
wire [512:0] u_ca_in_486;
wire [512:0] u_ca_in_487;
wire [512:0] u_ca_in_488;
wire [512:0] u_ca_in_489;
wire [512:0] u_ca_in_490;
wire [512:0] u_ca_in_491;
wire [512:0] u_ca_in_492;
wire [512:0] u_ca_in_493;
wire [512:0] u_ca_in_494;
wire [512:0] u_ca_in_495;
wire [512:0] u_ca_in_496;
wire [512:0] u_ca_in_497;
wire [512:0] u_ca_in_498;
wire [512:0] u_ca_in_499;
wire [512:0] u_ca_in_500;
wire [512:0] u_ca_in_501;
wire [512:0] u_ca_in_502;
wire [512:0] u_ca_in_503;
wire [512:0] u_ca_in_504;
wire [512:0] u_ca_in_505;
wire [512:0] u_ca_in_506;
wire [512:0] u_ca_in_507;
wire [512:0] u_ca_in_508;
wire [512:0] u_ca_in_509;
wire [512:0] u_ca_in_510;
wire [512:0] u_ca_in_511;
wire [512:0] u_ca_in_512;
wire [512:0] u_ca_in_513;
wire [512:0] u_ca_in_514;
wire [512:0] u_ca_in_515;
wire [512:0] u_ca_in_516;
wire [512:0] u_ca_in_517;
wire [512:0] u_ca_in_518;
wire [512:0] u_ca_in_519;
wire [512:0] u_ca_in_520;
wire [512:0] u_ca_in_521;
wire [512:0] u_ca_in_522;
wire [512:0] u_ca_in_523;
wire [512:0] u_ca_in_524;
wire [512:0] u_ca_in_525;
wire [512:0] u_ca_in_526;
wire [512:0] u_ca_in_527;
wire [512:0] u_ca_in_528;
wire [512:0] u_ca_in_529;
wire [512:0] u_ca_in_530;
wire [512:0] u_ca_in_531;
wire [512:0] u_ca_in_532;
wire [512:0] u_ca_in_533;
wire [512:0] u_ca_in_534;
wire [512:0] u_ca_in_535;
wire [512:0] u_ca_in_536;
wire [512:0] u_ca_in_537;
wire [512:0] u_ca_in_538;
wire [512:0] u_ca_in_539;
wire [512:0] u_ca_in_540;
wire [512:0] u_ca_in_541;
wire [512:0] u_ca_in_542;
wire [512:0] u_ca_in_543;
wire [512:0] u_ca_in_544;
wire [512:0] u_ca_in_545;
wire [512:0] u_ca_in_546;
wire [512:0] u_ca_in_547;
wire [512:0] u_ca_in_548;
wire [512:0] u_ca_in_549;
wire [512:0] u_ca_in_550;
wire [512:0] u_ca_in_551;
wire [512:0] u_ca_in_552;
wire [512:0] u_ca_in_553;
wire [512:0] u_ca_in_554;
wire [512:0] u_ca_in_555;
wire [512:0] u_ca_in_556;
wire [512:0] u_ca_in_557;
wire [512:0] u_ca_in_558;
wire [512:0] u_ca_in_559;
wire [512:0] u_ca_in_560;
wire [512:0] u_ca_in_561;
wire [512:0] u_ca_in_562;
wire [512:0] u_ca_in_563;
wire [512:0] u_ca_in_564;
wire [512:0] u_ca_in_565;
wire [512:0] u_ca_in_566;
wire [512:0] u_ca_in_567;
wire [512:0] u_ca_in_568;
wire [512:0] u_ca_in_569;
wire [512:0] u_ca_in_570;
wire [512:0] u_ca_in_571;
wire [512:0] u_ca_in_572;
wire [512:0] u_ca_in_573;
wire [512:0] u_ca_in_574;
wire [512:0] u_ca_in_575;
wire [512:0] u_ca_in_576;
wire [512:0] u_ca_in_577;
wire [512:0] u_ca_in_578;
wire [512:0] u_ca_in_579;
wire [512:0] u_ca_in_580;
wire [512:0] u_ca_in_581;
wire [512:0] u_ca_in_582;
wire [512:0] u_ca_in_583;
wire [512:0] u_ca_in_584;
wire [512:0] u_ca_in_585;
wire [512:0] u_ca_in_586;
wire [512:0] u_ca_in_587;
wire [512:0] u_ca_in_588;
wire [512:0] u_ca_in_589;
wire [512:0] u_ca_in_590;
wire [512:0] u_ca_in_591;
wire [512:0] u_ca_in_592;
wire [512:0] u_ca_in_593;
wire [512:0] u_ca_in_594;
wire [512:0] u_ca_in_595;
wire [512:0] u_ca_in_596;
wire [512:0] u_ca_in_597;
wire [512:0] u_ca_in_598;
wire [512:0] u_ca_in_599;
wire [512:0] u_ca_in_600;
wire [512:0] u_ca_in_601;
wire [512:0] u_ca_in_602;
wire [512:0] u_ca_in_603;
wire [512:0] u_ca_in_604;
wire [512:0] u_ca_in_605;
wire [512:0] u_ca_in_606;
wire [512:0] u_ca_in_607;
wire [512:0] u_ca_in_608;
wire [512:0] u_ca_in_609;
wire [512:0] u_ca_in_610;
wire [512:0] u_ca_in_611;
wire [512:0] u_ca_in_612;
wire [512:0] u_ca_in_613;
wire [512:0] u_ca_in_614;
wire [512:0] u_ca_in_615;
wire [512:0] u_ca_in_616;
wire [512:0] u_ca_in_617;
wire [512:0] u_ca_in_618;
wire [512:0] u_ca_in_619;
wire [512:0] u_ca_in_620;
wire [512:0] u_ca_in_621;
wire [512:0] u_ca_in_622;
wire [512:0] u_ca_in_623;
wire [512:0] u_ca_in_624;
wire [512:0] u_ca_in_625;
wire [512:0] u_ca_in_626;
wire [512:0] u_ca_in_627;
wire [512:0] u_ca_in_628;
wire [512:0] u_ca_in_629;
wire [512:0] u_ca_in_630;
wire [512:0] u_ca_in_631;
wire [512:0] u_ca_in_632;
wire [512:0] u_ca_in_633;
wire [512:0] u_ca_in_634;
wire [512:0] u_ca_in_635;
wire [512:0] u_ca_in_636;
wire [512:0] u_ca_in_637;
wire [512:0] u_ca_in_638;
wire [512:0] u_ca_in_639;
wire [512:0] u_ca_in_640;
wire [512:0] u_ca_in_641;
wire [512:0] u_ca_in_642;
wire [512:0] u_ca_in_643;
wire [512:0] u_ca_in_644;
wire [512:0] u_ca_in_645;
wire [512:0] u_ca_in_646;
wire [512:0] u_ca_in_647;
wire [512:0] u_ca_in_648;
wire [512:0] u_ca_in_649;
wire [512:0] u_ca_in_650;
wire [512:0] u_ca_in_651;
wire [512:0] u_ca_in_652;
wire [512:0] u_ca_in_653;
wire [512:0] u_ca_in_654;
wire [512:0] u_ca_in_655;
wire [512:0] u_ca_in_656;
wire [512:0] u_ca_in_657;
wire [512:0] u_ca_in_658;
wire [512:0] u_ca_in_659;
wire [512:0] u_ca_in_660;
wire [512:0] u_ca_in_661;
wire [512:0] u_ca_in_662;
wire [512:0] u_ca_in_663;
wire [512:0] u_ca_in_664;
wire [512:0] u_ca_in_665;
wire [512:0] u_ca_in_666;
wire [512:0] u_ca_in_667;
wire [512:0] u_ca_in_668;
wire [512:0] u_ca_in_669;
wire [512:0] u_ca_in_670;
wire [512:0] u_ca_in_671;
wire [512:0] u_ca_in_672;
wire [512:0] u_ca_in_673;
wire [512:0] u_ca_in_674;
wire [512:0] u_ca_in_675;
wire [512:0] u_ca_in_676;
wire [512:0] u_ca_in_677;
wire [512:0] u_ca_in_678;
wire [512:0] u_ca_in_679;
wire [512:0] u_ca_in_680;
wire [512:0] u_ca_in_681;
wire [512:0] u_ca_in_682;
wire [512:0] u_ca_in_683;
wire [512:0] u_ca_in_684;
wire [512:0] u_ca_in_685;
wire [512:0] u_ca_in_686;
wire [512:0] u_ca_in_687;
wire [512:0] u_ca_in_688;
wire [512:0] u_ca_in_689;
wire [512:0] u_ca_in_690;
wire [512:0] u_ca_in_691;
wire [512:0] u_ca_in_692;
wire [512:0] u_ca_in_693;
wire [512:0] u_ca_in_694;
wire [512:0] u_ca_in_695;
wire [512:0] u_ca_in_696;
wire [512:0] u_ca_in_697;
wire [512:0] u_ca_in_698;
wire [512:0] u_ca_in_699;
wire [512:0] u_ca_in_700;
wire [512:0] u_ca_in_701;
wire [512:0] u_ca_in_702;
wire [512:0] u_ca_in_703;
wire [512:0] u_ca_in_704;
wire [512:0] u_ca_in_705;
wire [512:0] u_ca_in_706;
wire [512:0] u_ca_in_707;
wire [512:0] u_ca_in_708;
wire [512:0] u_ca_in_709;
wire [512:0] u_ca_in_710;
wire [512:0] u_ca_in_711;
wire [512:0] u_ca_in_712;
wire [512:0] u_ca_in_713;
wire [512:0] u_ca_in_714;
wire [512:0] u_ca_in_715;
wire [512:0] u_ca_in_716;
wire [512:0] u_ca_in_717;
wire [512:0] u_ca_in_718;
wire [512:0] u_ca_in_719;
wire [512:0] u_ca_in_720;
wire [512:0] u_ca_in_721;
wire [512:0] u_ca_in_722;
wire [512:0] u_ca_in_723;
wire [512:0] u_ca_in_724;
wire [512:0] u_ca_in_725;
wire [512:0] u_ca_in_726;
wire [512:0] u_ca_in_727;
wire [512:0] u_ca_in_728;
wire [512:0] u_ca_in_729;
wire [512:0] u_ca_in_730;
wire [512:0] u_ca_in_731;
wire [512:0] u_ca_in_732;
wire [512:0] u_ca_in_733;
wire [512:0] u_ca_in_734;
wire [512:0] u_ca_in_735;
wire [512:0] u_ca_in_736;
wire [512:0] u_ca_in_737;
wire [512:0] u_ca_in_738;
wire [512:0] u_ca_in_739;
wire [512:0] u_ca_in_740;
wire [512:0] u_ca_in_741;
wire [512:0] u_ca_in_742;
wire [512:0] u_ca_in_743;
wire [512:0] u_ca_in_744;
wire [512:0] u_ca_in_745;
wire [512:0] u_ca_in_746;
wire [512:0] u_ca_in_747;
wire [512:0] u_ca_in_748;
wire [512:0] u_ca_in_749;
wire [512:0] u_ca_in_750;
wire [512:0] u_ca_in_751;
wire [512:0] u_ca_in_752;
wire [512:0] u_ca_in_753;
wire [512:0] u_ca_in_754;
wire [512:0] u_ca_in_755;
wire [512:0] u_ca_in_756;
wire [512:0] u_ca_in_757;
wire [512:0] u_ca_in_758;
wire [512:0] u_ca_in_759;
wire [512:0] u_ca_in_760;
wire [512:0] u_ca_in_761;
wire [512:0] u_ca_in_762;
wire [512:0] u_ca_in_763;
wire [512:0] u_ca_in_764;
wire [512:0] u_ca_in_765;
wire [512:0] u_ca_in_766;
wire [512:0] u_ca_in_767;
wire [512:0] u_ca_in_768;
wire [512:0] u_ca_in_769;
wire [512:0] u_ca_in_770;
wire [512:0] u_ca_in_771;
wire [512:0] u_ca_in_772;
wire [512:0] u_ca_in_773;
wire [512:0] u_ca_in_774;
wire [512:0] u_ca_in_775;
wire [512:0] u_ca_in_776;
wire [512:0] u_ca_in_777;
wire [512:0] u_ca_in_778;
wire [512:0] u_ca_in_779;
wire [512:0] u_ca_in_780;
wire [512:0] u_ca_in_781;
wire [512:0] u_ca_in_782;
wire [512:0] u_ca_in_783;
wire [512:0] u_ca_in_784;
wire [512:0] u_ca_in_785;
wire [512:0] u_ca_in_786;
wire [512:0] u_ca_in_787;
wire [512:0] u_ca_in_788;
wire [512:0] u_ca_in_789;
wire [512:0] u_ca_in_790;
wire [512:0] u_ca_in_791;
wire [512:0] u_ca_in_792;
wire [512:0] u_ca_in_793;
wire [512:0] u_ca_in_794;
wire [512:0] u_ca_in_795;
wire [512:0] u_ca_in_796;
wire [512:0] u_ca_in_797;
wire [512:0] u_ca_in_798;
wire [512:0] u_ca_in_799;
wire [512:0] u_ca_in_800;
wire [512:0] u_ca_in_801;
wire [512:0] u_ca_in_802;
wire [512:0] u_ca_in_803;
wire [512:0] u_ca_in_804;
wire [512:0] u_ca_in_805;
wire [512:0] u_ca_in_806;
wire [512:0] u_ca_in_807;
wire [512:0] u_ca_in_808;
wire [512:0] u_ca_in_809;
wire [512:0] u_ca_in_810;
wire [512:0] u_ca_in_811;
wire [512:0] u_ca_in_812;
wire [512:0] u_ca_in_813;
wire [512:0] u_ca_in_814;
wire [512:0] u_ca_in_815;
wire [512:0] u_ca_in_816;
wire [512:0] u_ca_in_817;
wire [512:0] u_ca_in_818;
wire [512:0] u_ca_in_819;
wire [512:0] u_ca_in_820;
wire [512:0] u_ca_in_821;
wire [512:0] u_ca_in_822;
wire [512:0] u_ca_in_823;
wire [512:0] u_ca_in_824;
wire [512:0] u_ca_in_825;
wire [512:0] u_ca_in_826;
wire [512:0] u_ca_in_827;
wire [512:0] u_ca_in_828;
wire [512:0] u_ca_in_829;
wire [512:0] u_ca_in_830;
wire [512:0] u_ca_in_831;
wire [512:0] u_ca_in_832;
wire [512:0] u_ca_in_833;
wire [512:0] u_ca_in_834;
wire [512:0] u_ca_in_835;
wire [512:0] u_ca_in_836;
wire [512:0] u_ca_in_837;
wire [512:0] u_ca_in_838;
wire [512:0] u_ca_in_839;
wire [512:0] u_ca_in_840;
wire [512:0] u_ca_in_841;
wire [512:0] u_ca_in_842;
wire [512:0] u_ca_in_843;
wire [512:0] u_ca_in_844;
wire [512:0] u_ca_in_845;
wire [512:0] u_ca_in_846;
wire [512:0] u_ca_in_847;
wire [512:0] u_ca_in_848;
wire [512:0] u_ca_in_849;
wire [512:0] u_ca_in_850;
wire [512:0] u_ca_in_851;
wire [512:0] u_ca_in_852;
wire [512:0] u_ca_in_853;
wire [512:0] u_ca_in_854;
wire [512:0] u_ca_in_855;
wire [512:0] u_ca_in_856;
wire [512:0] u_ca_in_857;
wire [512:0] u_ca_in_858;
wire [512:0] u_ca_in_859;
wire [512:0] u_ca_in_860;
wire [512:0] u_ca_in_861;
wire [512:0] u_ca_in_862;
wire [512:0] u_ca_in_863;
wire [512:0] u_ca_in_864;
wire [512:0] u_ca_in_865;
wire [512:0] u_ca_in_866;
wire [512:0] u_ca_in_867;
wire [512:0] u_ca_in_868;
wire [512:0] u_ca_in_869;
wire [512:0] u_ca_in_870;
wire [512:0] u_ca_in_871;
wire [512:0] u_ca_in_872;
wire [512:0] u_ca_in_873;
wire [512:0] u_ca_in_874;
wire [512:0] u_ca_in_875;
wire [512:0] u_ca_in_876;
wire [512:0] u_ca_in_877;
wire [512:0] u_ca_in_878;
wire [512:0] u_ca_in_879;
wire [512:0] u_ca_in_880;
wire [512:0] u_ca_in_881;
wire [512:0] u_ca_in_882;
wire [512:0] u_ca_in_883;
wire [512:0] u_ca_in_884;
wire [512:0] u_ca_in_885;
wire [512:0] u_ca_in_886;
wire [512:0] u_ca_in_887;
wire [512:0] u_ca_in_888;
wire [512:0] u_ca_in_889;
wire [512:0] u_ca_in_890;
wire [512:0] u_ca_in_891;
wire [512:0] u_ca_in_892;
wire [512:0] u_ca_in_893;
wire [512:0] u_ca_in_894;
wire [512:0] u_ca_in_895;
wire [512:0] u_ca_in_896;
wire [512:0] u_ca_in_897;
wire [512:0] u_ca_in_898;
wire [512:0] u_ca_in_899;
wire [512:0] u_ca_in_900;
wire [512:0] u_ca_in_901;
wire [512:0] u_ca_in_902;
wire [512:0] u_ca_in_903;
wire [512:0] u_ca_in_904;
wire [512:0] u_ca_in_905;
wire [512:0] u_ca_in_906;
wire [512:0] u_ca_in_907;
wire [512:0] u_ca_in_908;
wire [512:0] u_ca_in_909;
wire [512:0] u_ca_in_910;
wire [512:0] u_ca_in_911;
wire [512:0] u_ca_in_912;
wire [512:0] u_ca_in_913;
wire [512:0] u_ca_in_914;
wire [512:0] u_ca_in_915;
wire [512:0] u_ca_in_916;
wire [512:0] u_ca_in_917;
wire [512:0] u_ca_in_918;
wire [512:0] u_ca_in_919;
wire [512:0] u_ca_in_920;
wire [512:0] u_ca_in_921;
wire [512:0] u_ca_in_922;
wire [512:0] u_ca_in_923;
wire [512:0] u_ca_in_924;
wire [512:0] u_ca_in_925;
wire [512:0] u_ca_in_926;
wire [512:0] u_ca_in_927;
wire [512:0] u_ca_in_928;
wire [512:0] u_ca_in_929;
wire [512:0] u_ca_in_930;
wire [512:0] u_ca_in_931;
wire [512:0] u_ca_in_932;
wire [512:0] u_ca_in_933;
wire [512:0] u_ca_in_934;
wire [512:0] u_ca_in_935;
wire [512:0] u_ca_in_936;
wire [512:0] u_ca_in_937;
wire [512:0] u_ca_in_938;
wire [512:0] u_ca_in_939;
wire [512:0] u_ca_in_940;
wire [512:0] u_ca_in_941;
wire [512:0] u_ca_in_942;
wire [512:0] u_ca_in_943;
wire [512:0] u_ca_in_944;
wire [512:0] u_ca_in_945;
wire [512:0] u_ca_in_946;
wire [512:0] u_ca_in_947;
wire [512:0] u_ca_in_948;
wire [512:0] u_ca_in_949;
wire [512:0] u_ca_in_950;
wire [512:0] u_ca_in_951;
wire [512:0] u_ca_in_952;
wire [512:0] u_ca_in_953;
wire [512:0] u_ca_in_954;
wire [512:0] u_ca_in_955;
wire [512:0] u_ca_in_956;
wire [512:0] u_ca_in_957;
wire [512:0] u_ca_in_958;
wire [512:0] u_ca_in_959;
wire [512:0] u_ca_in_960;
wire [512:0] u_ca_in_961;
wire [512:0] u_ca_in_962;
wire [512:0] u_ca_in_963;
wire [512:0] u_ca_in_964;
wire [512:0] u_ca_in_965;
wire [512:0] u_ca_in_966;
wire [512:0] u_ca_in_967;
wire [512:0] u_ca_in_968;
wire [512:0] u_ca_in_969;
wire [512:0] u_ca_in_970;
wire [512:0] u_ca_in_971;
wire [512:0] u_ca_in_972;
wire [512:0] u_ca_in_973;
wire [512:0] u_ca_in_974;
wire [512:0] u_ca_in_975;
wire [512:0] u_ca_in_976;
wire [512:0] u_ca_in_977;
wire [512:0] u_ca_in_978;
wire [512:0] u_ca_in_979;
wire [512:0] u_ca_in_980;
wire [512:0] u_ca_in_981;
wire [512:0] u_ca_in_982;
wire [512:0] u_ca_in_983;
wire [512:0] u_ca_in_984;
wire [512:0] u_ca_in_985;
wire [512:0] u_ca_in_986;
wire [512:0] u_ca_in_987;
wire [512:0] u_ca_in_988;
wire [512:0] u_ca_in_989;
wire [512:0] u_ca_in_990;
wire [512:0] u_ca_in_991;
wire [512:0] u_ca_in_992;
wire [512:0] u_ca_in_993;
wire [512:0] u_ca_in_994;
wire [512:0] u_ca_in_995;
wire [512:0] u_ca_in_996;
wire [512:0] u_ca_in_997;
wire [512:0] u_ca_in_998;
wire [512:0] u_ca_in_999;
wire [512:0] u_ca_in_1000;
wire [512:0] u_ca_in_1001;
wire [512:0] u_ca_in_1002;
wire [512:0] u_ca_in_1003;
wire [512:0] u_ca_in_1004;
wire [512:0] u_ca_in_1005;
wire [512:0] u_ca_in_1006;
wire [512:0] u_ca_in_1007;
wire [512:0] u_ca_in_1008;
wire [512:0] u_ca_in_1009;
wire [512:0] u_ca_in_1010;
wire [512:0] u_ca_in_1011;
wire [512:0] u_ca_in_1012;
wire [512:0] u_ca_in_1013;
wire [512:0] u_ca_in_1014;
wire [512:0] u_ca_in_1015;
wire [512:0] u_ca_in_1016;
wire [512:0] u_ca_in_1017;
wire [512:0] u_ca_in_1018;
wire [512:0] u_ca_in_1019;
wire [512:0] u_ca_in_1020;
wire [512:0] u_ca_in_1021;
wire [512:0] u_ca_in_1022;
wire [512:0] u_ca_in_1023;
wire [151:0] u_ca_out_0;
wire [151:0] u_ca_out_1;
wire [151:0] u_ca_out_2;
wire [151:0] u_ca_out_3;
wire [151:0] u_ca_out_4;
wire [151:0] u_ca_out_5;
wire [151:0] u_ca_out_6;
wire [151:0] u_ca_out_7;
wire [151:0] u_ca_out_8;
wire [151:0] u_ca_out_9;
wire [151:0] u_ca_out_10;
wire [151:0] u_ca_out_11;
wire [151:0] u_ca_out_12;
wire [151:0] u_ca_out_13;
wire [151:0] u_ca_out_14;
wire [151:0] u_ca_out_15;
wire [151:0] u_ca_out_16;
wire [151:0] u_ca_out_17;
wire [151:0] u_ca_out_18;
wire [151:0] u_ca_out_19;
wire [151:0] u_ca_out_20;
wire [151:0] u_ca_out_21;
wire [151:0] u_ca_out_22;
wire [151:0] u_ca_out_23;
wire [151:0] u_ca_out_24;
wire [151:0] u_ca_out_25;
wire [151:0] u_ca_out_26;
wire [151:0] u_ca_out_27;
wire [151:0] u_ca_out_28;
wire [151:0] u_ca_out_29;
wire [151:0] u_ca_out_30;
wire [151:0] u_ca_out_31;
wire [151:0] u_ca_out_32;
wire [151:0] u_ca_out_33;
wire [151:0] u_ca_out_34;
wire [151:0] u_ca_out_35;
wire [151:0] u_ca_out_36;
wire [151:0] u_ca_out_37;
wire [151:0] u_ca_out_38;
wire [151:0] u_ca_out_39;
wire [151:0] u_ca_out_40;
wire [151:0] u_ca_out_41;
wire [151:0] u_ca_out_42;
wire [151:0] u_ca_out_43;
wire [151:0] u_ca_out_44;
wire [151:0] u_ca_out_45;
wire [151:0] u_ca_out_46;
wire [151:0] u_ca_out_47;
wire [151:0] u_ca_out_48;
wire [151:0] u_ca_out_49;
wire [151:0] u_ca_out_50;
wire [151:0] u_ca_out_51;
wire [151:0] u_ca_out_52;
wire [151:0] u_ca_out_53;
wire [151:0] u_ca_out_54;
wire [151:0] u_ca_out_55;
wire [151:0] u_ca_out_56;
wire [151:0] u_ca_out_57;
wire [151:0] u_ca_out_58;
wire [151:0] u_ca_out_59;
wire [151:0] u_ca_out_60;
wire [151:0] u_ca_out_61;
wire [151:0] u_ca_out_62;
wire [151:0] u_ca_out_63;
wire [151:0] u_ca_out_64;
wire [151:0] u_ca_out_65;
wire [151:0] u_ca_out_66;
wire [151:0] u_ca_out_67;
wire [151:0] u_ca_out_68;
wire [151:0] u_ca_out_69;
wire [151:0] u_ca_out_70;
wire [151:0] u_ca_out_71;
wire [151:0] u_ca_out_72;
wire [151:0] u_ca_out_73;
wire [151:0] u_ca_out_74;
wire [151:0] u_ca_out_75;
wire [151:0] u_ca_out_76;
wire [151:0] u_ca_out_77;
wire [151:0] u_ca_out_78;
wire [151:0] u_ca_out_79;
wire [151:0] u_ca_out_80;
wire [151:0] u_ca_out_81;
wire [151:0] u_ca_out_82;
wire [151:0] u_ca_out_83;
wire [151:0] u_ca_out_84;
wire [151:0] u_ca_out_85;
wire [151:0] u_ca_out_86;
wire [151:0] u_ca_out_87;
wire [151:0] u_ca_out_88;
wire [151:0] u_ca_out_89;
wire [151:0] u_ca_out_90;
wire [151:0] u_ca_out_91;
wire [151:0] u_ca_out_92;
wire [151:0] u_ca_out_93;
wire [151:0] u_ca_out_94;
wire [151:0] u_ca_out_95;
wire [151:0] u_ca_out_96;
wire [151:0] u_ca_out_97;
wire [151:0] u_ca_out_98;
wire [151:0] u_ca_out_99;
wire [151:0] u_ca_out_100;
wire [151:0] u_ca_out_101;
wire [151:0] u_ca_out_102;
wire [151:0] u_ca_out_103;
wire [151:0] u_ca_out_104;
wire [151:0] u_ca_out_105;
wire [151:0] u_ca_out_106;
wire [151:0] u_ca_out_107;
wire [151:0] u_ca_out_108;
wire [151:0] u_ca_out_109;
wire [151:0] u_ca_out_110;
wire [151:0] u_ca_out_111;
wire [151:0] u_ca_out_112;
wire [151:0] u_ca_out_113;
wire [151:0] u_ca_out_114;
wire [151:0] u_ca_out_115;
wire [151:0] u_ca_out_116;
wire [151:0] u_ca_out_117;
wire [151:0] u_ca_out_118;
wire [151:0] u_ca_out_119;
wire [151:0] u_ca_out_120;
wire [151:0] u_ca_out_121;
wire [151:0] u_ca_out_122;
wire [151:0] u_ca_out_123;
wire [151:0] u_ca_out_124;
wire [151:0] u_ca_out_125;
wire [151:0] u_ca_out_126;
wire [151:0] u_ca_out_127;
wire [151:0] u_ca_out_128;
wire [151:0] u_ca_out_129;
wire [151:0] u_ca_out_130;
wire [151:0] u_ca_out_131;
wire [151:0] u_ca_out_132;
wire [151:0] u_ca_out_133;
wire [151:0] u_ca_out_134;
wire [151:0] u_ca_out_135;
wire [151:0] u_ca_out_136;
wire [151:0] u_ca_out_137;
wire [151:0] u_ca_out_138;
wire [151:0] u_ca_out_139;
wire [151:0] u_ca_out_140;
wire [151:0] u_ca_out_141;
wire [151:0] u_ca_out_142;
wire [151:0] u_ca_out_143;
wire [151:0] u_ca_out_144;
wire [151:0] u_ca_out_145;
wire [151:0] u_ca_out_146;
wire [151:0] u_ca_out_147;
wire [151:0] u_ca_out_148;
wire [151:0] u_ca_out_149;
wire [151:0] u_ca_out_150;
wire [151:0] u_ca_out_151;
wire [151:0] u_ca_out_152;
wire [151:0] u_ca_out_153;
wire [151:0] u_ca_out_154;
wire [151:0] u_ca_out_155;
wire [151:0] u_ca_out_156;
wire [151:0] u_ca_out_157;
wire [151:0] u_ca_out_158;
wire [151:0] u_ca_out_159;
wire [151:0] u_ca_out_160;
wire [151:0] u_ca_out_161;
wire [151:0] u_ca_out_162;
wire [151:0] u_ca_out_163;
wire [151:0] u_ca_out_164;
wire [151:0] u_ca_out_165;
wire [151:0] u_ca_out_166;
wire [151:0] u_ca_out_167;
wire [151:0] u_ca_out_168;
wire [151:0] u_ca_out_169;
wire [151:0] u_ca_out_170;
wire [151:0] u_ca_out_171;
wire [151:0] u_ca_out_172;
wire [151:0] u_ca_out_173;
wire [151:0] u_ca_out_174;
wire [151:0] u_ca_out_175;
wire [151:0] u_ca_out_176;
wire [151:0] u_ca_out_177;
wire [151:0] u_ca_out_178;
wire [151:0] u_ca_out_179;
wire [151:0] u_ca_out_180;
wire [151:0] u_ca_out_181;
wire [151:0] u_ca_out_182;
wire [151:0] u_ca_out_183;
wire [151:0] u_ca_out_184;
wire [151:0] u_ca_out_185;
wire [151:0] u_ca_out_186;
wire [151:0] u_ca_out_187;
wire [151:0] u_ca_out_188;
wire [151:0] u_ca_out_189;
wire [151:0] u_ca_out_190;
wire [151:0] u_ca_out_191;
wire [151:0] u_ca_out_192;
wire [151:0] u_ca_out_193;
wire [151:0] u_ca_out_194;
wire [151:0] u_ca_out_195;
wire [151:0] u_ca_out_196;
wire [151:0] u_ca_out_197;
wire [151:0] u_ca_out_198;
wire [151:0] u_ca_out_199;
wire [151:0] u_ca_out_200;
wire [151:0] u_ca_out_201;
wire [151:0] u_ca_out_202;
wire [151:0] u_ca_out_203;
wire [151:0] u_ca_out_204;
wire [151:0] u_ca_out_205;
wire [151:0] u_ca_out_206;
wire [151:0] u_ca_out_207;
wire [151:0] u_ca_out_208;
wire [151:0] u_ca_out_209;
wire [151:0] u_ca_out_210;
wire [151:0] u_ca_out_211;
wire [151:0] u_ca_out_212;
wire [151:0] u_ca_out_213;
wire [151:0] u_ca_out_214;
wire [151:0] u_ca_out_215;
wire [151:0] u_ca_out_216;
wire [151:0] u_ca_out_217;
wire [151:0] u_ca_out_218;
wire [151:0] u_ca_out_219;
wire [151:0] u_ca_out_220;
wire [151:0] u_ca_out_221;
wire [151:0] u_ca_out_222;
wire [151:0] u_ca_out_223;
wire [151:0] u_ca_out_224;
wire [151:0] u_ca_out_225;
wire [151:0] u_ca_out_226;
wire [151:0] u_ca_out_227;
wire [151:0] u_ca_out_228;
wire [151:0] u_ca_out_229;
wire [151:0] u_ca_out_230;
wire [151:0] u_ca_out_231;
wire [151:0] u_ca_out_232;
wire [151:0] u_ca_out_233;
wire [151:0] u_ca_out_234;
wire [151:0] u_ca_out_235;
wire [151:0] u_ca_out_236;
wire [151:0] u_ca_out_237;
wire [151:0] u_ca_out_238;
wire [151:0] u_ca_out_239;
wire [151:0] u_ca_out_240;
wire [151:0] u_ca_out_241;
wire [151:0] u_ca_out_242;
wire [151:0] u_ca_out_243;
wire [151:0] u_ca_out_244;
wire [151:0] u_ca_out_245;
wire [151:0] u_ca_out_246;
wire [151:0] u_ca_out_247;
wire [151:0] u_ca_out_248;
wire [151:0] u_ca_out_249;
wire [151:0] u_ca_out_250;
wire [151:0] u_ca_out_251;
wire [151:0] u_ca_out_252;
wire [151:0] u_ca_out_253;
wire [151:0] u_ca_out_254;
wire [151:0] u_ca_out_255;
wire [151:0] u_ca_out_256;
wire [151:0] u_ca_out_257;
wire [151:0] u_ca_out_258;
wire [151:0] u_ca_out_259;
wire [151:0] u_ca_out_260;
wire [151:0] u_ca_out_261;
wire [151:0] u_ca_out_262;
wire [151:0] u_ca_out_263;
wire [151:0] u_ca_out_264;
wire [151:0] u_ca_out_265;
wire [151:0] u_ca_out_266;
wire [151:0] u_ca_out_267;
wire [151:0] u_ca_out_268;
wire [151:0] u_ca_out_269;
wire [151:0] u_ca_out_270;
wire [151:0] u_ca_out_271;
wire [151:0] u_ca_out_272;
wire [151:0] u_ca_out_273;
wire [151:0] u_ca_out_274;
wire [151:0] u_ca_out_275;
wire [151:0] u_ca_out_276;
wire [151:0] u_ca_out_277;
wire [151:0] u_ca_out_278;
wire [151:0] u_ca_out_279;
wire [151:0] u_ca_out_280;
wire [151:0] u_ca_out_281;
wire [151:0] u_ca_out_282;
wire [151:0] u_ca_out_283;
wire [151:0] u_ca_out_284;
wire [151:0] u_ca_out_285;
wire [151:0] u_ca_out_286;
wire [151:0] u_ca_out_287;
wire [151:0] u_ca_out_288;
wire [151:0] u_ca_out_289;
wire [151:0] u_ca_out_290;
wire [151:0] u_ca_out_291;
wire [151:0] u_ca_out_292;
wire [151:0] u_ca_out_293;
wire [151:0] u_ca_out_294;
wire [151:0] u_ca_out_295;
wire [151:0] u_ca_out_296;
wire [151:0] u_ca_out_297;
wire [151:0] u_ca_out_298;
wire [151:0] u_ca_out_299;
wire [151:0] u_ca_out_300;
wire [151:0] u_ca_out_301;
wire [151:0] u_ca_out_302;
wire [151:0] u_ca_out_303;
wire [151:0] u_ca_out_304;
wire [151:0] u_ca_out_305;
wire [151:0] u_ca_out_306;
wire [151:0] u_ca_out_307;
wire [151:0] u_ca_out_308;
wire [151:0] u_ca_out_309;
wire [151:0] u_ca_out_310;
wire [151:0] u_ca_out_311;
wire [151:0] u_ca_out_312;
wire [151:0] u_ca_out_313;
wire [151:0] u_ca_out_314;
wire [151:0] u_ca_out_315;
wire [151:0] u_ca_out_316;
wire [151:0] u_ca_out_317;
wire [151:0] u_ca_out_318;
wire [151:0] u_ca_out_319;
wire [151:0] u_ca_out_320;
wire [151:0] u_ca_out_321;
wire [151:0] u_ca_out_322;
wire [151:0] u_ca_out_323;
wire [151:0] u_ca_out_324;
wire [151:0] u_ca_out_325;
wire [151:0] u_ca_out_326;
wire [151:0] u_ca_out_327;
wire [151:0] u_ca_out_328;
wire [151:0] u_ca_out_329;
wire [151:0] u_ca_out_330;
wire [151:0] u_ca_out_331;
wire [151:0] u_ca_out_332;
wire [151:0] u_ca_out_333;
wire [151:0] u_ca_out_334;
wire [151:0] u_ca_out_335;
wire [151:0] u_ca_out_336;
wire [151:0] u_ca_out_337;
wire [151:0] u_ca_out_338;
wire [151:0] u_ca_out_339;
wire [151:0] u_ca_out_340;
wire [151:0] u_ca_out_341;
wire [151:0] u_ca_out_342;
wire [151:0] u_ca_out_343;
wire [151:0] u_ca_out_344;
wire [151:0] u_ca_out_345;
wire [151:0] u_ca_out_346;
wire [151:0] u_ca_out_347;
wire [151:0] u_ca_out_348;
wire [151:0] u_ca_out_349;
wire [151:0] u_ca_out_350;
wire [151:0] u_ca_out_351;
wire [151:0] u_ca_out_352;
wire [151:0] u_ca_out_353;
wire [151:0] u_ca_out_354;
wire [151:0] u_ca_out_355;
wire [151:0] u_ca_out_356;
wire [151:0] u_ca_out_357;
wire [151:0] u_ca_out_358;
wire [151:0] u_ca_out_359;
wire [151:0] u_ca_out_360;
wire [151:0] u_ca_out_361;
wire [151:0] u_ca_out_362;
wire [151:0] u_ca_out_363;
wire [151:0] u_ca_out_364;
wire [151:0] u_ca_out_365;
wire [151:0] u_ca_out_366;
wire [151:0] u_ca_out_367;
wire [151:0] u_ca_out_368;
wire [151:0] u_ca_out_369;
wire [151:0] u_ca_out_370;
wire [151:0] u_ca_out_371;
wire [151:0] u_ca_out_372;
wire [151:0] u_ca_out_373;
wire [151:0] u_ca_out_374;
wire [151:0] u_ca_out_375;
wire [151:0] u_ca_out_376;
wire [151:0] u_ca_out_377;
wire [151:0] u_ca_out_378;
wire [151:0] u_ca_out_379;
wire [151:0] u_ca_out_380;
wire [151:0] u_ca_out_381;
wire [151:0] u_ca_out_382;
wire [151:0] u_ca_out_383;
wire [151:0] u_ca_out_384;
wire [151:0] u_ca_out_385;
wire [151:0] u_ca_out_386;
wire [151:0] u_ca_out_387;
wire [151:0] u_ca_out_388;
wire [151:0] u_ca_out_389;
wire [151:0] u_ca_out_390;
wire [151:0] u_ca_out_391;
wire [151:0] u_ca_out_392;
wire [151:0] u_ca_out_393;
wire [151:0] u_ca_out_394;
wire [151:0] u_ca_out_395;
wire [151:0] u_ca_out_396;
wire [151:0] u_ca_out_397;
wire [151:0] u_ca_out_398;
wire [151:0] u_ca_out_399;
wire [151:0] u_ca_out_400;
wire [151:0] u_ca_out_401;
wire [151:0] u_ca_out_402;
wire [151:0] u_ca_out_403;
wire [151:0] u_ca_out_404;
wire [151:0] u_ca_out_405;
wire [151:0] u_ca_out_406;
wire [151:0] u_ca_out_407;
wire [151:0] u_ca_out_408;
wire [151:0] u_ca_out_409;
wire [151:0] u_ca_out_410;
wire [151:0] u_ca_out_411;
wire [151:0] u_ca_out_412;
wire [151:0] u_ca_out_413;
wire [151:0] u_ca_out_414;
wire [151:0] u_ca_out_415;
wire [151:0] u_ca_out_416;
wire [151:0] u_ca_out_417;
wire [151:0] u_ca_out_418;
wire [151:0] u_ca_out_419;
wire [151:0] u_ca_out_420;
wire [151:0] u_ca_out_421;
wire [151:0] u_ca_out_422;
wire [151:0] u_ca_out_423;
wire [151:0] u_ca_out_424;
wire [151:0] u_ca_out_425;
wire [151:0] u_ca_out_426;
wire [151:0] u_ca_out_427;
wire [151:0] u_ca_out_428;
wire [151:0] u_ca_out_429;
wire [151:0] u_ca_out_430;
wire [151:0] u_ca_out_431;
wire [151:0] u_ca_out_432;
wire [151:0] u_ca_out_433;
wire [151:0] u_ca_out_434;
wire [151:0] u_ca_out_435;
wire [151:0] u_ca_out_436;
wire [151:0] u_ca_out_437;
wire [151:0] u_ca_out_438;
wire [151:0] u_ca_out_439;
wire [151:0] u_ca_out_440;
wire [151:0] u_ca_out_441;
wire [151:0] u_ca_out_442;
wire [151:0] u_ca_out_443;
wire [151:0] u_ca_out_444;
wire [151:0] u_ca_out_445;
wire [151:0] u_ca_out_446;
wire [151:0] u_ca_out_447;
wire [151:0] u_ca_out_448;
wire [151:0] u_ca_out_449;
wire [151:0] u_ca_out_450;
wire [151:0] u_ca_out_451;
wire [151:0] u_ca_out_452;
wire [151:0] u_ca_out_453;
wire [151:0] u_ca_out_454;
wire [151:0] u_ca_out_455;
wire [151:0] u_ca_out_456;
wire [151:0] u_ca_out_457;
wire [151:0] u_ca_out_458;
wire [151:0] u_ca_out_459;
wire [151:0] u_ca_out_460;
wire [151:0] u_ca_out_461;
wire [151:0] u_ca_out_462;
wire [151:0] u_ca_out_463;
wire [151:0] u_ca_out_464;
wire [151:0] u_ca_out_465;
wire [151:0] u_ca_out_466;
wire [151:0] u_ca_out_467;
wire [151:0] u_ca_out_468;
wire [151:0] u_ca_out_469;
wire [151:0] u_ca_out_470;
wire [151:0] u_ca_out_471;
wire [151:0] u_ca_out_472;
wire [151:0] u_ca_out_473;
wire [151:0] u_ca_out_474;
wire [151:0] u_ca_out_475;
wire [151:0] u_ca_out_476;
wire [151:0] u_ca_out_477;
wire [151:0] u_ca_out_478;
wire [151:0] u_ca_out_479;
wire [151:0] u_ca_out_480;
wire [151:0] u_ca_out_481;
wire [151:0] u_ca_out_482;
wire [151:0] u_ca_out_483;
wire [151:0] u_ca_out_484;
wire [151:0] u_ca_out_485;
wire [151:0] u_ca_out_486;
wire [151:0] u_ca_out_487;
wire [151:0] u_ca_out_488;
wire [151:0] u_ca_out_489;
wire [151:0] u_ca_out_490;
wire [151:0] u_ca_out_491;
wire [151:0] u_ca_out_492;
wire [151:0] u_ca_out_493;
wire [151:0] u_ca_out_494;
wire [151:0] u_ca_out_495;
wire [151:0] u_ca_out_496;
wire [151:0] u_ca_out_497;
wire [151:0] u_ca_out_498;
wire [151:0] u_ca_out_499;
wire [151:0] u_ca_out_500;
wire [151:0] u_ca_out_501;
wire [151:0] u_ca_out_502;
wire [151:0] u_ca_out_503;
wire [151:0] u_ca_out_504;
wire [151:0] u_ca_out_505;
wire [151:0] u_ca_out_506;
wire [151:0] u_ca_out_507;
wire [151:0] u_ca_out_508;
wire [151:0] u_ca_out_509;
wire [151:0] u_ca_out_510;
wire [151:0] u_ca_out_511;
wire [151:0] u_ca_out_512;
wire [151:0] u_ca_out_513;
wire [151:0] u_ca_out_514;
wire [151:0] u_ca_out_515;
wire [151:0] u_ca_out_516;
wire [151:0] u_ca_out_517;
wire [151:0] u_ca_out_518;
wire [151:0] u_ca_out_519;
wire [151:0] u_ca_out_520;
wire [151:0] u_ca_out_521;
wire [151:0] u_ca_out_522;
wire [151:0] u_ca_out_523;
wire [151:0] u_ca_out_524;
wire [151:0] u_ca_out_525;
wire [151:0] u_ca_out_526;
wire [151:0] u_ca_out_527;
wire [151:0] u_ca_out_528;
wire [151:0] u_ca_out_529;
wire [151:0] u_ca_out_530;
wire [151:0] u_ca_out_531;
wire [151:0] u_ca_out_532;
wire [151:0] u_ca_out_533;
wire [151:0] u_ca_out_534;
wire [151:0] u_ca_out_535;
wire [151:0] u_ca_out_536;
wire [151:0] u_ca_out_537;
wire [151:0] u_ca_out_538;
wire [151:0] u_ca_out_539;
wire [151:0] u_ca_out_540;
wire [151:0] u_ca_out_541;
wire [151:0] u_ca_out_542;
wire [151:0] u_ca_out_543;
wire [151:0] u_ca_out_544;
wire [151:0] u_ca_out_545;
wire [151:0] u_ca_out_546;
wire [151:0] u_ca_out_547;
wire [151:0] u_ca_out_548;
wire [151:0] u_ca_out_549;
wire [151:0] u_ca_out_550;
wire [151:0] u_ca_out_551;
wire [151:0] u_ca_out_552;
wire [151:0] u_ca_out_553;
wire [151:0] u_ca_out_554;
wire [151:0] u_ca_out_555;
wire [151:0] u_ca_out_556;
wire [151:0] u_ca_out_557;
wire [151:0] u_ca_out_558;
wire [151:0] u_ca_out_559;
wire [151:0] u_ca_out_560;
wire [151:0] u_ca_out_561;
wire [151:0] u_ca_out_562;
wire [151:0] u_ca_out_563;
wire [151:0] u_ca_out_564;
wire [151:0] u_ca_out_565;
wire [151:0] u_ca_out_566;
wire [151:0] u_ca_out_567;
wire [151:0] u_ca_out_568;
wire [151:0] u_ca_out_569;
wire [151:0] u_ca_out_570;
wire [151:0] u_ca_out_571;
wire [151:0] u_ca_out_572;
wire [151:0] u_ca_out_573;
wire [151:0] u_ca_out_574;
wire [151:0] u_ca_out_575;
wire [151:0] u_ca_out_576;
wire [151:0] u_ca_out_577;
wire [151:0] u_ca_out_578;
wire [151:0] u_ca_out_579;
wire [151:0] u_ca_out_580;
wire [151:0] u_ca_out_581;
wire [151:0] u_ca_out_582;
wire [151:0] u_ca_out_583;
wire [151:0] u_ca_out_584;
wire [151:0] u_ca_out_585;
wire [151:0] u_ca_out_586;
wire [151:0] u_ca_out_587;
wire [151:0] u_ca_out_588;
wire [151:0] u_ca_out_589;
wire [151:0] u_ca_out_590;
wire [151:0] u_ca_out_591;
wire [151:0] u_ca_out_592;
wire [151:0] u_ca_out_593;
wire [151:0] u_ca_out_594;
wire [151:0] u_ca_out_595;
wire [151:0] u_ca_out_596;
wire [151:0] u_ca_out_597;
wire [151:0] u_ca_out_598;
wire [151:0] u_ca_out_599;
wire [151:0] u_ca_out_600;
wire [151:0] u_ca_out_601;
wire [151:0] u_ca_out_602;
wire [151:0] u_ca_out_603;
wire [151:0] u_ca_out_604;
wire [151:0] u_ca_out_605;
wire [151:0] u_ca_out_606;
wire [151:0] u_ca_out_607;
wire [151:0] u_ca_out_608;
wire [151:0] u_ca_out_609;
wire [151:0] u_ca_out_610;
wire [151:0] u_ca_out_611;
wire [151:0] u_ca_out_612;
wire [151:0] u_ca_out_613;
wire [151:0] u_ca_out_614;
wire [151:0] u_ca_out_615;
wire [151:0] u_ca_out_616;
wire [151:0] u_ca_out_617;
wire [151:0] u_ca_out_618;
wire [151:0] u_ca_out_619;
wire [151:0] u_ca_out_620;
wire [151:0] u_ca_out_621;
wire [151:0] u_ca_out_622;
wire [151:0] u_ca_out_623;
wire [151:0] u_ca_out_624;
wire [151:0] u_ca_out_625;
wire [151:0] u_ca_out_626;
wire [151:0] u_ca_out_627;
wire [151:0] u_ca_out_628;
wire [151:0] u_ca_out_629;
wire [151:0] u_ca_out_630;
wire [151:0] u_ca_out_631;
wire [151:0] u_ca_out_632;
wire [151:0] u_ca_out_633;
wire [151:0] u_ca_out_634;
wire [151:0] u_ca_out_635;
wire [151:0] u_ca_out_636;
wire [151:0] u_ca_out_637;
wire [151:0] u_ca_out_638;
wire [151:0] u_ca_out_639;
wire [151:0] u_ca_out_640;
wire [151:0] u_ca_out_641;
wire [151:0] u_ca_out_642;
wire [151:0] u_ca_out_643;
wire [151:0] u_ca_out_644;
wire [151:0] u_ca_out_645;
wire [151:0] u_ca_out_646;
wire [151:0] u_ca_out_647;
wire [151:0] u_ca_out_648;
wire [151:0] u_ca_out_649;
wire [151:0] u_ca_out_650;
wire [151:0] u_ca_out_651;
wire [151:0] u_ca_out_652;
wire [151:0] u_ca_out_653;
wire [151:0] u_ca_out_654;
wire [151:0] u_ca_out_655;
wire [151:0] u_ca_out_656;
wire [151:0] u_ca_out_657;
wire [151:0] u_ca_out_658;
wire [151:0] u_ca_out_659;
wire [151:0] u_ca_out_660;
wire [151:0] u_ca_out_661;
wire [151:0] u_ca_out_662;
wire [151:0] u_ca_out_663;
wire [151:0] u_ca_out_664;
wire [151:0] u_ca_out_665;
wire [151:0] u_ca_out_666;
wire [151:0] u_ca_out_667;
wire [151:0] u_ca_out_668;
wire [151:0] u_ca_out_669;
wire [151:0] u_ca_out_670;
wire [151:0] u_ca_out_671;
wire [151:0] u_ca_out_672;
wire [151:0] u_ca_out_673;
wire [151:0] u_ca_out_674;
wire [151:0] u_ca_out_675;
wire [151:0] u_ca_out_676;
wire [151:0] u_ca_out_677;
wire [151:0] u_ca_out_678;
wire [151:0] u_ca_out_679;
wire [151:0] u_ca_out_680;
wire [151:0] u_ca_out_681;
wire [151:0] u_ca_out_682;
wire [151:0] u_ca_out_683;
wire [151:0] u_ca_out_684;
wire [151:0] u_ca_out_685;
wire [151:0] u_ca_out_686;
wire [151:0] u_ca_out_687;
wire [151:0] u_ca_out_688;
wire [151:0] u_ca_out_689;
wire [151:0] u_ca_out_690;
wire [151:0] u_ca_out_691;
wire [151:0] u_ca_out_692;
wire [151:0] u_ca_out_693;
wire [151:0] u_ca_out_694;
wire [151:0] u_ca_out_695;
wire [151:0] u_ca_out_696;
wire [151:0] u_ca_out_697;
wire [151:0] u_ca_out_698;
wire [151:0] u_ca_out_699;
wire [151:0] u_ca_out_700;
wire [151:0] u_ca_out_701;
wire [151:0] u_ca_out_702;
wire [151:0] u_ca_out_703;
wire [151:0] u_ca_out_704;
wire [151:0] u_ca_out_705;
wire [151:0] u_ca_out_706;
wire [151:0] u_ca_out_707;
wire [151:0] u_ca_out_708;
wire [151:0] u_ca_out_709;
wire [151:0] u_ca_out_710;
wire [151:0] u_ca_out_711;
wire [151:0] u_ca_out_712;
wire [151:0] u_ca_out_713;
wire [151:0] u_ca_out_714;
wire [151:0] u_ca_out_715;
wire [151:0] u_ca_out_716;
wire [151:0] u_ca_out_717;
wire [151:0] u_ca_out_718;
wire [151:0] u_ca_out_719;
wire [151:0] u_ca_out_720;
wire [151:0] u_ca_out_721;
wire [151:0] u_ca_out_722;
wire [151:0] u_ca_out_723;
wire [151:0] u_ca_out_724;
wire [151:0] u_ca_out_725;
wire [151:0] u_ca_out_726;
wire [151:0] u_ca_out_727;
wire [151:0] u_ca_out_728;
wire [151:0] u_ca_out_729;
wire [151:0] u_ca_out_730;
wire [151:0] u_ca_out_731;
wire [151:0] u_ca_out_732;
wire [151:0] u_ca_out_733;
wire [151:0] u_ca_out_734;
wire [151:0] u_ca_out_735;
wire [151:0] u_ca_out_736;
wire [151:0] u_ca_out_737;
wire [151:0] u_ca_out_738;
wire [151:0] u_ca_out_739;
wire [151:0] u_ca_out_740;
wire [151:0] u_ca_out_741;
wire [151:0] u_ca_out_742;
wire [151:0] u_ca_out_743;
wire [151:0] u_ca_out_744;
wire [151:0] u_ca_out_745;
wire [151:0] u_ca_out_746;
wire [151:0] u_ca_out_747;
wire [151:0] u_ca_out_748;
wire [151:0] u_ca_out_749;
wire [151:0] u_ca_out_750;
wire [151:0] u_ca_out_751;
wire [151:0] u_ca_out_752;
wire [151:0] u_ca_out_753;
wire [151:0] u_ca_out_754;
wire [151:0] u_ca_out_755;
wire [151:0] u_ca_out_756;
wire [151:0] u_ca_out_757;
wire [151:0] u_ca_out_758;
wire [151:0] u_ca_out_759;
wire [151:0] u_ca_out_760;
wire [151:0] u_ca_out_761;
wire [151:0] u_ca_out_762;
wire [151:0] u_ca_out_763;
wire [151:0] u_ca_out_764;
wire [151:0] u_ca_out_765;
wire [151:0] u_ca_out_766;
wire [151:0] u_ca_out_767;
wire [151:0] u_ca_out_768;
wire [151:0] u_ca_out_769;
wire [151:0] u_ca_out_770;
wire [151:0] u_ca_out_771;
wire [151:0] u_ca_out_772;
wire [151:0] u_ca_out_773;
wire [151:0] u_ca_out_774;
wire [151:0] u_ca_out_775;
wire [151:0] u_ca_out_776;
wire [151:0] u_ca_out_777;
wire [151:0] u_ca_out_778;
wire [151:0] u_ca_out_779;
wire [151:0] u_ca_out_780;
wire [151:0] u_ca_out_781;
wire [151:0] u_ca_out_782;
wire [151:0] u_ca_out_783;
wire [151:0] u_ca_out_784;
wire [151:0] u_ca_out_785;
wire [151:0] u_ca_out_786;
wire [151:0] u_ca_out_787;
wire [151:0] u_ca_out_788;
wire [151:0] u_ca_out_789;
wire [151:0] u_ca_out_790;
wire [151:0] u_ca_out_791;
wire [151:0] u_ca_out_792;
wire [151:0] u_ca_out_793;
wire [151:0] u_ca_out_794;
wire [151:0] u_ca_out_795;
wire [151:0] u_ca_out_796;
wire [151:0] u_ca_out_797;
wire [151:0] u_ca_out_798;
wire [151:0] u_ca_out_799;
wire [151:0] u_ca_out_800;
wire [151:0] u_ca_out_801;
wire [151:0] u_ca_out_802;
wire [151:0] u_ca_out_803;
wire [151:0] u_ca_out_804;
wire [151:0] u_ca_out_805;
wire [151:0] u_ca_out_806;
wire [151:0] u_ca_out_807;
wire [151:0] u_ca_out_808;
wire [151:0] u_ca_out_809;
wire [151:0] u_ca_out_810;
wire [151:0] u_ca_out_811;
wire [151:0] u_ca_out_812;
wire [151:0] u_ca_out_813;
wire [151:0] u_ca_out_814;
wire [151:0] u_ca_out_815;
wire [151:0] u_ca_out_816;
wire [151:0] u_ca_out_817;
wire [151:0] u_ca_out_818;
wire [151:0] u_ca_out_819;
wire [151:0] u_ca_out_820;
wire [151:0] u_ca_out_821;
wire [151:0] u_ca_out_822;
wire [151:0] u_ca_out_823;
wire [151:0] u_ca_out_824;
wire [151:0] u_ca_out_825;
wire [151:0] u_ca_out_826;
wire [151:0] u_ca_out_827;
wire [151:0] u_ca_out_828;
wire [151:0] u_ca_out_829;
wire [151:0] u_ca_out_830;
wire [151:0] u_ca_out_831;
wire [151:0] u_ca_out_832;
wire [151:0] u_ca_out_833;
wire [151:0] u_ca_out_834;
wire [151:0] u_ca_out_835;
wire [151:0] u_ca_out_836;
wire [151:0] u_ca_out_837;
wire [151:0] u_ca_out_838;
wire [151:0] u_ca_out_839;
wire [151:0] u_ca_out_840;
wire [151:0] u_ca_out_841;
wire [151:0] u_ca_out_842;
wire [151:0] u_ca_out_843;
wire [151:0] u_ca_out_844;
wire [151:0] u_ca_out_845;
wire [151:0] u_ca_out_846;
wire [151:0] u_ca_out_847;
wire [151:0] u_ca_out_848;
wire [151:0] u_ca_out_849;
wire [151:0] u_ca_out_850;
wire [151:0] u_ca_out_851;
wire [151:0] u_ca_out_852;
wire [151:0] u_ca_out_853;
wire [151:0] u_ca_out_854;
wire [151:0] u_ca_out_855;
wire [151:0] u_ca_out_856;
wire [151:0] u_ca_out_857;
wire [151:0] u_ca_out_858;
wire [151:0] u_ca_out_859;
wire [151:0] u_ca_out_860;
wire [151:0] u_ca_out_861;
wire [151:0] u_ca_out_862;
wire [151:0] u_ca_out_863;
wire [151:0] u_ca_out_864;
wire [151:0] u_ca_out_865;
wire [151:0] u_ca_out_866;
wire [151:0] u_ca_out_867;
wire [151:0] u_ca_out_868;
wire [151:0] u_ca_out_869;
wire [151:0] u_ca_out_870;
wire [151:0] u_ca_out_871;
wire [151:0] u_ca_out_872;
wire [151:0] u_ca_out_873;
wire [151:0] u_ca_out_874;
wire [151:0] u_ca_out_875;
wire [151:0] u_ca_out_876;
wire [151:0] u_ca_out_877;
wire [151:0] u_ca_out_878;
wire [151:0] u_ca_out_879;
wire [151:0] u_ca_out_880;
wire [151:0] u_ca_out_881;
wire [151:0] u_ca_out_882;
wire [151:0] u_ca_out_883;
wire [151:0] u_ca_out_884;
wire [151:0] u_ca_out_885;
wire [151:0] u_ca_out_886;
wire [151:0] u_ca_out_887;
wire [151:0] u_ca_out_888;
wire [151:0] u_ca_out_889;
wire [151:0] u_ca_out_890;
wire [151:0] u_ca_out_891;
wire [151:0] u_ca_out_892;
wire [151:0] u_ca_out_893;
wire [151:0] u_ca_out_894;
wire [151:0] u_ca_out_895;
wire [151:0] u_ca_out_896;
wire [151:0] u_ca_out_897;
wire [151:0] u_ca_out_898;
wire [151:0] u_ca_out_899;
wire [151:0] u_ca_out_900;
wire [151:0] u_ca_out_901;
wire [151:0] u_ca_out_902;
wire [151:0] u_ca_out_903;
wire [151:0] u_ca_out_904;
wire [151:0] u_ca_out_905;
wire [151:0] u_ca_out_906;
wire [151:0] u_ca_out_907;
wire [151:0] u_ca_out_908;
wire [151:0] u_ca_out_909;
wire [151:0] u_ca_out_910;
wire [151:0] u_ca_out_911;
wire [151:0] u_ca_out_912;
wire [151:0] u_ca_out_913;
wire [151:0] u_ca_out_914;
wire [151:0] u_ca_out_915;
wire [151:0] u_ca_out_916;
wire [151:0] u_ca_out_917;
wire [151:0] u_ca_out_918;
wire [151:0] u_ca_out_919;
wire [151:0] u_ca_out_920;
wire [151:0] u_ca_out_921;
wire [151:0] u_ca_out_922;
wire [151:0] u_ca_out_923;
wire [151:0] u_ca_out_924;
wire [151:0] u_ca_out_925;
wire [151:0] u_ca_out_926;
wire [151:0] u_ca_out_927;
wire [151:0] u_ca_out_928;
wire [151:0] u_ca_out_929;
wire [151:0] u_ca_out_930;
wire [151:0] u_ca_out_931;
wire [151:0] u_ca_out_932;
wire [151:0] u_ca_out_933;
wire [151:0] u_ca_out_934;
wire [151:0] u_ca_out_935;
wire [151:0] u_ca_out_936;
wire [151:0] u_ca_out_937;
wire [151:0] u_ca_out_938;
wire [151:0] u_ca_out_939;
wire [151:0] u_ca_out_940;
wire [151:0] u_ca_out_941;
wire [151:0] u_ca_out_942;
wire [151:0] u_ca_out_943;
wire [151:0] u_ca_out_944;
wire [151:0] u_ca_out_945;
wire [151:0] u_ca_out_946;
wire [151:0] u_ca_out_947;
wire [151:0] u_ca_out_948;
wire [151:0] u_ca_out_949;
wire [151:0] u_ca_out_950;
wire [151:0] u_ca_out_951;
wire [151:0] u_ca_out_952;
wire [151:0] u_ca_out_953;
wire [151:0] u_ca_out_954;
wire [151:0] u_ca_out_955;
wire [151:0] u_ca_out_956;
wire [151:0] u_ca_out_957;
wire [151:0] u_ca_out_958;
wire [151:0] u_ca_out_959;
wire [151:0] u_ca_out_960;
wire [151:0] u_ca_out_961;
wire [151:0] u_ca_out_962;
wire [151:0] u_ca_out_963;
wire [151:0] u_ca_out_964;
wire [151:0] u_ca_out_965;
wire [151:0] u_ca_out_966;
wire [151:0] u_ca_out_967;
wire [151:0] u_ca_out_968;
wire [151:0] u_ca_out_969;
wire [151:0] u_ca_out_970;
wire [151:0] u_ca_out_971;
wire [151:0] u_ca_out_972;
wire [151:0] u_ca_out_973;
wire [151:0] u_ca_out_974;
wire [151:0] u_ca_out_975;
wire [151:0] u_ca_out_976;
wire [151:0] u_ca_out_977;
wire [151:0] u_ca_out_978;
wire [151:0] u_ca_out_979;
wire [151:0] u_ca_out_980;
wire [151:0] u_ca_out_981;
wire [151:0] u_ca_out_982;
wire [151:0] u_ca_out_983;
wire [151:0] u_ca_out_984;
wire [151:0] u_ca_out_985;
wire [151:0] u_ca_out_986;
wire [151:0] u_ca_out_987;
wire [151:0] u_ca_out_988;
wire [151:0] u_ca_out_989;
wire [151:0] u_ca_out_990;
wire [151:0] u_ca_out_991;
wire [151:0] u_ca_out_992;
wire [151:0] u_ca_out_993;
wire [151:0] u_ca_out_994;
wire [151:0] u_ca_out_995;
wire [151:0] u_ca_out_996;
wire [151:0] u_ca_out_997;
wire [151:0] u_ca_out_998;
wire [151:0] u_ca_out_999;
wire [151:0] u_ca_out_1000;
wire [151:0] u_ca_out_1001;
wire [151:0] u_ca_out_1002;
wire [151:0] u_ca_out_1003;
wire [151:0] u_ca_out_1004;
wire [151:0] u_ca_out_1005;
wire [151:0] u_ca_out_1006;
wire [151:0] u_ca_out_1007;
wire [151:0] u_ca_out_1008;
wire [151:0] u_ca_out_1009;
wire [151:0] u_ca_out_1010;
wire [151:0] u_ca_out_1011;
wire [151:0] u_ca_out_1012;
wire [151:0] u_ca_out_1013;
wire [151:0] u_ca_out_1014;
wire [151:0] u_ca_out_1015;
wire [151:0] u_ca_out_1016;
wire [151:0] u_ca_out_1017;
wire [151:0] u_ca_out_1018;
wire [151:0] u_ca_out_1019;
wire [151:0] u_ca_out_1020;
wire [151:0] u_ca_out_1021;
wire [151:0] u_ca_out_1022;
wire [151:0] u_ca_out_1023;

assign u_ca_in_0 = {{1{1'b0}}, col_in_0};
assign u_ca_in_1 = {{1{1'b0}}, col_in_1};
assign u_ca_in_2 = {{1{1'b0}}, col_in_2};
assign u_ca_in_3 = {{1{1'b0}}, col_in_3};
assign u_ca_in_4 = {{1{1'b0}}, col_in_4};
assign u_ca_in_5 = {{1{1'b0}}, col_in_5};
assign u_ca_in_6 = {{1{1'b0}}, col_in_6};
assign u_ca_in_7 = {{1{1'b0}}, col_in_7};
assign u_ca_in_8 = {{1{1'b0}}, col_in_8};
assign u_ca_in_9 = {{1{1'b0}}, col_in_9};
assign u_ca_in_10 = {{1{1'b0}}, col_in_10};
assign u_ca_in_11 = {{1{1'b0}}, col_in_11};
assign u_ca_in_12 = {{1{1'b0}}, col_in_12};
assign u_ca_in_13 = {{1{1'b0}}, col_in_13};
assign u_ca_in_14 = {{1{1'b0}}, col_in_14};
assign u_ca_in_15 = {{1{1'b0}}, col_in_15};
assign u_ca_in_16 = {{1{1'b0}}, col_in_16};
assign u_ca_in_17 = {{1{1'b0}}, col_in_17};
assign u_ca_in_18 = {{1{1'b0}}, col_in_18};
assign u_ca_in_19 = {{1{1'b0}}, col_in_19};
assign u_ca_in_20 = {{1{1'b0}}, col_in_20};
assign u_ca_in_21 = {{1{1'b0}}, col_in_21};
assign u_ca_in_22 = {{1{1'b0}}, col_in_22};
assign u_ca_in_23 = {{1{1'b0}}, col_in_23};
assign u_ca_in_24 = {{1{1'b0}}, col_in_24};
assign u_ca_in_25 = {{1{1'b0}}, col_in_25};
assign u_ca_in_26 = {{1{1'b0}}, col_in_26};
assign u_ca_in_27 = {{1{1'b0}}, col_in_27};
assign u_ca_in_28 = {{1{1'b0}}, col_in_28};
assign u_ca_in_29 = {{1{1'b0}}, col_in_29};
assign u_ca_in_30 = {{1{1'b0}}, col_in_30};
assign u_ca_in_31 = {{1{1'b0}}, col_in_31};
assign u_ca_in_32 = {{1{1'b0}}, col_in_32};
assign u_ca_in_33 = {{1{1'b0}}, col_in_33};
assign u_ca_in_34 = {{1{1'b0}}, col_in_34};
assign u_ca_in_35 = {{1{1'b0}}, col_in_35};
assign u_ca_in_36 = {{1{1'b0}}, col_in_36};
assign u_ca_in_37 = {{1{1'b0}}, col_in_37};
assign u_ca_in_38 = {{1{1'b0}}, col_in_38};
assign u_ca_in_39 = {{1{1'b0}}, col_in_39};
assign u_ca_in_40 = {{1{1'b0}}, col_in_40};
assign u_ca_in_41 = {{1{1'b0}}, col_in_41};
assign u_ca_in_42 = {{1{1'b0}}, col_in_42};
assign u_ca_in_43 = {{1{1'b0}}, col_in_43};
assign u_ca_in_44 = {{1{1'b0}}, col_in_44};
assign u_ca_in_45 = {{1{1'b0}}, col_in_45};
assign u_ca_in_46 = {{1{1'b0}}, col_in_46};
assign u_ca_in_47 = {{1{1'b0}}, col_in_47};
assign u_ca_in_48 = {{1{1'b0}}, col_in_48};
assign u_ca_in_49 = {{1{1'b0}}, col_in_49};
assign u_ca_in_50 = {{1{1'b0}}, col_in_50};
assign u_ca_in_51 = {{1{1'b0}}, col_in_51};
assign u_ca_in_52 = {{1{1'b0}}, col_in_52};
assign u_ca_in_53 = {{1{1'b0}}, col_in_53};
assign u_ca_in_54 = {{1{1'b0}}, col_in_54};
assign u_ca_in_55 = {{1{1'b0}}, col_in_55};
assign u_ca_in_56 = {{1{1'b0}}, col_in_56};
assign u_ca_in_57 = {{1{1'b0}}, col_in_57};
assign u_ca_in_58 = {{1{1'b0}}, col_in_58};
assign u_ca_in_59 = {{1{1'b0}}, col_in_59};
assign u_ca_in_60 = {{1{1'b0}}, col_in_60};
assign u_ca_in_61 = {{1{1'b0}}, col_in_61};
assign u_ca_in_62 = {{1{1'b0}}, col_in_62};
assign u_ca_in_63 = {{1{1'b0}}, col_in_63};
assign u_ca_in_64 = {{1{1'b0}}, col_in_64};
assign u_ca_in_65 = {{1{1'b0}}, col_in_65};
assign u_ca_in_66 = {{1{1'b0}}, col_in_66};
assign u_ca_in_67 = {{1{1'b0}}, col_in_67};
assign u_ca_in_68 = {{1{1'b0}}, col_in_68};
assign u_ca_in_69 = {{1{1'b0}}, col_in_69};
assign u_ca_in_70 = {{1{1'b0}}, col_in_70};
assign u_ca_in_71 = {{1{1'b0}}, col_in_71};
assign u_ca_in_72 = {{1{1'b0}}, col_in_72};
assign u_ca_in_73 = {{1{1'b0}}, col_in_73};
assign u_ca_in_74 = {{1{1'b0}}, col_in_74};
assign u_ca_in_75 = {{1{1'b0}}, col_in_75};
assign u_ca_in_76 = {{1{1'b0}}, col_in_76};
assign u_ca_in_77 = {{1{1'b0}}, col_in_77};
assign u_ca_in_78 = {{1{1'b0}}, col_in_78};
assign u_ca_in_79 = {{1{1'b0}}, col_in_79};
assign u_ca_in_80 = {{1{1'b0}}, col_in_80};
assign u_ca_in_81 = {{1{1'b0}}, col_in_81};
assign u_ca_in_82 = {{1{1'b0}}, col_in_82};
assign u_ca_in_83 = {{1{1'b0}}, col_in_83};
assign u_ca_in_84 = {{1{1'b0}}, col_in_84};
assign u_ca_in_85 = {{1{1'b0}}, col_in_85};
assign u_ca_in_86 = {{1{1'b0}}, col_in_86};
assign u_ca_in_87 = {{1{1'b0}}, col_in_87};
assign u_ca_in_88 = {{1{1'b0}}, col_in_88};
assign u_ca_in_89 = {{1{1'b0}}, col_in_89};
assign u_ca_in_90 = {{1{1'b0}}, col_in_90};
assign u_ca_in_91 = {{1{1'b0}}, col_in_91};
assign u_ca_in_92 = {{1{1'b0}}, col_in_92};
assign u_ca_in_93 = {{1{1'b0}}, col_in_93};
assign u_ca_in_94 = {{1{1'b0}}, col_in_94};
assign u_ca_in_95 = {{1{1'b0}}, col_in_95};
assign u_ca_in_96 = {{1{1'b0}}, col_in_96};
assign u_ca_in_97 = {{1{1'b0}}, col_in_97};
assign u_ca_in_98 = {{1{1'b0}}, col_in_98};
assign u_ca_in_99 = {{1{1'b0}}, col_in_99};
assign u_ca_in_100 = {{1{1'b0}}, col_in_100};
assign u_ca_in_101 = {{1{1'b0}}, col_in_101};
assign u_ca_in_102 = {{1{1'b0}}, col_in_102};
assign u_ca_in_103 = {{1{1'b0}}, col_in_103};
assign u_ca_in_104 = {{1{1'b0}}, col_in_104};
assign u_ca_in_105 = {{1{1'b0}}, col_in_105};
assign u_ca_in_106 = {{1{1'b0}}, col_in_106};
assign u_ca_in_107 = {{1{1'b0}}, col_in_107};
assign u_ca_in_108 = {{1{1'b0}}, col_in_108};
assign u_ca_in_109 = {{1{1'b0}}, col_in_109};
assign u_ca_in_110 = {{1{1'b0}}, col_in_110};
assign u_ca_in_111 = {{1{1'b0}}, col_in_111};
assign u_ca_in_112 = {{1{1'b0}}, col_in_112};
assign u_ca_in_113 = {{1{1'b0}}, col_in_113};
assign u_ca_in_114 = {{1{1'b0}}, col_in_114};
assign u_ca_in_115 = {{1{1'b0}}, col_in_115};
assign u_ca_in_116 = {{1{1'b0}}, col_in_116};
assign u_ca_in_117 = {{1{1'b0}}, col_in_117};
assign u_ca_in_118 = {{1{1'b0}}, col_in_118};
assign u_ca_in_119 = {{1{1'b0}}, col_in_119};
assign u_ca_in_120 = {{1{1'b0}}, col_in_120};
assign u_ca_in_121 = {{1{1'b0}}, col_in_121};
assign u_ca_in_122 = {{1{1'b0}}, col_in_122};
assign u_ca_in_123 = {{1{1'b0}}, col_in_123};
assign u_ca_in_124 = {{1{1'b0}}, col_in_124};
assign u_ca_in_125 = {{1{1'b0}}, col_in_125};
assign u_ca_in_126 = {{1{1'b0}}, col_in_126};
assign u_ca_in_127 = {{1{1'b0}}, col_in_127};
assign u_ca_in_128 = {{1{1'b0}}, col_in_128};
assign u_ca_in_129 = {{1{1'b0}}, col_in_129};
assign u_ca_in_130 = {{1{1'b0}}, col_in_130};
assign u_ca_in_131 = {{1{1'b0}}, col_in_131};
assign u_ca_in_132 = {{1{1'b0}}, col_in_132};
assign u_ca_in_133 = {{1{1'b0}}, col_in_133};
assign u_ca_in_134 = {{1{1'b0}}, col_in_134};
assign u_ca_in_135 = {{1{1'b0}}, col_in_135};
assign u_ca_in_136 = {{1{1'b0}}, col_in_136};
assign u_ca_in_137 = {{1{1'b0}}, col_in_137};
assign u_ca_in_138 = {{1{1'b0}}, col_in_138};
assign u_ca_in_139 = {{1{1'b0}}, col_in_139};
assign u_ca_in_140 = {{1{1'b0}}, col_in_140};
assign u_ca_in_141 = {{1{1'b0}}, col_in_141};
assign u_ca_in_142 = {{1{1'b0}}, col_in_142};
assign u_ca_in_143 = {{1{1'b0}}, col_in_143};
assign u_ca_in_144 = {{1{1'b0}}, col_in_144};
assign u_ca_in_145 = {{1{1'b0}}, col_in_145};
assign u_ca_in_146 = {{1{1'b0}}, col_in_146};
assign u_ca_in_147 = {{1{1'b0}}, col_in_147};
assign u_ca_in_148 = {{1{1'b0}}, col_in_148};
assign u_ca_in_149 = {{1{1'b0}}, col_in_149};
assign u_ca_in_150 = {{1{1'b0}}, col_in_150};
assign u_ca_in_151 = {{1{1'b0}}, col_in_151};
assign u_ca_in_152 = {{1{1'b0}}, col_in_152};
assign u_ca_in_153 = {{1{1'b0}}, col_in_153};
assign u_ca_in_154 = {{1{1'b0}}, col_in_154};
assign u_ca_in_155 = {{1{1'b0}}, col_in_155};
assign u_ca_in_156 = {{1{1'b0}}, col_in_156};
assign u_ca_in_157 = {{1{1'b0}}, col_in_157};
assign u_ca_in_158 = {{1{1'b0}}, col_in_158};
assign u_ca_in_159 = {{1{1'b0}}, col_in_159};
assign u_ca_in_160 = {{1{1'b0}}, col_in_160};
assign u_ca_in_161 = {{1{1'b0}}, col_in_161};
assign u_ca_in_162 = {{1{1'b0}}, col_in_162};
assign u_ca_in_163 = {{1{1'b0}}, col_in_163};
assign u_ca_in_164 = {{1{1'b0}}, col_in_164};
assign u_ca_in_165 = {{1{1'b0}}, col_in_165};
assign u_ca_in_166 = {{1{1'b0}}, col_in_166};
assign u_ca_in_167 = {{1{1'b0}}, col_in_167};
assign u_ca_in_168 = {{1{1'b0}}, col_in_168};
assign u_ca_in_169 = {{1{1'b0}}, col_in_169};
assign u_ca_in_170 = {{1{1'b0}}, col_in_170};
assign u_ca_in_171 = {{1{1'b0}}, col_in_171};
assign u_ca_in_172 = {{1{1'b0}}, col_in_172};
assign u_ca_in_173 = {{1{1'b0}}, col_in_173};
assign u_ca_in_174 = {{1{1'b0}}, col_in_174};
assign u_ca_in_175 = {{1{1'b0}}, col_in_175};
assign u_ca_in_176 = {{1{1'b0}}, col_in_176};
assign u_ca_in_177 = {{1{1'b0}}, col_in_177};
assign u_ca_in_178 = {{1{1'b0}}, col_in_178};
assign u_ca_in_179 = {{1{1'b0}}, col_in_179};
assign u_ca_in_180 = {{1{1'b0}}, col_in_180};
assign u_ca_in_181 = {{1{1'b0}}, col_in_181};
assign u_ca_in_182 = {{1{1'b0}}, col_in_182};
assign u_ca_in_183 = {{1{1'b0}}, col_in_183};
assign u_ca_in_184 = {{1{1'b0}}, col_in_184};
assign u_ca_in_185 = {{1{1'b0}}, col_in_185};
assign u_ca_in_186 = {{1{1'b0}}, col_in_186};
assign u_ca_in_187 = {{1{1'b0}}, col_in_187};
assign u_ca_in_188 = {{1{1'b0}}, col_in_188};
assign u_ca_in_189 = {{1{1'b0}}, col_in_189};
assign u_ca_in_190 = {{1{1'b0}}, col_in_190};
assign u_ca_in_191 = {{1{1'b0}}, col_in_191};
assign u_ca_in_192 = {{1{1'b0}}, col_in_192};
assign u_ca_in_193 = {{1{1'b0}}, col_in_193};
assign u_ca_in_194 = {{1{1'b0}}, col_in_194};
assign u_ca_in_195 = {{1{1'b0}}, col_in_195};
assign u_ca_in_196 = {{1{1'b0}}, col_in_196};
assign u_ca_in_197 = {{1{1'b0}}, col_in_197};
assign u_ca_in_198 = {{1{1'b0}}, col_in_198};
assign u_ca_in_199 = {{1{1'b0}}, col_in_199};
assign u_ca_in_200 = {{1{1'b0}}, col_in_200};
assign u_ca_in_201 = {{1{1'b0}}, col_in_201};
assign u_ca_in_202 = {{1{1'b0}}, col_in_202};
assign u_ca_in_203 = {{1{1'b0}}, col_in_203};
assign u_ca_in_204 = {{1{1'b0}}, col_in_204};
assign u_ca_in_205 = {{1{1'b0}}, col_in_205};
assign u_ca_in_206 = {{1{1'b0}}, col_in_206};
assign u_ca_in_207 = {{1{1'b0}}, col_in_207};
assign u_ca_in_208 = {{1{1'b0}}, col_in_208};
assign u_ca_in_209 = {{1{1'b0}}, col_in_209};
assign u_ca_in_210 = {{1{1'b0}}, col_in_210};
assign u_ca_in_211 = {{1{1'b0}}, col_in_211};
assign u_ca_in_212 = {{1{1'b0}}, col_in_212};
assign u_ca_in_213 = {{1{1'b0}}, col_in_213};
assign u_ca_in_214 = {{1{1'b0}}, col_in_214};
assign u_ca_in_215 = {{1{1'b0}}, col_in_215};
assign u_ca_in_216 = {{1{1'b0}}, col_in_216};
assign u_ca_in_217 = {{1{1'b0}}, col_in_217};
assign u_ca_in_218 = {{1{1'b0}}, col_in_218};
assign u_ca_in_219 = {{1{1'b0}}, col_in_219};
assign u_ca_in_220 = {{1{1'b0}}, col_in_220};
assign u_ca_in_221 = {{1{1'b0}}, col_in_221};
assign u_ca_in_222 = {{1{1'b0}}, col_in_222};
assign u_ca_in_223 = {{1{1'b0}}, col_in_223};
assign u_ca_in_224 = {{1{1'b0}}, col_in_224};
assign u_ca_in_225 = {{1{1'b0}}, col_in_225};
assign u_ca_in_226 = {{1{1'b0}}, col_in_226};
assign u_ca_in_227 = {{1{1'b0}}, col_in_227};
assign u_ca_in_228 = {{1{1'b0}}, col_in_228};
assign u_ca_in_229 = {{1{1'b0}}, col_in_229};
assign u_ca_in_230 = {{1{1'b0}}, col_in_230};
assign u_ca_in_231 = {{1{1'b0}}, col_in_231};
assign u_ca_in_232 = {{1{1'b0}}, col_in_232};
assign u_ca_in_233 = {{1{1'b0}}, col_in_233};
assign u_ca_in_234 = {{1{1'b0}}, col_in_234};
assign u_ca_in_235 = {{1{1'b0}}, col_in_235};
assign u_ca_in_236 = {{1{1'b0}}, col_in_236};
assign u_ca_in_237 = {{1{1'b0}}, col_in_237};
assign u_ca_in_238 = {{1{1'b0}}, col_in_238};
assign u_ca_in_239 = {{1{1'b0}}, col_in_239};
assign u_ca_in_240 = {{1{1'b0}}, col_in_240};
assign u_ca_in_241 = {{1{1'b0}}, col_in_241};
assign u_ca_in_242 = {{1{1'b0}}, col_in_242};
assign u_ca_in_243 = {{1{1'b0}}, col_in_243};
assign u_ca_in_244 = {{1{1'b0}}, col_in_244};
assign u_ca_in_245 = {{1{1'b0}}, col_in_245};
assign u_ca_in_246 = {{1{1'b0}}, col_in_246};
assign u_ca_in_247 = {{1{1'b0}}, col_in_247};
assign u_ca_in_248 = {{1{1'b0}}, col_in_248};
assign u_ca_in_249 = {{1{1'b0}}, col_in_249};
assign u_ca_in_250 = {{1{1'b0}}, col_in_250};
assign u_ca_in_251 = {{1{1'b0}}, col_in_251};
assign u_ca_in_252 = {{1{1'b0}}, col_in_252};
assign u_ca_in_253 = {{1{1'b0}}, col_in_253};
assign u_ca_in_254 = {{1{1'b0}}, col_in_254};
assign u_ca_in_255 = {{1{1'b0}}, col_in_255};
assign u_ca_in_256 = {{1{1'b0}}, col_in_256};
assign u_ca_in_257 = {{1{1'b0}}, col_in_257};
assign u_ca_in_258 = {{1{1'b0}}, col_in_258};
assign u_ca_in_259 = {{1{1'b0}}, col_in_259};
assign u_ca_in_260 = {{1{1'b0}}, col_in_260};
assign u_ca_in_261 = {{1{1'b0}}, col_in_261};
assign u_ca_in_262 = {{1{1'b0}}, col_in_262};
assign u_ca_in_263 = {{1{1'b0}}, col_in_263};
assign u_ca_in_264 = {{1{1'b0}}, col_in_264};
assign u_ca_in_265 = {{1{1'b0}}, col_in_265};
assign u_ca_in_266 = {{1{1'b0}}, col_in_266};
assign u_ca_in_267 = {{1{1'b0}}, col_in_267};
assign u_ca_in_268 = {{1{1'b0}}, col_in_268};
assign u_ca_in_269 = {{1{1'b0}}, col_in_269};
assign u_ca_in_270 = {{1{1'b0}}, col_in_270};
assign u_ca_in_271 = {{1{1'b0}}, col_in_271};
assign u_ca_in_272 = {{1{1'b0}}, col_in_272};
assign u_ca_in_273 = {{1{1'b0}}, col_in_273};
assign u_ca_in_274 = {{1{1'b0}}, col_in_274};
assign u_ca_in_275 = {{1{1'b0}}, col_in_275};
assign u_ca_in_276 = {{1{1'b0}}, col_in_276};
assign u_ca_in_277 = {{1{1'b0}}, col_in_277};
assign u_ca_in_278 = {{1{1'b0}}, col_in_278};
assign u_ca_in_279 = {{1{1'b0}}, col_in_279};
assign u_ca_in_280 = {{1{1'b0}}, col_in_280};
assign u_ca_in_281 = {{1{1'b0}}, col_in_281};
assign u_ca_in_282 = {{1{1'b0}}, col_in_282};
assign u_ca_in_283 = {{1{1'b0}}, col_in_283};
assign u_ca_in_284 = {{1{1'b0}}, col_in_284};
assign u_ca_in_285 = {{1{1'b0}}, col_in_285};
assign u_ca_in_286 = {{1{1'b0}}, col_in_286};
assign u_ca_in_287 = {{1{1'b0}}, col_in_287};
assign u_ca_in_288 = {{1{1'b0}}, col_in_288};
assign u_ca_in_289 = {{1{1'b0}}, col_in_289};
assign u_ca_in_290 = {{1{1'b0}}, col_in_290};
assign u_ca_in_291 = {{1{1'b0}}, col_in_291};
assign u_ca_in_292 = {{1{1'b0}}, col_in_292};
assign u_ca_in_293 = {{1{1'b0}}, col_in_293};
assign u_ca_in_294 = {{1{1'b0}}, col_in_294};
assign u_ca_in_295 = {{1{1'b0}}, col_in_295};
assign u_ca_in_296 = {{1{1'b0}}, col_in_296};
assign u_ca_in_297 = {{1{1'b0}}, col_in_297};
assign u_ca_in_298 = {{1{1'b0}}, col_in_298};
assign u_ca_in_299 = {{1{1'b0}}, col_in_299};
assign u_ca_in_300 = {{1{1'b0}}, col_in_300};
assign u_ca_in_301 = {{1{1'b0}}, col_in_301};
assign u_ca_in_302 = {{1{1'b0}}, col_in_302};
assign u_ca_in_303 = {{1{1'b0}}, col_in_303};
assign u_ca_in_304 = {{1{1'b0}}, col_in_304};
assign u_ca_in_305 = {{1{1'b0}}, col_in_305};
assign u_ca_in_306 = {{1{1'b0}}, col_in_306};
assign u_ca_in_307 = {{1{1'b0}}, col_in_307};
assign u_ca_in_308 = {{1{1'b0}}, col_in_308};
assign u_ca_in_309 = {{1{1'b0}}, col_in_309};
assign u_ca_in_310 = {{1{1'b0}}, col_in_310};
assign u_ca_in_311 = {{1{1'b0}}, col_in_311};
assign u_ca_in_312 = {{1{1'b0}}, col_in_312};
assign u_ca_in_313 = {{1{1'b0}}, col_in_313};
assign u_ca_in_314 = {{1{1'b0}}, col_in_314};
assign u_ca_in_315 = {{1{1'b0}}, col_in_315};
assign u_ca_in_316 = {{1{1'b0}}, col_in_316};
assign u_ca_in_317 = {{1{1'b0}}, col_in_317};
assign u_ca_in_318 = {{1{1'b0}}, col_in_318};
assign u_ca_in_319 = {{1{1'b0}}, col_in_319};
assign u_ca_in_320 = {{1{1'b0}}, col_in_320};
assign u_ca_in_321 = {{1{1'b0}}, col_in_321};
assign u_ca_in_322 = {{1{1'b0}}, col_in_322};
assign u_ca_in_323 = {{1{1'b0}}, col_in_323};
assign u_ca_in_324 = {{1{1'b0}}, col_in_324};
assign u_ca_in_325 = {{1{1'b0}}, col_in_325};
assign u_ca_in_326 = {{1{1'b0}}, col_in_326};
assign u_ca_in_327 = {{1{1'b0}}, col_in_327};
assign u_ca_in_328 = {{1{1'b0}}, col_in_328};
assign u_ca_in_329 = {{1{1'b0}}, col_in_329};
assign u_ca_in_330 = {{1{1'b0}}, col_in_330};
assign u_ca_in_331 = {{1{1'b0}}, col_in_331};
assign u_ca_in_332 = {{1{1'b0}}, col_in_332};
assign u_ca_in_333 = {{1{1'b0}}, col_in_333};
assign u_ca_in_334 = {{1{1'b0}}, col_in_334};
assign u_ca_in_335 = {{1{1'b0}}, col_in_335};
assign u_ca_in_336 = {{1{1'b0}}, col_in_336};
assign u_ca_in_337 = {{1{1'b0}}, col_in_337};
assign u_ca_in_338 = {{1{1'b0}}, col_in_338};
assign u_ca_in_339 = {{1{1'b0}}, col_in_339};
assign u_ca_in_340 = {{1{1'b0}}, col_in_340};
assign u_ca_in_341 = {{1{1'b0}}, col_in_341};
assign u_ca_in_342 = {{1{1'b0}}, col_in_342};
assign u_ca_in_343 = {{1{1'b0}}, col_in_343};
assign u_ca_in_344 = {{1{1'b0}}, col_in_344};
assign u_ca_in_345 = {{1{1'b0}}, col_in_345};
assign u_ca_in_346 = {{1{1'b0}}, col_in_346};
assign u_ca_in_347 = {{1{1'b0}}, col_in_347};
assign u_ca_in_348 = {{1{1'b0}}, col_in_348};
assign u_ca_in_349 = {{1{1'b0}}, col_in_349};
assign u_ca_in_350 = {{1{1'b0}}, col_in_350};
assign u_ca_in_351 = {{1{1'b0}}, col_in_351};
assign u_ca_in_352 = {{1{1'b0}}, col_in_352};
assign u_ca_in_353 = {{1{1'b0}}, col_in_353};
assign u_ca_in_354 = {{1{1'b0}}, col_in_354};
assign u_ca_in_355 = {{1{1'b0}}, col_in_355};
assign u_ca_in_356 = {{1{1'b0}}, col_in_356};
assign u_ca_in_357 = {{1{1'b0}}, col_in_357};
assign u_ca_in_358 = {{1{1'b0}}, col_in_358};
assign u_ca_in_359 = {{1{1'b0}}, col_in_359};
assign u_ca_in_360 = {{1{1'b0}}, col_in_360};
assign u_ca_in_361 = {{1{1'b0}}, col_in_361};
assign u_ca_in_362 = {{1{1'b0}}, col_in_362};
assign u_ca_in_363 = {{1{1'b0}}, col_in_363};
assign u_ca_in_364 = {{1{1'b0}}, col_in_364};
assign u_ca_in_365 = {{1{1'b0}}, col_in_365};
assign u_ca_in_366 = {{1{1'b0}}, col_in_366};
assign u_ca_in_367 = {{1{1'b0}}, col_in_367};
assign u_ca_in_368 = {{1{1'b0}}, col_in_368};
assign u_ca_in_369 = {{1{1'b0}}, col_in_369};
assign u_ca_in_370 = {{1{1'b0}}, col_in_370};
assign u_ca_in_371 = {{1{1'b0}}, col_in_371};
assign u_ca_in_372 = {{1{1'b0}}, col_in_372};
assign u_ca_in_373 = {{1{1'b0}}, col_in_373};
assign u_ca_in_374 = {{1{1'b0}}, col_in_374};
assign u_ca_in_375 = {{1{1'b0}}, col_in_375};
assign u_ca_in_376 = {{1{1'b0}}, col_in_376};
assign u_ca_in_377 = {{1{1'b0}}, col_in_377};
assign u_ca_in_378 = {{1{1'b0}}, col_in_378};
assign u_ca_in_379 = {{1{1'b0}}, col_in_379};
assign u_ca_in_380 = {{1{1'b0}}, col_in_380};
assign u_ca_in_381 = {{1{1'b0}}, col_in_381};
assign u_ca_in_382 = {{1{1'b0}}, col_in_382};
assign u_ca_in_383 = {{1{1'b0}}, col_in_383};
assign u_ca_in_384 = {{1{1'b0}}, col_in_384};
assign u_ca_in_385 = {{1{1'b0}}, col_in_385};
assign u_ca_in_386 = {{1{1'b0}}, col_in_386};
assign u_ca_in_387 = {{1{1'b0}}, col_in_387};
assign u_ca_in_388 = {{1{1'b0}}, col_in_388};
assign u_ca_in_389 = {{1{1'b0}}, col_in_389};
assign u_ca_in_390 = {{1{1'b0}}, col_in_390};
assign u_ca_in_391 = {{1{1'b0}}, col_in_391};
assign u_ca_in_392 = {{1{1'b0}}, col_in_392};
assign u_ca_in_393 = {{1{1'b0}}, col_in_393};
assign u_ca_in_394 = {{1{1'b0}}, col_in_394};
assign u_ca_in_395 = {{1{1'b0}}, col_in_395};
assign u_ca_in_396 = {{1{1'b0}}, col_in_396};
assign u_ca_in_397 = {{1{1'b0}}, col_in_397};
assign u_ca_in_398 = {{1{1'b0}}, col_in_398};
assign u_ca_in_399 = {{1{1'b0}}, col_in_399};
assign u_ca_in_400 = {{1{1'b0}}, col_in_400};
assign u_ca_in_401 = {{1{1'b0}}, col_in_401};
assign u_ca_in_402 = {{1{1'b0}}, col_in_402};
assign u_ca_in_403 = {{1{1'b0}}, col_in_403};
assign u_ca_in_404 = {{1{1'b0}}, col_in_404};
assign u_ca_in_405 = {{1{1'b0}}, col_in_405};
assign u_ca_in_406 = {{1{1'b0}}, col_in_406};
assign u_ca_in_407 = {{1{1'b0}}, col_in_407};
assign u_ca_in_408 = {{1{1'b0}}, col_in_408};
assign u_ca_in_409 = {{1{1'b0}}, col_in_409};
assign u_ca_in_410 = {{1{1'b0}}, col_in_410};
assign u_ca_in_411 = {{1{1'b0}}, col_in_411};
assign u_ca_in_412 = {{1{1'b0}}, col_in_412};
assign u_ca_in_413 = {{1{1'b0}}, col_in_413};
assign u_ca_in_414 = {{1{1'b0}}, col_in_414};
assign u_ca_in_415 = {{1{1'b0}}, col_in_415};
assign u_ca_in_416 = {{1{1'b0}}, col_in_416};
assign u_ca_in_417 = {{1{1'b0}}, col_in_417};
assign u_ca_in_418 = {{1{1'b0}}, col_in_418};
assign u_ca_in_419 = {{1{1'b0}}, col_in_419};
assign u_ca_in_420 = {{1{1'b0}}, col_in_420};
assign u_ca_in_421 = {{1{1'b0}}, col_in_421};
assign u_ca_in_422 = {{1{1'b0}}, col_in_422};
assign u_ca_in_423 = {{1{1'b0}}, col_in_423};
assign u_ca_in_424 = {{1{1'b0}}, col_in_424};
assign u_ca_in_425 = {{1{1'b0}}, col_in_425};
assign u_ca_in_426 = {{1{1'b0}}, col_in_426};
assign u_ca_in_427 = {{1{1'b0}}, col_in_427};
assign u_ca_in_428 = {{1{1'b0}}, col_in_428};
assign u_ca_in_429 = {{1{1'b0}}, col_in_429};
assign u_ca_in_430 = {{1{1'b0}}, col_in_430};
assign u_ca_in_431 = {{1{1'b0}}, col_in_431};
assign u_ca_in_432 = {{1{1'b0}}, col_in_432};
assign u_ca_in_433 = {{1{1'b0}}, col_in_433};
assign u_ca_in_434 = {{1{1'b0}}, col_in_434};
assign u_ca_in_435 = {{1{1'b0}}, col_in_435};
assign u_ca_in_436 = {{1{1'b0}}, col_in_436};
assign u_ca_in_437 = {{1{1'b0}}, col_in_437};
assign u_ca_in_438 = {{1{1'b0}}, col_in_438};
assign u_ca_in_439 = {{1{1'b0}}, col_in_439};
assign u_ca_in_440 = {{1{1'b0}}, col_in_440};
assign u_ca_in_441 = {{1{1'b0}}, col_in_441};
assign u_ca_in_442 = {{1{1'b0}}, col_in_442};
assign u_ca_in_443 = {{1{1'b0}}, col_in_443};
assign u_ca_in_444 = {{1{1'b0}}, col_in_444};
assign u_ca_in_445 = {{1{1'b0}}, col_in_445};
assign u_ca_in_446 = {{1{1'b0}}, col_in_446};
assign u_ca_in_447 = {{1{1'b0}}, col_in_447};
assign u_ca_in_448 = {{1{1'b0}}, col_in_448};
assign u_ca_in_449 = {{1{1'b0}}, col_in_449};
assign u_ca_in_450 = {{1{1'b0}}, col_in_450};
assign u_ca_in_451 = {{1{1'b0}}, col_in_451};
assign u_ca_in_452 = {{1{1'b0}}, col_in_452};
assign u_ca_in_453 = {{1{1'b0}}, col_in_453};
assign u_ca_in_454 = {{1{1'b0}}, col_in_454};
assign u_ca_in_455 = {{1{1'b0}}, col_in_455};
assign u_ca_in_456 = {{1{1'b0}}, col_in_456};
assign u_ca_in_457 = {{1{1'b0}}, col_in_457};
assign u_ca_in_458 = {{1{1'b0}}, col_in_458};
assign u_ca_in_459 = {{1{1'b0}}, col_in_459};
assign u_ca_in_460 = {{1{1'b0}}, col_in_460};
assign u_ca_in_461 = {{1{1'b0}}, col_in_461};
assign u_ca_in_462 = {{1{1'b0}}, col_in_462};
assign u_ca_in_463 = {{1{1'b0}}, col_in_463};
assign u_ca_in_464 = {{1{1'b0}}, col_in_464};
assign u_ca_in_465 = {{1{1'b0}}, col_in_465};
assign u_ca_in_466 = {{1{1'b0}}, col_in_466};
assign u_ca_in_467 = {{1{1'b0}}, col_in_467};
assign u_ca_in_468 = {{1{1'b0}}, col_in_468};
assign u_ca_in_469 = {{1{1'b0}}, col_in_469};
assign u_ca_in_470 = {{1{1'b0}}, col_in_470};
assign u_ca_in_471 = {{1{1'b0}}, col_in_471};
assign u_ca_in_472 = {{1{1'b0}}, col_in_472};
assign u_ca_in_473 = {{1{1'b0}}, col_in_473};
assign u_ca_in_474 = {{1{1'b0}}, col_in_474};
assign u_ca_in_475 = {{1{1'b0}}, col_in_475};
assign u_ca_in_476 = {{1{1'b0}}, col_in_476};
assign u_ca_in_477 = {{1{1'b0}}, col_in_477};
assign u_ca_in_478 = {{1{1'b0}}, col_in_478};
assign u_ca_in_479 = {{1{1'b0}}, col_in_479};
assign u_ca_in_480 = {{1{1'b0}}, col_in_480};
assign u_ca_in_481 = {{1{1'b0}}, col_in_481};
assign u_ca_in_482 = {{1{1'b0}}, col_in_482};
assign u_ca_in_483 = {{1{1'b0}}, col_in_483};
assign u_ca_in_484 = {{1{1'b0}}, col_in_484};
assign u_ca_in_485 = {{1{1'b0}}, col_in_485};
assign u_ca_in_486 = {{1{1'b0}}, col_in_486};
assign u_ca_in_487 = {{1{1'b0}}, col_in_487};
assign u_ca_in_488 = {{1{1'b0}}, col_in_488};
assign u_ca_in_489 = {{1{1'b0}}, col_in_489};
assign u_ca_in_490 = {{1{1'b0}}, col_in_490};
assign u_ca_in_491 = {{1{1'b0}}, col_in_491};
assign u_ca_in_492 = {{1{1'b0}}, col_in_492};
assign u_ca_in_493 = {{1{1'b0}}, col_in_493};
assign u_ca_in_494 = {{1{1'b0}}, col_in_494};
assign u_ca_in_495 = {{1{1'b0}}, col_in_495};
assign u_ca_in_496 = {{1{1'b0}}, col_in_496};
assign u_ca_in_497 = {{1{1'b0}}, col_in_497};
assign u_ca_in_498 = {{1{1'b0}}, col_in_498};
assign u_ca_in_499 = {{1{1'b0}}, col_in_499};
assign u_ca_in_500 = {{1{1'b0}}, col_in_500};
assign u_ca_in_501 = {{1{1'b0}}, col_in_501};
assign u_ca_in_502 = {{1{1'b0}}, col_in_502};
assign u_ca_in_503 = {{1{1'b0}}, col_in_503};
assign u_ca_in_504 = {{1{1'b0}}, col_in_504};
assign u_ca_in_505 = {{1{1'b0}}, col_in_505};
assign u_ca_in_506 = {{1{1'b0}}, col_in_506};
assign u_ca_in_507 = {{1{1'b0}}, col_in_507};
assign u_ca_in_508 = {{1{1'b0}}, col_in_508};
assign u_ca_in_509 = {{1{1'b0}}, col_in_509};
assign u_ca_in_510 = {{1{1'b0}}, col_in_510};
assign u_ca_in_511 = {{1{1'b0}}, col_in_511};
assign u_ca_in_512 = {{1{1'b0}}, col_in_512};
assign u_ca_in_513 = {{1{1'b0}}, col_in_513};
assign u_ca_in_514 = {{1{1'b0}}, col_in_514};
assign u_ca_in_515 = {{1{1'b0}}, col_in_515};
assign u_ca_in_516 = {{1{1'b0}}, col_in_516};
assign u_ca_in_517 = {{1{1'b0}}, col_in_517};
assign u_ca_in_518 = {{1{1'b0}}, col_in_518};
assign u_ca_in_519 = {{1{1'b0}}, col_in_519};
assign u_ca_in_520 = {{1{1'b0}}, col_in_520};
assign u_ca_in_521 = {{1{1'b0}}, col_in_521};
assign u_ca_in_522 = {{1{1'b0}}, col_in_522};
assign u_ca_in_523 = {{1{1'b0}}, col_in_523};
assign u_ca_in_524 = {{1{1'b0}}, col_in_524};
assign u_ca_in_525 = {{1{1'b0}}, col_in_525};
assign u_ca_in_526 = {{1{1'b0}}, col_in_526};
assign u_ca_in_527 = {{1{1'b0}}, col_in_527};
assign u_ca_in_528 = {{1{1'b0}}, col_in_528};
assign u_ca_in_529 = {{1{1'b0}}, col_in_529};
assign u_ca_in_530 = {{1{1'b0}}, col_in_530};
assign u_ca_in_531 = {{1{1'b0}}, col_in_531};
assign u_ca_in_532 = {{1{1'b0}}, col_in_532};
assign u_ca_in_533 = {{1{1'b0}}, col_in_533};
assign u_ca_in_534 = {{1{1'b0}}, col_in_534};
assign u_ca_in_535 = {{1{1'b0}}, col_in_535};
assign u_ca_in_536 = {{1{1'b0}}, col_in_536};
assign u_ca_in_537 = {{1{1'b0}}, col_in_537};
assign u_ca_in_538 = {{1{1'b0}}, col_in_538};
assign u_ca_in_539 = {{1{1'b0}}, col_in_539};
assign u_ca_in_540 = {{1{1'b0}}, col_in_540};
assign u_ca_in_541 = {{1{1'b0}}, col_in_541};
assign u_ca_in_542 = {{1{1'b0}}, col_in_542};
assign u_ca_in_543 = {{1{1'b0}}, col_in_543};
assign u_ca_in_544 = {{1{1'b0}}, col_in_544};
assign u_ca_in_545 = {{1{1'b0}}, col_in_545};
assign u_ca_in_546 = {{1{1'b0}}, col_in_546};
assign u_ca_in_547 = {{1{1'b0}}, col_in_547};
assign u_ca_in_548 = {{1{1'b0}}, col_in_548};
assign u_ca_in_549 = {{1{1'b0}}, col_in_549};
assign u_ca_in_550 = {{1{1'b0}}, col_in_550};
assign u_ca_in_551 = {{1{1'b0}}, col_in_551};
assign u_ca_in_552 = {{1{1'b0}}, col_in_552};
assign u_ca_in_553 = {{1{1'b0}}, col_in_553};
assign u_ca_in_554 = {{1{1'b0}}, col_in_554};
assign u_ca_in_555 = {{1{1'b0}}, col_in_555};
assign u_ca_in_556 = {{1{1'b0}}, col_in_556};
assign u_ca_in_557 = {{1{1'b0}}, col_in_557};
assign u_ca_in_558 = {{1{1'b0}}, col_in_558};
assign u_ca_in_559 = {{1{1'b0}}, col_in_559};
assign u_ca_in_560 = {{1{1'b0}}, col_in_560};
assign u_ca_in_561 = {{1{1'b0}}, col_in_561};
assign u_ca_in_562 = {{1{1'b0}}, col_in_562};
assign u_ca_in_563 = {{1{1'b0}}, col_in_563};
assign u_ca_in_564 = {{1{1'b0}}, col_in_564};
assign u_ca_in_565 = {{1{1'b0}}, col_in_565};
assign u_ca_in_566 = {{1{1'b0}}, col_in_566};
assign u_ca_in_567 = {{1{1'b0}}, col_in_567};
assign u_ca_in_568 = {{1{1'b0}}, col_in_568};
assign u_ca_in_569 = {{1{1'b0}}, col_in_569};
assign u_ca_in_570 = {{1{1'b0}}, col_in_570};
assign u_ca_in_571 = {{1{1'b0}}, col_in_571};
assign u_ca_in_572 = {{1{1'b0}}, col_in_572};
assign u_ca_in_573 = {{1{1'b0}}, col_in_573};
assign u_ca_in_574 = {{1{1'b0}}, col_in_574};
assign u_ca_in_575 = {{1{1'b0}}, col_in_575};
assign u_ca_in_576 = {{1{1'b0}}, col_in_576};
assign u_ca_in_577 = {{1{1'b0}}, col_in_577};
assign u_ca_in_578 = {{1{1'b0}}, col_in_578};
assign u_ca_in_579 = {{1{1'b0}}, col_in_579};
assign u_ca_in_580 = {{1{1'b0}}, col_in_580};
assign u_ca_in_581 = {{1{1'b0}}, col_in_581};
assign u_ca_in_582 = {{1{1'b0}}, col_in_582};
assign u_ca_in_583 = {{1{1'b0}}, col_in_583};
assign u_ca_in_584 = {{1{1'b0}}, col_in_584};
assign u_ca_in_585 = {{1{1'b0}}, col_in_585};
assign u_ca_in_586 = {{1{1'b0}}, col_in_586};
assign u_ca_in_587 = {{1{1'b0}}, col_in_587};
assign u_ca_in_588 = {{1{1'b0}}, col_in_588};
assign u_ca_in_589 = {{1{1'b0}}, col_in_589};
assign u_ca_in_590 = {{1{1'b0}}, col_in_590};
assign u_ca_in_591 = {{1{1'b0}}, col_in_591};
assign u_ca_in_592 = {{1{1'b0}}, col_in_592};
assign u_ca_in_593 = {{1{1'b0}}, col_in_593};
assign u_ca_in_594 = {{1{1'b0}}, col_in_594};
assign u_ca_in_595 = {{1{1'b0}}, col_in_595};
assign u_ca_in_596 = {{1{1'b0}}, col_in_596};
assign u_ca_in_597 = {{1{1'b0}}, col_in_597};
assign u_ca_in_598 = {{1{1'b0}}, col_in_598};
assign u_ca_in_599 = {{1{1'b0}}, col_in_599};
assign u_ca_in_600 = {{1{1'b0}}, col_in_600};
assign u_ca_in_601 = {{1{1'b0}}, col_in_601};
assign u_ca_in_602 = {{1{1'b0}}, col_in_602};
assign u_ca_in_603 = {{1{1'b0}}, col_in_603};
assign u_ca_in_604 = {{1{1'b0}}, col_in_604};
assign u_ca_in_605 = {{1{1'b0}}, col_in_605};
assign u_ca_in_606 = {{1{1'b0}}, col_in_606};
assign u_ca_in_607 = {{1{1'b0}}, col_in_607};
assign u_ca_in_608 = {{1{1'b0}}, col_in_608};
assign u_ca_in_609 = {{1{1'b0}}, col_in_609};
assign u_ca_in_610 = {{1{1'b0}}, col_in_610};
assign u_ca_in_611 = {{1{1'b0}}, col_in_611};
assign u_ca_in_612 = {{1{1'b0}}, col_in_612};
assign u_ca_in_613 = {{1{1'b0}}, col_in_613};
assign u_ca_in_614 = {{1{1'b0}}, col_in_614};
assign u_ca_in_615 = {{1{1'b0}}, col_in_615};
assign u_ca_in_616 = {{1{1'b0}}, col_in_616};
assign u_ca_in_617 = {{1{1'b0}}, col_in_617};
assign u_ca_in_618 = {{1{1'b0}}, col_in_618};
assign u_ca_in_619 = {{1{1'b0}}, col_in_619};
assign u_ca_in_620 = {{1{1'b0}}, col_in_620};
assign u_ca_in_621 = {{1{1'b0}}, col_in_621};
assign u_ca_in_622 = {{1{1'b0}}, col_in_622};
assign u_ca_in_623 = {{1{1'b0}}, col_in_623};
assign u_ca_in_624 = {{1{1'b0}}, col_in_624};
assign u_ca_in_625 = {{1{1'b0}}, col_in_625};
assign u_ca_in_626 = {{1{1'b0}}, col_in_626};
assign u_ca_in_627 = {{1{1'b0}}, col_in_627};
assign u_ca_in_628 = {{1{1'b0}}, col_in_628};
assign u_ca_in_629 = {{1{1'b0}}, col_in_629};
assign u_ca_in_630 = {{1{1'b0}}, col_in_630};
assign u_ca_in_631 = {{1{1'b0}}, col_in_631};
assign u_ca_in_632 = {{1{1'b0}}, col_in_632};
assign u_ca_in_633 = {{1{1'b0}}, col_in_633};
assign u_ca_in_634 = {{1{1'b0}}, col_in_634};
assign u_ca_in_635 = {{1{1'b0}}, col_in_635};
assign u_ca_in_636 = {{1{1'b0}}, col_in_636};
assign u_ca_in_637 = {{1{1'b0}}, col_in_637};
assign u_ca_in_638 = {{1{1'b0}}, col_in_638};
assign u_ca_in_639 = {{1{1'b0}}, col_in_639};
assign u_ca_in_640 = {{1{1'b0}}, col_in_640};
assign u_ca_in_641 = {{1{1'b0}}, col_in_641};
assign u_ca_in_642 = {{1{1'b0}}, col_in_642};
assign u_ca_in_643 = {{1{1'b0}}, col_in_643};
assign u_ca_in_644 = {{1{1'b0}}, col_in_644};
assign u_ca_in_645 = {{1{1'b0}}, col_in_645};
assign u_ca_in_646 = {{1{1'b0}}, col_in_646};
assign u_ca_in_647 = {{1{1'b0}}, col_in_647};
assign u_ca_in_648 = {{1{1'b0}}, col_in_648};
assign u_ca_in_649 = {{1{1'b0}}, col_in_649};
assign u_ca_in_650 = {{1{1'b0}}, col_in_650};
assign u_ca_in_651 = {{1{1'b0}}, col_in_651};
assign u_ca_in_652 = {{1{1'b0}}, col_in_652};
assign u_ca_in_653 = {{1{1'b0}}, col_in_653};
assign u_ca_in_654 = {{1{1'b0}}, col_in_654};
assign u_ca_in_655 = {{1{1'b0}}, col_in_655};
assign u_ca_in_656 = {{1{1'b0}}, col_in_656};
assign u_ca_in_657 = {{1{1'b0}}, col_in_657};
assign u_ca_in_658 = {{1{1'b0}}, col_in_658};
assign u_ca_in_659 = {{1{1'b0}}, col_in_659};
assign u_ca_in_660 = {{1{1'b0}}, col_in_660};
assign u_ca_in_661 = {{1{1'b0}}, col_in_661};
assign u_ca_in_662 = {{1{1'b0}}, col_in_662};
assign u_ca_in_663 = {{1{1'b0}}, col_in_663};
assign u_ca_in_664 = {{1{1'b0}}, col_in_664};
assign u_ca_in_665 = {{1{1'b0}}, col_in_665};
assign u_ca_in_666 = {{1{1'b0}}, col_in_666};
assign u_ca_in_667 = {{1{1'b0}}, col_in_667};
assign u_ca_in_668 = {{1{1'b0}}, col_in_668};
assign u_ca_in_669 = {{1{1'b0}}, col_in_669};
assign u_ca_in_670 = {{1{1'b0}}, col_in_670};
assign u_ca_in_671 = {{1{1'b0}}, col_in_671};
assign u_ca_in_672 = {{1{1'b0}}, col_in_672};
assign u_ca_in_673 = {{1{1'b0}}, col_in_673};
assign u_ca_in_674 = {{1{1'b0}}, col_in_674};
assign u_ca_in_675 = {{1{1'b0}}, col_in_675};
assign u_ca_in_676 = {{1{1'b0}}, col_in_676};
assign u_ca_in_677 = {{1{1'b0}}, col_in_677};
assign u_ca_in_678 = {{1{1'b0}}, col_in_678};
assign u_ca_in_679 = {{1{1'b0}}, col_in_679};
assign u_ca_in_680 = {{1{1'b0}}, col_in_680};
assign u_ca_in_681 = {{1{1'b0}}, col_in_681};
assign u_ca_in_682 = {{1{1'b0}}, col_in_682};
assign u_ca_in_683 = {{1{1'b0}}, col_in_683};
assign u_ca_in_684 = {{1{1'b0}}, col_in_684};
assign u_ca_in_685 = {{1{1'b0}}, col_in_685};
assign u_ca_in_686 = {{1{1'b0}}, col_in_686};
assign u_ca_in_687 = {{1{1'b0}}, col_in_687};
assign u_ca_in_688 = {{1{1'b0}}, col_in_688};
assign u_ca_in_689 = {{1{1'b0}}, col_in_689};
assign u_ca_in_690 = {{1{1'b0}}, col_in_690};
assign u_ca_in_691 = {{1{1'b0}}, col_in_691};
assign u_ca_in_692 = {{1{1'b0}}, col_in_692};
assign u_ca_in_693 = {{1{1'b0}}, col_in_693};
assign u_ca_in_694 = {{1{1'b0}}, col_in_694};
assign u_ca_in_695 = {{1{1'b0}}, col_in_695};
assign u_ca_in_696 = {{1{1'b0}}, col_in_696};
assign u_ca_in_697 = {{1{1'b0}}, col_in_697};
assign u_ca_in_698 = {{1{1'b0}}, col_in_698};
assign u_ca_in_699 = {{1{1'b0}}, col_in_699};
assign u_ca_in_700 = {{1{1'b0}}, col_in_700};
assign u_ca_in_701 = {{1{1'b0}}, col_in_701};
assign u_ca_in_702 = {{1{1'b0}}, col_in_702};
assign u_ca_in_703 = {{1{1'b0}}, col_in_703};
assign u_ca_in_704 = {{1{1'b0}}, col_in_704};
assign u_ca_in_705 = {{1{1'b0}}, col_in_705};
assign u_ca_in_706 = {{1{1'b0}}, col_in_706};
assign u_ca_in_707 = {{1{1'b0}}, col_in_707};
assign u_ca_in_708 = {{1{1'b0}}, col_in_708};
assign u_ca_in_709 = {{1{1'b0}}, col_in_709};
assign u_ca_in_710 = {{1{1'b0}}, col_in_710};
assign u_ca_in_711 = {{1{1'b0}}, col_in_711};
assign u_ca_in_712 = {{1{1'b0}}, col_in_712};
assign u_ca_in_713 = {{1{1'b0}}, col_in_713};
assign u_ca_in_714 = {{1{1'b0}}, col_in_714};
assign u_ca_in_715 = {{1{1'b0}}, col_in_715};
assign u_ca_in_716 = {{1{1'b0}}, col_in_716};
assign u_ca_in_717 = {{1{1'b0}}, col_in_717};
assign u_ca_in_718 = {{1{1'b0}}, col_in_718};
assign u_ca_in_719 = {{1{1'b0}}, col_in_719};
assign u_ca_in_720 = {{1{1'b0}}, col_in_720};
assign u_ca_in_721 = {{1{1'b0}}, col_in_721};
assign u_ca_in_722 = {{1{1'b0}}, col_in_722};
assign u_ca_in_723 = {{1{1'b0}}, col_in_723};
assign u_ca_in_724 = {{1{1'b0}}, col_in_724};
assign u_ca_in_725 = {{1{1'b0}}, col_in_725};
assign u_ca_in_726 = {{1{1'b0}}, col_in_726};
assign u_ca_in_727 = {{1{1'b0}}, col_in_727};
assign u_ca_in_728 = {{1{1'b0}}, col_in_728};
assign u_ca_in_729 = {{1{1'b0}}, col_in_729};
assign u_ca_in_730 = {{1{1'b0}}, col_in_730};
assign u_ca_in_731 = {{1{1'b0}}, col_in_731};
assign u_ca_in_732 = {{1{1'b0}}, col_in_732};
assign u_ca_in_733 = {{1{1'b0}}, col_in_733};
assign u_ca_in_734 = {{1{1'b0}}, col_in_734};
assign u_ca_in_735 = {{1{1'b0}}, col_in_735};
assign u_ca_in_736 = {{1{1'b0}}, col_in_736};
assign u_ca_in_737 = {{1{1'b0}}, col_in_737};
assign u_ca_in_738 = {{1{1'b0}}, col_in_738};
assign u_ca_in_739 = {{1{1'b0}}, col_in_739};
assign u_ca_in_740 = {{1{1'b0}}, col_in_740};
assign u_ca_in_741 = {{1{1'b0}}, col_in_741};
assign u_ca_in_742 = {{1{1'b0}}, col_in_742};
assign u_ca_in_743 = {{1{1'b0}}, col_in_743};
assign u_ca_in_744 = {{1{1'b0}}, col_in_744};
assign u_ca_in_745 = {{1{1'b0}}, col_in_745};
assign u_ca_in_746 = {{1{1'b0}}, col_in_746};
assign u_ca_in_747 = {{1{1'b0}}, col_in_747};
assign u_ca_in_748 = {{1{1'b0}}, col_in_748};
assign u_ca_in_749 = {{1{1'b0}}, col_in_749};
assign u_ca_in_750 = {{1{1'b0}}, col_in_750};
assign u_ca_in_751 = {{1{1'b0}}, col_in_751};
assign u_ca_in_752 = {{1{1'b0}}, col_in_752};
assign u_ca_in_753 = {{1{1'b0}}, col_in_753};
assign u_ca_in_754 = {{1{1'b0}}, col_in_754};
assign u_ca_in_755 = {{1{1'b0}}, col_in_755};
assign u_ca_in_756 = {{1{1'b0}}, col_in_756};
assign u_ca_in_757 = {{1{1'b0}}, col_in_757};
assign u_ca_in_758 = {{1{1'b0}}, col_in_758};
assign u_ca_in_759 = {{1{1'b0}}, col_in_759};
assign u_ca_in_760 = {{1{1'b0}}, col_in_760};
assign u_ca_in_761 = {{1{1'b0}}, col_in_761};
assign u_ca_in_762 = {{1{1'b0}}, col_in_762};
assign u_ca_in_763 = {{1{1'b0}}, col_in_763};
assign u_ca_in_764 = {{1{1'b0}}, col_in_764};
assign u_ca_in_765 = {{1{1'b0}}, col_in_765};
assign u_ca_in_766 = {{1{1'b0}}, col_in_766};
assign u_ca_in_767 = {{1{1'b0}}, col_in_767};
assign u_ca_in_768 = {{1{1'b0}}, col_in_768};
assign u_ca_in_769 = {{1{1'b0}}, col_in_769};
assign u_ca_in_770 = {{1{1'b0}}, col_in_770};
assign u_ca_in_771 = {{1{1'b0}}, col_in_771};
assign u_ca_in_772 = {{1{1'b0}}, col_in_772};
assign u_ca_in_773 = {{1{1'b0}}, col_in_773};
assign u_ca_in_774 = {{1{1'b0}}, col_in_774};
assign u_ca_in_775 = {{1{1'b0}}, col_in_775};
assign u_ca_in_776 = {{1{1'b0}}, col_in_776};
assign u_ca_in_777 = {{1{1'b0}}, col_in_777};
assign u_ca_in_778 = {{1{1'b0}}, col_in_778};
assign u_ca_in_779 = {{1{1'b0}}, col_in_779};
assign u_ca_in_780 = {{1{1'b0}}, col_in_780};
assign u_ca_in_781 = {{1{1'b0}}, col_in_781};
assign u_ca_in_782 = {{1{1'b0}}, col_in_782};
assign u_ca_in_783 = {{1{1'b0}}, col_in_783};
assign u_ca_in_784 = {{1{1'b0}}, col_in_784};
assign u_ca_in_785 = {{1{1'b0}}, col_in_785};
assign u_ca_in_786 = {{1{1'b0}}, col_in_786};
assign u_ca_in_787 = {{1{1'b0}}, col_in_787};
assign u_ca_in_788 = {{1{1'b0}}, col_in_788};
assign u_ca_in_789 = {{1{1'b0}}, col_in_789};
assign u_ca_in_790 = {{1{1'b0}}, col_in_790};
assign u_ca_in_791 = {{1{1'b0}}, col_in_791};
assign u_ca_in_792 = {{1{1'b0}}, col_in_792};
assign u_ca_in_793 = {{1{1'b0}}, col_in_793};
assign u_ca_in_794 = {{1{1'b0}}, col_in_794};
assign u_ca_in_795 = {{1{1'b0}}, col_in_795};
assign u_ca_in_796 = {{1{1'b0}}, col_in_796};
assign u_ca_in_797 = {{1{1'b0}}, col_in_797};
assign u_ca_in_798 = {{1{1'b0}}, col_in_798};
assign u_ca_in_799 = {{1{1'b0}}, col_in_799};
assign u_ca_in_800 = {{1{1'b0}}, col_in_800};
assign u_ca_in_801 = {{1{1'b0}}, col_in_801};
assign u_ca_in_802 = {{1{1'b0}}, col_in_802};
assign u_ca_in_803 = {{1{1'b0}}, col_in_803};
assign u_ca_in_804 = {{1{1'b0}}, col_in_804};
assign u_ca_in_805 = {{1{1'b0}}, col_in_805};
assign u_ca_in_806 = {{1{1'b0}}, col_in_806};
assign u_ca_in_807 = {{1{1'b0}}, col_in_807};
assign u_ca_in_808 = {{1{1'b0}}, col_in_808};
assign u_ca_in_809 = {{1{1'b0}}, col_in_809};
assign u_ca_in_810 = {{1{1'b0}}, col_in_810};
assign u_ca_in_811 = {{1{1'b0}}, col_in_811};
assign u_ca_in_812 = {{1{1'b0}}, col_in_812};
assign u_ca_in_813 = {{1{1'b0}}, col_in_813};
assign u_ca_in_814 = {{1{1'b0}}, col_in_814};
assign u_ca_in_815 = {{1{1'b0}}, col_in_815};
assign u_ca_in_816 = {{1{1'b0}}, col_in_816};
assign u_ca_in_817 = {{1{1'b0}}, col_in_817};
assign u_ca_in_818 = {{1{1'b0}}, col_in_818};
assign u_ca_in_819 = {{1{1'b0}}, col_in_819};
assign u_ca_in_820 = {{1{1'b0}}, col_in_820};
assign u_ca_in_821 = {{1{1'b0}}, col_in_821};
assign u_ca_in_822 = {{1{1'b0}}, col_in_822};
assign u_ca_in_823 = {{1{1'b0}}, col_in_823};
assign u_ca_in_824 = {{1{1'b0}}, col_in_824};
assign u_ca_in_825 = {{1{1'b0}}, col_in_825};
assign u_ca_in_826 = {{1{1'b0}}, col_in_826};
assign u_ca_in_827 = {{1{1'b0}}, col_in_827};
assign u_ca_in_828 = {{1{1'b0}}, col_in_828};
assign u_ca_in_829 = {{1{1'b0}}, col_in_829};
assign u_ca_in_830 = {{1{1'b0}}, col_in_830};
assign u_ca_in_831 = {{1{1'b0}}, col_in_831};
assign u_ca_in_832 = {{1{1'b0}}, col_in_832};
assign u_ca_in_833 = {{1{1'b0}}, col_in_833};
assign u_ca_in_834 = {{1{1'b0}}, col_in_834};
assign u_ca_in_835 = {{1{1'b0}}, col_in_835};
assign u_ca_in_836 = {{1{1'b0}}, col_in_836};
assign u_ca_in_837 = {{1{1'b0}}, col_in_837};
assign u_ca_in_838 = {{1{1'b0}}, col_in_838};
assign u_ca_in_839 = {{1{1'b0}}, col_in_839};
assign u_ca_in_840 = {{1{1'b0}}, col_in_840};
assign u_ca_in_841 = {{1{1'b0}}, col_in_841};
assign u_ca_in_842 = {{1{1'b0}}, col_in_842};
assign u_ca_in_843 = {{1{1'b0}}, col_in_843};
assign u_ca_in_844 = {{1{1'b0}}, col_in_844};
assign u_ca_in_845 = {{1{1'b0}}, col_in_845};
assign u_ca_in_846 = {{1{1'b0}}, col_in_846};
assign u_ca_in_847 = {{1{1'b0}}, col_in_847};
assign u_ca_in_848 = {{1{1'b0}}, col_in_848};
assign u_ca_in_849 = {{1{1'b0}}, col_in_849};
assign u_ca_in_850 = {{1{1'b0}}, col_in_850};
assign u_ca_in_851 = {{1{1'b0}}, col_in_851};
assign u_ca_in_852 = {{1{1'b0}}, col_in_852};
assign u_ca_in_853 = {{1{1'b0}}, col_in_853};
assign u_ca_in_854 = {{1{1'b0}}, col_in_854};
assign u_ca_in_855 = {{1{1'b0}}, col_in_855};
assign u_ca_in_856 = {{1{1'b0}}, col_in_856};
assign u_ca_in_857 = {{1{1'b0}}, col_in_857};
assign u_ca_in_858 = {{1{1'b0}}, col_in_858};
assign u_ca_in_859 = {{1{1'b0}}, col_in_859};
assign u_ca_in_860 = {{1{1'b0}}, col_in_860};
assign u_ca_in_861 = {{1{1'b0}}, col_in_861};
assign u_ca_in_862 = {{1{1'b0}}, col_in_862};
assign u_ca_in_863 = {{1{1'b0}}, col_in_863};
assign u_ca_in_864 = {{1{1'b0}}, col_in_864};
assign u_ca_in_865 = {{1{1'b0}}, col_in_865};
assign u_ca_in_866 = {{1{1'b0}}, col_in_866};
assign u_ca_in_867 = {{1{1'b0}}, col_in_867};
assign u_ca_in_868 = {{1{1'b0}}, col_in_868};
assign u_ca_in_869 = {{1{1'b0}}, col_in_869};
assign u_ca_in_870 = {{1{1'b0}}, col_in_870};
assign u_ca_in_871 = {{1{1'b0}}, col_in_871};
assign u_ca_in_872 = {{1{1'b0}}, col_in_872};
assign u_ca_in_873 = {{1{1'b0}}, col_in_873};
assign u_ca_in_874 = {{1{1'b0}}, col_in_874};
assign u_ca_in_875 = {{1{1'b0}}, col_in_875};
assign u_ca_in_876 = {{1{1'b0}}, col_in_876};
assign u_ca_in_877 = {{1{1'b0}}, col_in_877};
assign u_ca_in_878 = {{1{1'b0}}, col_in_878};
assign u_ca_in_879 = {{1{1'b0}}, col_in_879};
assign u_ca_in_880 = {{1{1'b0}}, col_in_880};
assign u_ca_in_881 = {{1{1'b0}}, col_in_881};
assign u_ca_in_882 = {{1{1'b0}}, col_in_882};
assign u_ca_in_883 = {{1{1'b0}}, col_in_883};
assign u_ca_in_884 = {{1{1'b0}}, col_in_884};
assign u_ca_in_885 = {{1{1'b0}}, col_in_885};
assign u_ca_in_886 = {{1{1'b0}}, col_in_886};
assign u_ca_in_887 = {{1{1'b0}}, col_in_887};
assign u_ca_in_888 = {{1{1'b0}}, col_in_888};
assign u_ca_in_889 = {{1{1'b0}}, col_in_889};
assign u_ca_in_890 = {{1{1'b0}}, col_in_890};
assign u_ca_in_891 = {{1{1'b0}}, col_in_891};
assign u_ca_in_892 = {{1{1'b0}}, col_in_892};
assign u_ca_in_893 = {{1{1'b0}}, col_in_893};
assign u_ca_in_894 = {{1{1'b0}}, col_in_894};
assign u_ca_in_895 = {{1{1'b0}}, col_in_895};
assign u_ca_in_896 = {{1{1'b0}}, col_in_896};
assign u_ca_in_897 = {{1{1'b0}}, col_in_897};
assign u_ca_in_898 = {{1{1'b0}}, col_in_898};
assign u_ca_in_899 = {{1{1'b0}}, col_in_899};
assign u_ca_in_900 = {{1{1'b0}}, col_in_900};
assign u_ca_in_901 = {{1{1'b0}}, col_in_901};
assign u_ca_in_902 = {{1{1'b0}}, col_in_902};
assign u_ca_in_903 = {{1{1'b0}}, col_in_903};
assign u_ca_in_904 = {{1{1'b0}}, col_in_904};
assign u_ca_in_905 = {{1{1'b0}}, col_in_905};
assign u_ca_in_906 = {{1{1'b0}}, col_in_906};
assign u_ca_in_907 = {{1{1'b0}}, col_in_907};
assign u_ca_in_908 = {{1{1'b0}}, col_in_908};
assign u_ca_in_909 = {{1{1'b0}}, col_in_909};
assign u_ca_in_910 = {{1{1'b0}}, col_in_910};
assign u_ca_in_911 = {{1{1'b0}}, col_in_911};
assign u_ca_in_912 = {{1{1'b0}}, col_in_912};
assign u_ca_in_913 = {{1{1'b0}}, col_in_913};
assign u_ca_in_914 = {{1{1'b0}}, col_in_914};
assign u_ca_in_915 = {{1{1'b0}}, col_in_915};
assign u_ca_in_916 = {{1{1'b0}}, col_in_916};
assign u_ca_in_917 = {{1{1'b0}}, col_in_917};
assign u_ca_in_918 = {{1{1'b0}}, col_in_918};
assign u_ca_in_919 = {{1{1'b0}}, col_in_919};
assign u_ca_in_920 = {{1{1'b0}}, col_in_920};
assign u_ca_in_921 = {{1{1'b0}}, col_in_921};
assign u_ca_in_922 = {{1{1'b0}}, col_in_922};
assign u_ca_in_923 = {{1{1'b0}}, col_in_923};
assign u_ca_in_924 = {{1{1'b0}}, col_in_924};
assign u_ca_in_925 = {{1{1'b0}}, col_in_925};
assign u_ca_in_926 = {{1{1'b0}}, col_in_926};
assign u_ca_in_927 = {{1{1'b0}}, col_in_927};
assign u_ca_in_928 = {{1{1'b0}}, col_in_928};
assign u_ca_in_929 = {{1{1'b0}}, col_in_929};
assign u_ca_in_930 = {{1{1'b0}}, col_in_930};
assign u_ca_in_931 = {{1{1'b0}}, col_in_931};
assign u_ca_in_932 = {{1{1'b0}}, col_in_932};
assign u_ca_in_933 = {{1{1'b0}}, col_in_933};
assign u_ca_in_934 = {{1{1'b0}}, col_in_934};
assign u_ca_in_935 = {{1{1'b0}}, col_in_935};
assign u_ca_in_936 = {{1{1'b0}}, col_in_936};
assign u_ca_in_937 = {{1{1'b0}}, col_in_937};
assign u_ca_in_938 = {{1{1'b0}}, col_in_938};
assign u_ca_in_939 = {{1{1'b0}}, col_in_939};
assign u_ca_in_940 = {{1{1'b0}}, col_in_940};
assign u_ca_in_941 = {{1{1'b0}}, col_in_941};
assign u_ca_in_942 = {{1{1'b0}}, col_in_942};
assign u_ca_in_943 = {{1{1'b0}}, col_in_943};
assign u_ca_in_944 = {{1{1'b0}}, col_in_944};
assign u_ca_in_945 = {{1{1'b0}}, col_in_945};
assign u_ca_in_946 = {{1{1'b0}}, col_in_946};
assign u_ca_in_947 = {{1{1'b0}}, col_in_947};
assign u_ca_in_948 = {{1{1'b0}}, col_in_948};
assign u_ca_in_949 = {{1{1'b0}}, col_in_949};
assign u_ca_in_950 = {{1{1'b0}}, col_in_950};
assign u_ca_in_951 = {{1{1'b0}}, col_in_951};
assign u_ca_in_952 = {{1{1'b0}}, col_in_952};
assign u_ca_in_953 = {{1{1'b0}}, col_in_953};
assign u_ca_in_954 = {{1{1'b0}}, col_in_954};
assign u_ca_in_955 = {{1{1'b0}}, col_in_955};
assign u_ca_in_956 = {{1{1'b0}}, col_in_956};
assign u_ca_in_957 = {{1{1'b0}}, col_in_957};
assign u_ca_in_958 = {{1{1'b0}}, col_in_958};
assign u_ca_in_959 = {{1{1'b0}}, col_in_959};
assign u_ca_in_960 = {{1{1'b0}}, col_in_960};
assign u_ca_in_961 = {{1{1'b0}}, col_in_961};
assign u_ca_in_962 = {{1{1'b0}}, col_in_962};
assign u_ca_in_963 = {{1{1'b0}}, col_in_963};
assign u_ca_in_964 = {{1{1'b0}}, col_in_964};
assign u_ca_in_965 = {{1{1'b0}}, col_in_965};
assign u_ca_in_966 = {{1{1'b0}}, col_in_966};
assign u_ca_in_967 = {{1{1'b0}}, col_in_967};
assign u_ca_in_968 = {{1{1'b0}}, col_in_968};
assign u_ca_in_969 = {{1{1'b0}}, col_in_969};
assign u_ca_in_970 = {{1{1'b0}}, col_in_970};
assign u_ca_in_971 = {{1{1'b0}}, col_in_971};
assign u_ca_in_972 = {{1{1'b0}}, col_in_972};
assign u_ca_in_973 = {{1{1'b0}}, col_in_973};
assign u_ca_in_974 = {{1{1'b0}}, col_in_974};
assign u_ca_in_975 = {{1{1'b0}}, col_in_975};
assign u_ca_in_976 = {{1{1'b0}}, col_in_976};
assign u_ca_in_977 = {{1{1'b0}}, col_in_977};
assign u_ca_in_978 = {{1{1'b0}}, col_in_978};
assign u_ca_in_979 = {{1{1'b0}}, col_in_979};
assign u_ca_in_980 = {{1{1'b0}}, col_in_980};
assign u_ca_in_981 = {{1{1'b0}}, col_in_981};
assign u_ca_in_982 = {{1{1'b0}}, col_in_982};
assign u_ca_in_983 = {{1{1'b0}}, col_in_983};
assign u_ca_in_984 = {{1{1'b0}}, col_in_984};
assign u_ca_in_985 = {{1{1'b0}}, col_in_985};
assign u_ca_in_986 = {{1{1'b0}}, col_in_986};
assign u_ca_in_987 = {{1{1'b0}}, col_in_987};
assign u_ca_in_988 = {{1{1'b0}}, col_in_988};
assign u_ca_in_989 = {{1{1'b0}}, col_in_989};
assign u_ca_in_990 = {{1{1'b0}}, col_in_990};
assign u_ca_in_991 = {{1{1'b0}}, col_in_991};
assign u_ca_in_992 = {{1{1'b0}}, col_in_992};
assign u_ca_in_993 = {{1{1'b0}}, col_in_993};
assign u_ca_in_994 = {{1{1'b0}}, col_in_994};
assign u_ca_in_995 = {{1{1'b0}}, col_in_995};
assign u_ca_in_996 = {{1{1'b0}}, col_in_996};
assign u_ca_in_997 = {{1{1'b0}}, col_in_997};
assign u_ca_in_998 = {{1{1'b0}}, col_in_998};
assign u_ca_in_999 = {{1{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{1{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{1{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{1{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{1{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{1{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{1{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{1{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{1{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{1{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{1{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{1{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{1{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{1{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{1{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{1{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{1{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{1{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{1{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{1{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{1{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{1{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{1{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{1{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{1{1'b0}}, col_in_1023};

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_513_152 u_ca_513_152_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_513_152 u_ca_513_152_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_513_152 u_ca_513_152_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_513_152 u_ca_513_152_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_513_152 u_ca_513_152_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_513_152 u_ca_513_152_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_513_152 u_ca_513_152_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_513_152 u_ca_513_152_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_513_152 u_ca_513_152_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_513_152 u_ca_513_152_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_513_152 u_ca_513_152_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_513_152 u_ca_513_152_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_513_152 u_ca_513_152_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_513_152 u_ca_513_152_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_513_152 u_ca_513_152_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_513_152 u_ca_513_152_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_513_152 u_ca_513_152_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_513_152 u_ca_513_152_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_513_152 u_ca_513_152_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_513_152 u_ca_513_152_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_513_152 u_ca_513_152_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_513_152 u_ca_513_152_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_513_152 u_ca_513_152_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_513_152 u_ca_513_152_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_513_152 u_ca_513_152_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_513_152 u_ca_513_152_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_513_152 u_ca_513_152_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_513_152 u_ca_513_152_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_513_152 u_ca_513_152_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_513_152 u_ca_513_152_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_513_152 u_ca_513_152_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_513_152 u_ca_513_152_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_513_152 u_ca_513_152_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_513_152 u_ca_513_152_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_513_152 u_ca_513_152_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_513_152 u_ca_513_152_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_513_152 u_ca_513_152_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_513_152 u_ca_513_152_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_513_152 u_ca_513_152_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_513_152 u_ca_513_152_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_513_152 u_ca_513_152_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_513_152 u_ca_513_152_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_513_152 u_ca_513_152_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_513_152 u_ca_513_152_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_513_152 u_ca_513_152_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_513_152 u_ca_513_152_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_513_152 u_ca_513_152_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_513_152 u_ca_513_152_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_513_152 u_ca_513_152_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_513_152 u_ca_513_152_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_513_152 u_ca_513_152_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_513_152 u_ca_513_152_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_513_152 u_ca_513_152_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_513_152 u_ca_513_152_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_513_152 u_ca_513_152_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_513_152 u_ca_513_152_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_513_152 u_ca_513_152_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_513_152 u_ca_513_152_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_513_152 u_ca_513_152_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_513_152 u_ca_513_152_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_513_152 u_ca_513_152_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_513_152 u_ca_513_152_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_513_152 u_ca_513_152_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_513_152 u_ca_513_152_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_513_152 u_ca_513_152_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_513_152 u_ca_513_152_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_513_152 u_ca_513_152_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_513_152 u_ca_513_152_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_513_152 u_ca_513_152_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_513_152 u_ca_513_152_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_513_152 u_ca_513_152_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_513_152 u_ca_513_152_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_513_152 u_ca_513_152_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_513_152 u_ca_513_152_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_513_152 u_ca_513_152_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_513_152 u_ca_513_152_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_513_152 u_ca_513_152_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_513_152 u_ca_513_152_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_513_152 u_ca_513_152_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_513_152 u_ca_513_152_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_513_152 u_ca_513_152_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_513_152 u_ca_513_152_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_513_152 u_ca_513_152_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_513_152 u_ca_513_152_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_513_152 u_ca_513_152_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_513_152 u_ca_513_152_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_513_152 u_ca_513_152_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_513_152 u_ca_513_152_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_513_152 u_ca_513_152_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_513_152 u_ca_513_152_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_513_152 u_ca_513_152_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_513_152 u_ca_513_152_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_513_152 u_ca_513_152_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_513_152 u_ca_513_152_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_513_152 u_ca_513_152_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_513_152 u_ca_513_152_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_513_152 u_ca_513_152_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_513_152 u_ca_513_152_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_513_152 u_ca_513_152_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_513_152 u_ca_513_152_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_513_152 u_ca_513_152_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_513_152 u_ca_513_152_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_513_152 u_ca_513_152_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_513_152 u_ca_513_152_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_513_152 u_ca_513_152_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_513_152 u_ca_513_152_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_513_152 u_ca_513_152_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_513_152 u_ca_513_152_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_513_152 u_ca_513_152_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_513_152 u_ca_513_152_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_513_152 u_ca_513_152_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_513_152 u_ca_513_152_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_513_152 u_ca_513_152_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_513_152 u_ca_513_152_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_513_152 u_ca_513_152_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_513_152 u_ca_513_152_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_513_152 u_ca_513_152_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_513_152 u_ca_513_152_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_513_152 u_ca_513_152_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_513_152 u_ca_513_152_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_513_152 u_ca_513_152_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_513_152 u_ca_513_152_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_513_152 u_ca_513_152_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_513_152 u_ca_513_152_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_513_152 u_ca_513_152_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_513_152 u_ca_513_152_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_513_152 u_ca_513_152_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_513_152 u_ca_513_152_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_513_152 u_ca_513_152_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_513_152 u_ca_513_152_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_513_152 u_ca_513_152_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_513_152 u_ca_513_152_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_513_152 u_ca_513_152_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_513_152 u_ca_513_152_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_513_152 u_ca_513_152_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_513_152 u_ca_513_152_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_513_152 u_ca_513_152_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_513_152 u_ca_513_152_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_513_152 u_ca_513_152_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_513_152 u_ca_513_152_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_513_152 u_ca_513_152_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_513_152 u_ca_513_152_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_513_152 u_ca_513_152_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_513_152 u_ca_513_152_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_513_152 u_ca_513_152_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_513_152 u_ca_513_152_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_513_152 u_ca_513_152_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_513_152 u_ca_513_152_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_513_152 u_ca_513_152_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_513_152 u_ca_513_152_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_513_152 u_ca_513_152_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_513_152 u_ca_513_152_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_513_152 u_ca_513_152_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_513_152 u_ca_513_152_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_513_152 u_ca_513_152_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_513_152 u_ca_513_152_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_513_152 u_ca_513_152_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_513_152 u_ca_513_152_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_513_152 u_ca_513_152_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_513_152 u_ca_513_152_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_513_152 u_ca_513_152_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_513_152 u_ca_513_152_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_513_152 u_ca_513_152_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_513_152 u_ca_513_152_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_513_152 u_ca_513_152_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_513_152 u_ca_513_152_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_513_152 u_ca_513_152_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_513_152 u_ca_513_152_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_513_152 u_ca_513_152_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_513_152 u_ca_513_152_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_513_152 u_ca_513_152_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_513_152 u_ca_513_152_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_513_152 u_ca_513_152_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_513_152 u_ca_513_152_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_513_152 u_ca_513_152_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_513_152 u_ca_513_152_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_513_152 u_ca_513_152_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_513_152 u_ca_513_152_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_513_152 u_ca_513_152_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_513_152 u_ca_513_152_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_513_152 u_ca_513_152_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_513_152 u_ca_513_152_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_513_152 u_ca_513_152_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_513_152 u_ca_513_152_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_513_152 u_ca_513_152_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_513_152 u_ca_513_152_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_513_152 u_ca_513_152_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_513_152 u_ca_513_152_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_513_152 u_ca_513_152_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_513_152 u_ca_513_152_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_513_152 u_ca_513_152_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_513_152 u_ca_513_152_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_513_152 u_ca_513_152_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_513_152 u_ca_513_152_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_513_152 u_ca_513_152_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_513_152 u_ca_513_152_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_513_152 u_ca_513_152_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_513_152 u_ca_513_152_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_513_152 u_ca_513_152_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_513_152 u_ca_513_152_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_513_152 u_ca_513_152_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_513_152 u_ca_513_152_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_513_152 u_ca_513_152_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_513_152 u_ca_513_152_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_513_152 u_ca_513_152_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_513_152 u_ca_513_152_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_513_152 u_ca_513_152_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_513_152 u_ca_513_152_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_513_152 u_ca_513_152_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_513_152 u_ca_513_152_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_513_152 u_ca_513_152_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_513_152 u_ca_513_152_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_513_152 u_ca_513_152_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_513_152 u_ca_513_152_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_513_152 u_ca_513_152_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_513_152 u_ca_513_152_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_513_152 u_ca_513_152_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_513_152 u_ca_513_152_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_513_152 u_ca_513_152_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_513_152 u_ca_513_152_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_513_152 u_ca_513_152_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_513_152 u_ca_513_152_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_513_152 u_ca_513_152_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_513_152 u_ca_513_152_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_513_152 u_ca_513_152_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_513_152 u_ca_513_152_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_513_152 u_ca_513_152_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_513_152 u_ca_513_152_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_513_152 u_ca_513_152_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_513_152 u_ca_513_152_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_513_152 u_ca_513_152_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_513_152 u_ca_513_152_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_513_152 u_ca_513_152_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_513_152 u_ca_513_152_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_513_152 u_ca_513_152_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_513_152 u_ca_513_152_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_513_152 u_ca_513_152_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_513_152 u_ca_513_152_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_513_152 u_ca_513_152_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_513_152 u_ca_513_152_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_513_152 u_ca_513_152_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_513_152 u_ca_513_152_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_513_152 u_ca_513_152_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_513_152 u_ca_513_152_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_513_152 u_ca_513_152_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_513_152 u_ca_513_152_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_513_152 u_ca_513_152_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_513_152 u_ca_513_152_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_513_152 u_ca_513_152_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_513_152 u_ca_513_152_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_513_152 u_ca_513_152_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_513_152 u_ca_513_152_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_513_152 u_ca_513_152_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_513_152 u_ca_513_152_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_513_152 u_ca_513_152_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_513_152 u_ca_513_152_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_513_152 u_ca_513_152_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_513_152 u_ca_513_152_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_513_152 u_ca_513_152_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_513_152 u_ca_513_152_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_513_152 u_ca_513_152_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_513_152 u_ca_513_152_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_513_152 u_ca_513_152_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_513_152 u_ca_513_152_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_513_152 u_ca_513_152_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_513_152 u_ca_513_152_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_513_152 u_ca_513_152_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_513_152 u_ca_513_152_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_513_152 u_ca_513_152_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_513_152 u_ca_513_152_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_513_152 u_ca_513_152_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_513_152 u_ca_513_152_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_513_152 u_ca_513_152_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_513_152 u_ca_513_152_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_513_152 u_ca_513_152_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_513_152 u_ca_513_152_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_513_152 u_ca_513_152_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_513_152 u_ca_513_152_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_513_152 u_ca_513_152_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_513_152 u_ca_513_152_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_513_152 u_ca_513_152_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_513_152 u_ca_513_152_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_513_152 u_ca_513_152_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_513_152 u_ca_513_152_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_513_152 u_ca_513_152_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_513_152 u_ca_513_152_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_513_152 u_ca_513_152_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_513_152 u_ca_513_152_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_513_152 u_ca_513_152_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_513_152 u_ca_513_152_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_513_152 u_ca_513_152_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_513_152 u_ca_513_152_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_513_152 u_ca_513_152_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_513_152 u_ca_513_152_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_513_152 u_ca_513_152_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_513_152 u_ca_513_152_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_513_152 u_ca_513_152_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_513_152 u_ca_513_152_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_513_152 u_ca_513_152_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_513_152 u_ca_513_152_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_513_152 u_ca_513_152_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_513_152 u_ca_513_152_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_513_152 u_ca_513_152_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_513_152 u_ca_513_152_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_513_152 u_ca_513_152_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_513_152 u_ca_513_152_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_513_152 u_ca_513_152_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_513_152 u_ca_513_152_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_513_152 u_ca_513_152_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_513_152 u_ca_513_152_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_513_152 u_ca_513_152_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_513_152 u_ca_513_152_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_513_152 u_ca_513_152_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_513_152 u_ca_513_152_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_513_152 u_ca_513_152_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_513_152 u_ca_513_152_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_513_152 u_ca_513_152_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_513_152 u_ca_513_152_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_513_152 u_ca_513_152_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_513_152 u_ca_513_152_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_513_152 u_ca_513_152_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_513_152 u_ca_513_152_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_513_152 u_ca_513_152_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_513_152 u_ca_513_152_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_513_152 u_ca_513_152_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_513_152 u_ca_513_152_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_513_152 u_ca_513_152_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_513_152 u_ca_513_152_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_513_152 u_ca_513_152_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_513_152 u_ca_513_152_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_513_152 u_ca_513_152_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_513_152 u_ca_513_152_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_513_152 u_ca_513_152_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_513_152 u_ca_513_152_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_513_152 u_ca_513_152_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_513_152 u_ca_513_152_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_513_152 u_ca_513_152_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_513_152 u_ca_513_152_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_513_152 u_ca_513_152_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_513_152 u_ca_513_152_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_513_152 u_ca_513_152_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_513_152 u_ca_513_152_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_513_152 u_ca_513_152_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_513_152 u_ca_513_152_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_513_152 u_ca_513_152_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_513_152 u_ca_513_152_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_513_152 u_ca_513_152_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_513_152 u_ca_513_152_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_513_152 u_ca_513_152_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_513_152 u_ca_513_152_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_513_152 u_ca_513_152_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_513_152 u_ca_513_152_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_513_152 u_ca_513_152_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_513_152 u_ca_513_152_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_513_152 u_ca_513_152_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_513_152 u_ca_513_152_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_513_152 u_ca_513_152_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_513_152 u_ca_513_152_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_513_152 u_ca_513_152_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_513_152 u_ca_513_152_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_513_152 u_ca_513_152_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_513_152 u_ca_513_152_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_513_152 u_ca_513_152_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_513_152 u_ca_513_152_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_513_152 u_ca_513_152_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_513_152 u_ca_513_152_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_513_152 u_ca_513_152_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_513_152 u_ca_513_152_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_513_152 u_ca_513_152_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_513_152 u_ca_513_152_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_513_152 u_ca_513_152_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_513_152 u_ca_513_152_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_513_152 u_ca_513_152_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_513_152 u_ca_513_152_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_513_152 u_ca_513_152_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_513_152 u_ca_513_152_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_513_152 u_ca_513_152_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_513_152 u_ca_513_152_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_513_152 u_ca_513_152_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_513_152 u_ca_513_152_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_513_152 u_ca_513_152_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_513_152 u_ca_513_152_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_513_152 u_ca_513_152_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_513_152 u_ca_513_152_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_513_152 u_ca_513_152_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_513_152 u_ca_513_152_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_513_152 u_ca_513_152_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_513_152 u_ca_513_152_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_513_152 u_ca_513_152_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_513_152 u_ca_513_152_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_513_152 u_ca_513_152_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_513_152 u_ca_513_152_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_513_152 u_ca_513_152_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_513_152 u_ca_513_152_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_513_152 u_ca_513_152_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_513_152 u_ca_513_152_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_513_152 u_ca_513_152_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_513_152 u_ca_513_152_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_513_152 u_ca_513_152_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_513_152 u_ca_513_152_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_513_152 u_ca_513_152_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_513_152 u_ca_513_152_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_513_152 u_ca_513_152_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_513_152 u_ca_513_152_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_513_152 u_ca_513_152_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_513_152 u_ca_513_152_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_513_152 u_ca_513_152_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_513_152 u_ca_513_152_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_513_152 u_ca_513_152_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_513_152 u_ca_513_152_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_513_152 u_ca_513_152_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_513_152 u_ca_513_152_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_513_152 u_ca_513_152_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_513_152 u_ca_513_152_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_513_152 u_ca_513_152_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_513_152 u_ca_513_152_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_513_152 u_ca_513_152_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_513_152 u_ca_513_152_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_513_152 u_ca_513_152_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_513_152 u_ca_513_152_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_513_152 u_ca_513_152_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_513_152 u_ca_513_152_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_513_152 u_ca_513_152_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_513_152 u_ca_513_152_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_513_152 u_ca_513_152_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_513_152 u_ca_513_152_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_513_152 u_ca_513_152_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_513_152 u_ca_513_152_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_513_152 u_ca_513_152_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_513_152 u_ca_513_152_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_513_152 u_ca_513_152_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_513_152 u_ca_513_152_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_513_152 u_ca_513_152_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_513_152 u_ca_513_152_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_513_152 u_ca_513_152_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_513_152 u_ca_513_152_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_513_152 u_ca_513_152_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_513_152 u_ca_513_152_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_513_152 u_ca_513_152_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_513_152 u_ca_513_152_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_513_152 u_ca_513_152_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_513_152 u_ca_513_152_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_513_152 u_ca_513_152_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_513_152 u_ca_513_152_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_513_152 u_ca_513_152_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_513_152 u_ca_513_152_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_513_152 u_ca_513_152_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_513_152 u_ca_513_152_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_513_152 u_ca_513_152_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_513_152 u_ca_513_152_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_513_152 u_ca_513_152_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_513_152 u_ca_513_152_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_513_152 u_ca_513_152_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_513_152 u_ca_513_152_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_513_152 u_ca_513_152_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_513_152 u_ca_513_152_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_513_152 u_ca_513_152_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_513_152 u_ca_513_152_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_513_152 u_ca_513_152_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_513_152 u_ca_513_152_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_513_152 u_ca_513_152_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_513_152 u_ca_513_152_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_513_152 u_ca_513_152_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_513_152 u_ca_513_152_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_513_152 u_ca_513_152_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_513_152 u_ca_513_152_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_513_152 u_ca_513_152_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_513_152 u_ca_513_152_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_513_152 u_ca_513_152_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_513_152 u_ca_513_152_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_513_152 u_ca_513_152_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_513_152 u_ca_513_152_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_513_152 u_ca_513_152_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_513_152 u_ca_513_152_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_513_152 u_ca_513_152_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_513_152 u_ca_513_152_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_513_152 u_ca_513_152_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_513_152 u_ca_513_152_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_513_152 u_ca_513_152_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_513_152 u_ca_513_152_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_513_152 u_ca_513_152_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_513_152 u_ca_513_152_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_513_152 u_ca_513_152_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_513_152 u_ca_513_152_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_513_152 u_ca_513_152_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_513_152 u_ca_513_152_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_513_152 u_ca_513_152_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_513_152 u_ca_513_152_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_513_152 u_ca_513_152_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_513_152 u_ca_513_152_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_513_152 u_ca_513_152_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_513_152 u_ca_513_152_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_513_152 u_ca_513_152_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_513_152 u_ca_513_152_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_513_152 u_ca_513_152_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_513_152 u_ca_513_152_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_513_152 u_ca_513_152_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_513_152 u_ca_513_152_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_513_152 u_ca_513_152_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_513_152 u_ca_513_152_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_513_152 u_ca_513_152_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_513_152 u_ca_513_152_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_513_152 u_ca_513_152_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_513_152 u_ca_513_152_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_513_152 u_ca_513_152_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_513_152 u_ca_513_152_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_513_152 u_ca_513_152_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_513_152 u_ca_513_152_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_513_152 u_ca_513_152_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_513_152 u_ca_513_152_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_513_152 u_ca_513_152_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_513_152 u_ca_513_152_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_513_152 u_ca_513_152_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_513_152 u_ca_513_152_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_513_152 u_ca_513_152_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_513_152 u_ca_513_152_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_513_152 u_ca_513_152_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_513_152 u_ca_513_152_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_513_152 u_ca_513_152_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_513_152 u_ca_513_152_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_513_152 u_ca_513_152_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_513_152 u_ca_513_152_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_513_152 u_ca_513_152_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_513_152 u_ca_513_152_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_513_152 u_ca_513_152_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_513_152 u_ca_513_152_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_513_152 u_ca_513_152_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_513_152 u_ca_513_152_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_513_152 u_ca_513_152_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_513_152 u_ca_513_152_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_513_152 u_ca_513_152_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_513_152 u_ca_513_152_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_513_152 u_ca_513_152_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_513_152 u_ca_513_152_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_513_152 u_ca_513_152_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_513_152 u_ca_513_152_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_513_152 u_ca_513_152_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_513_152 u_ca_513_152_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_513_152 u_ca_513_152_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_513_152 u_ca_513_152_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_513_152 u_ca_513_152_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_513_152 u_ca_513_152_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_513_152 u_ca_513_152_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_513_152 u_ca_513_152_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_513_152 u_ca_513_152_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_513_152 u_ca_513_152_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_513_152 u_ca_513_152_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_513_152 u_ca_513_152_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_513_152 u_ca_513_152_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_513_152 u_ca_513_152_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_513_152 u_ca_513_152_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_513_152 u_ca_513_152_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_513_152 u_ca_513_152_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_513_152 u_ca_513_152_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_513_152 u_ca_513_152_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_513_152 u_ca_513_152_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_513_152 u_ca_513_152_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_513_152 u_ca_513_152_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_513_152 u_ca_513_152_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_513_152 u_ca_513_152_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_513_152 u_ca_513_152_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_513_152 u_ca_513_152_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_513_152 u_ca_513_152_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_513_152 u_ca_513_152_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_513_152 u_ca_513_152_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_513_152 u_ca_513_152_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_513_152 u_ca_513_152_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_513_152 u_ca_513_152_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_513_152 u_ca_513_152_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_513_152 u_ca_513_152_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_513_152 u_ca_513_152_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_513_152 u_ca_513_152_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_513_152 u_ca_513_152_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_513_152 u_ca_513_152_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_513_152 u_ca_513_152_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_513_152 u_ca_513_152_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_513_152 u_ca_513_152_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_513_152 u_ca_513_152_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_513_152 u_ca_513_152_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_513_152 u_ca_513_152_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_513_152 u_ca_513_152_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_513_152 u_ca_513_152_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_513_152 u_ca_513_152_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_513_152 u_ca_513_152_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_513_152 u_ca_513_152_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_513_152 u_ca_513_152_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_513_152 u_ca_513_152_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_513_152 u_ca_513_152_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_513_152 u_ca_513_152_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_513_152 u_ca_513_152_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_513_152 u_ca_513_152_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_513_152 u_ca_513_152_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_513_152 u_ca_513_152_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_513_152 u_ca_513_152_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_513_152 u_ca_513_152_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_513_152 u_ca_513_152_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_513_152 u_ca_513_152_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_513_152 u_ca_513_152_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_513_152 u_ca_513_152_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_513_152 u_ca_513_152_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_513_152 u_ca_513_152_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_513_152 u_ca_513_152_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_513_152 u_ca_513_152_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_513_152 u_ca_513_152_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_513_152 u_ca_513_152_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_513_152 u_ca_513_152_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_513_152 u_ca_513_152_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_513_152 u_ca_513_152_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_513_152 u_ca_513_152_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_513_152 u_ca_513_152_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_513_152 u_ca_513_152_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_513_152 u_ca_513_152_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_513_152 u_ca_513_152_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_513_152 u_ca_513_152_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_513_152 u_ca_513_152_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_513_152 u_ca_513_152_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_513_152 u_ca_513_152_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_513_152 u_ca_513_152_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_513_152 u_ca_513_152_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_513_152 u_ca_513_152_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_513_152 u_ca_513_152_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_513_152 u_ca_513_152_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_513_152 u_ca_513_152_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_513_152 u_ca_513_152_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_513_152 u_ca_513_152_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_513_152 u_ca_513_152_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_513_152 u_ca_513_152_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_513_152 u_ca_513_152_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_513_152 u_ca_513_152_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_513_152 u_ca_513_152_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_513_152 u_ca_513_152_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_513_152 u_ca_513_152_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_513_152 u_ca_513_152_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_513_152 u_ca_513_152_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_513_152 u_ca_513_152_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_513_152 u_ca_513_152_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_513_152 u_ca_513_152_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_513_152 u_ca_513_152_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_513_152 u_ca_513_152_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_513_152 u_ca_513_152_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_513_152 u_ca_513_152_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_513_152 u_ca_513_152_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_513_152 u_ca_513_152_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_513_152 u_ca_513_152_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_513_152 u_ca_513_152_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_513_152 u_ca_513_152_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_513_152 u_ca_513_152_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_513_152 u_ca_513_152_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_513_152 u_ca_513_152_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_513_152 u_ca_513_152_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_513_152 u_ca_513_152_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_513_152 u_ca_513_152_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_513_152 u_ca_513_152_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_513_152 u_ca_513_152_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_513_152 u_ca_513_152_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_513_152 u_ca_513_152_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_513_152 u_ca_513_152_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_513_152 u_ca_513_152_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_513_152 u_ca_513_152_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_513_152 u_ca_513_152_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_513_152 u_ca_513_152_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_513_152 u_ca_513_152_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_513_152 u_ca_513_152_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_513_152 u_ca_513_152_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_513_152 u_ca_513_152_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_513_152 u_ca_513_152_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_513_152 u_ca_513_152_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_513_152 u_ca_513_152_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_513_152 u_ca_513_152_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_513_152 u_ca_513_152_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_513_152 u_ca_513_152_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_513_152 u_ca_513_152_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_513_152 u_ca_513_152_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_513_152 u_ca_513_152_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_513_152 u_ca_513_152_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_513_152 u_ca_513_152_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_513_152 u_ca_513_152_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_513_152 u_ca_513_152_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_513_152 u_ca_513_152_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_513_152 u_ca_513_152_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_513_152 u_ca_513_152_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_513_152 u_ca_513_152_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_513_152 u_ca_513_152_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_513_152 u_ca_513_152_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_513_152 u_ca_513_152_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_513_152 u_ca_513_152_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_513_152 u_ca_513_152_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_513_152 u_ca_513_152_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_513_152 u_ca_513_152_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_513_152 u_ca_513_152_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_513_152 u_ca_513_152_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_513_152 u_ca_513_152_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_513_152 u_ca_513_152_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_513_152 u_ca_513_152_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_513_152 u_ca_513_152_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_513_152 u_ca_513_152_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_513_152 u_ca_513_152_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_513_152 u_ca_513_152_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_513_152 u_ca_513_152_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_513_152 u_ca_513_152_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_513_152 u_ca_513_152_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_513_152 u_ca_513_152_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_513_152 u_ca_513_152_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_513_152 u_ca_513_152_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_513_152 u_ca_513_152_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_513_152 u_ca_513_152_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_513_152 u_ca_513_152_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_513_152 u_ca_513_152_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_513_152 u_ca_513_152_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_513_152 u_ca_513_152_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_513_152 u_ca_513_152_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_513_152 u_ca_513_152_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_513_152 u_ca_513_152_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_513_152 u_ca_513_152_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_513_152 u_ca_513_152_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_513_152 u_ca_513_152_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_513_152 u_ca_513_152_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_513_152 u_ca_513_152_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_513_152 u_ca_513_152_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_513_152 u_ca_513_152_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_513_152 u_ca_513_152_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_513_152 u_ca_513_152_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_513_152 u_ca_513_152_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_513_152 u_ca_513_152_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_513_152 u_ca_513_152_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_513_152 u_ca_513_152_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_513_152 u_ca_513_152_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_513_152 u_ca_513_152_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_513_152 u_ca_513_152_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_513_152 u_ca_513_152_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_513_152 u_ca_513_152_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_513_152 u_ca_513_152_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_513_152 u_ca_513_152_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_513_152 u_ca_513_152_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_513_152 u_ca_513_152_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_513_152 u_ca_513_152_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_513_152 u_ca_513_152_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_513_152 u_ca_513_152_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_513_152 u_ca_513_152_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_513_152 u_ca_513_152_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_513_152 u_ca_513_152_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_513_152 u_ca_513_152_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_513_152 u_ca_513_152_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_513_152 u_ca_513_152_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_513_152 u_ca_513_152_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_513_152 u_ca_513_152_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_513_152 u_ca_513_152_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_513_152 u_ca_513_152_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_513_152 u_ca_513_152_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_513_152 u_ca_513_152_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_513_152 u_ca_513_152_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_513_152 u_ca_513_152_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_513_152 u_ca_513_152_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_513_152 u_ca_513_152_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_513_152 u_ca_513_152_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_513_152 u_ca_513_152_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_513_152 u_ca_513_152_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_513_152 u_ca_513_152_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_513_152 u_ca_513_152_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_513_152 u_ca_513_152_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_513_152 u_ca_513_152_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_513_152 u_ca_513_152_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_513_152 u_ca_513_152_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_513_152 u_ca_513_152_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_513_152 u_ca_513_152_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_513_152 u_ca_513_152_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_513_152 u_ca_513_152_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_513_152 u_ca_513_152_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_513_152 u_ca_513_152_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_513_152 u_ca_513_152_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_513_152 u_ca_513_152_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_513_152 u_ca_513_152_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_513_152 u_ca_513_152_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_513_152 u_ca_513_152_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_513_152 u_ca_513_152_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_513_152 u_ca_513_152_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_513_152 u_ca_513_152_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_513_152 u_ca_513_152_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_513_152 u_ca_513_152_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_513_152 u_ca_513_152_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_513_152 u_ca_513_152_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_513_152 u_ca_513_152_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_513_152 u_ca_513_152_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_513_152 u_ca_513_152_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_513_152 u_ca_513_152_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_513_152 u_ca_513_152_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_513_152 u_ca_513_152_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_513_152 u_ca_513_152_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_513_152 u_ca_513_152_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_513_152 u_ca_513_152_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_513_152 u_ca_513_152_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_513_152 u_ca_513_152_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_513_152 u_ca_513_152_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_513_152 u_ca_513_152_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_513_152 u_ca_513_152_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_513_152 u_ca_513_152_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_513_152 u_ca_513_152_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_513_152 u_ca_513_152_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_513_152 u_ca_513_152_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_513_152 u_ca_513_152_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_513_152 u_ca_513_152_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_513_152 u_ca_513_152_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_513_152 u_ca_513_152_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_513_152 u_ca_513_152_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_513_152 u_ca_513_152_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_513_152 u_ca_513_152_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_513_152 u_ca_513_152_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_513_152 u_ca_513_152_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_513_152 u_ca_513_152_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_513_152 u_ca_513_152_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_513_152 u_ca_513_152_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_513_152 u_ca_513_152_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_513_152 u_ca_513_152_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_513_152 u_ca_513_152_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_513_152 u_ca_513_152_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_513_152 u_ca_513_152_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_513_152 u_ca_513_152_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_513_152 u_ca_513_152_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_513_152 u_ca_513_152_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_513_152 u_ca_513_152_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_513_152 u_ca_513_152_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_513_152 u_ca_513_152_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_513_152 u_ca_513_152_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_513_152 u_ca_513_152_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_513_152 u_ca_513_152_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_513_152 u_ca_513_152_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_513_152 u_ca_513_152_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_513_152 u_ca_513_152_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_513_152 u_ca_513_152_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_513_152 u_ca_513_152_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_513_152 u_ca_513_152_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_513_152 u_ca_513_152_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_513_152 u_ca_513_152_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_513_152 u_ca_513_152_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_513_152 u_ca_513_152_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_513_152 u_ca_513_152_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_513_152 u_ca_513_152_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_513_152 u_ca_513_152_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_513_152 u_ca_513_152_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_513_152 u_ca_513_152_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_513_152 u_ca_513_152_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_513_152 u_ca_513_152_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_513_152 u_ca_513_152_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_513_152 u_ca_513_152_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_513_152 u_ca_513_152_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_513_152 u_ca_513_152_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_513_152 u_ca_513_152_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_513_152 u_ca_513_152_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_513_152 u_ca_513_152_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_513_152 u_ca_513_152_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_513_152 u_ca_513_152_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_513_152 u_ca_513_152_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_513_152 u_ca_513_152_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_513_152 u_ca_513_152_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_513_152 u_ca_513_152_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_513_152 u_ca_513_152_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_513_152 u_ca_513_152_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_513_152 u_ca_513_152_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_513_152 u_ca_513_152_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_513_152 u_ca_513_152_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_513_152 u_ca_513_152_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_513_152 u_ca_513_152_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_513_152 u_ca_513_152_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_513_152 u_ca_513_152_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_513_152 u_ca_513_152_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_513_152 u_ca_513_152_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_513_152 u_ca_513_152_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_513_152 u_ca_513_152_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_513_152 u_ca_513_152_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_513_152 u_ca_513_152_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_513_152 u_ca_513_152_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_513_152 u_ca_513_152_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_513_152 u_ca_513_152_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_513_152 u_ca_513_152_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_513_152 u_ca_513_152_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_513_152 u_ca_513_152_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_513_152 u_ca_513_152_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_513_152 u_ca_513_152_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_513_152 u_ca_513_152_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_513_152 u_ca_513_152_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_513_152 u_ca_513_152_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_513_152 u_ca_513_152_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_513_152 u_ca_513_152_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_513_152 u_ca_513_152_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_513_152 u_ca_513_152_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_513_152 u_ca_513_152_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_513_152 u_ca_513_152_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_513_152 u_ca_513_152_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_513_152 u_ca_513_152_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_513_152 u_ca_513_152_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_513_152 u_ca_513_152_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_513_152 u_ca_513_152_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_513_152 u_ca_513_152_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_513_152 u_ca_513_152_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_513_152 u_ca_513_152_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_513_152 u_ca_513_152_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_513_152 u_ca_513_152_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_513_152 u_ca_513_152_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_513_152 u_ca_513_152_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_513_152 u_ca_513_152_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_513_152 u_ca_513_152_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_513_152 u_ca_513_152_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_513_152 u_ca_513_152_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_513_152 u_ca_513_152_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_513_152 u_ca_513_152_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_513_152 u_ca_513_152_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_513_152 u_ca_513_152_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_513_152 u_ca_513_152_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_513_152 u_ca_513_152_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_513_152 u_ca_513_152_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_513_152 u_ca_513_152_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_513_152 u_ca_513_152_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_513_152 u_ca_513_152_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_513_152 u_ca_513_152_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_513_152 u_ca_513_152_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_513_152 u_ca_513_152_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_513_152 u_ca_513_152_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_513_152 u_ca_513_152_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_513_152 u_ca_513_152_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_513_152 u_ca_513_152_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_513_152 u_ca_513_152_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_513_152 u_ca_513_152_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_513_152 u_ca_513_152_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_513_152 u_ca_513_152_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_513_152 u_ca_513_152_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_513_152 u_ca_513_152_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_513_152 u_ca_513_152_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_513_152 u_ca_513_152_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_513_152 u_ca_513_152_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_513_152 u_ca_513_152_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_513_152 u_ca_513_152_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_513_152 u_ca_513_152_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_513_152 u_ca_513_152_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_513_152 u_ca_513_152_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_513_152 u_ca_513_152_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_513_152 u_ca_513_152_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_513_152 u_ca_513_152_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_513_152 u_ca_513_152_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_513_152 u_ca_513_152_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_513_152 u_ca_513_152_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_513_152 u_ca_513_152_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_513_152 u_ca_513_152_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_513_152 u_ca_513_152_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_513_152 u_ca_513_152_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_513_152 u_ca_513_152_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_513_152 u_ca_513_152_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_513_152 u_ca_513_152_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_513_152 u_ca_513_152_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_513_152 u_ca_513_152_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_513_152 u_ca_513_152_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_513_152 u_ca_513_152_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_513_152 u_ca_513_152_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_513_152 u_ca_513_152_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_513_152 u_ca_513_152_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_513_152 u_ca_513_152_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_513_152 u_ca_513_152_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_513_152 u_ca_513_152_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_513_152 u_ca_513_152_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_513_152 u_ca_513_152_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_513_152 u_ca_513_152_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_513_152 u_ca_513_152_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_513_152 u_ca_513_152_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_513_152 u_ca_513_152_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_513_152 u_ca_513_152_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_513_152 u_ca_513_152_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_513_152 u_ca_513_152_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_513_152 u_ca_513_152_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_513_152 u_ca_513_152_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_513_152 u_ca_513_152_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_513_152 u_ca_513_152_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_513_152 u_ca_513_152_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_513_152 u_ca_513_152_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_513_152 u_ca_513_152_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_513_152 u_ca_513_152_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_513_152 u_ca_513_152_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_513_152 u_ca_513_152_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_513_152 u_ca_513_152_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_513_152 u_ca_513_152_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_513_152 u_ca_513_152_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_513_152 u_ca_513_152_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_513_152 u_ca_513_152_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_513_152 u_ca_513_152_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_513_152 u_ca_513_152_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_513_152 u_ca_513_152_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_513_152 u_ca_513_152_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_513_152 u_ca_513_152_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_513_152 u_ca_513_152_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_513_152 u_ca_513_152_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_513_152 u_ca_513_152_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_513_152 u_ca_513_152_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_513_152 u_ca_513_152_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_513_152 u_ca_513_152_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_513_152 u_ca_513_152_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_513_152 u_ca_513_152_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_513_152 u_ca_513_152_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_513_152 u_ca_513_152_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_513_152 u_ca_513_152_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_513_152 u_ca_513_152_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_513_152 u_ca_513_152_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_513_152 u_ca_513_152_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_513_152 u_ca_513_152_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_513_152 u_ca_513_152_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_513_152 u_ca_513_152_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_513_152 u_ca_513_152_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_513_152 u_ca_513_152_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_513_152 u_ca_513_152_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_513_152 u_ca_513_152_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_513_152 u_ca_513_152_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_513_152 u_ca_513_152_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_513_152 u_ca_513_152_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_513_152 u_ca_513_152_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_513_152 u_ca_513_152_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_513_152 u_ca_513_152_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_513_152 u_ca_513_152_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_513_152 u_ca_513_152_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_513_152 u_ca_513_152_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_513_152 u_ca_513_152_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_513_152 u_ca_513_152_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_513_152 u_ca_513_152_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_513_152 u_ca_513_152_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_513_152 u_ca_513_152_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_513_152 u_ca_513_152_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_513_152 u_ca_513_152_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_513_152 u_ca_513_152_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{133{1'b0}}, u_ca_out_0[18:0]};
assign col_out_1 = {{76{1'b0}}, u_ca_out_1[18:0], u_ca_out_0[75:19]};
assign col_out_2 = {{19{1'b0}}, u_ca_out_2[18:0], u_ca_out_1[75:19], u_ca_out_0[132:76]};
assign col_out_3 = {u_ca_out_3[18:0],u_ca_out_2[75:19], u_ca_out_1[132:76], u_ca_out_0[151:133]};
assign col_out_4 = {u_ca_out_4[18:0],u_ca_out_3[75:19], u_ca_out_2[132:76], u_ca_out_1[151:133]};
assign col_out_5 = {u_ca_out_5[18:0],u_ca_out_4[75:19], u_ca_out_3[132:76], u_ca_out_2[151:133]};
assign col_out_6 = {u_ca_out_6[18:0],u_ca_out_5[75:19], u_ca_out_4[132:76], u_ca_out_3[151:133]};
assign col_out_7 = {u_ca_out_7[18:0],u_ca_out_6[75:19], u_ca_out_5[132:76], u_ca_out_4[151:133]};
assign col_out_8 = {u_ca_out_8[18:0],u_ca_out_7[75:19], u_ca_out_6[132:76], u_ca_out_5[151:133]};
assign col_out_9 = {u_ca_out_9[18:0],u_ca_out_8[75:19], u_ca_out_7[132:76], u_ca_out_6[151:133]};
assign col_out_10 = {u_ca_out_10[18:0],u_ca_out_9[75:19], u_ca_out_8[132:76], u_ca_out_7[151:133]};
assign col_out_11 = {u_ca_out_11[18:0],u_ca_out_10[75:19], u_ca_out_9[132:76], u_ca_out_8[151:133]};
assign col_out_12 = {u_ca_out_12[18:0],u_ca_out_11[75:19], u_ca_out_10[132:76], u_ca_out_9[151:133]};
assign col_out_13 = {u_ca_out_13[18:0],u_ca_out_12[75:19], u_ca_out_11[132:76], u_ca_out_10[151:133]};
assign col_out_14 = {u_ca_out_14[18:0],u_ca_out_13[75:19], u_ca_out_12[132:76], u_ca_out_11[151:133]};
assign col_out_15 = {u_ca_out_15[18:0],u_ca_out_14[75:19], u_ca_out_13[132:76], u_ca_out_12[151:133]};
assign col_out_16 = {u_ca_out_16[18:0],u_ca_out_15[75:19], u_ca_out_14[132:76], u_ca_out_13[151:133]};
assign col_out_17 = {u_ca_out_17[18:0],u_ca_out_16[75:19], u_ca_out_15[132:76], u_ca_out_14[151:133]};
assign col_out_18 = {u_ca_out_18[18:0],u_ca_out_17[75:19], u_ca_out_16[132:76], u_ca_out_15[151:133]};
assign col_out_19 = {u_ca_out_19[18:0],u_ca_out_18[75:19], u_ca_out_17[132:76], u_ca_out_16[151:133]};
assign col_out_20 = {u_ca_out_20[18:0],u_ca_out_19[75:19], u_ca_out_18[132:76], u_ca_out_17[151:133]};
assign col_out_21 = {u_ca_out_21[18:0],u_ca_out_20[75:19], u_ca_out_19[132:76], u_ca_out_18[151:133]};
assign col_out_22 = {u_ca_out_22[18:0],u_ca_out_21[75:19], u_ca_out_20[132:76], u_ca_out_19[151:133]};
assign col_out_23 = {u_ca_out_23[18:0],u_ca_out_22[75:19], u_ca_out_21[132:76], u_ca_out_20[151:133]};
assign col_out_24 = {u_ca_out_24[18:0],u_ca_out_23[75:19], u_ca_out_22[132:76], u_ca_out_21[151:133]};
assign col_out_25 = {u_ca_out_25[18:0],u_ca_out_24[75:19], u_ca_out_23[132:76], u_ca_out_22[151:133]};
assign col_out_26 = {u_ca_out_26[18:0],u_ca_out_25[75:19], u_ca_out_24[132:76], u_ca_out_23[151:133]};
assign col_out_27 = {u_ca_out_27[18:0],u_ca_out_26[75:19], u_ca_out_25[132:76], u_ca_out_24[151:133]};
assign col_out_28 = {u_ca_out_28[18:0],u_ca_out_27[75:19], u_ca_out_26[132:76], u_ca_out_25[151:133]};
assign col_out_29 = {u_ca_out_29[18:0],u_ca_out_28[75:19], u_ca_out_27[132:76], u_ca_out_26[151:133]};
assign col_out_30 = {u_ca_out_30[18:0],u_ca_out_29[75:19], u_ca_out_28[132:76], u_ca_out_27[151:133]};
assign col_out_31 = {u_ca_out_31[18:0],u_ca_out_30[75:19], u_ca_out_29[132:76], u_ca_out_28[151:133]};
assign col_out_32 = {u_ca_out_32[18:0],u_ca_out_31[75:19], u_ca_out_30[132:76], u_ca_out_29[151:133]};
assign col_out_33 = {u_ca_out_33[18:0],u_ca_out_32[75:19], u_ca_out_31[132:76], u_ca_out_30[151:133]};
assign col_out_34 = {u_ca_out_34[18:0],u_ca_out_33[75:19], u_ca_out_32[132:76], u_ca_out_31[151:133]};
assign col_out_35 = {u_ca_out_35[18:0],u_ca_out_34[75:19], u_ca_out_33[132:76], u_ca_out_32[151:133]};
assign col_out_36 = {u_ca_out_36[18:0],u_ca_out_35[75:19], u_ca_out_34[132:76], u_ca_out_33[151:133]};
assign col_out_37 = {u_ca_out_37[18:0],u_ca_out_36[75:19], u_ca_out_35[132:76], u_ca_out_34[151:133]};
assign col_out_38 = {u_ca_out_38[18:0],u_ca_out_37[75:19], u_ca_out_36[132:76], u_ca_out_35[151:133]};
assign col_out_39 = {u_ca_out_39[18:0],u_ca_out_38[75:19], u_ca_out_37[132:76], u_ca_out_36[151:133]};
assign col_out_40 = {u_ca_out_40[18:0],u_ca_out_39[75:19], u_ca_out_38[132:76], u_ca_out_37[151:133]};
assign col_out_41 = {u_ca_out_41[18:0],u_ca_out_40[75:19], u_ca_out_39[132:76], u_ca_out_38[151:133]};
assign col_out_42 = {u_ca_out_42[18:0],u_ca_out_41[75:19], u_ca_out_40[132:76], u_ca_out_39[151:133]};
assign col_out_43 = {u_ca_out_43[18:0],u_ca_out_42[75:19], u_ca_out_41[132:76], u_ca_out_40[151:133]};
assign col_out_44 = {u_ca_out_44[18:0],u_ca_out_43[75:19], u_ca_out_42[132:76], u_ca_out_41[151:133]};
assign col_out_45 = {u_ca_out_45[18:0],u_ca_out_44[75:19], u_ca_out_43[132:76], u_ca_out_42[151:133]};
assign col_out_46 = {u_ca_out_46[18:0],u_ca_out_45[75:19], u_ca_out_44[132:76], u_ca_out_43[151:133]};
assign col_out_47 = {u_ca_out_47[18:0],u_ca_out_46[75:19], u_ca_out_45[132:76], u_ca_out_44[151:133]};
assign col_out_48 = {u_ca_out_48[18:0],u_ca_out_47[75:19], u_ca_out_46[132:76], u_ca_out_45[151:133]};
assign col_out_49 = {u_ca_out_49[18:0],u_ca_out_48[75:19], u_ca_out_47[132:76], u_ca_out_46[151:133]};
assign col_out_50 = {u_ca_out_50[18:0],u_ca_out_49[75:19], u_ca_out_48[132:76], u_ca_out_47[151:133]};
assign col_out_51 = {u_ca_out_51[18:0],u_ca_out_50[75:19], u_ca_out_49[132:76], u_ca_out_48[151:133]};
assign col_out_52 = {u_ca_out_52[18:0],u_ca_out_51[75:19], u_ca_out_50[132:76], u_ca_out_49[151:133]};
assign col_out_53 = {u_ca_out_53[18:0],u_ca_out_52[75:19], u_ca_out_51[132:76], u_ca_out_50[151:133]};
assign col_out_54 = {u_ca_out_54[18:0],u_ca_out_53[75:19], u_ca_out_52[132:76], u_ca_out_51[151:133]};
assign col_out_55 = {u_ca_out_55[18:0],u_ca_out_54[75:19], u_ca_out_53[132:76], u_ca_out_52[151:133]};
assign col_out_56 = {u_ca_out_56[18:0],u_ca_out_55[75:19], u_ca_out_54[132:76], u_ca_out_53[151:133]};
assign col_out_57 = {u_ca_out_57[18:0],u_ca_out_56[75:19], u_ca_out_55[132:76], u_ca_out_54[151:133]};
assign col_out_58 = {u_ca_out_58[18:0],u_ca_out_57[75:19], u_ca_out_56[132:76], u_ca_out_55[151:133]};
assign col_out_59 = {u_ca_out_59[18:0],u_ca_out_58[75:19], u_ca_out_57[132:76], u_ca_out_56[151:133]};
assign col_out_60 = {u_ca_out_60[18:0],u_ca_out_59[75:19], u_ca_out_58[132:76], u_ca_out_57[151:133]};
assign col_out_61 = {u_ca_out_61[18:0],u_ca_out_60[75:19], u_ca_out_59[132:76], u_ca_out_58[151:133]};
assign col_out_62 = {u_ca_out_62[18:0],u_ca_out_61[75:19], u_ca_out_60[132:76], u_ca_out_59[151:133]};
assign col_out_63 = {u_ca_out_63[18:0],u_ca_out_62[75:19], u_ca_out_61[132:76], u_ca_out_60[151:133]};
assign col_out_64 = {u_ca_out_64[18:0],u_ca_out_63[75:19], u_ca_out_62[132:76], u_ca_out_61[151:133]};
assign col_out_65 = {u_ca_out_65[18:0],u_ca_out_64[75:19], u_ca_out_63[132:76], u_ca_out_62[151:133]};
assign col_out_66 = {u_ca_out_66[18:0],u_ca_out_65[75:19], u_ca_out_64[132:76], u_ca_out_63[151:133]};
assign col_out_67 = {u_ca_out_67[18:0],u_ca_out_66[75:19], u_ca_out_65[132:76], u_ca_out_64[151:133]};
assign col_out_68 = {u_ca_out_68[18:0],u_ca_out_67[75:19], u_ca_out_66[132:76], u_ca_out_65[151:133]};
assign col_out_69 = {u_ca_out_69[18:0],u_ca_out_68[75:19], u_ca_out_67[132:76], u_ca_out_66[151:133]};
assign col_out_70 = {u_ca_out_70[18:0],u_ca_out_69[75:19], u_ca_out_68[132:76], u_ca_out_67[151:133]};
assign col_out_71 = {u_ca_out_71[18:0],u_ca_out_70[75:19], u_ca_out_69[132:76], u_ca_out_68[151:133]};
assign col_out_72 = {u_ca_out_72[18:0],u_ca_out_71[75:19], u_ca_out_70[132:76], u_ca_out_69[151:133]};
assign col_out_73 = {u_ca_out_73[18:0],u_ca_out_72[75:19], u_ca_out_71[132:76], u_ca_out_70[151:133]};
assign col_out_74 = {u_ca_out_74[18:0],u_ca_out_73[75:19], u_ca_out_72[132:76], u_ca_out_71[151:133]};
assign col_out_75 = {u_ca_out_75[18:0],u_ca_out_74[75:19], u_ca_out_73[132:76], u_ca_out_72[151:133]};
assign col_out_76 = {u_ca_out_76[18:0],u_ca_out_75[75:19], u_ca_out_74[132:76], u_ca_out_73[151:133]};
assign col_out_77 = {u_ca_out_77[18:0],u_ca_out_76[75:19], u_ca_out_75[132:76], u_ca_out_74[151:133]};
assign col_out_78 = {u_ca_out_78[18:0],u_ca_out_77[75:19], u_ca_out_76[132:76], u_ca_out_75[151:133]};
assign col_out_79 = {u_ca_out_79[18:0],u_ca_out_78[75:19], u_ca_out_77[132:76], u_ca_out_76[151:133]};
assign col_out_80 = {u_ca_out_80[18:0],u_ca_out_79[75:19], u_ca_out_78[132:76], u_ca_out_77[151:133]};
assign col_out_81 = {u_ca_out_81[18:0],u_ca_out_80[75:19], u_ca_out_79[132:76], u_ca_out_78[151:133]};
assign col_out_82 = {u_ca_out_82[18:0],u_ca_out_81[75:19], u_ca_out_80[132:76], u_ca_out_79[151:133]};
assign col_out_83 = {u_ca_out_83[18:0],u_ca_out_82[75:19], u_ca_out_81[132:76], u_ca_out_80[151:133]};
assign col_out_84 = {u_ca_out_84[18:0],u_ca_out_83[75:19], u_ca_out_82[132:76], u_ca_out_81[151:133]};
assign col_out_85 = {u_ca_out_85[18:0],u_ca_out_84[75:19], u_ca_out_83[132:76], u_ca_out_82[151:133]};
assign col_out_86 = {u_ca_out_86[18:0],u_ca_out_85[75:19], u_ca_out_84[132:76], u_ca_out_83[151:133]};
assign col_out_87 = {u_ca_out_87[18:0],u_ca_out_86[75:19], u_ca_out_85[132:76], u_ca_out_84[151:133]};
assign col_out_88 = {u_ca_out_88[18:0],u_ca_out_87[75:19], u_ca_out_86[132:76], u_ca_out_85[151:133]};
assign col_out_89 = {u_ca_out_89[18:0],u_ca_out_88[75:19], u_ca_out_87[132:76], u_ca_out_86[151:133]};
assign col_out_90 = {u_ca_out_90[18:0],u_ca_out_89[75:19], u_ca_out_88[132:76], u_ca_out_87[151:133]};
assign col_out_91 = {u_ca_out_91[18:0],u_ca_out_90[75:19], u_ca_out_89[132:76], u_ca_out_88[151:133]};
assign col_out_92 = {u_ca_out_92[18:0],u_ca_out_91[75:19], u_ca_out_90[132:76], u_ca_out_89[151:133]};
assign col_out_93 = {u_ca_out_93[18:0],u_ca_out_92[75:19], u_ca_out_91[132:76], u_ca_out_90[151:133]};
assign col_out_94 = {u_ca_out_94[18:0],u_ca_out_93[75:19], u_ca_out_92[132:76], u_ca_out_91[151:133]};
assign col_out_95 = {u_ca_out_95[18:0],u_ca_out_94[75:19], u_ca_out_93[132:76], u_ca_out_92[151:133]};
assign col_out_96 = {u_ca_out_96[18:0],u_ca_out_95[75:19], u_ca_out_94[132:76], u_ca_out_93[151:133]};
assign col_out_97 = {u_ca_out_97[18:0],u_ca_out_96[75:19], u_ca_out_95[132:76], u_ca_out_94[151:133]};
assign col_out_98 = {u_ca_out_98[18:0],u_ca_out_97[75:19], u_ca_out_96[132:76], u_ca_out_95[151:133]};
assign col_out_99 = {u_ca_out_99[18:0],u_ca_out_98[75:19], u_ca_out_97[132:76], u_ca_out_96[151:133]};
assign col_out_100 = {u_ca_out_100[18:0],u_ca_out_99[75:19], u_ca_out_98[132:76], u_ca_out_97[151:133]};
assign col_out_101 = {u_ca_out_101[18:0],u_ca_out_100[75:19], u_ca_out_99[132:76], u_ca_out_98[151:133]};
assign col_out_102 = {u_ca_out_102[18:0],u_ca_out_101[75:19], u_ca_out_100[132:76], u_ca_out_99[151:133]};
assign col_out_103 = {u_ca_out_103[18:0],u_ca_out_102[75:19], u_ca_out_101[132:76], u_ca_out_100[151:133]};
assign col_out_104 = {u_ca_out_104[18:0],u_ca_out_103[75:19], u_ca_out_102[132:76], u_ca_out_101[151:133]};
assign col_out_105 = {u_ca_out_105[18:0],u_ca_out_104[75:19], u_ca_out_103[132:76], u_ca_out_102[151:133]};
assign col_out_106 = {u_ca_out_106[18:0],u_ca_out_105[75:19], u_ca_out_104[132:76], u_ca_out_103[151:133]};
assign col_out_107 = {u_ca_out_107[18:0],u_ca_out_106[75:19], u_ca_out_105[132:76], u_ca_out_104[151:133]};
assign col_out_108 = {u_ca_out_108[18:0],u_ca_out_107[75:19], u_ca_out_106[132:76], u_ca_out_105[151:133]};
assign col_out_109 = {u_ca_out_109[18:0],u_ca_out_108[75:19], u_ca_out_107[132:76], u_ca_out_106[151:133]};
assign col_out_110 = {u_ca_out_110[18:0],u_ca_out_109[75:19], u_ca_out_108[132:76], u_ca_out_107[151:133]};
assign col_out_111 = {u_ca_out_111[18:0],u_ca_out_110[75:19], u_ca_out_109[132:76], u_ca_out_108[151:133]};
assign col_out_112 = {u_ca_out_112[18:0],u_ca_out_111[75:19], u_ca_out_110[132:76], u_ca_out_109[151:133]};
assign col_out_113 = {u_ca_out_113[18:0],u_ca_out_112[75:19], u_ca_out_111[132:76], u_ca_out_110[151:133]};
assign col_out_114 = {u_ca_out_114[18:0],u_ca_out_113[75:19], u_ca_out_112[132:76], u_ca_out_111[151:133]};
assign col_out_115 = {u_ca_out_115[18:0],u_ca_out_114[75:19], u_ca_out_113[132:76], u_ca_out_112[151:133]};
assign col_out_116 = {u_ca_out_116[18:0],u_ca_out_115[75:19], u_ca_out_114[132:76], u_ca_out_113[151:133]};
assign col_out_117 = {u_ca_out_117[18:0],u_ca_out_116[75:19], u_ca_out_115[132:76], u_ca_out_114[151:133]};
assign col_out_118 = {u_ca_out_118[18:0],u_ca_out_117[75:19], u_ca_out_116[132:76], u_ca_out_115[151:133]};
assign col_out_119 = {u_ca_out_119[18:0],u_ca_out_118[75:19], u_ca_out_117[132:76], u_ca_out_116[151:133]};
assign col_out_120 = {u_ca_out_120[18:0],u_ca_out_119[75:19], u_ca_out_118[132:76], u_ca_out_117[151:133]};
assign col_out_121 = {u_ca_out_121[18:0],u_ca_out_120[75:19], u_ca_out_119[132:76], u_ca_out_118[151:133]};
assign col_out_122 = {u_ca_out_122[18:0],u_ca_out_121[75:19], u_ca_out_120[132:76], u_ca_out_119[151:133]};
assign col_out_123 = {u_ca_out_123[18:0],u_ca_out_122[75:19], u_ca_out_121[132:76], u_ca_out_120[151:133]};
assign col_out_124 = {u_ca_out_124[18:0],u_ca_out_123[75:19], u_ca_out_122[132:76], u_ca_out_121[151:133]};
assign col_out_125 = {u_ca_out_125[18:0],u_ca_out_124[75:19], u_ca_out_123[132:76], u_ca_out_122[151:133]};
assign col_out_126 = {u_ca_out_126[18:0],u_ca_out_125[75:19], u_ca_out_124[132:76], u_ca_out_123[151:133]};
assign col_out_127 = {u_ca_out_127[18:0],u_ca_out_126[75:19], u_ca_out_125[132:76], u_ca_out_124[151:133]};
assign col_out_128 = {u_ca_out_128[18:0],u_ca_out_127[75:19], u_ca_out_126[132:76], u_ca_out_125[151:133]};
assign col_out_129 = {u_ca_out_129[18:0],u_ca_out_128[75:19], u_ca_out_127[132:76], u_ca_out_126[151:133]};
assign col_out_130 = {u_ca_out_130[18:0],u_ca_out_129[75:19], u_ca_out_128[132:76], u_ca_out_127[151:133]};
assign col_out_131 = {u_ca_out_131[18:0],u_ca_out_130[75:19], u_ca_out_129[132:76], u_ca_out_128[151:133]};
assign col_out_132 = {u_ca_out_132[18:0],u_ca_out_131[75:19], u_ca_out_130[132:76], u_ca_out_129[151:133]};
assign col_out_133 = {u_ca_out_133[18:0],u_ca_out_132[75:19], u_ca_out_131[132:76], u_ca_out_130[151:133]};
assign col_out_134 = {u_ca_out_134[18:0],u_ca_out_133[75:19], u_ca_out_132[132:76], u_ca_out_131[151:133]};
assign col_out_135 = {u_ca_out_135[18:0],u_ca_out_134[75:19], u_ca_out_133[132:76], u_ca_out_132[151:133]};
assign col_out_136 = {u_ca_out_136[18:0],u_ca_out_135[75:19], u_ca_out_134[132:76], u_ca_out_133[151:133]};
assign col_out_137 = {u_ca_out_137[18:0],u_ca_out_136[75:19], u_ca_out_135[132:76], u_ca_out_134[151:133]};
assign col_out_138 = {u_ca_out_138[18:0],u_ca_out_137[75:19], u_ca_out_136[132:76], u_ca_out_135[151:133]};
assign col_out_139 = {u_ca_out_139[18:0],u_ca_out_138[75:19], u_ca_out_137[132:76], u_ca_out_136[151:133]};
assign col_out_140 = {u_ca_out_140[18:0],u_ca_out_139[75:19], u_ca_out_138[132:76], u_ca_out_137[151:133]};
assign col_out_141 = {u_ca_out_141[18:0],u_ca_out_140[75:19], u_ca_out_139[132:76], u_ca_out_138[151:133]};
assign col_out_142 = {u_ca_out_142[18:0],u_ca_out_141[75:19], u_ca_out_140[132:76], u_ca_out_139[151:133]};
assign col_out_143 = {u_ca_out_143[18:0],u_ca_out_142[75:19], u_ca_out_141[132:76], u_ca_out_140[151:133]};
assign col_out_144 = {u_ca_out_144[18:0],u_ca_out_143[75:19], u_ca_out_142[132:76], u_ca_out_141[151:133]};
assign col_out_145 = {u_ca_out_145[18:0],u_ca_out_144[75:19], u_ca_out_143[132:76], u_ca_out_142[151:133]};
assign col_out_146 = {u_ca_out_146[18:0],u_ca_out_145[75:19], u_ca_out_144[132:76], u_ca_out_143[151:133]};
assign col_out_147 = {u_ca_out_147[18:0],u_ca_out_146[75:19], u_ca_out_145[132:76], u_ca_out_144[151:133]};
assign col_out_148 = {u_ca_out_148[18:0],u_ca_out_147[75:19], u_ca_out_146[132:76], u_ca_out_145[151:133]};
assign col_out_149 = {u_ca_out_149[18:0],u_ca_out_148[75:19], u_ca_out_147[132:76], u_ca_out_146[151:133]};
assign col_out_150 = {u_ca_out_150[18:0],u_ca_out_149[75:19], u_ca_out_148[132:76], u_ca_out_147[151:133]};
assign col_out_151 = {u_ca_out_151[18:0],u_ca_out_150[75:19], u_ca_out_149[132:76], u_ca_out_148[151:133]};
assign col_out_152 = {u_ca_out_152[18:0],u_ca_out_151[75:19], u_ca_out_150[132:76], u_ca_out_149[151:133]};
assign col_out_153 = {u_ca_out_153[18:0],u_ca_out_152[75:19], u_ca_out_151[132:76], u_ca_out_150[151:133]};
assign col_out_154 = {u_ca_out_154[18:0],u_ca_out_153[75:19], u_ca_out_152[132:76], u_ca_out_151[151:133]};
assign col_out_155 = {u_ca_out_155[18:0],u_ca_out_154[75:19], u_ca_out_153[132:76], u_ca_out_152[151:133]};
assign col_out_156 = {u_ca_out_156[18:0],u_ca_out_155[75:19], u_ca_out_154[132:76], u_ca_out_153[151:133]};
assign col_out_157 = {u_ca_out_157[18:0],u_ca_out_156[75:19], u_ca_out_155[132:76], u_ca_out_154[151:133]};
assign col_out_158 = {u_ca_out_158[18:0],u_ca_out_157[75:19], u_ca_out_156[132:76], u_ca_out_155[151:133]};
assign col_out_159 = {u_ca_out_159[18:0],u_ca_out_158[75:19], u_ca_out_157[132:76], u_ca_out_156[151:133]};
assign col_out_160 = {u_ca_out_160[18:0],u_ca_out_159[75:19], u_ca_out_158[132:76], u_ca_out_157[151:133]};
assign col_out_161 = {u_ca_out_161[18:0],u_ca_out_160[75:19], u_ca_out_159[132:76], u_ca_out_158[151:133]};
assign col_out_162 = {u_ca_out_162[18:0],u_ca_out_161[75:19], u_ca_out_160[132:76], u_ca_out_159[151:133]};
assign col_out_163 = {u_ca_out_163[18:0],u_ca_out_162[75:19], u_ca_out_161[132:76], u_ca_out_160[151:133]};
assign col_out_164 = {u_ca_out_164[18:0],u_ca_out_163[75:19], u_ca_out_162[132:76], u_ca_out_161[151:133]};
assign col_out_165 = {u_ca_out_165[18:0],u_ca_out_164[75:19], u_ca_out_163[132:76], u_ca_out_162[151:133]};
assign col_out_166 = {u_ca_out_166[18:0],u_ca_out_165[75:19], u_ca_out_164[132:76], u_ca_out_163[151:133]};
assign col_out_167 = {u_ca_out_167[18:0],u_ca_out_166[75:19], u_ca_out_165[132:76], u_ca_out_164[151:133]};
assign col_out_168 = {u_ca_out_168[18:0],u_ca_out_167[75:19], u_ca_out_166[132:76], u_ca_out_165[151:133]};
assign col_out_169 = {u_ca_out_169[18:0],u_ca_out_168[75:19], u_ca_out_167[132:76], u_ca_out_166[151:133]};
assign col_out_170 = {u_ca_out_170[18:0],u_ca_out_169[75:19], u_ca_out_168[132:76], u_ca_out_167[151:133]};
assign col_out_171 = {u_ca_out_171[18:0],u_ca_out_170[75:19], u_ca_out_169[132:76], u_ca_out_168[151:133]};
assign col_out_172 = {u_ca_out_172[18:0],u_ca_out_171[75:19], u_ca_out_170[132:76], u_ca_out_169[151:133]};
assign col_out_173 = {u_ca_out_173[18:0],u_ca_out_172[75:19], u_ca_out_171[132:76], u_ca_out_170[151:133]};
assign col_out_174 = {u_ca_out_174[18:0],u_ca_out_173[75:19], u_ca_out_172[132:76], u_ca_out_171[151:133]};
assign col_out_175 = {u_ca_out_175[18:0],u_ca_out_174[75:19], u_ca_out_173[132:76], u_ca_out_172[151:133]};
assign col_out_176 = {u_ca_out_176[18:0],u_ca_out_175[75:19], u_ca_out_174[132:76], u_ca_out_173[151:133]};
assign col_out_177 = {u_ca_out_177[18:0],u_ca_out_176[75:19], u_ca_out_175[132:76], u_ca_out_174[151:133]};
assign col_out_178 = {u_ca_out_178[18:0],u_ca_out_177[75:19], u_ca_out_176[132:76], u_ca_out_175[151:133]};
assign col_out_179 = {u_ca_out_179[18:0],u_ca_out_178[75:19], u_ca_out_177[132:76], u_ca_out_176[151:133]};
assign col_out_180 = {u_ca_out_180[18:0],u_ca_out_179[75:19], u_ca_out_178[132:76], u_ca_out_177[151:133]};
assign col_out_181 = {u_ca_out_181[18:0],u_ca_out_180[75:19], u_ca_out_179[132:76], u_ca_out_178[151:133]};
assign col_out_182 = {u_ca_out_182[18:0],u_ca_out_181[75:19], u_ca_out_180[132:76], u_ca_out_179[151:133]};
assign col_out_183 = {u_ca_out_183[18:0],u_ca_out_182[75:19], u_ca_out_181[132:76], u_ca_out_180[151:133]};
assign col_out_184 = {u_ca_out_184[18:0],u_ca_out_183[75:19], u_ca_out_182[132:76], u_ca_out_181[151:133]};
assign col_out_185 = {u_ca_out_185[18:0],u_ca_out_184[75:19], u_ca_out_183[132:76], u_ca_out_182[151:133]};
assign col_out_186 = {u_ca_out_186[18:0],u_ca_out_185[75:19], u_ca_out_184[132:76], u_ca_out_183[151:133]};
assign col_out_187 = {u_ca_out_187[18:0],u_ca_out_186[75:19], u_ca_out_185[132:76], u_ca_out_184[151:133]};
assign col_out_188 = {u_ca_out_188[18:0],u_ca_out_187[75:19], u_ca_out_186[132:76], u_ca_out_185[151:133]};
assign col_out_189 = {u_ca_out_189[18:0],u_ca_out_188[75:19], u_ca_out_187[132:76], u_ca_out_186[151:133]};
assign col_out_190 = {u_ca_out_190[18:0],u_ca_out_189[75:19], u_ca_out_188[132:76], u_ca_out_187[151:133]};
assign col_out_191 = {u_ca_out_191[18:0],u_ca_out_190[75:19], u_ca_out_189[132:76], u_ca_out_188[151:133]};
assign col_out_192 = {u_ca_out_192[18:0],u_ca_out_191[75:19], u_ca_out_190[132:76], u_ca_out_189[151:133]};
assign col_out_193 = {u_ca_out_193[18:0],u_ca_out_192[75:19], u_ca_out_191[132:76], u_ca_out_190[151:133]};
assign col_out_194 = {u_ca_out_194[18:0],u_ca_out_193[75:19], u_ca_out_192[132:76], u_ca_out_191[151:133]};
assign col_out_195 = {u_ca_out_195[18:0],u_ca_out_194[75:19], u_ca_out_193[132:76], u_ca_out_192[151:133]};
assign col_out_196 = {u_ca_out_196[18:0],u_ca_out_195[75:19], u_ca_out_194[132:76], u_ca_out_193[151:133]};
assign col_out_197 = {u_ca_out_197[18:0],u_ca_out_196[75:19], u_ca_out_195[132:76], u_ca_out_194[151:133]};
assign col_out_198 = {u_ca_out_198[18:0],u_ca_out_197[75:19], u_ca_out_196[132:76], u_ca_out_195[151:133]};
assign col_out_199 = {u_ca_out_199[18:0],u_ca_out_198[75:19], u_ca_out_197[132:76], u_ca_out_196[151:133]};
assign col_out_200 = {u_ca_out_200[18:0],u_ca_out_199[75:19], u_ca_out_198[132:76], u_ca_out_197[151:133]};
assign col_out_201 = {u_ca_out_201[18:0],u_ca_out_200[75:19], u_ca_out_199[132:76], u_ca_out_198[151:133]};
assign col_out_202 = {u_ca_out_202[18:0],u_ca_out_201[75:19], u_ca_out_200[132:76], u_ca_out_199[151:133]};
assign col_out_203 = {u_ca_out_203[18:0],u_ca_out_202[75:19], u_ca_out_201[132:76], u_ca_out_200[151:133]};
assign col_out_204 = {u_ca_out_204[18:0],u_ca_out_203[75:19], u_ca_out_202[132:76], u_ca_out_201[151:133]};
assign col_out_205 = {u_ca_out_205[18:0],u_ca_out_204[75:19], u_ca_out_203[132:76], u_ca_out_202[151:133]};
assign col_out_206 = {u_ca_out_206[18:0],u_ca_out_205[75:19], u_ca_out_204[132:76], u_ca_out_203[151:133]};
assign col_out_207 = {u_ca_out_207[18:0],u_ca_out_206[75:19], u_ca_out_205[132:76], u_ca_out_204[151:133]};
assign col_out_208 = {u_ca_out_208[18:0],u_ca_out_207[75:19], u_ca_out_206[132:76], u_ca_out_205[151:133]};
assign col_out_209 = {u_ca_out_209[18:0],u_ca_out_208[75:19], u_ca_out_207[132:76], u_ca_out_206[151:133]};
assign col_out_210 = {u_ca_out_210[18:0],u_ca_out_209[75:19], u_ca_out_208[132:76], u_ca_out_207[151:133]};
assign col_out_211 = {u_ca_out_211[18:0],u_ca_out_210[75:19], u_ca_out_209[132:76], u_ca_out_208[151:133]};
assign col_out_212 = {u_ca_out_212[18:0],u_ca_out_211[75:19], u_ca_out_210[132:76], u_ca_out_209[151:133]};
assign col_out_213 = {u_ca_out_213[18:0],u_ca_out_212[75:19], u_ca_out_211[132:76], u_ca_out_210[151:133]};
assign col_out_214 = {u_ca_out_214[18:0],u_ca_out_213[75:19], u_ca_out_212[132:76], u_ca_out_211[151:133]};
assign col_out_215 = {u_ca_out_215[18:0],u_ca_out_214[75:19], u_ca_out_213[132:76], u_ca_out_212[151:133]};
assign col_out_216 = {u_ca_out_216[18:0],u_ca_out_215[75:19], u_ca_out_214[132:76], u_ca_out_213[151:133]};
assign col_out_217 = {u_ca_out_217[18:0],u_ca_out_216[75:19], u_ca_out_215[132:76], u_ca_out_214[151:133]};
assign col_out_218 = {u_ca_out_218[18:0],u_ca_out_217[75:19], u_ca_out_216[132:76], u_ca_out_215[151:133]};
assign col_out_219 = {u_ca_out_219[18:0],u_ca_out_218[75:19], u_ca_out_217[132:76], u_ca_out_216[151:133]};
assign col_out_220 = {u_ca_out_220[18:0],u_ca_out_219[75:19], u_ca_out_218[132:76], u_ca_out_217[151:133]};
assign col_out_221 = {u_ca_out_221[18:0],u_ca_out_220[75:19], u_ca_out_219[132:76], u_ca_out_218[151:133]};
assign col_out_222 = {u_ca_out_222[18:0],u_ca_out_221[75:19], u_ca_out_220[132:76], u_ca_out_219[151:133]};
assign col_out_223 = {u_ca_out_223[18:0],u_ca_out_222[75:19], u_ca_out_221[132:76], u_ca_out_220[151:133]};
assign col_out_224 = {u_ca_out_224[18:0],u_ca_out_223[75:19], u_ca_out_222[132:76], u_ca_out_221[151:133]};
assign col_out_225 = {u_ca_out_225[18:0],u_ca_out_224[75:19], u_ca_out_223[132:76], u_ca_out_222[151:133]};
assign col_out_226 = {u_ca_out_226[18:0],u_ca_out_225[75:19], u_ca_out_224[132:76], u_ca_out_223[151:133]};
assign col_out_227 = {u_ca_out_227[18:0],u_ca_out_226[75:19], u_ca_out_225[132:76], u_ca_out_224[151:133]};
assign col_out_228 = {u_ca_out_228[18:0],u_ca_out_227[75:19], u_ca_out_226[132:76], u_ca_out_225[151:133]};
assign col_out_229 = {u_ca_out_229[18:0],u_ca_out_228[75:19], u_ca_out_227[132:76], u_ca_out_226[151:133]};
assign col_out_230 = {u_ca_out_230[18:0],u_ca_out_229[75:19], u_ca_out_228[132:76], u_ca_out_227[151:133]};
assign col_out_231 = {u_ca_out_231[18:0],u_ca_out_230[75:19], u_ca_out_229[132:76], u_ca_out_228[151:133]};
assign col_out_232 = {u_ca_out_232[18:0],u_ca_out_231[75:19], u_ca_out_230[132:76], u_ca_out_229[151:133]};
assign col_out_233 = {u_ca_out_233[18:0],u_ca_out_232[75:19], u_ca_out_231[132:76], u_ca_out_230[151:133]};
assign col_out_234 = {u_ca_out_234[18:0],u_ca_out_233[75:19], u_ca_out_232[132:76], u_ca_out_231[151:133]};
assign col_out_235 = {u_ca_out_235[18:0],u_ca_out_234[75:19], u_ca_out_233[132:76], u_ca_out_232[151:133]};
assign col_out_236 = {u_ca_out_236[18:0],u_ca_out_235[75:19], u_ca_out_234[132:76], u_ca_out_233[151:133]};
assign col_out_237 = {u_ca_out_237[18:0],u_ca_out_236[75:19], u_ca_out_235[132:76], u_ca_out_234[151:133]};
assign col_out_238 = {u_ca_out_238[18:0],u_ca_out_237[75:19], u_ca_out_236[132:76], u_ca_out_235[151:133]};
assign col_out_239 = {u_ca_out_239[18:0],u_ca_out_238[75:19], u_ca_out_237[132:76], u_ca_out_236[151:133]};
assign col_out_240 = {u_ca_out_240[18:0],u_ca_out_239[75:19], u_ca_out_238[132:76], u_ca_out_237[151:133]};
assign col_out_241 = {u_ca_out_241[18:0],u_ca_out_240[75:19], u_ca_out_239[132:76], u_ca_out_238[151:133]};
assign col_out_242 = {u_ca_out_242[18:0],u_ca_out_241[75:19], u_ca_out_240[132:76], u_ca_out_239[151:133]};
assign col_out_243 = {u_ca_out_243[18:0],u_ca_out_242[75:19], u_ca_out_241[132:76], u_ca_out_240[151:133]};
assign col_out_244 = {u_ca_out_244[18:0],u_ca_out_243[75:19], u_ca_out_242[132:76], u_ca_out_241[151:133]};
assign col_out_245 = {u_ca_out_245[18:0],u_ca_out_244[75:19], u_ca_out_243[132:76], u_ca_out_242[151:133]};
assign col_out_246 = {u_ca_out_246[18:0],u_ca_out_245[75:19], u_ca_out_244[132:76], u_ca_out_243[151:133]};
assign col_out_247 = {u_ca_out_247[18:0],u_ca_out_246[75:19], u_ca_out_245[132:76], u_ca_out_244[151:133]};
assign col_out_248 = {u_ca_out_248[18:0],u_ca_out_247[75:19], u_ca_out_246[132:76], u_ca_out_245[151:133]};
assign col_out_249 = {u_ca_out_249[18:0],u_ca_out_248[75:19], u_ca_out_247[132:76], u_ca_out_246[151:133]};
assign col_out_250 = {u_ca_out_250[18:0],u_ca_out_249[75:19], u_ca_out_248[132:76], u_ca_out_247[151:133]};
assign col_out_251 = {u_ca_out_251[18:0],u_ca_out_250[75:19], u_ca_out_249[132:76], u_ca_out_248[151:133]};
assign col_out_252 = {u_ca_out_252[18:0],u_ca_out_251[75:19], u_ca_out_250[132:76], u_ca_out_249[151:133]};
assign col_out_253 = {u_ca_out_253[18:0],u_ca_out_252[75:19], u_ca_out_251[132:76], u_ca_out_250[151:133]};
assign col_out_254 = {u_ca_out_254[18:0],u_ca_out_253[75:19], u_ca_out_252[132:76], u_ca_out_251[151:133]};
assign col_out_255 = {u_ca_out_255[18:0],u_ca_out_254[75:19], u_ca_out_253[132:76], u_ca_out_252[151:133]};
assign col_out_256 = {u_ca_out_256[18:0],u_ca_out_255[75:19], u_ca_out_254[132:76], u_ca_out_253[151:133]};
assign col_out_257 = {u_ca_out_257[18:0],u_ca_out_256[75:19], u_ca_out_255[132:76], u_ca_out_254[151:133]};
assign col_out_258 = {u_ca_out_258[18:0],u_ca_out_257[75:19], u_ca_out_256[132:76], u_ca_out_255[151:133]};
assign col_out_259 = {u_ca_out_259[18:0],u_ca_out_258[75:19], u_ca_out_257[132:76], u_ca_out_256[151:133]};
assign col_out_260 = {u_ca_out_260[18:0],u_ca_out_259[75:19], u_ca_out_258[132:76], u_ca_out_257[151:133]};
assign col_out_261 = {u_ca_out_261[18:0],u_ca_out_260[75:19], u_ca_out_259[132:76], u_ca_out_258[151:133]};
assign col_out_262 = {u_ca_out_262[18:0],u_ca_out_261[75:19], u_ca_out_260[132:76], u_ca_out_259[151:133]};
assign col_out_263 = {u_ca_out_263[18:0],u_ca_out_262[75:19], u_ca_out_261[132:76], u_ca_out_260[151:133]};
assign col_out_264 = {u_ca_out_264[18:0],u_ca_out_263[75:19], u_ca_out_262[132:76], u_ca_out_261[151:133]};
assign col_out_265 = {u_ca_out_265[18:0],u_ca_out_264[75:19], u_ca_out_263[132:76], u_ca_out_262[151:133]};
assign col_out_266 = {u_ca_out_266[18:0],u_ca_out_265[75:19], u_ca_out_264[132:76], u_ca_out_263[151:133]};
assign col_out_267 = {u_ca_out_267[18:0],u_ca_out_266[75:19], u_ca_out_265[132:76], u_ca_out_264[151:133]};
assign col_out_268 = {u_ca_out_268[18:0],u_ca_out_267[75:19], u_ca_out_266[132:76], u_ca_out_265[151:133]};
assign col_out_269 = {u_ca_out_269[18:0],u_ca_out_268[75:19], u_ca_out_267[132:76], u_ca_out_266[151:133]};
assign col_out_270 = {u_ca_out_270[18:0],u_ca_out_269[75:19], u_ca_out_268[132:76], u_ca_out_267[151:133]};
assign col_out_271 = {u_ca_out_271[18:0],u_ca_out_270[75:19], u_ca_out_269[132:76], u_ca_out_268[151:133]};
assign col_out_272 = {u_ca_out_272[18:0],u_ca_out_271[75:19], u_ca_out_270[132:76], u_ca_out_269[151:133]};
assign col_out_273 = {u_ca_out_273[18:0],u_ca_out_272[75:19], u_ca_out_271[132:76], u_ca_out_270[151:133]};
assign col_out_274 = {u_ca_out_274[18:0],u_ca_out_273[75:19], u_ca_out_272[132:76], u_ca_out_271[151:133]};
assign col_out_275 = {u_ca_out_275[18:0],u_ca_out_274[75:19], u_ca_out_273[132:76], u_ca_out_272[151:133]};
assign col_out_276 = {u_ca_out_276[18:0],u_ca_out_275[75:19], u_ca_out_274[132:76], u_ca_out_273[151:133]};
assign col_out_277 = {u_ca_out_277[18:0],u_ca_out_276[75:19], u_ca_out_275[132:76], u_ca_out_274[151:133]};
assign col_out_278 = {u_ca_out_278[18:0],u_ca_out_277[75:19], u_ca_out_276[132:76], u_ca_out_275[151:133]};
assign col_out_279 = {u_ca_out_279[18:0],u_ca_out_278[75:19], u_ca_out_277[132:76], u_ca_out_276[151:133]};
assign col_out_280 = {u_ca_out_280[18:0],u_ca_out_279[75:19], u_ca_out_278[132:76], u_ca_out_277[151:133]};
assign col_out_281 = {u_ca_out_281[18:0],u_ca_out_280[75:19], u_ca_out_279[132:76], u_ca_out_278[151:133]};
assign col_out_282 = {u_ca_out_282[18:0],u_ca_out_281[75:19], u_ca_out_280[132:76], u_ca_out_279[151:133]};
assign col_out_283 = {u_ca_out_283[18:0],u_ca_out_282[75:19], u_ca_out_281[132:76], u_ca_out_280[151:133]};
assign col_out_284 = {u_ca_out_284[18:0],u_ca_out_283[75:19], u_ca_out_282[132:76], u_ca_out_281[151:133]};
assign col_out_285 = {u_ca_out_285[18:0],u_ca_out_284[75:19], u_ca_out_283[132:76], u_ca_out_282[151:133]};
assign col_out_286 = {u_ca_out_286[18:0],u_ca_out_285[75:19], u_ca_out_284[132:76], u_ca_out_283[151:133]};
assign col_out_287 = {u_ca_out_287[18:0],u_ca_out_286[75:19], u_ca_out_285[132:76], u_ca_out_284[151:133]};
assign col_out_288 = {u_ca_out_288[18:0],u_ca_out_287[75:19], u_ca_out_286[132:76], u_ca_out_285[151:133]};
assign col_out_289 = {u_ca_out_289[18:0],u_ca_out_288[75:19], u_ca_out_287[132:76], u_ca_out_286[151:133]};
assign col_out_290 = {u_ca_out_290[18:0],u_ca_out_289[75:19], u_ca_out_288[132:76], u_ca_out_287[151:133]};
assign col_out_291 = {u_ca_out_291[18:0],u_ca_out_290[75:19], u_ca_out_289[132:76], u_ca_out_288[151:133]};
assign col_out_292 = {u_ca_out_292[18:0],u_ca_out_291[75:19], u_ca_out_290[132:76], u_ca_out_289[151:133]};
assign col_out_293 = {u_ca_out_293[18:0],u_ca_out_292[75:19], u_ca_out_291[132:76], u_ca_out_290[151:133]};
assign col_out_294 = {u_ca_out_294[18:0],u_ca_out_293[75:19], u_ca_out_292[132:76], u_ca_out_291[151:133]};
assign col_out_295 = {u_ca_out_295[18:0],u_ca_out_294[75:19], u_ca_out_293[132:76], u_ca_out_292[151:133]};
assign col_out_296 = {u_ca_out_296[18:0],u_ca_out_295[75:19], u_ca_out_294[132:76], u_ca_out_293[151:133]};
assign col_out_297 = {u_ca_out_297[18:0],u_ca_out_296[75:19], u_ca_out_295[132:76], u_ca_out_294[151:133]};
assign col_out_298 = {u_ca_out_298[18:0],u_ca_out_297[75:19], u_ca_out_296[132:76], u_ca_out_295[151:133]};
assign col_out_299 = {u_ca_out_299[18:0],u_ca_out_298[75:19], u_ca_out_297[132:76], u_ca_out_296[151:133]};
assign col_out_300 = {u_ca_out_300[18:0],u_ca_out_299[75:19], u_ca_out_298[132:76], u_ca_out_297[151:133]};
assign col_out_301 = {u_ca_out_301[18:0],u_ca_out_300[75:19], u_ca_out_299[132:76], u_ca_out_298[151:133]};
assign col_out_302 = {u_ca_out_302[18:0],u_ca_out_301[75:19], u_ca_out_300[132:76], u_ca_out_299[151:133]};
assign col_out_303 = {u_ca_out_303[18:0],u_ca_out_302[75:19], u_ca_out_301[132:76], u_ca_out_300[151:133]};
assign col_out_304 = {u_ca_out_304[18:0],u_ca_out_303[75:19], u_ca_out_302[132:76], u_ca_out_301[151:133]};
assign col_out_305 = {u_ca_out_305[18:0],u_ca_out_304[75:19], u_ca_out_303[132:76], u_ca_out_302[151:133]};
assign col_out_306 = {u_ca_out_306[18:0],u_ca_out_305[75:19], u_ca_out_304[132:76], u_ca_out_303[151:133]};
assign col_out_307 = {u_ca_out_307[18:0],u_ca_out_306[75:19], u_ca_out_305[132:76], u_ca_out_304[151:133]};
assign col_out_308 = {u_ca_out_308[18:0],u_ca_out_307[75:19], u_ca_out_306[132:76], u_ca_out_305[151:133]};
assign col_out_309 = {u_ca_out_309[18:0],u_ca_out_308[75:19], u_ca_out_307[132:76], u_ca_out_306[151:133]};
assign col_out_310 = {u_ca_out_310[18:0],u_ca_out_309[75:19], u_ca_out_308[132:76], u_ca_out_307[151:133]};
assign col_out_311 = {u_ca_out_311[18:0],u_ca_out_310[75:19], u_ca_out_309[132:76], u_ca_out_308[151:133]};
assign col_out_312 = {u_ca_out_312[18:0],u_ca_out_311[75:19], u_ca_out_310[132:76], u_ca_out_309[151:133]};
assign col_out_313 = {u_ca_out_313[18:0],u_ca_out_312[75:19], u_ca_out_311[132:76], u_ca_out_310[151:133]};
assign col_out_314 = {u_ca_out_314[18:0],u_ca_out_313[75:19], u_ca_out_312[132:76], u_ca_out_311[151:133]};
assign col_out_315 = {u_ca_out_315[18:0],u_ca_out_314[75:19], u_ca_out_313[132:76], u_ca_out_312[151:133]};
assign col_out_316 = {u_ca_out_316[18:0],u_ca_out_315[75:19], u_ca_out_314[132:76], u_ca_out_313[151:133]};
assign col_out_317 = {u_ca_out_317[18:0],u_ca_out_316[75:19], u_ca_out_315[132:76], u_ca_out_314[151:133]};
assign col_out_318 = {u_ca_out_318[18:0],u_ca_out_317[75:19], u_ca_out_316[132:76], u_ca_out_315[151:133]};
assign col_out_319 = {u_ca_out_319[18:0],u_ca_out_318[75:19], u_ca_out_317[132:76], u_ca_out_316[151:133]};
assign col_out_320 = {u_ca_out_320[18:0],u_ca_out_319[75:19], u_ca_out_318[132:76], u_ca_out_317[151:133]};
assign col_out_321 = {u_ca_out_321[18:0],u_ca_out_320[75:19], u_ca_out_319[132:76], u_ca_out_318[151:133]};
assign col_out_322 = {u_ca_out_322[18:0],u_ca_out_321[75:19], u_ca_out_320[132:76], u_ca_out_319[151:133]};
assign col_out_323 = {u_ca_out_323[18:0],u_ca_out_322[75:19], u_ca_out_321[132:76], u_ca_out_320[151:133]};
assign col_out_324 = {u_ca_out_324[18:0],u_ca_out_323[75:19], u_ca_out_322[132:76], u_ca_out_321[151:133]};
assign col_out_325 = {u_ca_out_325[18:0],u_ca_out_324[75:19], u_ca_out_323[132:76], u_ca_out_322[151:133]};
assign col_out_326 = {u_ca_out_326[18:0],u_ca_out_325[75:19], u_ca_out_324[132:76], u_ca_out_323[151:133]};
assign col_out_327 = {u_ca_out_327[18:0],u_ca_out_326[75:19], u_ca_out_325[132:76], u_ca_out_324[151:133]};
assign col_out_328 = {u_ca_out_328[18:0],u_ca_out_327[75:19], u_ca_out_326[132:76], u_ca_out_325[151:133]};
assign col_out_329 = {u_ca_out_329[18:0],u_ca_out_328[75:19], u_ca_out_327[132:76], u_ca_out_326[151:133]};
assign col_out_330 = {u_ca_out_330[18:0],u_ca_out_329[75:19], u_ca_out_328[132:76], u_ca_out_327[151:133]};
assign col_out_331 = {u_ca_out_331[18:0],u_ca_out_330[75:19], u_ca_out_329[132:76], u_ca_out_328[151:133]};
assign col_out_332 = {u_ca_out_332[18:0],u_ca_out_331[75:19], u_ca_out_330[132:76], u_ca_out_329[151:133]};
assign col_out_333 = {u_ca_out_333[18:0],u_ca_out_332[75:19], u_ca_out_331[132:76], u_ca_out_330[151:133]};
assign col_out_334 = {u_ca_out_334[18:0],u_ca_out_333[75:19], u_ca_out_332[132:76], u_ca_out_331[151:133]};
assign col_out_335 = {u_ca_out_335[18:0],u_ca_out_334[75:19], u_ca_out_333[132:76], u_ca_out_332[151:133]};
assign col_out_336 = {u_ca_out_336[18:0],u_ca_out_335[75:19], u_ca_out_334[132:76], u_ca_out_333[151:133]};
assign col_out_337 = {u_ca_out_337[18:0],u_ca_out_336[75:19], u_ca_out_335[132:76], u_ca_out_334[151:133]};
assign col_out_338 = {u_ca_out_338[18:0],u_ca_out_337[75:19], u_ca_out_336[132:76], u_ca_out_335[151:133]};
assign col_out_339 = {u_ca_out_339[18:0],u_ca_out_338[75:19], u_ca_out_337[132:76], u_ca_out_336[151:133]};
assign col_out_340 = {u_ca_out_340[18:0],u_ca_out_339[75:19], u_ca_out_338[132:76], u_ca_out_337[151:133]};
assign col_out_341 = {u_ca_out_341[18:0],u_ca_out_340[75:19], u_ca_out_339[132:76], u_ca_out_338[151:133]};
assign col_out_342 = {u_ca_out_342[18:0],u_ca_out_341[75:19], u_ca_out_340[132:76], u_ca_out_339[151:133]};
assign col_out_343 = {u_ca_out_343[18:0],u_ca_out_342[75:19], u_ca_out_341[132:76], u_ca_out_340[151:133]};
assign col_out_344 = {u_ca_out_344[18:0],u_ca_out_343[75:19], u_ca_out_342[132:76], u_ca_out_341[151:133]};
assign col_out_345 = {u_ca_out_345[18:0],u_ca_out_344[75:19], u_ca_out_343[132:76], u_ca_out_342[151:133]};
assign col_out_346 = {u_ca_out_346[18:0],u_ca_out_345[75:19], u_ca_out_344[132:76], u_ca_out_343[151:133]};
assign col_out_347 = {u_ca_out_347[18:0],u_ca_out_346[75:19], u_ca_out_345[132:76], u_ca_out_344[151:133]};
assign col_out_348 = {u_ca_out_348[18:0],u_ca_out_347[75:19], u_ca_out_346[132:76], u_ca_out_345[151:133]};
assign col_out_349 = {u_ca_out_349[18:0],u_ca_out_348[75:19], u_ca_out_347[132:76], u_ca_out_346[151:133]};
assign col_out_350 = {u_ca_out_350[18:0],u_ca_out_349[75:19], u_ca_out_348[132:76], u_ca_out_347[151:133]};
assign col_out_351 = {u_ca_out_351[18:0],u_ca_out_350[75:19], u_ca_out_349[132:76], u_ca_out_348[151:133]};
assign col_out_352 = {u_ca_out_352[18:0],u_ca_out_351[75:19], u_ca_out_350[132:76], u_ca_out_349[151:133]};
assign col_out_353 = {u_ca_out_353[18:0],u_ca_out_352[75:19], u_ca_out_351[132:76], u_ca_out_350[151:133]};
assign col_out_354 = {u_ca_out_354[18:0],u_ca_out_353[75:19], u_ca_out_352[132:76], u_ca_out_351[151:133]};
assign col_out_355 = {u_ca_out_355[18:0],u_ca_out_354[75:19], u_ca_out_353[132:76], u_ca_out_352[151:133]};
assign col_out_356 = {u_ca_out_356[18:0],u_ca_out_355[75:19], u_ca_out_354[132:76], u_ca_out_353[151:133]};
assign col_out_357 = {u_ca_out_357[18:0],u_ca_out_356[75:19], u_ca_out_355[132:76], u_ca_out_354[151:133]};
assign col_out_358 = {u_ca_out_358[18:0],u_ca_out_357[75:19], u_ca_out_356[132:76], u_ca_out_355[151:133]};
assign col_out_359 = {u_ca_out_359[18:0],u_ca_out_358[75:19], u_ca_out_357[132:76], u_ca_out_356[151:133]};
assign col_out_360 = {u_ca_out_360[18:0],u_ca_out_359[75:19], u_ca_out_358[132:76], u_ca_out_357[151:133]};
assign col_out_361 = {u_ca_out_361[18:0],u_ca_out_360[75:19], u_ca_out_359[132:76], u_ca_out_358[151:133]};
assign col_out_362 = {u_ca_out_362[18:0],u_ca_out_361[75:19], u_ca_out_360[132:76], u_ca_out_359[151:133]};
assign col_out_363 = {u_ca_out_363[18:0],u_ca_out_362[75:19], u_ca_out_361[132:76], u_ca_out_360[151:133]};
assign col_out_364 = {u_ca_out_364[18:0],u_ca_out_363[75:19], u_ca_out_362[132:76], u_ca_out_361[151:133]};
assign col_out_365 = {u_ca_out_365[18:0],u_ca_out_364[75:19], u_ca_out_363[132:76], u_ca_out_362[151:133]};
assign col_out_366 = {u_ca_out_366[18:0],u_ca_out_365[75:19], u_ca_out_364[132:76], u_ca_out_363[151:133]};
assign col_out_367 = {u_ca_out_367[18:0],u_ca_out_366[75:19], u_ca_out_365[132:76], u_ca_out_364[151:133]};
assign col_out_368 = {u_ca_out_368[18:0],u_ca_out_367[75:19], u_ca_out_366[132:76], u_ca_out_365[151:133]};
assign col_out_369 = {u_ca_out_369[18:0],u_ca_out_368[75:19], u_ca_out_367[132:76], u_ca_out_366[151:133]};
assign col_out_370 = {u_ca_out_370[18:0],u_ca_out_369[75:19], u_ca_out_368[132:76], u_ca_out_367[151:133]};
assign col_out_371 = {u_ca_out_371[18:0],u_ca_out_370[75:19], u_ca_out_369[132:76], u_ca_out_368[151:133]};
assign col_out_372 = {u_ca_out_372[18:0],u_ca_out_371[75:19], u_ca_out_370[132:76], u_ca_out_369[151:133]};
assign col_out_373 = {u_ca_out_373[18:0],u_ca_out_372[75:19], u_ca_out_371[132:76], u_ca_out_370[151:133]};
assign col_out_374 = {u_ca_out_374[18:0],u_ca_out_373[75:19], u_ca_out_372[132:76], u_ca_out_371[151:133]};
assign col_out_375 = {u_ca_out_375[18:0],u_ca_out_374[75:19], u_ca_out_373[132:76], u_ca_out_372[151:133]};
assign col_out_376 = {u_ca_out_376[18:0],u_ca_out_375[75:19], u_ca_out_374[132:76], u_ca_out_373[151:133]};
assign col_out_377 = {u_ca_out_377[18:0],u_ca_out_376[75:19], u_ca_out_375[132:76], u_ca_out_374[151:133]};
assign col_out_378 = {u_ca_out_378[18:0],u_ca_out_377[75:19], u_ca_out_376[132:76], u_ca_out_375[151:133]};
assign col_out_379 = {u_ca_out_379[18:0],u_ca_out_378[75:19], u_ca_out_377[132:76], u_ca_out_376[151:133]};
assign col_out_380 = {u_ca_out_380[18:0],u_ca_out_379[75:19], u_ca_out_378[132:76], u_ca_out_377[151:133]};
assign col_out_381 = {u_ca_out_381[18:0],u_ca_out_380[75:19], u_ca_out_379[132:76], u_ca_out_378[151:133]};
assign col_out_382 = {u_ca_out_382[18:0],u_ca_out_381[75:19], u_ca_out_380[132:76], u_ca_out_379[151:133]};
assign col_out_383 = {u_ca_out_383[18:0],u_ca_out_382[75:19], u_ca_out_381[132:76], u_ca_out_380[151:133]};
assign col_out_384 = {u_ca_out_384[18:0],u_ca_out_383[75:19], u_ca_out_382[132:76], u_ca_out_381[151:133]};
assign col_out_385 = {u_ca_out_385[18:0],u_ca_out_384[75:19], u_ca_out_383[132:76], u_ca_out_382[151:133]};
assign col_out_386 = {u_ca_out_386[18:0],u_ca_out_385[75:19], u_ca_out_384[132:76], u_ca_out_383[151:133]};
assign col_out_387 = {u_ca_out_387[18:0],u_ca_out_386[75:19], u_ca_out_385[132:76], u_ca_out_384[151:133]};
assign col_out_388 = {u_ca_out_388[18:0],u_ca_out_387[75:19], u_ca_out_386[132:76], u_ca_out_385[151:133]};
assign col_out_389 = {u_ca_out_389[18:0],u_ca_out_388[75:19], u_ca_out_387[132:76], u_ca_out_386[151:133]};
assign col_out_390 = {u_ca_out_390[18:0],u_ca_out_389[75:19], u_ca_out_388[132:76], u_ca_out_387[151:133]};
assign col_out_391 = {u_ca_out_391[18:0],u_ca_out_390[75:19], u_ca_out_389[132:76], u_ca_out_388[151:133]};
assign col_out_392 = {u_ca_out_392[18:0],u_ca_out_391[75:19], u_ca_out_390[132:76], u_ca_out_389[151:133]};
assign col_out_393 = {u_ca_out_393[18:0],u_ca_out_392[75:19], u_ca_out_391[132:76], u_ca_out_390[151:133]};
assign col_out_394 = {u_ca_out_394[18:0],u_ca_out_393[75:19], u_ca_out_392[132:76], u_ca_out_391[151:133]};
assign col_out_395 = {u_ca_out_395[18:0],u_ca_out_394[75:19], u_ca_out_393[132:76], u_ca_out_392[151:133]};
assign col_out_396 = {u_ca_out_396[18:0],u_ca_out_395[75:19], u_ca_out_394[132:76], u_ca_out_393[151:133]};
assign col_out_397 = {u_ca_out_397[18:0],u_ca_out_396[75:19], u_ca_out_395[132:76], u_ca_out_394[151:133]};
assign col_out_398 = {u_ca_out_398[18:0],u_ca_out_397[75:19], u_ca_out_396[132:76], u_ca_out_395[151:133]};
assign col_out_399 = {u_ca_out_399[18:0],u_ca_out_398[75:19], u_ca_out_397[132:76], u_ca_out_396[151:133]};
assign col_out_400 = {u_ca_out_400[18:0],u_ca_out_399[75:19], u_ca_out_398[132:76], u_ca_out_397[151:133]};
assign col_out_401 = {u_ca_out_401[18:0],u_ca_out_400[75:19], u_ca_out_399[132:76], u_ca_out_398[151:133]};
assign col_out_402 = {u_ca_out_402[18:0],u_ca_out_401[75:19], u_ca_out_400[132:76], u_ca_out_399[151:133]};
assign col_out_403 = {u_ca_out_403[18:0],u_ca_out_402[75:19], u_ca_out_401[132:76], u_ca_out_400[151:133]};
assign col_out_404 = {u_ca_out_404[18:0],u_ca_out_403[75:19], u_ca_out_402[132:76], u_ca_out_401[151:133]};
assign col_out_405 = {u_ca_out_405[18:0],u_ca_out_404[75:19], u_ca_out_403[132:76], u_ca_out_402[151:133]};
assign col_out_406 = {u_ca_out_406[18:0],u_ca_out_405[75:19], u_ca_out_404[132:76], u_ca_out_403[151:133]};
assign col_out_407 = {u_ca_out_407[18:0],u_ca_out_406[75:19], u_ca_out_405[132:76], u_ca_out_404[151:133]};
assign col_out_408 = {u_ca_out_408[18:0],u_ca_out_407[75:19], u_ca_out_406[132:76], u_ca_out_405[151:133]};
assign col_out_409 = {u_ca_out_409[18:0],u_ca_out_408[75:19], u_ca_out_407[132:76], u_ca_out_406[151:133]};
assign col_out_410 = {u_ca_out_410[18:0],u_ca_out_409[75:19], u_ca_out_408[132:76], u_ca_out_407[151:133]};
assign col_out_411 = {u_ca_out_411[18:0],u_ca_out_410[75:19], u_ca_out_409[132:76], u_ca_out_408[151:133]};
assign col_out_412 = {u_ca_out_412[18:0],u_ca_out_411[75:19], u_ca_out_410[132:76], u_ca_out_409[151:133]};
assign col_out_413 = {u_ca_out_413[18:0],u_ca_out_412[75:19], u_ca_out_411[132:76], u_ca_out_410[151:133]};
assign col_out_414 = {u_ca_out_414[18:0],u_ca_out_413[75:19], u_ca_out_412[132:76], u_ca_out_411[151:133]};
assign col_out_415 = {u_ca_out_415[18:0],u_ca_out_414[75:19], u_ca_out_413[132:76], u_ca_out_412[151:133]};
assign col_out_416 = {u_ca_out_416[18:0],u_ca_out_415[75:19], u_ca_out_414[132:76], u_ca_out_413[151:133]};
assign col_out_417 = {u_ca_out_417[18:0],u_ca_out_416[75:19], u_ca_out_415[132:76], u_ca_out_414[151:133]};
assign col_out_418 = {u_ca_out_418[18:0],u_ca_out_417[75:19], u_ca_out_416[132:76], u_ca_out_415[151:133]};
assign col_out_419 = {u_ca_out_419[18:0],u_ca_out_418[75:19], u_ca_out_417[132:76], u_ca_out_416[151:133]};
assign col_out_420 = {u_ca_out_420[18:0],u_ca_out_419[75:19], u_ca_out_418[132:76], u_ca_out_417[151:133]};
assign col_out_421 = {u_ca_out_421[18:0],u_ca_out_420[75:19], u_ca_out_419[132:76], u_ca_out_418[151:133]};
assign col_out_422 = {u_ca_out_422[18:0],u_ca_out_421[75:19], u_ca_out_420[132:76], u_ca_out_419[151:133]};
assign col_out_423 = {u_ca_out_423[18:0],u_ca_out_422[75:19], u_ca_out_421[132:76], u_ca_out_420[151:133]};
assign col_out_424 = {u_ca_out_424[18:0],u_ca_out_423[75:19], u_ca_out_422[132:76], u_ca_out_421[151:133]};
assign col_out_425 = {u_ca_out_425[18:0],u_ca_out_424[75:19], u_ca_out_423[132:76], u_ca_out_422[151:133]};
assign col_out_426 = {u_ca_out_426[18:0],u_ca_out_425[75:19], u_ca_out_424[132:76], u_ca_out_423[151:133]};
assign col_out_427 = {u_ca_out_427[18:0],u_ca_out_426[75:19], u_ca_out_425[132:76], u_ca_out_424[151:133]};
assign col_out_428 = {u_ca_out_428[18:0],u_ca_out_427[75:19], u_ca_out_426[132:76], u_ca_out_425[151:133]};
assign col_out_429 = {u_ca_out_429[18:0],u_ca_out_428[75:19], u_ca_out_427[132:76], u_ca_out_426[151:133]};
assign col_out_430 = {u_ca_out_430[18:0],u_ca_out_429[75:19], u_ca_out_428[132:76], u_ca_out_427[151:133]};
assign col_out_431 = {u_ca_out_431[18:0],u_ca_out_430[75:19], u_ca_out_429[132:76], u_ca_out_428[151:133]};
assign col_out_432 = {u_ca_out_432[18:0],u_ca_out_431[75:19], u_ca_out_430[132:76], u_ca_out_429[151:133]};
assign col_out_433 = {u_ca_out_433[18:0],u_ca_out_432[75:19], u_ca_out_431[132:76], u_ca_out_430[151:133]};
assign col_out_434 = {u_ca_out_434[18:0],u_ca_out_433[75:19], u_ca_out_432[132:76], u_ca_out_431[151:133]};
assign col_out_435 = {u_ca_out_435[18:0],u_ca_out_434[75:19], u_ca_out_433[132:76], u_ca_out_432[151:133]};
assign col_out_436 = {u_ca_out_436[18:0],u_ca_out_435[75:19], u_ca_out_434[132:76], u_ca_out_433[151:133]};
assign col_out_437 = {u_ca_out_437[18:0],u_ca_out_436[75:19], u_ca_out_435[132:76], u_ca_out_434[151:133]};
assign col_out_438 = {u_ca_out_438[18:0],u_ca_out_437[75:19], u_ca_out_436[132:76], u_ca_out_435[151:133]};
assign col_out_439 = {u_ca_out_439[18:0],u_ca_out_438[75:19], u_ca_out_437[132:76], u_ca_out_436[151:133]};
assign col_out_440 = {u_ca_out_440[18:0],u_ca_out_439[75:19], u_ca_out_438[132:76], u_ca_out_437[151:133]};
assign col_out_441 = {u_ca_out_441[18:0],u_ca_out_440[75:19], u_ca_out_439[132:76], u_ca_out_438[151:133]};
assign col_out_442 = {u_ca_out_442[18:0],u_ca_out_441[75:19], u_ca_out_440[132:76], u_ca_out_439[151:133]};
assign col_out_443 = {u_ca_out_443[18:0],u_ca_out_442[75:19], u_ca_out_441[132:76], u_ca_out_440[151:133]};
assign col_out_444 = {u_ca_out_444[18:0],u_ca_out_443[75:19], u_ca_out_442[132:76], u_ca_out_441[151:133]};
assign col_out_445 = {u_ca_out_445[18:0],u_ca_out_444[75:19], u_ca_out_443[132:76], u_ca_out_442[151:133]};
assign col_out_446 = {u_ca_out_446[18:0],u_ca_out_445[75:19], u_ca_out_444[132:76], u_ca_out_443[151:133]};
assign col_out_447 = {u_ca_out_447[18:0],u_ca_out_446[75:19], u_ca_out_445[132:76], u_ca_out_444[151:133]};
assign col_out_448 = {u_ca_out_448[18:0],u_ca_out_447[75:19], u_ca_out_446[132:76], u_ca_out_445[151:133]};
assign col_out_449 = {u_ca_out_449[18:0],u_ca_out_448[75:19], u_ca_out_447[132:76], u_ca_out_446[151:133]};
assign col_out_450 = {u_ca_out_450[18:0],u_ca_out_449[75:19], u_ca_out_448[132:76], u_ca_out_447[151:133]};
assign col_out_451 = {u_ca_out_451[18:0],u_ca_out_450[75:19], u_ca_out_449[132:76], u_ca_out_448[151:133]};
assign col_out_452 = {u_ca_out_452[18:0],u_ca_out_451[75:19], u_ca_out_450[132:76], u_ca_out_449[151:133]};
assign col_out_453 = {u_ca_out_453[18:0],u_ca_out_452[75:19], u_ca_out_451[132:76], u_ca_out_450[151:133]};
assign col_out_454 = {u_ca_out_454[18:0],u_ca_out_453[75:19], u_ca_out_452[132:76], u_ca_out_451[151:133]};
assign col_out_455 = {u_ca_out_455[18:0],u_ca_out_454[75:19], u_ca_out_453[132:76], u_ca_out_452[151:133]};
assign col_out_456 = {u_ca_out_456[18:0],u_ca_out_455[75:19], u_ca_out_454[132:76], u_ca_out_453[151:133]};
assign col_out_457 = {u_ca_out_457[18:0],u_ca_out_456[75:19], u_ca_out_455[132:76], u_ca_out_454[151:133]};
assign col_out_458 = {u_ca_out_458[18:0],u_ca_out_457[75:19], u_ca_out_456[132:76], u_ca_out_455[151:133]};
assign col_out_459 = {u_ca_out_459[18:0],u_ca_out_458[75:19], u_ca_out_457[132:76], u_ca_out_456[151:133]};
assign col_out_460 = {u_ca_out_460[18:0],u_ca_out_459[75:19], u_ca_out_458[132:76], u_ca_out_457[151:133]};
assign col_out_461 = {u_ca_out_461[18:0],u_ca_out_460[75:19], u_ca_out_459[132:76], u_ca_out_458[151:133]};
assign col_out_462 = {u_ca_out_462[18:0],u_ca_out_461[75:19], u_ca_out_460[132:76], u_ca_out_459[151:133]};
assign col_out_463 = {u_ca_out_463[18:0],u_ca_out_462[75:19], u_ca_out_461[132:76], u_ca_out_460[151:133]};
assign col_out_464 = {u_ca_out_464[18:0],u_ca_out_463[75:19], u_ca_out_462[132:76], u_ca_out_461[151:133]};
assign col_out_465 = {u_ca_out_465[18:0],u_ca_out_464[75:19], u_ca_out_463[132:76], u_ca_out_462[151:133]};
assign col_out_466 = {u_ca_out_466[18:0],u_ca_out_465[75:19], u_ca_out_464[132:76], u_ca_out_463[151:133]};
assign col_out_467 = {u_ca_out_467[18:0],u_ca_out_466[75:19], u_ca_out_465[132:76], u_ca_out_464[151:133]};
assign col_out_468 = {u_ca_out_468[18:0],u_ca_out_467[75:19], u_ca_out_466[132:76], u_ca_out_465[151:133]};
assign col_out_469 = {u_ca_out_469[18:0],u_ca_out_468[75:19], u_ca_out_467[132:76], u_ca_out_466[151:133]};
assign col_out_470 = {u_ca_out_470[18:0],u_ca_out_469[75:19], u_ca_out_468[132:76], u_ca_out_467[151:133]};
assign col_out_471 = {u_ca_out_471[18:0],u_ca_out_470[75:19], u_ca_out_469[132:76], u_ca_out_468[151:133]};
assign col_out_472 = {u_ca_out_472[18:0],u_ca_out_471[75:19], u_ca_out_470[132:76], u_ca_out_469[151:133]};
assign col_out_473 = {u_ca_out_473[18:0],u_ca_out_472[75:19], u_ca_out_471[132:76], u_ca_out_470[151:133]};
assign col_out_474 = {u_ca_out_474[18:0],u_ca_out_473[75:19], u_ca_out_472[132:76], u_ca_out_471[151:133]};
assign col_out_475 = {u_ca_out_475[18:0],u_ca_out_474[75:19], u_ca_out_473[132:76], u_ca_out_472[151:133]};
assign col_out_476 = {u_ca_out_476[18:0],u_ca_out_475[75:19], u_ca_out_474[132:76], u_ca_out_473[151:133]};
assign col_out_477 = {u_ca_out_477[18:0],u_ca_out_476[75:19], u_ca_out_475[132:76], u_ca_out_474[151:133]};
assign col_out_478 = {u_ca_out_478[18:0],u_ca_out_477[75:19], u_ca_out_476[132:76], u_ca_out_475[151:133]};
assign col_out_479 = {u_ca_out_479[18:0],u_ca_out_478[75:19], u_ca_out_477[132:76], u_ca_out_476[151:133]};
assign col_out_480 = {u_ca_out_480[18:0],u_ca_out_479[75:19], u_ca_out_478[132:76], u_ca_out_477[151:133]};
assign col_out_481 = {u_ca_out_481[18:0],u_ca_out_480[75:19], u_ca_out_479[132:76], u_ca_out_478[151:133]};
assign col_out_482 = {u_ca_out_482[18:0],u_ca_out_481[75:19], u_ca_out_480[132:76], u_ca_out_479[151:133]};
assign col_out_483 = {u_ca_out_483[18:0],u_ca_out_482[75:19], u_ca_out_481[132:76], u_ca_out_480[151:133]};
assign col_out_484 = {u_ca_out_484[18:0],u_ca_out_483[75:19], u_ca_out_482[132:76], u_ca_out_481[151:133]};
assign col_out_485 = {u_ca_out_485[18:0],u_ca_out_484[75:19], u_ca_out_483[132:76], u_ca_out_482[151:133]};
assign col_out_486 = {u_ca_out_486[18:0],u_ca_out_485[75:19], u_ca_out_484[132:76], u_ca_out_483[151:133]};
assign col_out_487 = {u_ca_out_487[18:0],u_ca_out_486[75:19], u_ca_out_485[132:76], u_ca_out_484[151:133]};
assign col_out_488 = {u_ca_out_488[18:0],u_ca_out_487[75:19], u_ca_out_486[132:76], u_ca_out_485[151:133]};
assign col_out_489 = {u_ca_out_489[18:0],u_ca_out_488[75:19], u_ca_out_487[132:76], u_ca_out_486[151:133]};
assign col_out_490 = {u_ca_out_490[18:0],u_ca_out_489[75:19], u_ca_out_488[132:76], u_ca_out_487[151:133]};
assign col_out_491 = {u_ca_out_491[18:0],u_ca_out_490[75:19], u_ca_out_489[132:76], u_ca_out_488[151:133]};
assign col_out_492 = {u_ca_out_492[18:0],u_ca_out_491[75:19], u_ca_out_490[132:76], u_ca_out_489[151:133]};
assign col_out_493 = {u_ca_out_493[18:0],u_ca_out_492[75:19], u_ca_out_491[132:76], u_ca_out_490[151:133]};
assign col_out_494 = {u_ca_out_494[18:0],u_ca_out_493[75:19], u_ca_out_492[132:76], u_ca_out_491[151:133]};
assign col_out_495 = {u_ca_out_495[18:0],u_ca_out_494[75:19], u_ca_out_493[132:76], u_ca_out_492[151:133]};
assign col_out_496 = {u_ca_out_496[18:0],u_ca_out_495[75:19], u_ca_out_494[132:76], u_ca_out_493[151:133]};
assign col_out_497 = {u_ca_out_497[18:0],u_ca_out_496[75:19], u_ca_out_495[132:76], u_ca_out_494[151:133]};
assign col_out_498 = {u_ca_out_498[18:0],u_ca_out_497[75:19], u_ca_out_496[132:76], u_ca_out_495[151:133]};
assign col_out_499 = {u_ca_out_499[18:0],u_ca_out_498[75:19], u_ca_out_497[132:76], u_ca_out_496[151:133]};
assign col_out_500 = {u_ca_out_500[18:0],u_ca_out_499[75:19], u_ca_out_498[132:76], u_ca_out_497[151:133]};
assign col_out_501 = {u_ca_out_501[18:0],u_ca_out_500[75:19], u_ca_out_499[132:76], u_ca_out_498[151:133]};
assign col_out_502 = {u_ca_out_502[18:0],u_ca_out_501[75:19], u_ca_out_500[132:76], u_ca_out_499[151:133]};
assign col_out_503 = {u_ca_out_503[18:0],u_ca_out_502[75:19], u_ca_out_501[132:76], u_ca_out_500[151:133]};
assign col_out_504 = {u_ca_out_504[18:0],u_ca_out_503[75:19], u_ca_out_502[132:76], u_ca_out_501[151:133]};
assign col_out_505 = {u_ca_out_505[18:0],u_ca_out_504[75:19], u_ca_out_503[132:76], u_ca_out_502[151:133]};
assign col_out_506 = {u_ca_out_506[18:0],u_ca_out_505[75:19], u_ca_out_504[132:76], u_ca_out_503[151:133]};
assign col_out_507 = {u_ca_out_507[18:0],u_ca_out_506[75:19], u_ca_out_505[132:76], u_ca_out_504[151:133]};
assign col_out_508 = {u_ca_out_508[18:0],u_ca_out_507[75:19], u_ca_out_506[132:76], u_ca_out_505[151:133]};
assign col_out_509 = {u_ca_out_509[18:0],u_ca_out_508[75:19], u_ca_out_507[132:76], u_ca_out_506[151:133]};
assign col_out_510 = {u_ca_out_510[18:0],u_ca_out_509[75:19], u_ca_out_508[132:76], u_ca_out_507[151:133]};
assign col_out_511 = {u_ca_out_511[18:0],u_ca_out_510[75:19], u_ca_out_509[132:76], u_ca_out_508[151:133]};
assign col_out_512 = {u_ca_out_512[18:0],u_ca_out_511[75:19], u_ca_out_510[132:76], u_ca_out_509[151:133]};
assign col_out_513 = {u_ca_out_513[18:0],u_ca_out_512[75:19], u_ca_out_511[132:76], u_ca_out_510[151:133]};
assign col_out_514 = {u_ca_out_514[18:0],u_ca_out_513[75:19], u_ca_out_512[132:76], u_ca_out_511[151:133]};
assign col_out_515 = {u_ca_out_515[18:0],u_ca_out_514[75:19], u_ca_out_513[132:76], u_ca_out_512[151:133]};
assign col_out_516 = {u_ca_out_516[18:0],u_ca_out_515[75:19], u_ca_out_514[132:76], u_ca_out_513[151:133]};
assign col_out_517 = {u_ca_out_517[18:0],u_ca_out_516[75:19], u_ca_out_515[132:76], u_ca_out_514[151:133]};
assign col_out_518 = {u_ca_out_518[18:0],u_ca_out_517[75:19], u_ca_out_516[132:76], u_ca_out_515[151:133]};
assign col_out_519 = {u_ca_out_519[18:0],u_ca_out_518[75:19], u_ca_out_517[132:76], u_ca_out_516[151:133]};
assign col_out_520 = {u_ca_out_520[18:0],u_ca_out_519[75:19], u_ca_out_518[132:76], u_ca_out_517[151:133]};
assign col_out_521 = {u_ca_out_521[18:0],u_ca_out_520[75:19], u_ca_out_519[132:76], u_ca_out_518[151:133]};
assign col_out_522 = {u_ca_out_522[18:0],u_ca_out_521[75:19], u_ca_out_520[132:76], u_ca_out_519[151:133]};
assign col_out_523 = {u_ca_out_523[18:0],u_ca_out_522[75:19], u_ca_out_521[132:76], u_ca_out_520[151:133]};
assign col_out_524 = {u_ca_out_524[18:0],u_ca_out_523[75:19], u_ca_out_522[132:76], u_ca_out_521[151:133]};
assign col_out_525 = {u_ca_out_525[18:0],u_ca_out_524[75:19], u_ca_out_523[132:76], u_ca_out_522[151:133]};
assign col_out_526 = {u_ca_out_526[18:0],u_ca_out_525[75:19], u_ca_out_524[132:76], u_ca_out_523[151:133]};
assign col_out_527 = {u_ca_out_527[18:0],u_ca_out_526[75:19], u_ca_out_525[132:76], u_ca_out_524[151:133]};
assign col_out_528 = {u_ca_out_528[18:0],u_ca_out_527[75:19], u_ca_out_526[132:76], u_ca_out_525[151:133]};
assign col_out_529 = {u_ca_out_529[18:0],u_ca_out_528[75:19], u_ca_out_527[132:76], u_ca_out_526[151:133]};
assign col_out_530 = {u_ca_out_530[18:0],u_ca_out_529[75:19], u_ca_out_528[132:76], u_ca_out_527[151:133]};
assign col_out_531 = {u_ca_out_531[18:0],u_ca_out_530[75:19], u_ca_out_529[132:76], u_ca_out_528[151:133]};
assign col_out_532 = {u_ca_out_532[18:0],u_ca_out_531[75:19], u_ca_out_530[132:76], u_ca_out_529[151:133]};
assign col_out_533 = {u_ca_out_533[18:0],u_ca_out_532[75:19], u_ca_out_531[132:76], u_ca_out_530[151:133]};
assign col_out_534 = {u_ca_out_534[18:0],u_ca_out_533[75:19], u_ca_out_532[132:76], u_ca_out_531[151:133]};
assign col_out_535 = {u_ca_out_535[18:0],u_ca_out_534[75:19], u_ca_out_533[132:76], u_ca_out_532[151:133]};
assign col_out_536 = {u_ca_out_536[18:0],u_ca_out_535[75:19], u_ca_out_534[132:76], u_ca_out_533[151:133]};
assign col_out_537 = {u_ca_out_537[18:0],u_ca_out_536[75:19], u_ca_out_535[132:76], u_ca_out_534[151:133]};
assign col_out_538 = {u_ca_out_538[18:0],u_ca_out_537[75:19], u_ca_out_536[132:76], u_ca_out_535[151:133]};
assign col_out_539 = {u_ca_out_539[18:0],u_ca_out_538[75:19], u_ca_out_537[132:76], u_ca_out_536[151:133]};
assign col_out_540 = {u_ca_out_540[18:0],u_ca_out_539[75:19], u_ca_out_538[132:76], u_ca_out_537[151:133]};
assign col_out_541 = {u_ca_out_541[18:0],u_ca_out_540[75:19], u_ca_out_539[132:76], u_ca_out_538[151:133]};
assign col_out_542 = {u_ca_out_542[18:0],u_ca_out_541[75:19], u_ca_out_540[132:76], u_ca_out_539[151:133]};
assign col_out_543 = {u_ca_out_543[18:0],u_ca_out_542[75:19], u_ca_out_541[132:76], u_ca_out_540[151:133]};
assign col_out_544 = {u_ca_out_544[18:0],u_ca_out_543[75:19], u_ca_out_542[132:76], u_ca_out_541[151:133]};
assign col_out_545 = {u_ca_out_545[18:0],u_ca_out_544[75:19], u_ca_out_543[132:76], u_ca_out_542[151:133]};
assign col_out_546 = {u_ca_out_546[18:0],u_ca_out_545[75:19], u_ca_out_544[132:76], u_ca_out_543[151:133]};
assign col_out_547 = {u_ca_out_547[18:0],u_ca_out_546[75:19], u_ca_out_545[132:76], u_ca_out_544[151:133]};
assign col_out_548 = {u_ca_out_548[18:0],u_ca_out_547[75:19], u_ca_out_546[132:76], u_ca_out_545[151:133]};
assign col_out_549 = {u_ca_out_549[18:0],u_ca_out_548[75:19], u_ca_out_547[132:76], u_ca_out_546[151:133]};
assign col_out_550 = {u_ca_out_550[18:0],u_ca_out_549[75:19], u_ca_out_548[132:76], u_ca_out_547[151:133]};
assign col_out_551 = {u_ca_out_551[18:0],u_ca_out_550[75:19], u_ca_out_549[132:76], u_ca_out_548[151:133]};
assign col_out_552 = {u_ca_out_552[18:0],u_ca_out_551[75:19], u_ca_out_550[132:76], u_ca_out_549[151:133]};
assign col_out_553 = {u_ca_out_553[18:0],u_ca_out_552[75:19], u_ca_out_551[132:76], u_ca_out_550[151:133]};
assign col_out_554 = {u_ca_out_554[18:0],u_ca_out_553[75:19], u_ca_out_552[132:76], u_ca_out_551[151:133]};
assign col_out_555 = {u_ca_out_555[18:0],u_ca_out_554[75:19], u_ca_out_553[132:76], u_ca_out_552[151:133]};
assign col_out_556 = {u_ca_out_556[18:0],u_ca_out_555[75:19], u_ca_out_554[132:76], u_ca_out_553[151:133]};
assign col_out_557 = {u_ca_out_557[18:0],u_ca_out_556[75:19], u_ca_out_555[132:76], u_ca_out_554[151:133]};
assign col_out_558 = {u_ca_out_558[18:0],u_ca_out_557[75:19], u_ca_out_556[132:76], u_ca_out_555[151:133]};
assign col_out_559 = {u_ca_out_559[18:0],u_ca_out_558[75:19], u_ca_out_557[132:76], u_ca_out_556[151:133]};
assign col_out_560 = {u_ca_out_560[18:0],u_ca_out_559[75:19], u_ca_out_558[132:76], u_ca_out_557[151:133]};
assign col_out_561 = {u_ca_out_561[18:0],u_ca_out_560[75:19], u_ca_out_559[132:76], u_ca_out_558[151:133]};
assign col_out_562 = {u_ca_out_562[18:0],u_ca_out_561[75:19], u_ca_out_560[132:76], u_ca_out_559[151:133]};
assign col_out_563 = {u_ca_out_563[18:0],u_ca_out_562[75:19], u_ca_out_561[132:76], u_ca_out_560[151:133]};
assign col_out_564 = {u_ca_out_564[18:0],u_ca_out_563[75:19], u_ca_out_562[132:76], u_ca_out_561[151:133]};
assign col_out_565 = {u_ca_out_565[18:0],u_ca_out_564[75:19], u_ca_out_563[132:76], u_ca_out_562[151:133]};
assign col_out_566 = {u_ca_out_566[18:0],u_ca_out_565[75:19], u_ca_out_564[132:76], u_ca_out_563[151:133]};
assign col_out_567 = {u_ca_out_567[18:0],u_ca_out_566[75:19], u_ca_out_565[132:76], u_ca_out_564[151:133]};
assign col_out_568 = {u_ca_out_568[18:0],u_ca_out_567[75:19], u_ca_out_566[132:76], u_ca_out_565[151:133]};
assign col_out_569 = {u_ca_out_569[18:0],u_ca_out_568[75:19], u_ca_out_567[132:76], u_ca_out_566[151:133]};
assign col_out_570 = {u_ca_out_570[18:0],u_ca_out_569[75:19], u_ca_out_568[132:76], u_ca_out_567[151:133]};
assign col_out_571 = {u_ca_out_571[18:0],u_ca_out_570[75:19], u_ca_out_569[132:76], u_ca_out_568[151:133]};
assign col_out_572 = {u_ca_out_572[18:0],u_ca_out_571[75:19], u_ca_out_570[132:76], u_ca_out_569[151:133]};
assign col_out_573 = {u_ca_out_573[18:0],u_ca_out_572[75:19], u_ca_out_571[132:76], u_ca_out_570[151:133]};
assign col_out_574 = {u_ca_out_574[18:0],u_ca_out_573[75:19], u_ca_out_572[132:76], u_ca_out_571[151:133]};
assign col_out_575 = {u_ca_out_575[18:0],u_ca_out_574[75:19], u_ca_out_573[132:76], u_ca_out_572[151:133]};
assign col_out_576 = {u_ca_out_576[18:0],u_ca_out_575[75:19], u_ca_out_574[132:76], u_ca_out_573[151:133]};
assign col_out_577 = {u_ca_out_577[18:0],u_ca_out_576[75:19], u_ca_out_575[132:76], u_ca_out_574[151:133]};
assign col_out_578 = {u_ca_out_578[18:0],u_ca_out_577[75:19], u_ca_out_576[132:76], u_ca_out_575[151:133]};
assign col_out_579 = {u_ca_out_579[18:0],u_ca_out_578[75:19], u_ca_out_577[132:76], u_ca_out_576[151:133]};
assign col_out_580 = {u_ca_out_580[18:0],u_ca_out_579[75:19], u_ca_out_578[132:76], u_ca_out_577[151:133]};
assign col_out_581 = {u_ca_out_581[18:0],u_ca_out_580[75:19], u_ca_out_579[132:76], u_ca_out_578[151:133]};
assign col_out_582 = {u_ca_out_582[18:0],u_ca_out_581[75:19], u_ca_out_580[132:76], u_ca_out_579[151:133]};
assign col_out_583 = {u_ca_out_583[18:0],u_ca_out_582[75:19], u_ca_out_581[132:76], u_ca_out_580[151:133]};
assign col_out_584 = {u_ca_out_584[18:0],u_ca_out_583[75:19], u_ca_out_582[132:76], u_ca_out_581[151:133]};
assign col_out_585 = {u_ca_out_585[18:0],u_ca_out_584[75:19], u_ca_out_583[132:76], u_ca_out_582[151:133]};
assign col_out_586 = {u_ca_out_586[18:0],u_ca_out_585[75:19], u_ca_out_584[132:76], u_ca_out_583[151:133]};
assign col_out_587 = {u_ca_out_587[18:0],u_ca_out_586[75:19], u_ca_out_585[132:76], u_ca_out_584[151:133]};
assign col_out_588 = {u_ca_out_588[18:0],u_ca_out_587[75:19], u_ca_out_586[132:76], u_ca_out_585[151:133]};
assign col_out_589 = {u_ca_out_589[18:0],u_ca_out_588[75:19], u_ca_out_587[132:76], u_ca_out_586[151:133]};
assign col_out_590 = {u_ca_out_590[18:0],u_ca_out_589[75:19], u_ca_out_588[132:76], u_ca_out_587[151:133]};
assign col_out_591 = {u_ca_out_591[18:0],u_ca_out_590[75:19], u_ca_out_589[132:76], u_ca_out_588[151:133]};
assign col_out_592 = {u_ca_out_592[18:0],u_ca_out_591[75:19], u_ca_out_590[132:76], u_ca_out_589[151:133]};
assign col_out_593 = {u_ca_out_593[18:0],u_ca_out_592[75:19], u_ca_out_591[132:76], u_ca_out_590[151:133]};
assign col_out_594 = {u_ca_out_594[18:0],u_ca_out_593[75:19], u_ca_out_592[132:76], u_ca_out_591[151:133]};
assign col_out_595 = {u_ca_out_595[18:0],u_ca_out_594[75:19], u_ca_out_593[132:76], u_ca_out_592[151:133]};
assign col_out_596 = {u_ca_out_596[18:0],u_ca_out_595[75:19], u_ca_out_594[132:76], u_ca_out_593[151:133]};
assign col_out_597 = {u_ca_out_597[18:0],u_ca_out_596[75:19], u_ca_out_595[132:76], u_ca_out_594[151:133]};
assign col_out_598 = {u_ca_out_598[18:0],u_ca_out_597[75:19], u_ca_out_596[132:76], u_ca_out_595[151:133]};
assign col_out_599 = {u_ca_out_599[18:0],u_ca_out_598[75:19], u_ca_out_597[132:76], u_ca_out_596[151:133]};
assign col_out_600 = {u_ca_out_600[18:0],u_ca_out_599[75:19], u_ca_out_598[132:76], u_ca_out_597[151:133]};
assign col_out_601 = {u_ca_out_601[18:0],u_ca_out_600[75:19], u_ca_out_599[132:76], u_ca_out_598[151:133]};
assign col_out_602 = {u_ca_out_602[18:0],u_ca_out_601[75:19], u_ca_out_600[132:76], u_ca_out_599[151:133]};
assign col_out_603 = {u_ca_out_603[18:0],u_ca_out_602[75:19], u_ca_out_601[132:76], u_ca_out_600[151:133]};
assign col_out_604 = {u_ca_out_604[18:0],u_ca_out_603[75:19], u_ca_out_602[132:76], u_ca_out_601[151:133]};
assign col_out_605 = {u_ca_out_605[18:0],u_ca_out_604[75:19], u_ca_out_603[132:76], u_ca_out_602[151:133]};
assign col_out_606 = {u_ca_out_606[18:0],u_ca_out_605[75:19], u_ca_out_604[132:76], u_ca_out_603[151:133]};
assign col_out_607 = {u_ca_out_607[18:0],u_ca_out_606[75:19], u_ca_out_605[132:76], u_ca_out_604[151:133]};
assign col_out_608 = {u_ca_out_608[18:0],u_ca_out_607[75:19], u_ca_out_606[132:76], u_ca_out_605[151:133]};
assign col_out_609 = {u_ca_out_609[18:0],u_ca_out_608[75:19], u_ca_out_607[132:76], u_ca_out_606[151:133]};
assign col_out_610 = {u_ca_out_610[18:0],u_ca_out_609[75:19], u_ca_out_608[132:76], u_ca_out_607[151:133]};
assign col_out_611 = {u_ca_out_611[18:0],u_ca_out_610[75:19], u_ca_out_609[132:76], u_ca_out_608[151:133]};
assign col_out_612 = {u_ca_out_612[18:0],u_ca_out_611[75:19], u_ca_out_610[132:76], u_ca_out_609[151:133]};
assign col_out_613 = {u_ca_out_613[18:0],u_ca_out_612[75:19], u_ca_out_611[132:76], u_ca_out_610[151:133]};
assign col_out_614 = {u_ca_out_614[18:0],u_ca_out_613[75:19], u_ca_out_612[132:76], u_ca_out_611[151:133]};
assign col_out_615 = {u_ca_out_615[18:0],u_ca_out_614[75:19], u_ca_out_613[132:76], u_ca_out_612[151:133]};
assign col_out_616 = {u_ca_out_616[18:0],u_ca_out_615[75:19], u_ca_out_614[132:76], u_ca_out_613[151:133]};
assign col_out_617 = {u_ca_out_617[18:0],u_ca_out_616[75:19], u_ca_out_615[132:76], u_ca_out_614[151:133]};
assign col_out_618 = {u_ca_out_618[18:0],u_ca_out_617[75:19], u_ca_out_616[132:76], u_ca_out_615[151:133]};
assign col_out_619 = {u_ca_out_619[18:0],u_ca_out_618[75:19], u_ca_out_617[132:76], u_ca_out_616[151:133]};
assign col_out_620 = {u_ca_out_620[18:0],u_ca_out_619[75:19], u_ca_out_618[132:76], u_ca_out_617[151:133]};
assign col_out_621 = {u_ca_out_621[18:0],u_ca_out_620[75:19], u_ca_out_619[132:76], u_ca_out_618[151:133]};
assign col_out_622 = {u_ca_out_622[18:0],u_ca_out_621[75:19], u_ca_out_620[132:76], u_ca_out_619[151:133]};
assign col_out_623 = {u_ca_out_623[18:0],u_ca_out_622[75:19], u_ca_out_621[132:76], u_ca_out_620[151:133]};
assign col_out_624 = {u_ca_out_624[18:0],u_ca_out_623[75:19], u_ca_out_622[132:76], u_ca_out_621[151:133]};
assign col_out_625 = {u_ca_out_625[18:0],u_ca_out_624[75:19], u_ca_out_623[132:76], u_ca_out_622[151:133]};
assign col_out_626 = {u_ca_out_626[18:0],u_ca_out_625[75:19], u_ca_out_624[132:76], u_ca_out_623[151:133]};
assign col_out_627 = {u_ca_out_627[18:0],u_ca_out_626[75:19], u_ca_out_625[132:76], u_ca_out_624[151:133]};
assign col_out_628 = {u_ca_out_628[18:0],u_ca_out_627[75:19], u_ca_out_626[132:76], u_ca_out_625[151:133]};
assign col_out_629 = {u_ca_out_629[18:0],u_ca_out_628[75:19], u_ca_out_627[132:76], u_ca_out_626[151:133]};
assign col_out_630 = {u_ca_out_630[18:0],u_ca_out_629[75:19], u_ca_out_628[132:76], u_ca_out_627[151:133]};
assign col_out_631 = {u_ca_out_631[18:0],u_ca_out_630[75:19], u_ca_out_629[132:76], u_ca_out_628[151:133]};
assign col_out_632 = {u_ca_out_632[18:0],u_ca_out_631[75:19], u_ca_out_630[132:76], u_ca_out_629[151:133]};
assign col_out_633 = {u_ca_out_633[18:0],u_ca_out_632[75:19], u_ca_out_631[132:76], u_ca_out_630[151:133]};
assign col_out_634 = {u_ca_out_634[18:0],u_ca_out_633[75:19], u_ca_out_632[132:76], u_ca_out_631[151:133]};
assign col_out_635 = {u_ca_out_635[18:0],u_ca_out_634[75:19], u_ca_out_633[132:76], u_ca_out_632[151:133]};
assign col_out_636 = {u_ca_out_636[18:0],u_ca_out_635[75:19], u_ca_out_634[132:76], u_ca_out_633[151:133]};
assign col_out_637 = {u_ca_out_637[18:0],u_ca_out_636[75:19], u_ca_out_635[132:76], u_ca_out_634[151:133]};
assign col_out_638 = {u_ca_out_638[18:0],u_ca_out_637[75:19], u_ca_out_636[132:76], u_ca_out_635[151:133]};
assign col_out_639 = {u_ca_out_639[18:0],u_ca_out_638[75:19], u_ca_out_637[132:76], u_ca_out_636[151:133]};
assign col_out_640 = {u_ca_out_640[18:0],u_ca_out_639[75:19], u_ca_out_638[132:76], u_ca_out_637[151:133]};
assign col_out_641 = {u_ca_out_641[18:0],u_ca_out_640[75:19], u_ca_out_639[132:76], u_ca_out_638[151:133]};
assign col_out_642 = {u_ca_out_642[18:0],u_ca_out_641[75:19], u_ca_out_640[132:76], u_ca_out_639[151:133]};
assign col_out_643 = {u_ca_out_643[18:0],u_ca_out_642[75:19], u_ca_out_641[132:76], u_ca_out_640[151:133]};
assign col_out_644 = {u_ca_out_644[18:0],u_ca_out_643[75:19], u_ca_out_642[132:76], u_ca_out_641[151:133]};
assign col_out_645 = {u_ca_out_645[18:0],u_ca_out_644[75:19], u_ca_out_643[132:76], u_ca_out_642[151:133]};
assign col_out_646 = {u_ca_out_646[18:0],u_ca_out_645[75:19], u_ca_out_644[132:76], u_ca_out_643[151:133]};
assign col_out_647 = {u_ca_out_647[18:0],u_ca_out_646[75:19], u_ca_out_645[132:76], u_ca_out_644[151:133]};
assign col_out_648 = {u_ca_out_648[18:0],u_ca_out_647[75:19], u_ca_out_646[132:76], u_ca_out_645[151:133]};
assign col_out_649 = {u_ca_out_649[18:0],u_ca_out_648[75:19], u_ca_out_647[132:76], u_ca_out_646[151:133]};
assign col_out_650 = {u_ca_out_650[18:0],u_ca_out_649[75:19], u_ca_out_648[132:76], u_ca_out_647[151:133]};
assign col_out_651 = {u_ca_out_651[18:0],u_ca_out_650[75:19], u_ca_out_649[132:76], u_ca_out_648[151:133]};
assign col_out_652 = {u_ca_out_652[18:0],u_ca_out_651[75:19], u_ca_out_650[132:76], u_ca_out_649[151:133]};
assign col_out_653 = {u_ca_out_653[18:0],u_ca_out_652[75:19], u_ca_out_651[132:76], u_ca_out_650[151:133]};
assign col_out_654 = {u_ca_out_654[18:0],u_ca_out_653[75:19], u_ca_out_652[132:76], u_ca_out_651[151:133]};
assign col_out_655 = {u_ca_out_655[18:0],u_ca_out_654[75:19], u_ca_out_653[132:76], u_ca_out_652[151:133]};
assign col_out_656 = {u_ca_out_656[18:0],u_ca_out_655[75:19], u_ca_out_654[132:76], u_ca_out_653[151:133]};
assign col_out_657 = {u_ca_out_657[18:0],u_ca_out_656[75:19], u_ca_out_655[132:76], u_ca_out_654[151:133]};
assign col_out_658 = {u_ca_out_658[18:0],u_ca_out_657[75:19], u_ca_out_656[132:76], u_ca_out_655[151:133]};
assign col_out_659 = {u_ca_out_659[18:0],u_ca_out_658[75:19], u_ca_out_657[132:76], u_ca_out_656[151:133]};
assign col_out_660 = {u_ca_out_660[18:0],u_ca_out_659[75:19], u_ca_out_658[132:76], u_ca_out_657[151:133]};
assign col_out_661 = {u_ca_out_661[18:0],u_ca_out_660[75:19], u_ca_out_659[132:76], u_ca_out_658[151:133]};
assign col_out_662 = {u_ca_out_662[18:0],u_ca_out_661[75:19], u_ca_out_660[132:76], u_ca_out_659[151:133]};
assign col_out_663 = {u_ca_out_663[18:0],u_ca_out_662[75:19], u_ca_out_661[132:76], u_ca_out_660[151:133]};
assign col_out_664 = {u_ca_out_664[18:0],u_ca_out_663[75:19], u_ca_out_662[132:76], u_ca_out_661[151:133]};
assign col_out_665 = {u_ca_out_665[18:0],u_ca_out_664[75:19], u_ca_out_663[132:76], u_ca_out_662[151:133]};
assign col_out_666 = {u_ca_out_666[18:0],u_ca_out_665[75:19], u_ca_out_664[132:76], u_ca_out_663[151:133]};
assign col_out_667 = {u_ca_out_667[18:0],u_ca_out_666[75:19], u_ca_out_665[132:76], u_ca_out_664[151:133]};
assign col_out_668 = {u_ca_out_668[18:0],u_ca_out_667[75:19], u_ca_out_666[132:76], u_ca_out_665[151:133]};
assign col_out_669 = {u_ca_out_669[18:0],u_ca_out_668[75:19], u_ca_out_667[132:76], u_ca_out_666[151:133]};
assign col_out_670 = {u_ca_out_670[18:0],u_ca_out_669[75:19], u_ca_out_668[132:76], u_ca_out_667[151:133]};
assign col_out_671 = {u_ca_out_671[18:0],u_ca_out_670[75:19], u_ca_out_669[132:76], u_ca_out_668[151:133]};
assign col_out_672 = {u_ca_out_672[18:0],u_ca_out_671[75:19], u_ca_out_670[132:76], u_ca_out_669[151:133]};
assign col_out_673 = {u_ca_out_673[18:0],u_ca_out_672[75:19], u_ca_out_671[132:76], u_ca_out_670[151:133]};
assign col_out_674 = {u_ca_out_674[18:0],u_ca_out_673[75:19], u_ca_out_672[132:76], u_ca_out_671[151:133]};
assign col_out_675 = {u_ca_out_675[18:0],u_ca_out_674[75:19], u_ca_out_673[132:76], u_ca_out_672[151:133]};
assign col_out_676 = {u_ca_out_676[18:0],u_ca_out_675[75:19], u_ca_out_674[132:76], u_ca_out_673[151:133]};
assign col_out_677 = {u_ca_out_677[18:0],u_ca_out_676[75:19], u_ca_out_675[132:76], u_ca_out_674[151:133]};
assign col_out_678 = {u_ca_out_678[18:0],u_ca_out_677[75:19], u_ca_out_676[132:76], u_ca_out_675[151:133]};
assign col_out_679 = {u_ca_out_679[18:0],u_ca_out_678[75:19], u_ca_out_677[132:76], u_ca_out_676[151:133]};
assign col_out_680 = {u_ca_out_680[18:0],u_ca_out_679[75:19], u_ca_out_678[132:76], u_ca_out_677[151:133]};
assign col_out_681 = {u_ca_out_681[18:0],u_ca_out_680[75:19], u_ca_out_679[132:76], u_ca_out_678[151:133]};
assign col_out_682 = {u_ca_out_682[18:0],u_ca_out_681[75:19], u_ca_out_680[132:76], u_ca_out_679[151:133]};
assign col_out_683 = {u_ca_out_683[18:0],u_ca_out_682[75:19], u_ca_out_681[132:76], u_ca_out_680[151:133]};
assign col_out_684 = {u_ca_out_684[18:0],u_ca_out_683[75:19], u_ca_out_682[132:76], u_ca_out_681[151:133]};
assign col_out_685 = {u_ca_out_685[18:0],u_ca_out_684[75:19], u_ca_out_683[132:76], u_ca_out_682[151:133]};
assign col_out_686 = {u_ca_out_686[18:0],u_ca_out_685[75:19], u_ca_out_684[132:76], u_ca_out_683[151:133]};
assign col_out_687 = {u_ca_out_687[18:0],u_ca_out_686[75:19], u_ca_out_685[132:76], u_ca_out_684[151:133]};
assign col_out_688 = {u_ca_out_688[18:0],u_ca_out_687[75:19], u_ca_out_686[132:76], u_ca_out_685[151:133]};
assign col_out_689 = {u_ca_out_689[18:0],u_ca_out_688[75:19], u_ca_out_687[132:76], u_ca_out_686[151:133]};
assign col_out_690 = {u_ca_out_690[18:0],u_ca_out_689[75:19], u_ca_out_688[132:76], u_ca_out_687[151:133]};
assign col_out_691 = {u_ca_out_691[18:0],u_ca_out_690[75:19], u_ca_out_689[132:76], u_ca_out_688[151:133]};
assign col_out_692 = {u_ca_out_692[18:0],u_ca_out_691[75:19], u_ca_out_690[132:76], u_ca_out_689[151:133]};
assign col_out_693 = {u_ca_out_693[18:0],u_ca_out_692[75:19], u_ca_out_691[132:76], u_ca_out_690[151:133]};
assign col_out_694 = {u_ca_out_694[18:0],u_ca_out_693[75:19], u_ca_out_692[132:76], u_ca_out_691[151:133]};
assign col_out_695 = {u_ca_out_695[18:0],u_ca_out_694[75:19], u_ca_out_693[132:76], u_ca_out_692[151:133]};
assign col_out_696 = {u_ca_out_696[18:0],u_ca_out_695[75:19], u_ca_out_694[132:76], u_ca_out_693[151:133]};
assign col_out_697 = {u_ca_out_697[18:0],u_ca_out_696[75:19], u_ca_out_695[132:76], u_ca_out_694[151:133]};
assign col_out_698 = {u_ca_out_698[18:0],u_ca_out_697[75:19], u_ca_out_696[132:76], u_ca_out_695[151:133]};
assign col_out_699 = {u_ca_out_699[18:0],u_ca_out_698[75:19], u_ca_out_697[132:76], u_ca_out_696[151:133]};
assign col_out_700 = {u_ca_out_700[18:0],u_ca_out_699[75:19], u_ca_out_698[132:76], u_ca_out_697[151:133]};
assign col_out_701 = {u_ca_out_701[18:0],u_ca_out_700[75:19], u_ca_out_699[132:76], u_ca_out_698[151:133]};
assign col_out_702 = {u_ca_out_702[18:0],u_ca_out_701[75:19], u_ca_out_700[132:76], u_ca_out_699[151:133]};
assign col_out_703 = {u_ca_out_703[18:0],u_ca_out_702[75:19], u_ca_out_701[132:76], u_ca_out_700[151:133]};
assign col_out_704 = {u_ca_out_704[18:0],u_ca_out_703[75:19], u_ca_out_702[132:76], u_ca_out_701[151:133]};
assign col_out_705 = {u_ca_out_705[18:0],u_ca_out_704[75:19], u_ca_out_703[132:76], u_ca_out_702[151:133]};
assign col_out_706 = {u_ca_out_706[18:0],u_ca_out_705[75:19], u_ca_out_704[132:76], u_ca_out_703[151:133]};
assign col_out_707 = {u_ca_out_707[18:0],u_ca_out_706[75:19], u_ca_out_705[132:76], u_ca_out_704[151:133]};
assign col_out_708 = {u_ca_out_708[18:0],u_ca_out_707[75:19], u_ca_out_706[132:76], u_ca_out_705[151:133]};
assign col_out_709 = {u_ca_out_709[18:0],u_ca_out_708[75:19], u_ca_out_707[132:76], u_ca_out_706[151:133]};
assign col_out_710 = {u_ca_out_710[18:0],u_ca_out_709[75:19], u_ca_out_708[132:76], u_ca_out_707[151:133]};
assign col_out_711 = {u_ca_out_711[18:0],u_ca_out_710[75:19], u_ca_out_709[132:76], u_ca_out_708[151:133]};
assign col_out_712 = {u_ca_out_712[18:0],u_ca_out_711[75:19], u_ca_out_710[132:76], u_ca_out_709[151:133]};
assign col_out_713 = {u_ca_out_713[18:0],u_ca_out_712[75:19], u_ca_out_711[132:76], u_ca_out_710[151:133]};
assign col_out_714 = {u_ca_out_714[18:0],u_ca_out_713[75:19], u_ca_out_712[132:76], u_ca_out_711[151:133]};
assign col_out_715 = {u_ca_out_715[18:0],u_ca_out_714[75:19], u_ca_out_713[132:76], u_ca_out_712[151:133]};
assign col_out_716 = {u_ca_out_716[18:0],u_ca_out_715[75:19], u_ca_out_714[132:76], u_ca_out_713[151:133]};
assign col_out_717 = {u_ca_out_717[18:0],u_ca_out_716[75:19], u_ca_out_715[132:76], u_ca_out_714[151:133]};
assign col_out_718 = {u_ca_out_718[18:0],u_ca_out_717[75:19], u_ca_out_716[132:76], u_ca_out_715[151:133]};
assign col_out_719 = {u_ca_out_719[18:0],u_ca_out_718[75:19], u_ca_out_717[132:76], u_ca_out_716[151:133]};
assign col_out_720 = {u_ca_out_720[18:0],u_ca_out_719[75:19], u_ca_out_718[132:76], u_ca_out_717[151:133]};
assign col_out_721 = {u_ca_out_721[18:0],u_ca_out_720[75:19], u_ca_out_719[132:76], u_ca_out_718[151:133]};
assign col_out_722 = {u_ca_out_722[18:0],u_ca_out_721[75:19], u_ca_out_720[132:76], u_ca_out_719[151:133]};
assign col_out_723 = {u_ca_out_723[18:0],u_ca_out_722[75:19], u_ca_out_721[132:76], u_ca_out_720[151:133]};
assign col_out_724 = {u_ca_out_724[18:0],u_ca_out_723[75:19], u_ca_out_722[132:76], u_ca_out_721[151:133]};
assign col_out_725 = {u_ca_out_725[18:0],u_ca_out_724[75:19], u_ca_out_723[132:76], u_ca_out_722[151:133]};
assign col_out_726 = {u_ca_out_726[18:0],u_ca_out_725[75:19], u_ca_out_724[132:76], u_ca_out_723[151:133]};
assign col_out_727 = {u_ca_out_727[18:0],u_ca_out_726[75:19], u_ca_out_725[132:76], u_ca_out_724[151:133]};
assign col_out_728 = {u_ca_out_728[18:0],u_ca_out_727[75:19], u_ca_out_726[132:76], u_ca_out_725[151:133]};
assign col_out_729 = {u_ca_out_729[18:0],u_ca_out_728[75:19], u_ca_out_727[132:76], u_ca_out_726[151:133]};
assign col_out_730 = {u_ca_out_730[18:0],u_ca_out_729[75:19], u_ca_out_728[132:76], u_ca_out_727[151:133]};
assign col_out_731 = {u_ca_out_731[18:0],u_ca_out_730[75:19], u_ca_out_729[132:76], u_ca_out_728[151:133]};
assign col_out_732 = {u_ca_out_732[18:0],u_ca_out_731[75:19], u_ca_out_730[132:76], u_ca_out_729[151:133]};
assign col_out_733 = {u_ca_out_733[18:0],u_ca_out_732[75:19], u_ca_out_731[132:76], u_ca_out_730[151:133]};
assign col_out_734 = {u_ca_out_734[18:0],u_ca_out_733[75:19], u_ca_out_732[132:76], u_ca_out_731[151:133]};
assign col_out_735 = {u_ca_out_735[18:0],u_ca_out_734[75:19], u_ca_out_733[132:76], u_ca_out_732[151:133]};
assign col_out_736 = {u_ca_out_736[18:0],u_ca_out_735[75:19], u_ca_out_734[132:76], u_ca_out_733[151:133]};
assign col_out_737 = {u_ca_out_737[18:0],u_ca_out_736[75:19], u_ca_out_735[132:76], u_ca_out_734[151:133]};
assign col_out_738 = {u_ca_out_738[18:0],u_ca_out_737[75:19], u_ca_out_736[132:76], u_ca_out_735[151:133]};
assign col_out_739 = {u_ca_out_739[18:0],u_ca_out_738[75:19], u_ca_out_737[132:76], u_ca_out_736[151:133]};
assign col_out_740 = {u_ca_out_740[18:0],u_ca_out_739[75:19], u_ca_out_738[132:76], u_ca_out_737[151:133]};
assign col_out_741 = {u_ca_out_741[18:0],u_ca_out_740[75:19], u_ca_out_739[132:76], u_ca_out_738[151:133]};
assign col_out_742 = {u_ca_out_742[18:0],u_ca_out_741[75:19], u_ca_out_740[132:76], u_ca_out_739[151:133]};
assign col_out_743 = {u_ca_out_743[18:0],u_ca_out_742[75:19], u_ca_out_741[132:76], u_ca_out_740[151:133]};
assign col_out_744 = {u_ca_out_744[18:0],u_ca_out_743[75:19], u_ca_out_742[132:76], u_ca_out_741[151:133]};
assign col_out_745 = {u_ca_out_745[18:0],u_ca_out_744[75:19], u_ca_out_743[132:76], u_ca_out_742[151:133]};
assign col_out_746 = {u_ca_out_746[18:0],u_ca_out_745[75:19], u_ca_out_744[132:76], u_ca_out_743[151:133]};
assign col_out_747 = {u_ca_out_747[18:0],u_ca_out_746[75:19], u_ca_out_745[132:76], u_ca_out_744[151:133]};
assign col_out_748 = {u_ca_out_748[18:0],u_ca_out_747[75:19], u_ca_out_746[132:76], u_ca_out_745[151:133]};
assign col_out_749 = {u_ca_out_749[18:0],u_ca_out_748[75:19], u_ca_out_747[132:76], u_ca_out_746[151:133]};
assign col_out_750 = {u_ca_out_750[18:0],u_ca_out_749[75:19], u_ca_out_748[132:76], u_ca_out_747[151:133]};
assign col_out_751 = {u_ca_out_751[18:0],u_ca_out_750[75:19], u_ca_out_749[132:76], u_ca_out_748[151:133]};
assign col_out_752 = {u_ca_out_752[18:0],u_ca_out_751[75:19], u_ca_out_750[132:76], u_ca_out_749[151:133]};
assign col_out_753 = {u_ca_out_753[18:0],u_ca_out_752[75:19], u_ca_out_751[132:76], u_ca_out_750[151:133]};
assign col_out_754 = {u_ca_out_754[18:0],u_ca_out_753[75:19], u_ca_out_752[132:76], u_ca_out_751[151:133]};
assign col_out_755 = {u_ca_out_755[18:0],u_ca_out_754[75:19], u_ca_out_753[132:76], u_ca_out_752[151:133]};
assign col_out_756 = {u_ca_out_756[18:0],u_ca_out_755[75:19], u_ca_out_754[132:76], u_ca_out_753[151:133]};
assign col_out_757 = {u_ca_out_757[18:0],u_ca_out_756[75:19], u_ca_out_755[132:76], u_ca_out_754[151:133]};
assign col_out_758 = {u_ca_out_758[18:0],u_ca_out_757[75:19], u_ca_out_756[132:76], u_ca_out_755[151:133]};
assign col_out_759 = {u_ca_out_759[18:0],u_ca_out_758[75:19], u_ca_out_757[132:76], u_ca_out_756[151:133]};
assign col_out_760 = {u_ca_out_760[18:0],u_ca_out_759[75:19], u_ca_out_758[132:76], u_ca_out_757[151:133]};
assign col_out_761 = {u_ca_out_761[18:0],u_ca_out_760[75:19], u_ca_out_759[132:76], u_ca_out_758[151:133]};
assign col_out_762 = {u_ca_out_762[18:0],u_ca_out_761[75:19], u_ca_out_760[132:76], u_ca_out_759[151:133]};
assign col_out_763 = {u_ca_out_763[18:0],u_ca_out_762[75:19], u_ca_out_761[132:76], u_ca_out_760[151:133]};
assign col_out_764 = {u_ca_out_764[18:0],u_ca_out_763[75:19], u_ca_out_762[132:76], u_ca_out_761[151:133]};
assign col_out_765 = {u_ca_out_765[18:0],u_ca_out_764[75:19], u_ca_out_763[132:76], u_ca_out_762[151:133]};
assign col_out_766 = {u_ca_out_766[18:0],u_ca_out_765[75:19], u_ca_out_764[132:76], u_ca_out_763[151:133]};
assign col_out_767 = {u_ca_out_767[18:0],u_ca_out_766[75:19], u_ca_out_765[132:76], u_ca_out_764[151:133]};
assign col_out_768 = {u_ca_out_768[18:0],u_ca_out_767[75:19], u_ca_out_766[132:76], u_ca_out_765[151:133]};
assign col_out_769 = {u_ca_out_769[18:0],u_ca_out_768[75:19], u_ca_out_767[132:76], u_ca_out_766[151:133]};
assign col_out_770 = {u_ca_out_770[18:0],u_ca_out_769[75:19], u_ca_out_768[132:76], u_ca_out_767[151:133]};
assign col_out_771 = {u_ca_out_771[18:0],u_ca_out_770[75:19], u_ca_out_769[132:76], u_ca_out_768[151:133]};
assign col_out_772 = {u_ca_out_772[18:0],u_ca_out_771[75:19], u_ca_out_770[132:76], u_ca_out_769[151:133]};
assign col_out_773 = {u_ca_out_773[18:0],u_ca_out_772[75:19], u_ca_out_771[132:76], u_ca_out_770[151:133]};
assign col_out_774 = {u_ca_out_774[18:0],u_ca_out_773[75:19], u_ca_out_772[132:76], u_ca_out_771[151:133]};
assign col_out_775 = {u_ca_out_775[18:0],u_ca_out_774[75:19], u_ca_out_773[132:76], u_ca_out_772[151:133]};
assign col_out_776 = {u_ca_out_776[18:0],u_ca_out_775[75:19], u_ca_out_774[132:76], u_ca_out_773[151:133]};
assign col_out_777 = {u_ca_out_777[18:0],u_ca_out_776[75:19], u_ca_out_775[132:76], u_ca_out_774[151:133]};
assign col_out_778 = {u_ca_out_778[18:0],u_ca_out_777[75:19], u_ca_out_776[132:76], u_ca_out_775[151:133]};
assign col_out_779 = {u_ca_out_779[18:0],u_ca_out_778[75:19], u_ca_out_777[132:76], u_ca_out_776[151:133]};
assign col_out_780 = {u_ca_out_780[18:0],u_ca_out_779[75:19], u_ca_out_778[132:76], u_ca_out_777[151:133]};
assign col_out_781 = {u_ca_out_781[18:0],u_ca_out_780[75:19], u_ca_out_779[132:76], u_ca_out_778[151:133]};
assign col_out_782 = {u_ca_out_782[18:0],u_ca_out_781[75:19], u_ca_out_780[132:76], u_ca_out_779[151:133]};
assign col_out_783 = {u_ca_out_783[18:0],u_ca_out_782[75:19], u_ca_out_781[132:76], u_ca_out_780[151:133]};
assign col_out_784 = {u_ca_out_784[18:0],u_ca_out_783[75:19], u_ca_out_782[132:76], u_ca_out_781[151:133]};
assign col_out_785 = {u_ca_out_785[18:0],u_ca_out_784[75:19], u_ca_out_783[132:76], u_ca_out_782[151:133]};
assign col_out_786 = {u_ca_out_786[18:0],u_ca_out_785[75:19], u_ca_out_784[132:76], u_ca_out_783[151:133]};
assign col_out_787 = {u_ca_out_787[18:0],u_ca_out_786[75:19], u_ca_out_785[132:76], u_ca_out_784[151:133]};
assign col_out_788 = {u_ca_out_788[18:0],u_ca_out_787[75:19], u_ca_out_786[132:76], u_ca_out_785[151:133]};
assign col_out_789 = {u_ca_out_789[18:0],u_ca_out_788[75:19], u_ca_out_787[132:76], u_ca_out_786[151:133]};
assign col_out_790 = {u_ca_out_790[18:0],u_ca_out_789[75:19], u_ca_out_788[132:76], u_ca_out_787[151:133]};
assign col_out_791 = {u_ca_out_791[18:0],u_ca_out_790[75:19], u_ca_out_789[132:76], u_ca_out_788[151:133]};
assign col_out_792 = {u_ca_out_792[18:0],u_ca_out_791[75:19], u_ca_out_790[132:76], u_ca_out_789[151:133]};
assign col_out_793 = {u_ca_out_793[18:0],u_ca_out_792[75:19], u_ca_out_791[132:76], u_ca_out_790[151:133]};
assign col_out_794 = {u_ca_out_794[18:0],u_ca_out_793[75:19], u_ca_out_792[132:76], u_ca_out_791[151:133]};
assign col_out_795 = {u_ca_out_795[18:0],u_ca_out_794[75:19], u_ca_out_793[132:76], u_ca_out_792[151:133]};
assign col_out_796 = {u_ca_out_796[18:0],u_ca_out_795[75:19], u_ca_out_794[132:76], u_ca_out_793[151:133]};
assign col_out_797 = {u_ca_out_797[18:0],u_ca_out_796[75:19], u_ca_out_795[132:76], u_ca_out_794[151:133]};
assign col_out_798 = {u_ca_out_798[18:0],u_ca_out_797[75:19], u_ca_out_796[132:76], u_ca_out_795[151:133]};
assign col_out_799 = {u_ca_out_799[18:0],u_ca_out_798[75:19], u_ca_out_797[132:76], u_ca_out_796[151:133]};
assign col_out_800 = {u_ca_out_800[18:0],u_ca_out_799[75:19], u_ca_out_798[132:76], u_ca_out_797[151:133]};
assign col_out_801 = {u_ca_out_801[18:0],u_ca_out_800[75:19], u_ca_out_799[132:76], u_ca_out_798[151:133]};
assign col_out_802 = {u_ca_out_802[18:0],u_ca_out_801[75:19], u_ca_out_800[132:76], u_ca_out_799[151:133]};
assign col_out_803 = {u_ca_out_803[18:0],u_ca_out_802[75:19], u_ca_out_801[132:76], u_ca_out_800[151:133]};
assign col_out_804 = {u_ca_out_804[18:0],u_ca_out_803[75:19], u_ca_out_802[132:76], u_ca_out_801[151:133]};
assign col_out_805 = {u_ca_out_805[18:0],u_ca_out_804[75:19], u_ca_out_803[132:76], u_ca_out_802[151:133]};
assign col_out_806 = {u_ca_out_806[18:0],u_ca_out_805[75:19], u_ca_out_804[132:76], u_ca_out_803[151:133]};
assign col_out_807 = {u_ca_out_807[18:0],u_ca_out_806[75:19], u_ca_out_805[132:76], u_ca_out_804[151:133]};
assign col_out_808 = {u_ca_out_808[18:0],u_ca_out_807[75:19], u_ca_out_806[132:76], u_ca_out_805[151:133]};
assign col_out_809 = {u_ca_out_809[18:0],u_ca_out_808[75:19], u_ca_out_807[132:76], u_ca_out_806[151:133]};
assign col_out_810 = {u_ca_out_810[18:0],u_ca_out_809[75:19], u_ca_out_808[132:76], u_ca_out_807[151:133]};
assign col_out_811 = {u_ca_out_811[18:0],u_ca_out_810[75:19], u_ca_out_809[132:76], u_ca_out_808[151:133]};
assign col_out_812 = {u_ca_out_812[18:0],u_ca_out_811[75:19], u_ca_out_810[132:76], u_ca_out_809[151:133]};
assign col_out_813 = {u_ca_out_813[18:0],u_ca_out_812[75:19], u_ca_out_811[132:76], u_ca_out_810[151:133]};
assign col_out_814 = {u_ca_out_814[18:0],u_ca_out_813[75:19], u_ca_out_812[132:76], u_ca_out_811[151:133]};
assign col_out_815 = {u_ca_out_815[18:0],u_ca_out_814[75:19], u_ca_out_813[132:76], u_ca_out_812[151:133]};
assign col_out_816 = {u_ca_out_816[18:0],u_ca_out_815[75:19], u_ca_out_814[132:76], u_ca_out_813[151:133]};
assign col_out_817 = {u_ca_out_817[18:0],u_ca_out_816[75:19], u_ca_out_815[132:76], u_ca_out_814[151:133]};
assign col_out_818 = {u_ca_out_818[18:0],u_ca_out_817[75:19], u_ca_out_816[132:76], u_ca_out_815[151:133]};
assign col_out_819 = {u_ca_out_819[18:0],u_ca_out_818[75:19], u_ca_out_817[132:76], u_ca_out_816[151:133]};
assign col_out_820 = {u_ca_out_820[18:0],u_ca_out_819[75:19], u_ca_out_818[132:76], u_ca_out_817[151:133]};
assign col_out_821 = {u_ca_out_821[18:0],u_ca_out_820[75:19], u_ca_out_819[132:76], u_ca_out_818[151:133]};
assign col_out_822 = {u_ca_out_822[18:0],u_ca_out_821[75:19], u_ca_out_820[132:76], u_ca_out_819[151:133]};
assign col_out_823 = {u_ca_out_823[18:0],u_ca_out_822[75:19], u_ca_out_821[132:76], u_ca_out_820[151:133]};
assign col_out_824 = {u_ca_out_824[18:0],u_ca_out_823[75:19], u_ca_out_822[132:76], u_ca_out_821[151:133]};
assign col_out_825 = {u_ca_out_825[18:0],u_ca_out_824[75:19], u_ca_out_823[132:76], u_ca_out_822[151:133]};
assign col_out_826 = {u_ca_out_826[18:0],u_ca_out_825[75:19], u_ca_out_824[132:76], u_ca_out_823[151:133]};
assign col_out_827 = {u_ca_out_827[18:0],u_ca_out_826[75:19], u_ca_out_825[132:76], u_ca_out_824[151:133]};
assign col_out_828 = {u_ca_out_828[18:0],u_ca_out_827[75:19], u_ca_out_826[132:76], u_ca_out_825[151:133]};
assign col_out_829 = {u_ca_out_829[18:0],u_ca_out_828[75:19], u_ca_out_827[132:76], u_ca_out_826[151:133]};
assign col_out_830 = {u_ca_out_830[18:0],u_ca_out_829[75:19], u_ca_out_828[132:76], u_ca_out_827[151:133]};
assign col_out_831 = {u_ca_out_831[18:0],u_ca_out_830[75:19], u_ca_out_829[132:76], u_ca_out_828[151:133]};
assign col_out_832 = {u_ca_out_832[18:0],u_ca_out_831[75:19], u_ca_out_830[132:76], u_ca_out_829[151:133]};
assign col_out_833 = {u_ca_out_833[18:0],u_ca_out_832[75:19], u_ca_out_831[132:76], u_ca_out_830[151:133]};
assign col_out_834 = {u_ca_out_834[18:0],u_ca_out_833[75:19], u_ca_out_832[132:76], u_ca_out_831[151:133]};
assign col_out_835 = {u_ca_out_835[18:0],u_ca_out_834[75:19], u_ca_out_833[132:76], u_ca_out_832[151:133]};
assign col_out_836 = {u_ca_out_836[18:0],u_ca_out_835[75:19], u_ca_out_834[132:76], u_ca_out_833[151:133]};
assign col_out_837 = {u_ca_out_837[18:0],u_ca_out_836[75:19], u_ca_out_835[132:76], u_ca_out_834[151:133]};
assign col_out_838 = {u_ca_out_838[18:0],u_ca_out_837[75:19], u_ca_out_836[132:76], u_ca_out_835[151:133]};
assign col_out_839 = {u_ca_out_839[18:0],u_ca_out_838[75:19], u_ca_out_837[132:76], u_ca_out_836[151:133]};
assign col_out_840 = {u_ca_out_840[18:0],u_ca_out_839[75:19], u_ca_out_838[132:76], u_ca_out_837[151:133]};
assign col_out_841 = {u_ca_out_841[18:0],u_ca_out_840[75:19], u_ca_out_839[132:76], u_ca_out_838[151:133]};
assign col_out_842 = {u_ca_out_842[18:0],u_ca_out_841[75:19], u_ca_out_840[132:76], u_ca_out_839[151:133]};
assign col_out_843 = {u_ca_out_843[18:0],u_ca_out_842[75:19], u_ca_out_841[132:76], u_ca_out_840[151:133]};
assign col_out_844 = {u_ca_out_844[18:0],u_ca_out_843[75:19], u_ca_out_842[132:76], u_ca_out_841[151:133]};
assign col_out_845 = {u_ca_out_845[18:0],u_ca_out_844[75:19], u_ca_out_843[132:76], u_ca_out_842[151:133]};
assign col_out_846 = {u_ca_out_846[18:0],u_ca_out_845[75:19], u_ca_out_844[132:76], u_ca_out_843[151:133]};
assign col_out_847 = {u_ca_out_847[18:0],u_ca_out_846[75:19], u_ca_out_845[132:76], u_ca_out_844[151:133]};
assign col_out_848 = {u_ca_out_848[18:0],u_ca_out_847[75:19], u_ca_out_846[132:76], u_ca_out_845[151:133]};
assign col_out_849 = {u_ca_out_849[18:0],u_ca_out_848[75:19], u_ca_out_847[132:76], u_ca_out_846[151:133]};
assign col_out_850 = {u_ca_out_850[18:0],u_ca_out_849[75:19], u_ca_out_848[132:76], u_ca_out_847[151:133]};
assign col_out_851 = {u_ca_out_851[18:0],u_ca_out_850[75:19], u_ca_out_849[132:76], u_ca_out_848[151:133]};
assign col_out_852 = {u_ca_out_852[18:0],u_ca_out_851[75:19], u_ca_out_850[132:76], u_ca_out_849[151:133]};
assign col_out_853 = {u_ca_out_853[18:0],u_ca_out_852[75:19], u_ca_out_851[132:76], u_ca_out_850[151:133]};
assign col_out_854 = {u_ca_out_854[18:0],u_ca_out_853[75:19], u_ca_out_852[132:76], u_ca_out_851[151:133]};
assign col_out_855 = {u_ca_out_855[18:0],u_ca_out_854[75:19], u_ca_out_853[132:76], u_ca_out_852[151:133]};
assign col_out_856 = {u_ca_out_856[18:0],u_ca_out_855[75:19], u_ca_out_854[132:76], u_ca_out_853[151:133]};
assign col_out_857 = {u_ca_out_857[18:0],u_ca_out_856[75:19], u_ca_out_855[132:76], u_ca_out_854[151:133]};
assign col_out_858 = {u_ca_out_858[18:0],u_ca_out_857[75:19], u_ca_out_856[132:76], u_ca_out_855[151:133]};
assign col_out_859 = {u_ca_out_859[18:0],u_ca_out_858[75:19], u_ca_out_857[132:76], u_ca_out_856[151:133]};
assign col_out_860 = {u_ca_out_860[18:0],u_ca_out_859[75:19], u_ca_out_858[132:76], u_ca_out_857[151:133]};
assign col_out_861 = {u_ca_out_861[18:0],u_ca_out_860[75:19], u_ca_out_859[132:76], u_ca_out_858[151:133]};
assign col_out_862 = {u_ca_out_862[18:0],u_ca_out_861[75:19], u_ca_out_860[132:76], u_ca_out_859[151:133]};
assign col_out_863 = {u_ca_out_863[18:0],u_ca_out_862[75:19], u_ca_out_861[132:76], u_ca_out_860[151:133]};
assign col_out_864 = {u_ca_out_864[18:0],u_ca_out_863[75:19], u_ca_out_862[132:76], u_ca_out_861[151:133]};
assign col_out_865 = {u_ca_out_865[18:0],u_ca_out_864[75:19], u_ca_out_863[132:76], u_ca_out_862[151:133]};
assign col_out_866 = {u_ca_out_866[18:0],u_ca_out_865[75:19], u_ca_out_864[132:76], u_ca_out_863[151:133]};
assign col_out_867 = {u_ca_out_867[18:0],u_ca_out_866[75:19], u_ca_out_865[132:76], u_ca_out_864[151:133]};
assign col_out_868 = {u_ca_out_868[18:0],u_ca_out_867[75:19], u_ca_out_866[132:76], u_ca_out_865[151:133]};
assign col_out_869 = {u_ca_out_869[18:0],u_ca_out_868[75:19], u_ca_out_867[132:76], u_ca_out_866[151:133]};
assign col_out_870 = {u_ca_out_870[18:0],u_ca_out_869[75:19], u_ca_out_868[132:76], u_ca_out_867[151:133]};
assign col_out_871 = {u_ca_out_871[18:0],u_ca_out_870[75:19], u_ca_out_869[132:76], u_ca_out_868[151:133]};
assign col_out_872 = {u_ca_out_872[18:0],u_ca_out_871[75:19], u_ca_out_870[132:76], u_ca_out_869[151:133]};
assign col_out_873 = {u_ca_out_873[18:0],u_ca_out_872[75:19], u_ca_out_871[132:76], u_ca_out_870[151:133]};
assign col_out_874 = {u_ca_out_874[18:0],u_ca_out_873[75:19], u_ca_out_872[132:76], u_ca_out_871[151:133]};
assign col_out_875 = {u_ca_out_875[18:0],u_ca_out_874[75:19], u_ca_out_873[132:76], u_ca_out_872[151:133]};
assign col_out_876 = {u_ca_out_876[18:0],u_ca_out_875[75:19], u_ca_out_874[132:76], u_ca_out_873[151:133]};
assign col_out_877 = {u_ca_out_877[18:0],u_ca_out_876[75:19], u_ca_out_875[132:76], u_ca_out_874[151:133]};
assign col_out_878 = {u_ca_out_878[18:0],u_ca_out_877[75:19], u_ca_out_876[132:76], u_ca_out_875[151:133]};
assign col_out_879 = {u_ca_out_879[18:0],u_ca_out_878[75:19], u_ca_out_877[132:76], u_ca_out_876[151:133]};
assign col_out_880 = {u_ca_out_880[18:0],u_ca_out_879[75:19], u_ca_out_878[132:76], u_ca_out_877[151:133]};
assign col_out_881 = {u_ca_out_881[18:0],u_ca_out_880[75:19], u_ca_out_879[132:76], u_ca_out_878[151:133]};
assign col_out_882 = {u_ca_out_882[18:0],u_ca_out_881[75:19], u_ca_out_880[132:76], u_ca_out_879[151:133]};
assign col_out_883 = {u_ca_out_883[18:0],u_ca_out_882[75:19], u_ca_out_881[132:76], u_ca_out_880[151:133]};
assign col_out_884 = {u_ca_out_884[18:0],u_ca_out_883[75:19], u_ca_out_882[132:76], u_ca_out_881[151:133]};
assign col_out_885 = {u_ca_out_885[18:0],u_ca_out_884[75:19], u_ca_out_883[132:76], u_ca_out_882[151:133]};
assign col_out_886 = {u_ca_out_886[18:0],u_ca_out_885[75:19], u_ca_out_884[132:76], u_ca_out_883[151:133]};
assign col_out_887 = {u_ca_out_887[18:0],u_ca_out_886[75:19], u_ca_out_885[132:76], u_ca_out_884[151:133]};
assign col_out_888 = {u_ca_out_888[18:0],u_ca_out_887[75:19], u_ca_out_886[132:76], u_ca_out_885[151:133]};
assign col_out_889 = {u_ca_out_889[18:0],u_ca_out_888[75:19], u_ca_out_887[132:76], u_ca_out_886[151:133]};
assign col_out_890 = {u_ca_out_890[18:0],u_ca_out_889[75:19], u_ca_out_888[132:76], u_ca_out_887[151:133]};
assign col_out_891 = {u_ca_out_891[18:0],u_ca_out_890[75:19], u_ca_out_889[132:76], u_ca_out_888[151:133]};
assign col_out_892 = {u_ca_out_892[18:0],u_ca_out_891[75:19], u_ca_out_890[132:76], u_ca_out_889[151:133]};
assign col_out_893 = {u_ca_out_893[18:0],u_ca_out_892[75:19], u_ca_out_891[132:76], u_ca_out_890[151:133]};
assign col_out_894 = {u_ca_out_894[18:0],u_ca_out_893[75:19], u_ca_out_892[132:76], u_ca_out_891[151:133]};
assign col_out_895 = {u_ca_out_895[18:0],u_ca_out_894[75:19], u_ca_out_893[132:76], u_ca_out_892[151:133]};
assign col_out_896 = {u_ca_out_896[18:0],u_ca_out_895[75:19], u_ca_out_894[132:76], u_ca_out_893[151:133]};
assign col_out_897 = {u_ca_out_897[18:0],u_ca_out_896[75:19], u_ca_out_895[132:76], u_ca_out_894[151:133]};
assign col_out_898 = {u_ca_out_898[18:0],u_ca_out_897[75:19], u_ca_out_896[132:76], u_ca_out_895[151:133]};
assign col_out_899 = {u_ca_out_899[18:0],u_ca_out_898[75:19], u_ca_out_897[132:76], u_ca_out_896[151:133]};
assign col_out_900 = {u_ca_out_900[18:0],u_ca_out_899[75:19], u_ca_out_898[132:76], u_ca_out_897[151:133]};
assign col_out_901 = {u_ca_out_901[18:0],u_ca_out_900[75:19], u_ca_out_899[132:76], u_ca_out_898[151:133]};
assign col_out_902 = {u_ca_out_902[18:0],u_ca_out_901[75:19], u_ca_out_900[132:76], u_ca_out_899[151:133]};
assign col_out_903 = {u_ca_out_903[18:0],u_ca_out_902[75:19], u_ca_out_901[132:76], u_ca_out_900[151:133]};
assign col_out_904 = {u_ca_out_904[18:0],u_ca_out_903[75:19], u_ca_out_902[132:76], u_ca_out_901[151:133]};
assign col_out_905 = {u_ca_out_905[18:0],u_ca_out_904[75:19], u_ca_out_903[132:76], u_ca_out_902[151:133]};
assign col_out_906 = {u_ca_out_906[18:0],u_ca_out_905[75:19], u_ca_out_904[132:76], u_ca_out_903[151:133]};
assign col_out_907 = {u_ca_out_907[18:0],u_ca_out_906[75:19], u_ca_out_905[132:76], u_ca_out_904[151:133]};
assign col_out_908 = {u_ca_out_908[18:0],u_ca_out_907[75:19], u_ca_out_906[132:76], u_ca_out_905[151:133]};
assign col_out_909 = {u_ca_out_909[18:0],u_ca_out_908[75:19], u_ca_out_907[132:76], u_ca_out_906[151:133]};
assign col_out_910 = {u_ca_out_910[18:0],u_ca_out_909[75:19], u_ca_out_908[132:76], u_ca_out_907[151:133]};
assign col_out_911 = {u_ca_out_911[18:0],u_ca_out_910[75:19], u_ca_out_909[132:76], u_ca_out_908[151:133]};
assign col_out_912 = {u_ca_out_912[18:0],u_ca_out_911[75:19], u_ca_out_910[132:76], u_ca_out_909[151:133]};
assign col_out_913 = {u_ca_out_913[18:0],u_ca_out_912[75:19], u_ca_out_911[132:76], u_ca_out_910[151:133]};
assign col_out_914 = {u_ca_out_914[18:0],u_ca_out_913[75:19], u_ca_out_912[132:76], u_ca_out_911[151:133]};
assign col_out_915 = {u_ca_out_915[18:0],u_ca_out_914[75:19], u_ca_out_913[132:76], u_ca_out_912[151:133]};
assign col_out_916 = {u_ca_out_916[18:0],u_ca_out_915[75:19], u_ca_out_914[132:76], u_ca_out_913[151:133]};
assign col_out_917 = {u_ca_out_917[18:0],u_ca_out_916[75:19], u_ca_out_915[132:76], u_ca_out_914[151:133]};
assign col_out_918 = {u_ca_out_918[18:0],u_ca_out_917[75:19], u_ca_out_916[132:76], u_ca_out_915[151:133]};
assign col_out_919 = {u_ca_out_919[18:0],u_ca_out_918[75:19], u_ca_out_917[132:76], u_ca_out_916[151:133]};
assign col_out_920 = {u_ca_out_920[18:0],u_ca_out_919[75:19], u_ca_out_918[132:76], u_ca_out_917[151:133]};
assign col_out_921 = {u_ca_out_921[18:0],u_ca_out_920[75:19], u_ca_out_919[132:76], u_ca_out_918[151:133]};
assign col_out_922 = {u_ca_out_922[18:0],u_ca_out_921[75:19], u_ca_out_920[132:76], u_ca_out_919[151:133]};
assign col_out_923 = {u_ca_out_923[18:0],u_ca_out_922[75:19], u_ca_out_921[132:76], u_ca_out_920[151:133]};
assign col_out_924 = {u_ca_out_924[18:0],u_ca_out_923[75:19], u_ca_out_922[132:76], u_ca_out_921[151:133]};
assign col_out_925 = {u_ca_out_925[18:0],u_ca_out_924[75:19], u_ca_out_923[132:76], u_ca_out_922[151:133]};
assign col_out_926 = {u_ca_out_926[18:0],u_ca_out_925[75:19], u_ca_out_924[132:76], u_ca_out_923[151:133]};
assign col_out_927 = {u_ca_out_927[18:0],u_ca_out_926[75:19], u_ca_out_925[132:76], u_ca_out_924[151:133]};
assign col_out_928 = {u_ca_out_928[18:0],u_ca_out_927[75:19], u_ca_out_926[132:76], u_ca_out_925[151:133]};
assign col_out_929 = {u_ca_out_929[18:0],u_ca_out_928[75:19], u_ca_out_927[132:76], u_ca_out_926[151:133]};
assign col_out_930 = {u_ca_out_930[18:0],u_ca_out_929[75:19], u_ca_out_928[132:76], u_ca_out_927[151:133]};
assign col_out_931 = {u_ca_out_931[18:0],u_ca_out_930[75:19], u_ca_out_929[132:76], u_ca_out_928[151:133]};
assign col_out_932 = {u_ca_out_932[18:0],u_ca_out_931[75:19], u_ca_out_930[132:76], u_ca_out_929[151:133]};
assign col_out_933 = {u_ca_out_933[18:0],u_ca_out_932[75:19], u_ca_out_931[132:76], u_ca_out_930[151:133]};
assign col_out_934 = {u_ca_out_934[18:0],u_ca_out_933[75:19], u_ca_out_932[132:76], u_ca_out_931[151:133]};
assign col_out_935 = {u_ca_out_935[18:0],u_ca_out_934[75:19], u_ca_out_933[132:76], u_ca_out_932[151:133]};
assign col_out_936 = {u_ca_out_936[18:0],u_ca_out_935[75:19], u_ca_out_934[132:76], u_ca_out_933[151:133]};
assign col_out_937 = {u_ca_out_937[18:0],u_ca_out_936[75:19], u_ca_out_935[132:76], u_ca_out_934[151:133]};
assign col_out_938 = {u_ca_out_938[18:0],u_ca_out_937[75:19], u_ca_out_936[132:76], u_ca_out_935[151:133]};
assign col_out_939 = {u_ca_out_939[18:0],u_ca_out_938[75:19], u_ca_out_937[132:76], u_ca_out_936[151:133]};
assign col_out_940 = {u_ca_out_940[18:0],u_ca_out_939[75:19], u_ca_out_938[132:76], u_ca_out_937[151:133]};
assign col_out_941 = {u_ca_out_941[18:0],u_ca_out_940[75:19], u_ca_out_939[132:76], u_ca_out_938[151:133]};
assign col_out_942 = {u_ca_out_942[18:0],u_ca_out_941[75:19], u_ca_out_940[132:76], u_ca_out_939[151:133]};
assign col_out_943 = {u_ca_out_943[18:0],u_ca_out_942[75:19], u_ca_out_941[132:76], u_ca_out_940[151:133]};
assign col_out_944 = {u_ca_out_944[18:0],u_ca_out_943[75:19], u_ca_out_942[132:76], u_ca_out_941[151:133]};
assign col_out_945 = {u_ca_out_945[18:0],u_ca_out_944[75:19], u_ca_out_943[132:76], u_ca_out_942[151:133]};
assign col_out_946 = {u_ca_out_946[18:0],u_ca_out_945[75:19], u_ca_out_944[132:76], u_ca_out_943[151:133]};
assign col_out_947 = {u_ca_out_947[18:0],u_ca_out_946[75:19], u_ca_out_945[132:76], u_ca_out_944[151:133]};
assign col_out_948 = {u_ca_out_948[18:0],u_ca_out_947[75:19], u_ca_out_946[132:76], u_ca_out_945[151:133]};
assign col_out_949 = {u_ca_out_949[18:0],u_ca_out_948[75:19], u_ca_out_947[132:76], u_ca_out_946[151:133]};
assign col_out_950 = {u_ca_out_950[18:0],u_ca_out_949[75:19], u_ca_out_948[132:76], u_ca_out_947[151:133]};
assign col_out_951 = {u_ca_out_951[18:0],u_ca_out_950[75:19], u_ca_out_949[132:76], u_ca_out_948[151:133]};
assign col_out_952 = {u_ca_out_952[18:0],u_ca_out_951[75:19], u_ca_out_950[132:76], u_ca_out_949[151:133]};
assign col_out_953 = {u_ca_out_953[18:0],u_ca_out_952[75:19], u_ca_out_951[132:76], u_ca_out_950[151:133]};
assign col_out_954 = {u_ca_out_954[18:0],u_ca_out_953[75:19], u_ca_out_952[132:76], u_ca_out_951[151:133]};
assign col_out_955 = {u_ca_out_955[18:0],u_ca_out_954[75:19], u_ca_out_953[132:76], u_ca_out_952[151:133]};
assign col_out_956 = {u_ca_out_956[18:0],u_ca_out_955[75:19], u_ca_out_954[132:76], u_ca_out_953[151:133]};
assign col_out_957 = {u_ca_out_957[18:0],u_ca_out_956[75:19], u_ca_out_955[132:76], u_ca_out_954[151:133]};
assign col_out_958 = {u_ca_out_958[18:0],u_ca_out_957[75:19], u_ca_out_956[132:76], u_ca_out_955[151:133]};
assign col_out_959 = {u_ca_out_959[18:0],u_ca_out_958[75:19], u_ca_out_957[132:76], u_ca_out_956[151:133]};
assign col_out_960 = {u_ca_out_960[18:0],u_ca_out_959[75:19], u_ca_out_958[132:76], u_ca_out_957[151:133]};
assign col_out_961 = {u_ca_out_961[18:0],u_ca_out_960[75:19], u_ca_out_959[132:76], u_ca_out_958[151:133]};
assign col_out_962 = {u_ca_out_962[18:0],u_ca_out_961[75:19], u_ca_out_960[132:76], u_ca_out_959[151:133]};
assign col_out_963 = {u_ca_out_963[18:0],u_ca_out_962[75:19], u_ca_out_961[132:76], u_ca_out_960[151:133]};
assign col_out_964 = {u_ca_out_964[18:0],u_ca_out_963[75:19], u_ca_out_962[132:76], u_ca_out_961[151:133]};
assign col_out_965 = {u_ca_out_965[18:0],u_ca_out_964[75:19], u_ca_out_963[132:76], u_ca_out_962[151:133]};
assign col_out_966 = {u_ca_out_966[18:0],u_ca_out_965[75:19], u_ca_out_964[132:76], u_ca_out_963[151:133]};
assign col_out_967 = {u_ca_out_967[18:0],u_ca_out_966[75:19], u_ca_out_965[132:76], u_ca_out_964[151:133]};
assign col_out_968 = {u_ca_out_968[18:0],u_ca_out_967[75:19], u_ca_out_966[132:76], u_ca_out_965[151:133]};
assign col_out_969 = {u_ca_out_969[18:0],u_ca_out_968[75:19], u_ca_out_967[132:76], u_ca_out_966[151:133]};
assign col_out_970 = {u_ca_out_970[18:0],u_ca_out_969[75:19], u_ca_out_968[132:76], u_ca_out_967[151:133]};
assign col_out_971 = {u_ca_out_971[18:0],u_ca_out_970[75:19], u_ca_out_969[132:76], u_ca_out_968[151:133]};
assign col_out_972 = {u_ca_out_972[18:0],u_ca_out_971[75:19], u_ca_out_970[132:76], u_ca_out_969[151:133]};
assign col_out_973 = {u_ca_out_973[18:0],u_ca_out_972[75:19], u_ca_out_971[132:76], u_ca_out_970[151:133]};
assign col_out_974 = {u_ca_out_974[18:0],u_ca_out_973[75:19], u_ca_out_972[132:76], u_ca_out_971[151:133]};
assign col_out_975 = {u_ca_out_975[18:0],u_ca_out_974[75:19], u_ca_out_973[132:76], u_ca_out_972[151:133]};
assign col_out_976 = {u_ca_out_976[18:0],u_ca_out_975[75:19], u_ca_out_974[132:76], u_ca_out_973[151:133]};
assign col_out_977 = {u_ca_out_977[18:0],u_ca_out_976[75:19], u_ca_out_975[132:76], u_ca_out_974[151:133]};
assign col_out_978 = {u_ca_out_978[18:0],u_ca_out_977[75:19], u_ca_out_976[132:76], u_ca_out_975[151:133]};
assign col_out_979 = {u_ca_out_979[18:0],u_ca_out_978[75:19], u_ca_out_977[132:76], u_ca_out_976[151:133]};
assign col_out_980 = {u_ca_out_980[18:0],u_ca_out_979[75:19], u_ca_out_978[132:76], u_ca_out_977[151:133]};
assign col_out_981 = {u_ca_out_981[18:0],u_ca_out_980[75:19], u_ca_out_979[132:76], u_ca_out_978[151:133]};
assign col_out_982 = {u_ca_out_982[18:0],u_ca_out_981[75:19], u_ca_out_980[132:76], u_ca_out_979[151:133]};
assign col_out_983 = {u_ca_out_983[18:0],u_ca_out_982[75:19], u_ca_out_981[132:76], u_ca_out_980[151:133]};
assign col_out_984 = {u_ca_out_984[18:0],u_ca_out_983[75:19], u_ca_out_982[132:76], u_ca_out_981[151:133]};
assign col_out_985 = {u_ca_out_985[18:0],u_ca_out_984[75:19], u_ca_out_983[132:76], u_ca_out_982[151:133]};
assign col_out_986 = {u_ca_out_986[18:0],u_ca_out_985[75:19], u_ca_out_984[132:76], u_ca_out_983[151:133]};
assign col_out_987 = {u_ca_out_987[18:0],u_ca_out_986[75:19], u_ca_out_985[132:76], u_ca_out_984[151:133]};
assign col_out_988 = {u_ca_out_988[18:0],u_ca_out_987[75:19], u_ca_out_986[132:76], u_ca_out_985[151:133]};
assign col_out_989 = {u_ca_out_989[18:0],u_ca_out_988[75:19], u_ca_out_987[132:76], u_ca_out_986[151:133]};
assign col_out_990 = {u_ca_out_990[18:0],u_ca_out_989[75:19], u_ca_out_988[132:76], u_ca_out_987[151:133]};
assign col_out_991 = {u_ca_out_991[18:0],u_ca_out_990[75:19], u_ca_out_989[132:76], u_ca_out_988[151:133]};
assign col_out_992 = {u_ca_out_992[18:0],u_ca_out_991[75:19], u_ca_out_990[132:76], u_ca_out_989[151:133]};
assign col_out_993 = {u_ca_out_993[18:0],u_ca_out_992[75:19], u_ca_out_991[132:76], u_ca_out_990[151:133]};
assign col_out_994 = {u_ca_out_994[18:0],u_ca_out_993[75:19], u_ca_out_992[132:76], u_ca_out_991[151:133]};
assign col_out_995 = {u_ca_out_995[18:0],u_ca_out_994[75:19], u_ca_out_993[132:76], u_ca_out_992[151:133]};
assign col_out_996 = {u_ca_out_996[18:0],u_ca_out_995[75:19], u_ca_out_994[132:76], u_ca_out_993[151:133]};
assign col_out_997 = {u_ca_out_997[18:0],u_ca_out_996[75:19], u_ca_out_995[132:76], u_ca_out_994[151:133]};
assign col_out_998 = {u_ca_out_998[18:0],u_ca_out_997[75:19], u_ca_out_996[132:76], u_ca_out_995[151:133]};
assign col_out_999 = {u_ca_out_999[18:0],u_ca_out_998[75:19], u_ca_out_997[132:76], u_ca_out_996[151:133]};
assign col_out_1000 = {u_ca_out_1000[18:0],u_ca_out_999[75:19], u_ca_out_998[132:76], u_ca_out_997[151:133]};
assign col_out_1001 = {u_ca_out_1001[18:0],u_ca_out_1000[75:19], u_ca_out_999[132:76], u_ca_out_998[151:133]};
assign col_out_1002 = {u_ca_out_1002[18:0],u_ca_out_1001[75:19], u_ca_out_1000[132:76], u_ca_out_999[151:133]};
assign col_out_1003 = {u_ca_out_1003[18:0],u_ca_out_1002[75:19], u_ca_out_1001[132:76], u_ca_out_1000[151:133]};
assign col_out_1004 = {u_ca_out_1004[18:0],u_ca_out_1003[75:19], u_ca_out_1002[132:76], u_ca_out_1001[151:133]};
assign col_out_1005 = {u_ca_out_1005[18:0],u_ca_out_1004[75:19], u_ca_out_1003[132:76], u_ca_out_1002[151:133]};
assign col_out_1006 = {u_ca_out_1006[18:0],u_ca_out_1005[75:19], u_ca_out_1004[132:76], u_ca_out_1003[151:133]};
assign col_out_1007 = {u_ca_out_1007[18:0],u_ca_out_1006[75:19], u_ca_out_1005[132:76], u_ca_out_1004[151:133]};
assign col_out_1008 = {u_ca_out_1008[18:0],u_ca_out_1007[75:19], u_ca_out_1006[132:76], u_ca_out_1005[151:133]};
assign col_out_1009 = {u_ca_out_1009[18:0],u_ca_out_1008[75:19], u_ca_out_1007[132:76], u_ca_out_1006[151:133]};
assign col_out_1010 = {u_ca_out_1010[18:0],u_ca_out_1009[75:19], u_ca_out_1008[132:76], u_ca_out_1007[151:133]};
assign col_out_1011 = {u_ca_out_1011[18:0],u_ca_out_1010[75:19], u_ca_out_1009[132:76], u_ca_out_1008[151:133]};
assign col_out_1012 = {u_ca_out_1012[18:0],u_ca_out_1011[75:19], u_ca_out_1010[132:76], u_ca_out_1009[151:133]};
assign col_out_1013 = {u_ca_out_1013[18:0],u_ca_out_1012[75:19], u_ca_out_1011[132:76], u_ca_out_1010[151:133]};
assign col_out_1014 = {u_ca_out_1014[18:0],u_ca_out_1013[75:19], u_ca_out_1012[132:76], u_ca_out_1011[151:133]};
assign col_out_1015 = {u_ca_out_1015[18:0],u_ca_out_1014[75:19], u_ca_out_1013[132:76], u_ca_out_1012[151:133]};
assign col_out_1016 = {u_ca_out_1016[18:0],u_ca_out_1015[75:19], u_ca_out_1014[132:76], u_ca_out_1013[151:133]};
assign col_out_1017 = {u_ca_out_1017[18:0],u_ca_out_1016[75:19], u_ca_out_1015[132:76], u_ca_out_1014[151:133]};
assign col_out_1018 = {u_ca_out_1018[18:0],u_ca_out_1017[75:19], u_ca_out_1016[132:76], u_ca_out_1015[151:133]};
assign col_out_1019 = {u_ca_out_1019[18:0],u_ca_out_1018[75:19], u_ca_out_1017[132:76], u_ca_out_1016[151:133]};
assign col_out_1020 = {u_ca_out_1020[18:0],u_ca_out_1019[75:19], u_ca_out_1018[132:76], u_ca_out_1017[151:133]};
assign col_out_1021 = {u_ca_out_1021[18:0],u_ca_out_1020[75:19], u_ca_out_1019[132:76], u_ca_out_1018[151:133]};
assign col_out_1022 = {u_ca_out_1022[18:0],u_ca_out_1021[75:19], u_ca_out_1020[132:76], u_ca_out_1019[151:133]};
assign col_out_1023 = {u_ca_out_1023[18:0],u_ca_out_1022[75:19], u_ca_out_1021[132:76], u_ca_out_1020[151:133]};
assign col_out_1024 = {{19{1'b0}}, u_ca_out_1023[75:19], u_ca_out_1022[132:76], u_ca_out_1021[151:133]};
assign col_out_1025 = {{76{1'b0}}, u_ca_out_1023[132:76], u_ca_out_1022[151:133]};
assign col_out_1026 = {{133{1'b0}}, u_ca_out_1023[151:133]};

//---------------------------------------------------------


endmodule
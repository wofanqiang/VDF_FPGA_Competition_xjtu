module xpb_5_300
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h49ffe5270b2843e57efc7ec13f77c0fc6156a2a8c05ab2f30ecb879d609a88371807df76a545520a12377a5451c1457da68dfd351f0143a8808c0a9fe8f0baae55b4a9a7d21d716c6208c7758c6c65229bd6711b39024b847c4a75abb8601abef52661a66e5d01fb14e96b50bd72c683e1f4b12c40aa315f357e95215e151282;
    5'b00010 : xpb = 1024'h93ffca4e165087cafdf8fd827eef81f8c2ad455180b565e61d970f3ac135106e300fbeed4a8aa414246ef4a8a3828afb4d1bfa6a3e0287510118153fd1e1755cab69534fa43ae2d8c4118eeb18d8ca4537ace23672049708f894eb5770c0357dea4cc34cdcba03f629d2d6a17ae58d07c3e96258815462be6afd2a42bc2a2504;
    5'b00011 : xpb = 1024'h2d526a1f5f8a96e7b1f0046cae0cfba3b28de4c96b987861ae85dd826ecceb9d44cf20eb25a9778f97482fb611e5bfae8f8fcfb93a50faadd104e0817fffbb598ccec848c6c75700138053be0c696b36df7e59b91e80b57cbf52cf086ef5adaab06b92c99a4e0d63b7fc5b1340882d62570434a271b336ed5a0c445f915cd11b;
    5'b00100 : xpb = 1024'h77524f466ab2dacd30ec832ded84bca013e487722bf32b54bd51651fcf6773d45cd70061caeec999a97faa0a63a7052c361dccee59523e565190eb2168f07607e28371f098e4c86c75891b3398d5d0597b54cad4578301013b9d44b42755c869a591f47008ab0f5ecce5c663fdfaf3e638f8e5ceb25d684c8f8ad980ef71e39d;
    5'b00101 : xpb = 1024'h10a4ef17b3ece9e9e4e38a181ca2364b03c526ea16d63dd04e4033677cff4f037196625fa60d9d151c58e517d20a39df7891a23d55a0b1b3217db663170ebc04c3e8e6e9bb713c93c4f7e0068c66714b2326425703ff1f75025b2865258b40966bb0c3ecc63f18cc5b0f4ad5c39d9440cc13b818a2bc3c7b7e99f39dc4a48fb4;
    5'b00110 : xpb = 1024'h5aa4d43ebf152dcf63e008d95c19f747651bc992d730f0c35d0bbb04dd99d73a899e41d64b52ef1f2e905f6c23cb7f5d1f1f9f7274a1f55ba209c102ffff76b3199d90918d8eae002700a77c18d2d66dbefcb3723d016af97ea59e10ddeb5b5560d72593349c1ac76ff8b62681105ac4ae086944e3666ddab41888bf22b9a236;
    5'b00111 : xpb = 1024'ha4a4b965ca3d71b4e2dc879a9b91b843c6726c3b978ba3b66bd742a23e345f71a1a6214cf098412940c7d9c0758cc4dac5ad9ca793a339042295cba2e8f031616f523a395fac1f6c89096ef1a53f3b905ad3248d7603b67dfaf013bc964b761455fd8739a2f91cc284e221773e8321488ffd1a7124109f39e9971de080ceb4b8;
    5'b01000 : xpb = 1024'h3df75937137780d196d38e84caaf31eeb6530bb3826eb631fcc610e9ebcc3aa0b665834acbb714a4b3a114cde3eff98e082171f68ff1ac60f28296e4970e775e50b7af3282389393d87833c498cfdc8202a49c10227fd4f1c1adf76d9480ee411c1c56b6608d2630130ba5e90425c1a32317ecbb146f7368d8a637fd560160cf;
    5'b01001 : xpb = 1024'h87f73e5e1e9fc4b715d00d460a26f2eb17a9ae5c42c969250b9198874c66c2d7ce6d62c170fc66aec5d88f2235b13f0baeaf6f2baef2f009730ea1847fff320ca66c58da545605003a80fb3a253c41a49e7b0d2b5b8220763df86d194ce109001142b85cceea282b27f51139c1988827050c9de75519a4c80e24cd1eb4167351;
    5'b01010 : xpb = 1024'h2149de2f67d9d3d3c9c7143039446c96078a4dd42dac7ba09c8066cef9fe9e06e32cc4bf4c1b3a2a38b1ca2fa41473bef123447aab41636642fb6cc62e1d780987d1cdd376e2792789efc00d18cce296464c84ae07fe3eea04b650ca4b16812cd76187d98c7e3198b61e95ab873b288198277031457878f6fd33e73b89491f68;
    5'b01011 : xpb = 1024'h6b49c356730217b948c392f178bc2d9268e0f07cee072e93ab4bee6c5a99263dfb34a435f1608c344ae94483f5d5b93c97b141afca42a70ec3877766170e32b7dd86777b48ffea93ebf88782a53947b8e222f5c941008a6e8100c67603769bebcc87e97ffadb3393cb0800fc44adef057a1c215d8622aa5632b27c5ce75e31ea;
    5'b01100 : xpb = 1024'h49c6327bc3c26d5fcba99dba7d9a73d58c18ff4d8ea410f3c3abcb40831016d0ff40633cc7f5fafbdc27f916438edefda2516fec6911a6b937442a7c52c78b4beebec746b8c5ebb3b674c5598c9e8aa89f46d4bed7ca8e247beaa2701ac141892a6b8fcb86f3d015931856e0a508f600d36f3a776817e8521c19679bc90de01;
    5'b01101 : xpb = 1024'h4e9c484ec7646abb7bb7189ce7516839ba18329d9944f4024b06445168cb89a427fbe5aa71c4b1b9cff9f9e5b5fa336d80b31433e5925e1414004d47ae1d336314a0961c3da9d0279d7013cb25364dcd25cade67267ef466c4091fd2ba0c2ed787cd1aa326cc3efc6e1af0bec7c355e3ef2ba4d3b72bafe457402b9b1aa5f083;
    5'b01110 : xpb = 1024'h989c2d75d28caea0fab3975e26c929361b6ed546599fa6f559d1cbeec96611db4003c521170a03c3e231743a07bb78eb274111690493a1bc948c57e7970dee116a553fc40fc74193ff78db40b1a2b2efc1a14f825f813feb4053957e726c49967cf37c49952940f783045c0f85361c67d12055fff7d5e1438cbec0bc78bb0305;
    5'b01111 : xpb = 1024'h31eecd471bc6bdbdaeaa9e4855e6a2e10b4f74be4482b970eac09a3676fded0a54c3271ef228d73f550aaf47761ead9e69b4e6b800e2151964792329452c340e4bbab4bd3253b5bb4ee7a013a53353e16972c7050bfd5e5f0711792f70a1c1c343124bc652bd4a65112de0814ad8bcc2643b2849e834b5727bcddad94dedaf1c;
    5'b10000 : xpb = 1024'h7beeb26e26ef01a32da71d09955e63dd6ca6176704dd6c63f98c21d3d79875416ccb0695976e29496742299bc7dff31c1042e3ed1fe358c1e5052dc92e1ceebca16f5e6504712727b0f06789319fb9040549382044ffa9e3835beedb2901dc823838ad6cc11a4c6026174bd2084b8346462fd97628dee6d1b14c6ffaac02c19e;
    5'b10001 : xpb = 1024'h1541523f702910bfe19e23f3c47bdd885c86b6deefc07edf8a7af01b85305070818a6893728cfcc4da1b64a9364327cf52b6b93c1c31cc1eb4f1f90adc3b34b982d4d35e26fd9b4f005f2c5c253059f5ad1aafa2f17bc8574a19d28c273754aefe577ce97eae55cdb440d043cdee23a0d94aabc0193dbb00a05b8a1781356db5;
    5'b10010 : xpb = 1024'h5f4137667b5154a5609aa2b503f39e84bddd5987b01b31d2994677b8e5cad8a79992480a17d24eceec52defd88046d4cf944b6713b330fc7357e03aac52bef67d8897d05f91b0cbb6267f3d1b19cbf1848f120be2a7e13dbc6644837df976f6df37dde8fed0b57c8c92a3b948b60ea24bb3f5cec59e7ec5fd5da1f38df4a8037;
    5'b10011 : xpb = 1024'ha9411c8d8679988adf972176436b5f811f33fc307075e4c5a811ff56466560deb19a2780bd17a0d8fe8a5951d9c5b2ca9fd2b3a65a34536fb60a0e4aae1caa162e3e26adcb387e27c470bb473e09243ae4c791d963805f6042aebde397f78a2ce8a440365b6859c3de13a6e548d3b0a89d340e189a921dbf0b58b45a3d5f92b9;
    5'b10100 : xpb = 1024'h4293bc5ecfb3a7a7938e28607288d92c0f149ba85b58f7413900cd9df3fd3c0dc659897e983674547163945f4828e77de24688f55682c6cc85f6d98c5c3af0130fa39ba6edc4f24f13df801a3199c52c8c99095c0ffc7dd4096ca194962d0259aec30fb318fc63316c3d2b570e765103304ee0628af0f1edfa67ce7712923ed0;
    5'b10101 : xpb = 1024'h8c93a185dadbeb8d128aa721b2009a28706b3e511bb3aa3447cc553b5497c444de6168f53d7bc65e839b0eb399ea2cfb88d4862a75840a750682e42c452baac16558454ebfe263bb75e8478fbe062a4f286f7a7748fec95885b717404e8d1d18a3e971598759652c812696a7cbe917871243918ecb9b234d2fe6639870a75152;
    5'b10110 : xpb = 1024'h25e641572415faa9c681ae0be11e13d3604bddc90696bcafd8bb2383022f9f73f320caf3189a99d9f67449c1084d61aecb485b7971d27dd1d66faf6df349f0be46bdba47e26ed7e2c5570c62b196cb40d040f1f9f57ae7cc4c74faf14cc295456a0840d644ed6e9a0f501b19918bb7e1a55e63d8bbf9f77c1ef57db545d9fd69;
    5'b10111 : xpb = 1024'h6fe6267e2f3e3e8f457e2ccd2095d4cfc1a28071c6f16fa2e786ab2062ca27ab0b28aa69bddfebe408abc4155a0ea72c71d658ae90d3c17a56fbba0ddc3aab6c9c7263efb48c494f275fd3d83e0330636c1763152e7d3350c8bf709d0522b0045f2ea27cb34a70952439866a4efe7e6587531504fca428db547412d6a3ef0feb;
    5'b11000 : xpb = 1024'h938c64f78784dabf97533b74fb34e7ab1831fe9b1d4821e78757968106202da1fe80c6798febf5f7b84ff22c871dbdfb44a2dfd8d2234d726e8854f8a58f1697dd7d8e8d718bd7676ce98ab3193d15513e8da97daf951c48f7d544e03582831254d71f970de7a02b2630adc14a11ec01a6de74eed02fd0a43832cf37921bc02;
    5'b11001 : xpb = 1024'h5338ab7683a091917871b2788f2b0f7712d9c292722f35118741010570fc8b1137efebde3e4411698dbc79771a33215d5ad82b32ac23787fa7748fef7349ac17d38c8290a9362ee2d8d76020be003677afbf4bb313fb9d490bc7c9f9bbb842f01a73d39fdf3b7bfdc74c762cd213e543fc62987b2dad2e697901c214d736ce84;
    5'b11010 : xpb = 1024'h9d38909d8ec8d576f76e3139cea2d0737430653b3289e804960c88a2d19713484ff7cb54e38963739ff3f3cb6bf466db01662867cb24bc2828009a8f5c3a66c629412c387b53a04f3ae027964a6c9b9a4b95bcce4cfde8cd88123fa574185daf0f9a35464d987df8dc35e17d8f86abc7de5749a76e575fc8ae805736354be106;
    5'b11011 : xpb = 1024'h368b306ed802e493ab653823fdc04a1e641104b31d6cfa8026fb56ea7f2eee7764b72d52bea836ef12cd2ed8da579b8e43d9fdb6c7732f84f7ed65d10a58acc30aa6a1319de014768a4eec693dfd3c8bf3673450f97a07414ed02356724dd5dbd5b904c30b2c87666a5f65ef55294c2271721bf15eb633f79d8f71530a7e8d1d;
    5'b11100 : xpb = 1024'h808b1595e32b28792a61b6e53d380b1ac567a75bddc7ad7335c6de87dfc976ae7cbf0cc963ed88f92504a92d2c18e10bea67faebe674732d78797070f3496771605b4ad96ffd85e2ec57b3deca69a1ae8f3da56c327c52c5cb1a99022aadf09acadf6669798989617f48d140129c12a65366cd1d9f606556d30e067468939f9f;
    5'b11101 : xpb = 1024'h19ddb5672c653795de58bdcf6c5584c5b54846d3c8aabfeec6b5accf8d6151dd917e6ec73f0c5c7497dde43a9a7c15bf2cdbd03ae2c2e68a48663bb2a167ad6e41c0bfd29289fa0a3bc678b1bdfa42a0370f1ceedef8713991d87cb328e368c790fe35e6371d92cf0d7255b1d83eb300e6819f678fbf3985c21d20913dc64bb6;
    5'b11110 : xpb = 1024'h63dd9a8e378d7b7b5d553c90abcd45c2169ee97c890572e1d581346cedfbda14a9864e3de451ae7eaa155e8eec3d5b3cd369cd7001c42a32c8f246528a58681c9775697a64a76b769dcf40274a66a7c2d2e58e0a17fabcbe0e22f25ee14383868624978ca57a94ca225bc10295b17984c8765093d0696ae4f79bb5b29bdb5e38;
    5'b11111 : xpb = 1024'haddd7fb542b5bf60dc51bb51eb4506be77f58c25496025d4e44cbc0a4e96624bc18e2db489970088bc4cd8e33dfea0ba79f7caa520c56ddb497e50f2734922caed2a132236c4dce2ffd8079cd6d30ce56ebbff2550fd08428a6d680a99a39e457b4af93313d796c537452c5353244008aa6b01c011139c442d1a4ad3f9f070ba;
    endcase
end

endmodule

module xpb_5_635
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8d3f1fe0c6f9b59271c3ff3fa34732858ff583dd2bb9614799c3ca49e2020b12b823f539a09d4ccd437c3e0cec99aed3bbd3601533ccdf71a20337179a0db765e0a8ce2b38e52cb1bcafd7e1855812a9f9ccbceb304bd53fdcb9324709cb718540157cfb692da812c9a49c80488f6c8cca40fe19448ec5202d6d81fd53029937;
    5'b00010 : xpb = 1024'h69d0fa6bcc05365c188286a836341db9ae75048981fb2217b5aadb3e1101691d6cff6cfa77141b0be79a3cd2f5d54cdd138c984444e6ee9793672ed0f948fa1a4d0267a7c2395c1e66c5ad2071d46122ff94803dd4117d6f03e5d293596c4078512367cd219257980c895221994eb2f045a81d5038d22d10146b88f61d22cc03;
    5'b00011 : xpb = 1024'h4662d4f6d110b725bf410e10c92108edccf48535d83ce2e7d191ec324000c72821dae4bb4d8ae94a8bb83b98ff10eae66b45d0735600fdbd84cb268a58843cceb95c01244b8d8b8b10db825f5e50af9c055c439077d7259e2b1272dfa90d0f6b6231529ed9f7071d4f6e07c2ea0df953c10f3c872d1594fffb698feee742fecf;
    5'b00100 : xpb = 1024'h22f4af81d61c37ef65ff95795c0df421eb7405e22e7ea3b7ed78fd266f002532d6b65c7c2401b7892fd63a5f084c88efc2ff08a2671b0ce3762f1e43b7bf7f8325b59aa0d4e1baf7baf1579e4accfe150b2406e31b9ccdcd523f132bf8adde5e733f3d70925bb6a29252bd643acd3fb73c765bbe2158fcefe26796e7b163319b;
    5'b00101 : xpb = 1024'hb033cf629d15ed81d7c394b8ff5526a77b6989bf5a3804ff873cc770510230458eda51b5c49f04567352786bf4e637c37ed268b79ae7ec551832555b51cd36e9065e68cc0dc6e7a977a12f7fd02510bf04f0c3ce4be8a30d2ef8457302794fe3b354ba6bfb895eb55bf759e4835cac4406b759d765e7c2100fd518e50465cad2;
    5'b00110 : xpb = 1024'h8cc5a9eda2216e4b7e821c21924211db99e90a6bb079c5cfa323d86480018e5043b5c9769b15d29517707731fe21d5ccd68ba0e6ac01fb7b09964d14b108799d72b80248971b171621b704bebca15f380ab88720efae4b3c5624e5bf521a1ed6c462a53db3ee0e3a9edc0f85d41bf2a7821e790e5a2b29fff6d31fddce85fd9e;
    5'b00111 : xpb = 1024'h69578478a72cef152540a38a252efd0fb8688b1806bb869fbf0ae958af00ec5af8914137718ca0d3bb8e75f8075d73d62e44d915bd1c0aa0fafa44ce1043bc51df119bc5206f4682cbccd9fda91dadb110804a739373f36b7d51860ba1baedc9d570900f6c52bdbfe1c0c52724db390afd8598454e6e91efddd126d698a6306a;
    5'b01000 : xpb = 1024'h45e95f03ac386fdecbff2af2b81be843d6e80bc45cfd476fdaf1fa4cde004a65ad6cb8f848036f125fac74be109911df85fe1144ce3619c6ec5e3c876f7eff064b6b3541a9c375ef75e2af3c9599fc2a16480dc637399b9aa47e2657f15bbcbce67e7ae124b76d4524a57ac8759a7f6e78ecb77c42b1f9dfc4cf2dcf62c66336;
    5'b01001 : xpb = 1024'h227b398eb143f0a872bdb25b4b08d377f5678c70b33f083ff6d90b410cffa870624830b91e7a3d5103ca738419d4afe8ddb74973df5028ecddc23440ceba41bab7c4cebe3317a55c1ff8847b82164aa31c0fd118daff43c9cbaac6a440fc8baff78c65b2dd1c1cca678a3069c659c5d1f453d6b336f561cfabcd34c82ce69602;
    5'b01010 : xpb = 1024'hafba596f783da63ae481b19aee5005fd855d104ddef86987909cd58aef01b3831a6c25f2bf178a1e4746b191066e5ebc998aa989131d085e7fc56b5868c7f920986d9ce96bfcd20ddca85c5d076e5d4d15dc8e040b4b1909a863f8eb4ac7fd3537a1e2ae4649c4dd312eccea0ee9325ebe94d4cc7b8426efd93ab6c57fe92f39;
    5'b01011 : xpb = 1024'h8c4c33fa7d4927048b403903813cf131a3dc90fa353a2a57ac83e67f1e01118dcf479db3958e585ceb64b0570fa9fcc5f143e1b82437178471296311c8033bd504c73665f551017a86be319bf3eaabc61ba45156af10c138cf9099379a68cc2848afcd7ffeae74627413828b5fa878c239fbf4036fc78edfc038bdbe4a096205;
    5'b01100 : xpb = 1024'h68de0e858254a7ce31fec06c1429dc65c25c11a68b7beb27c86af7734d006f98842315746c05269b8f82af1d18e59acf48fd19e7355126aa628d5acb273e7e897120cfe27ea530e730d406dae066fa3f216c14a952d66967f6bd3983ea099b1b59bdb851b71323e7b6f8382cb067bf25b563133a640af6cfa736c4b7142994d1;
    5'b01101 : xpb = 1024'h456fe91087602897d8bd47d4a716c799e0db9252e1bdabf7e45208677bffcda338fe8d35427bf4da33a0ade3222138d8a0b65216466b35d053f152848679c13ddd7a695f07f96053dae9dc19cce348b82733d7fbf69c11971de9d9d039aa6a0e6acba3236f77d36cf9dcedce0127058930ca3271584e5ebf8e34cbafde49c79d;
    5'b01110 : xpb = 1024'h2201c39b8c6ba9617f7bcf3d3a03b2cdff5b12ff37ff6cc80039195baaff2badedda04f618f2c318d7beaca92b5cd6e1f86f8a45578544f645554a3de5b503f249d402db914d8fc084ffb158b95f97312cfb9b4e9a61b9c645167a1c894b39017bd98df527dc82f23cc1a36f51e64becac3151a84c91c6af7532d2a8a869fa69;
    5'b01111 : xpb = 1024'haf40e37c53655ef3f13fce7cdd4ae5538f5096dc63b8ce0f99fce3a58d0136c0a5fdfa2fb9900fe61b3aeab617f685b5b442ea5a8b522467e75881557fc2bb582a7cd106ca32bc7241af893a3eb7a9db26c85839caad8f0621cfac639316aa86bbef0af0910a2b0506663fef9a75b87976724fc191208bcfa2a054a5fb6c93a0;
    5'b10000 : xpb = 1024'h8bd2be075870dfbd97fe55e57037d087add01788b9fa8edfb5e3f499bc0094cb5ad971f09006de24bf58e97c213223bf0bfc22899c6c338dd8bc790edefdfe0c96d66a835386ebdeebc55e792b33f8542c901b8c6e73373548fc4cafe2b77979ccfcf5c2496eda8a494af590eb34fedcf1d96ef88563f3bf899e5b9ec58cc66c;
    5'b10001 : xpb = 1024'h686498925d7c60873ebcdd4e0324bbbbcc4f9835103c4fafd1cb058deafff2d60fb4e9b1667dac636376e8422a6dc1c863b55ab8ad8642b3ca2070c83e3940c1033003ffdcdb1b4b95db33b817b046cd3257dedf1238df647028ecfc3258486cde0ae09401d38a0f8c2fab323bf445406d408e2f79a75baf709c62978facf938;
    5'b10010 : xpb = 1024'h44f6731d6287e150e57b64b69611a6efeacf18e1667e107fedb2168219ff50e0c49061723cf47aa20794e70833a95fd1bb6e92e7bea051d9bb8468819d7483756f899d7c662f4ab83ff108f7042c9546381fa231b5fe879397558d4881f9175fef18cb65ba383994cf1460d38cb38ba3e8a7ad666deac39f579a699059cd2c04;
    5'b10011 : xpb = 1024'h21884da86793621a8c39ec1f28fe9224094e998dbcbfd1500999277648feaeeb796bd933136b48e0abb2e5ce3ce4fddb1327cb16cfba60fface8603afcafc629dbe336f8ef837a24ea06de35f0a8e3bf3de7658459c42fc2be822d94d199e6530026b637729ce91a11f91674dd72d207640ecc9d622e2b8f3e98708923ed5ed0;
    5'b10100 : xpb = 1024'haec76d892e8d17acfdfdeb5ecc45c4a999441d6ae8793297a35cf1c02b00b9fe318fce6cb40895adef2f23db297eacaecefb2b2c038740714eeb975296bd7d8fbc8c05242868a6d6a6b6b6177600f66937b4226f8a1005029b3b5fdbdb6557d8403c3332dbca912cdb9db2f526023e942e4fcab6a6bcf0af6c05f28676eff807;
    5'b10101 : xpb = 1024'h8b59481433989876a4bc72c75f32afddb7c39e173ebaf367bf4402b45a001808e66b462d8a7f63ec934d22a132ba4ab826b4635b14a14f97404f8f0bf5f8c04428e59ea0b1bcd64350cc8b56627d44e23d7be5c22dd5ad31c26800282b0626cb514a1e04942f40b21e82689676c184f7a9b6e9ed9b00589f5303f97f41102ad3;
    5'b10110 : xpb = 1024'h67eb229f38a419404b7afa2ff21f9b11d6431ec394fcb437db2b13a888ff76139b46bdee60f6322b376b21673bf5e8c17e6d9b8a25bb5ebd31b386c5553402f8953f381d3b1105affae260954ef9935b4343a914d19b5560e994a0747aa6f5be625808d64c93f03761671e37c780cb5b251e09248f43c08f3a0200780b305d9f;
    5'b10111 : xpb = 1024'h447cfd2a3daf9a09f2398198850c8645f4c29f6feb3e7507f712249cb7fed41e502235af376d0069db89202d453186cad626d3b936d56de323177e7eb46f45ad0198d199c465351ca4f835d43b75e1d4490b6c677560fd9010c140c0ca47c4b17365f3a804f89fbca44bd3d9184011bea085285b8387287f21000770d550906b;
    5'b11000 : xpb = 1024'h210ed7b542bb1ad398f8090117f9717a1342201c418035d812f93590e6fe322904fdad700de3cea87fa71ef34e6d24d42de00be847ef7d09147b763813aa88616df26b164db964894f0e0b1327f2304d4ed32fba1926a5bf37ede10d19e893a48473de79bd5d4f41e730897a68ff58221bec479277ca906f07fe0e699f70c337;
    5'b11001 : xpb = 1024'hae4df79609b4d0660abc0840bb40a3ffa337a3f96d39971facbcffdac9003d3bbd21a2a9ae811b75c3235d003b06d3a7e9b36bfd7bbc5c7ab67ead4fadb83fc74e9b3941869e913b0bbde2f4ad4a42f7489feca549727aff14a7135423b40529c4895b75268af754b0d525fab18ec4aee62d45abbc59558f356b9066f2735c6e;
    5'b11010 : xpb = 1024'h8adfd2210ec0512fb17a8fa94e2d8f33c1b724a5c37b57efc8a410cef7ff9b4671fd1a6a84f7e9b467415bc6444271b1416ca42c8cd66ba0a7e2a5090cf3827bbaf4d2be0ff2c0a7b5d3b83399c691704e67aff7ed38232e3bd3b3a07354d41cd5974646deefa6d9f3b9db9c024e0b12619464e2b09cbd7f1c69975fbc938f3a;
    5'b11011 : xpb = 1024'h6771acac13cbd1f958391711e11a7a67e036a55219bd18bfe48b21c326fef95126d8922b5b6eb7f30b5f5a8c4d7e0fba9925dc5b9df07ac699469cc26c2ec530274e6c3a9946f0145fe98d728642dfe9542f734a90fdcb5d630053ecc2f5a30fe6a531189754565f369e913d530d5175dcfb8419a4e0256f03679e5886b3c206;
    5'b11100 : xpb = 1024'h4403873718d752c2fef79e7a7407659bfeb625fe6ffed990007232b755fe575bdbb409ec31e58631af7d595256b9adc3f0df148aaf0a89ec8aaa947bcb6a07e493a805b7229b1f8109ff62b172bf2e6259f7369d34c3738c8a2cf43912967202f7b31bea4fb905e4798346dea3cc97d95862a35099238d5eea65a55150d3f4d2;
    5'b11101 : xpb = 1024'h209561c21de2d38ca5b625e306f450d01d35a6aac6409a601c5943ab84fdb566908f81ad085c5470539b58185ff54bcd48984cb9c02499127c0e8c352aa54a9900019f33abef4eedb41537f05f3b7cdb5fbef9efd8891bbbb1599485623740f608c106bc081db569bc67fc7ff48bde3cd3c9c2878d66f54ed163ac4a1af4279e;
    5'b11110 : xpb = 1024'hadd481a2e4dc891f177a2522aa3b8355ad2b2a87f1f9fba7b61d0df566ffc07948b376e6a8f9a13d971796254c8efaa1046baccef3f178841e11c34cc4b301fee0aa6d5ee4d47b9f70c50fd1e4938f85598bb6db08d4f0fb8e12c6cc6c02b27b48d683b7714b5d7c860c99003d1b4ac99e0ac0a0d1f5ba6efed12e476df6c0d5;
    5'b11111 : xpb = 1024'h8a665c2de9e809e8be38ac8b3d286e89cbaaab34483bbc77d2041ee995ff1e83fd8eeea77f706f7c3b3594eb55ca98aa5c24e4fe050b87aa0f75bb0623ee44b34d0406db6e28ab0c1adae510d10fddfe5f537a2dac9a992ab53f6718bba3816e59e46e8929b00d01c8f14ea18dda912d1971dfd7c639225ee5cf35403816f3a1;
    endcase
end

endmodule

module xpb_5_625
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1ae18a06b34c8ceac95784e39da27c1835509a5c9b9ac9e268339a004b512833bb2d41fb57017afb49f063237e25a3765795ea621b0d843f51649ba5494dde97b5d3276cfbe16ba160fffbdc150499f7136e33f71211624797723565457066f801ee6abf0e5cb70970d7f5596014e5a1e3e20abc47f88c0c56b4bb3f6f0d05a7;
    5'b00010 : xpb = 1024'h35c3140d669919d592af09c73b44f8306aa134b9373593c4d067340096a25067765a83f6ae02f5f693e0c646fc4b46ecaf2bd4c4361b087ea2c9374a929bbd2f6ba64ed9f7c2d742c1fff7b82a0933ee26dc67ee2422c48f2ee46aca8ae0cdf003dcd57e1cb96e12e1afeab2c029cb43c7c415788ff11818ad69767ede1a0b4e;
    5'b00011 : xpb = 1024'h50a49e1419e5a6c05c068eaad8e774489ff1cf15d2d05da7389ace00e1f3789b3187c5f2050470f1ddd1296a7a70ea6306c1bf2651288cbdf42dd2efdbe99bc721797646f3a442e422fff3943f0dcde53a4a9be5363426d6c656a02fd05134e805cb403d2b16251c5287e00c203eb0e5aba62034d7e9a425041e31be4d2710f5;
    5'b00100 : xpb = 1024'h6b86281acd3233ab255e138e7689f060d54269726e6b2789a0ce68012d44a0ceecb507ed5c05ebed27c18c8df8968dd95e57a9886c3610fd45926e9525377a5ed74c9db3ef85ae8583ffef70541267dc4db8cfdc4845891e5dc8d59515c19be007b9aafc3972dc25c35fd565805396878f882af11fe230315ad2ecfdbc34169c;
    5'b00101 : xpb = 1024'h8667b221807ec095eeb59872142c6c790a9303cf0a05f16c090202017895c902a7e249e8b30766e871b1efb176bc314fb5ed93ea8743953c96f70a3a6e8558f68d1fc520eb671a26e4ffeb4c691701d3612703d35a56eb65f53b0afa5b3202d809a815bb47cf932f3437cabee0687c29736a35ad67dabc3db187a83d2b411c43;
    5'b00110 : xpb = 1024'ha1493c2833cb4d80b80d1d55b1cee8913fe39e2ba5a0bb4e71359c01c3e6f136630f8be40a08e1e3bba252d4f4e1d4c60d837e4ca251197be85ba5dfb7d3378e42f2ec8de74885c845ffe7287e1b9bca749537ca6c684dad8cad405fa0a269d00b96807a562c4a38a50fc018407d61cb574c4069afd3484a083c637c9a4e21ea;
    5'b00111 : xpb = 1024'hb7d80d92529a5a2b65f2a623f171d5803be35576bc3e4b95b8c7cac5c356c621af4506696e3de50663476b18fa9677200ff40c89aabcd6f89210226c64ea1748476df4c3398f4249465e061fa44719093fe7228f1f382e46e92e3ca2be82e35de7d590fb3c008b48f27ce92a8c22143ec546c43a78077261881a3b78078c126;
    5'b01000 : xpb = 1024'h265f0adfd876328d7fb6af45dcb99970390ecfb4075eae9bc3c016aca7869495d6219261ede5594bb024d9d50dcf0ae858952b2ab5b951aeda859dcc0f9c800c3a4a06b92f7a5fc5f565dc3e0f490b87a76ca6200404e52c0605192f7158952de06bc3cec21cbfbdffffc3ec08d706e5d03676ffef7903326f365ef6ef85c6cd;
    5'b01001 : xpb = 1024'h414094e68bc2bf78490e34297a5c15886e5f6a10a2f9787e2bf3b0acf2d7bcc9914ed45d44e6d446fa153cf88bf4ae5eb02b158cd0c6d5ee2bea397158ea5ea3f01d2e262b5bcb675665d81a244da57ebadada17161647739d774e94b6c8fc25e25a2e8dd07976c770d7b94568ebec87b41881bc37718f3ec5eb1a365e92cc74;
    5'b01010 : xpb = 1024'h5c221eed3f0f4c631265b90d17fe91a0a3b0046d3e94426094274aad3e28e4fd4c7c16589be84f424405a01c0a1a51d507c0ffeeebd45a2d7d4ed516a2383d3ba5f05593273d3708b765d3f639523f75ce490e0e2827a9bb34e983f9fc39631de448994cded62dd0e1afae9ec900d22997fa8c787f6a1b4b1c9fd575cd9fd21b;
    5'b01011 : xpb = 1024'h7703a8f3f25bd94ddbbd3df0b5a10db8d9009ec9da2f0c42fc5ae4ad897a0d3107a95853f2e9ca3d8df6033f883ff54b5f56ea5106e1de6cceb370bbeb861bd35bc37d00231ea2aa1865cfd24e56d96ce1b742053a390c02cc5bb95f41a9ca15e637040bed32e4da5287a3f82915b7cb7bdc9734c762a757735490b53cacd7c2;
    5'b01100 : xpb = 1024'h91e532faa5a86638a514c2d4534389d10e51392675c9d625648e7eadd4cb3564c2d69a4f49eb4538d7e66663066598c1b6ecd4b321ef62ac20180c6134d3fa6b1196a46d1f000e4b7965cbae635b7363f52575fc4c4a6e4a63cdeec4871a310de8256ecafb8f9be3c35f9951892a9d6d5fbea1f10f5b3363ca094bf4abb9dd69;
    5'b01101 : xpb = 1024'hacc6bd0158f4f3236e6c47b7f0e605e943a1d3831164a007ccc218ae201c5d987e03dc4aa0ecc03421d6c986848b3c380e82bf153cfce6eb717ca8067e21d902c769cbda1ae179ecda65c78a78600d5b0893a9f35e5bd091fb402429cc8a9805ea13d98a09ec52ed34378eaae93f830f43a0acad5753bf7020be07341ac6e310;
    5'b01110 : xpb = 1024'h16fb01b24a534b456cbe54c47e2e3ab0077c6aaed787c972b718f958b86ad8c435e8a0cd2dc7bca0cc68ed631f52cee401fe819135579adf1242044d8c9d42e908edbe986731e84928cbc0c3f488e32127fce451e3e705c8dd25c79457d05c6bbcfab21f678011691e4f9d2551844287d8a8d8874f00ee4c3103476f00f1824c;
    5'b01111 : xpb = 1024'h31dc8bb8fd9fd8303615d9a81bd0b6c83ccd050b732293551f4c935903bc00f7f115e2c884c9379c165950869d78725a59946bf350651f1e63a69ff2d5eb2180bec0e605631353ea89cbbca0098d7d183b6b1848f5f868107497fcf99d40c363bee91cde75dcc8728f27927eb1992829bc8ae34396f97a5887b802ae6ffe87f3;
    5'b10000 : xpb = 1024'h4cbe15bfb0ec651aff6d5e8bb97332e0721d9f680ebd5d3787802d594f0d292bac4324c3dbcab2976049b3aa1b9e15d0b12a56556b72a35db50b3b981f39001874940d725ef4bf8beacbb87c1e92170f4ed94c400809ca580c0a325ee2b12a5bc0d7879d84397f7bffff87d811ae0dcba06cedffdef20664de6cbdeddf0b8d9a;
    5'b10001 : xpb = 1024'h679f9fc66438f205c8c4e36f5715aef8a76e39c4aa582719efb3c7599a5e515f677066bf32cc2d92aa3a16cd99c3b94708c040b78680279d066fd73d6886deb02a6734df5ad62b2d4bcbb4583396b106624780371a1b2c9fa37c67c428219153c2c5f25c9296368570d77d3171c2f36d844ef8bc26ea92713521792d4e189341;
    5'b10010 : xpb = 1024'h828129cd17857ef0921c6852f4b82b10dcbed42145f2f0fc57e76159e5af7993229da8ba89cda88df42a79f117e95cbd60562b19a18dabdc57d472e2b1d4bd47e03a5c4c56b796ceaccbb034489b4afd75b5b42e2c2c8ee73aee9d296d91f84bc4b45d1ba0f2ed8ee1af728ad1d7d90f683103786ee31e7d8bd6346cbd2598e8;
    5'b10011 : xpb = 1024'h9d62b3d3cad20bdb5b73ed36925aa729120f6e7de18dbadec01afb5a3100a1c6ddcaeab5e0cf23893e1add14960f0033b7ec157bbc9b301ba9390e87fb229bdf960d83b9529902700dcbac105d9fe4f48923e8253e3df12ed260d28eb3025f43c6a2c7daaf4fa498528767e431ecbeb14c130e34b6dbaa89e28aefac2c329e8f;
    5'b10100 : xpb = 1024'h796f884bc3063fd59c5fa431fa2dbefd5ea05a9a7b0e449aa71dc04c94f1cf295afaf386daa1ff5e8ad00f130d692dfab67d7f7b4f5e40f49fe6acf099e05c5d79176779ee970cc5c31a549d9c8babaa88d2283c3c92665b44675f93e4823a99989a0700ce363143c9f765e9a317e29e11b3a0eae88d965f2d02fe7125d3dcb;
    5'b10101 : xpb = 1024'h2278828b6f7cf0e8231d7f26bd4558080b3aa006434bae2c12a5760514a0452650dcf133c4ab9af1329d6414aefc365602fdc259d003684e9b63067452ebe45d8d649de49acadc6dbd31a125eecd54b1bbfb567ad5da88ad4bb8ab5e83b88aa19b780b2f1b401a1dad776bb7fa4663cbc4fd44caf68165724984eb26816a4372;
    5'b10110 : xpb = 1024'h3d5a0c9222c97dd2ec75040a5ae7d420408b3a62dee6780e7ad910055ff16d5a0c0a332f1bad15ec7c8dc7382d21d9cc5a93acbbeb10ec8decc7a2199c39c2f54337c55196ac480f1e319d0203d1eea8cf698a71e7ebeaf4e32ae0c3c928f1999d6675ee299cd1271e4f61115a5b496da8df4f873e79f17ea039a665f0774919;
    5'b10111 : xpb = 1024'h583b9698d6160abdb5cc88edf88a503875dbd4bf7a8141f0e30caa05ab42958dc737752a72ae90e7c67e2a5bab477d42b229971e061e70cd3e2c3dbee587a18cf90aecbe928db3b07f3198de18d6889fe2d7be68f9fd4d3c7a9d16290e9958919f54e0ad37f988308f27566aba702f0f8cc15a4386727d8af6ee61a55f844ec0;
    5'b11000 : xpb = 1024'h731d209f896297a87f240dd1962ccc50ab2c6f1c161c0bd34b404405f693bdc18264b725c9b00be3106e8d7f296d20b909bf8180212bf50c8f90d9642ed58024aede142b8e6f1f51e03194ba2ddb2296f645f2600c0eaf84120f4b8e5409bf89a1434b6c46563f39ffff4bc41a8514b170a364ffce6b09974da31ce4ce915467;
    5'b11001 : xpb = 1024'h8dfeaaa63caf2493487b92b533cf4868e07d0978b1b6d5b5b373de0641e4e5f53d91f92120b186de5a5ef0a2a792c42f61556be23c39794be0f5750978235ebc64b13b988a508af34131909642dfbc8e09b426571e2011cba98180f3997a2681a331b62b54b2f64370d7411d7a99fa5354856fbc166395a3a457d8243d9e5a0e;
    5'b11010 : xpb = 1024'ha8e034aceffbb17e11d31798d171c48115cda3d54d519f981ba778068d360e28f8bf3b1c77b301d9a44f53c625b867a5b8eb56445746fd8b325a10aec1713d541a8463058631f694a2318c7257e456851d225a4e3031741340f3b658deea8d79a52020ea630fad4ce1af3676daaedff538677a785e5c21affb0c9363acab5fb5;
    5'b11011 : xpb = 1024'h1314795de15a09a0102524a55eb9f947d9a83b011374c90305fe58b125848954b0a3ff9f048dfe464ee177a2c07ffa51ac6718c04fa1b17ed31f6cf5cfeca73a5c0855c3d28264f0f09785abd40d2c4b3c8b94acb5bca94a22d959c36a3051df7806f97fc0a36bc8cbc744f142f39f6dcd6fa6525609508c0b51d39e92d5fef1;
    5'b11100 : xpb = 1024'h2df6036494a6968ad97ca988fc5c75600ef8d55daf0f92e56e31f2b170d5b1886bd1419a5b8f794198d1dac63ea59dc803fd03226aaf35be2484089b193a85d211db7d30ce63d09251978187e911c6424ff9c8a3c7ce0b91ba4b8f28afa0b8d779f5643ecf0022d23c9f3a4aa308850fb151b10e9e01dc9862068ede01e30498;
    5'b11101 : xpb = 1024'h48d78d6b47f32375a2d42e6c99fef17844496fba4aaa5cc7d6658cb1bc26d9bc26fe8395b290f43ce2c23de9bccb413e5b92ed8485bcb9fd75e8a44062886469c7aea49dca453c33b2977d63fe1660396367fc9ad9df6dd951bdc48df5111fcf7be3cefddd5cd9dbad772fa4031d6ab19533bbcae5fa68a4b8bb4a1d70f00a3f;
    5'b11110 : xpb = 1024'h63b91771fb3fb0606c2bb35037a16d90799a0a16e64526aa3e9926b2077801efe22bc59109926f382cb2a10d3af0e4b4b328d7e6a0ca3e3cc74d3fe5abd643017d81cc0ac626a7d513977940131afa3076d63091ebf0d020e92ff9f33a8186c77dd239bcebb990e51e4f24fd633250537915c6872df2f4b10f70055cdffd0fe6;
    5'b11111 : xpb = 1024'h7e9aa178ae8c3d4b35833833d543e9a8aeeaa47381dff08ca6ccc0b252c92a239d59078c6093ea3376a30430b916882b0abec248bbd7c27c18b1db8af52421993354f377c20813767497751c281f94278a446488fe02326880a22f587ff1edbf7fc0a47bfa1647ee8f271a56c34735f55cf7d14375eb80bd6624c09c4f0a158d;
    endcase
end

endmodule

module xpb_5_785
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'habcb4c0972ab81b8723dd44edcdf0bbad78889fb9c7fe8c153423fa21667873be97acb8ec7ea29ffcfb568bf8cc75fb3ad042c11efd63500d987e1d4fb9ef88e0ef9d88ea5fb1a777aa4e2977d46917642ee41acc4b7813e8f0e20db373815dcd58eea54140b5f45eeacf771ba86a67a3d122098b734e47c114a23981a1e13ff;
    5'b00010 : xpb = 1024'ha6e952bd2368cea8197630c6a963d0243d9b10c66388310b28a7c5ee79cc616fcfad19a4c5add571000c92383630ae9cf5ee303dbcf999b60270844bbc6b7c6aa9a47c6e9c6537a9e2afc28c61b15ebb91d789c0fce8d56c688fafbbb44589277c16427e774dc5fe569a08047d3d26cb2b4a624f1e1e6bc7dc24cc2bab59c193;
    5'b00011 : xpb = 1024'ha2075970d4261b97c0ae8d3e75e8948da3ad97912a907954fe0d4c3add313ba3b5df67bac37180e23063bbb0df99fd863ed834698a1cfe6b2b5926c27d380047444f204e92cf54dc4abaa281461c2c00e0c0d1d5351a299a42113e9c3152fc72229d9aa8da902cb6be8718973ff3a71c1982a4058507f313a6ff74bf3c956f27;
    5'b00100 : xpb = 1024'h9d25602484e3688767e6e9b6426d58f709c01e5bf198c19ed372d287409615d79c11b5d0c1352c5360bae52989034c6f87c23895574063205441c9393e048423def9c42e8939720eb2c582762a86f9462faa19e96d4b7dc81b92cd7cae606fbcc924f2d33dd2936f2674292a02aa276d07bae5bbebf17a5f71da1d52cdd11cbb;
    5'b00101 : xpb = 1024'h984366d835a0b5770f1f462e0ef21d606fd2a526b8a109e8a8d858d3a3faf00b824403e6bef8d7c491120ea2326c9b58d0ac3cc12463c7d57d2a6baffed1080079a4680e7fa38f411ad0626b0ef1c68b7e9361fda57cd1f5f5145c5d2b6de3076fac4afda114fa278e6139bcc560a7bdf5f3277252db01ab3cb4c5e65f0cca4f;
    5'b00110 : xpb = 1024'h93616d8be65e0266b657a2a5db76e1c9d5e52bf17fa952327e3ddf20075fca3f687651fcbcbc8335c169381adbd5ea42199640ecf1872c8aa6130e26bf9d8bdd144f0bee760dac7382db425ff35c93d0cd7caa11ddae2623ce95eb3da87b56521633a328045760dff64e4a4f8817280ee42b6928b9c488f7078f6e79f04877e3;
    5'b00111 : xpb = 1024'h8e7f743f971b4f565d8fff1da7fba6333bf7b2bc46b19a7c53a3656c6ac4a4734ea8a012ba802ea6f1c06193853f392b62804518beaa913fcefbb09d806a0fb9aef9afce6c77c9a5eae62254d7c761161c65f22615df7a51a8177a1e2588c99cbcbafb526799c7985e3b5ae24acda85fd263aadf20ae1042d26a170d81842577;
    5'b01000 : xpb = 1024'h899d7af347d89c4604c85b9574806a9ca20a39870db9e2c62908ebb8ce297ea734daee28b843da1822178b0c2ea88814ab6a49448bcdf5f4f7e453144136939649a453ae62e1e6d852f10249bc322e5b6b4f3a3a4e10ce7f819908fea2963ce76342537ccadc2e50c6286b750d8428b0c09bec958797978e9d44bfa112bfd30b;
    5'b01001 : xpb = 1024'h84bb81a6f895e935ac00b80d41052f06081cc051d4c22b0ffe6e7205318e58db1b0d3c3eb6078589526eb484d811d6fdf4544d7058f15aaa20ccf58b02031772e44ef78e594c040abafbe23ea09cfba0ba38824e864222ad5b1a97df1fa3b03209c9aba72e1e95092e157c07d03aa901aed42e4bee811eda681f6834a3fb809f;
    5'b01010 : xpb = 1024'h7fd9885aa9533625533914850d89f36f6e2f471c9bca7359d3d3f85194f3330f013f8a54b3cb30fa82c5ddfd817b25e73d3e519c2614bf5f49b59801c2cf9b4f7ef99b6e4fb6213d2306c2338507c8e60921ca62be7376db349c26bf9cb1237cb05103d19160fbc196028c9a92f129529d0c7002556aa62632fa10c835372e33;
    5'b01011 : xpb = 1024'h7af78f0e5a108314fa7170fcda0eb7d8d441cde762d2bba3a9397e9df8580d42e771d86ab18edc6bb31d07762ae474d0862855c7f3382414729e3a78839c1f2c19a43f4e46203e6f8b11a2286972962b580b1276f6a4cb090e1db5a019be96c756d85bfbf4a36279fdef9d2d55a7a9a38b44b1b8bc542d71fdd4b95bc672dbc7;
    5'b01100 : xpb = 1024'h761595c20acdd004a1a9cd74a6937c423a5454b229db03ed7e9f04ea5bbce776cda42680af5287dce37430eed44dc3b9cf1259f3c05b88c99b86dcef4468a308b44ee32e3c8a5ba1f31c821d4ddd6370a6f45a8b2ed61f36e79f448096cc0a11fd5fb42657e5c93265dcadc0185e29f4797cf36f233db4bdc8af61ef57ae895b;
    5'b01101 : xpb = 1024'h71339c75bb8b1cf448e229ec731840aba066db7cf0e34c3754048b36bf21c1aab3d67496ad16334e13cb5a677db712a317fc5e1f8d7eed7ec46f7f66053526e54ef9870e32f478d45b276212324830b5f5dda29f67077364c120d36113d97d5ca3e70c50bb282feacdc9be52db14aa4567b535258a273c09938a0a82e8ea36ef;
    5'b01110 : xpb = 1024'h6c51a3296c4869e3f01a86643f9d051506796247b7eb9481296a118322869bde9a08c2acaad9debf442283e02720618c60e6624b5aa25233ed5821dcc601aac1e9a42aee295e9606c332420716b2fdfb44c6eab39f38c7929aa2624190e6f0a74a6e647b1e6a96a335b6cee59dcb2a9655ed76dbf110c3555e64b3167a25e483;
    5'b01111 : xpb = 1024'h676fa9dd1d05b6d39752e2dc0c21c97e6c8be9127ef3dccafecf97cf85eb7612803b10c2a89d8a307479ad58d089b075a9d0667727c5b6e91640c45386ce2e9e844ecece1fc8b3392b3d21fbfb1dcb4093b032c7d76a1bc07423f1220df463f1f0f5bca581acfd5b9da3df786081aae74425b89257fa4aa1293f5baa0b619217;
    5'b10000 : xpb = 1024'h628db090cdc303c33e8b3f53d8a68de7d29e6fdd45fc2514d4351e1be9505046666d5ed8a66135a1a4d0d6d179f2ff5ef2ba6aa2f4e91b9e3f2966ca479ab27b1ef972ae1632d06b934801f0df889885e2997adc0f9b6fee4da580028b01d73c977d14cfe4ef64140590f00b23382b38325dfa48bee3d1ecf41a043d9c9d3fab;
    5'b10001 : xpb = 1024'h5dabb7447e8050b2e5c39bcba52b525138b0f6a80d046d5ea99aa4684cb52a7a4c9faceea424e112d528004a235c4e483ba46ecec20c80536812094108673657b9a4168e0c9ced9dfb52e1e5c3f365cb3182c2f047ccc41c27270ee3080f4a873e046cfa4831cacc6d7e009de5eeab8920963bff25cd5938bef4acd12dd8ed3f;
    5'b10010 : xpb = 1024'h58c9bdf82f3d9da28cfbf84371b016ba9ec37d72d40cb5a87f002ab4b01a04ae32d1fb04a1e88c84057f29c2ccc59d31848e72fa8f2fe50890faabb7c933ba34544eba6e03070ad0635dc1daa85e3310806c0b047ffe184a00a89dc3851cbdd1e48bc524ab743184d56b1130a8a52bda0ece7db58cb6e08489cf5564bf149ad3;
    5'b10011 : xpb = 1024'h53e7c4abdffaea92343454bb3e34db2404d6043d9b14fdf25465b101137edee21904491a9fac37f535d6533b762eec1acd7877265c5349bdb9e34e2e8a003e10eef95e4df9712802cb68a1cf8cc90055cf555318b82f6c77da2a2ca4022a311c8b131d4f0eb6983d3d5821c36b5bac2afd06bf6bf3a067d054a9fdf850504867;
    5'b10100 : xpb = 1024'h4f05cb5f90b83781db6cb1330ab99f8d6ae88b08621d463c29cb374d76e3b915ff3697309d6fe366662d7cb41f983b0416627b522976ae72e2cbf0a54accc1ed89a4022defdb4535337381c47133cd9b1e3e9b2cf060c0a5b3abbb847f37a467319a757971f8fef5a54532562e122c7beb3f01225a89ef1c1f84a68be18bf5fb;
    5'b10101 : xpb = 1024'h4a23d2134175847182a50daad73e63f6d0fb11d329258e85ff30bd99da489349e568e5469b338ed79684a62cc90189ed5f4c7f7df69a13280bb4931c0b9945ca244ea60de64562679b7e61b9559e9ae06d27e341289214d38d2d4a64fc4517b1d821cda3d53b65ae0d3242e8f0c8acccd97742d8c1737667ea5f4f1f72c7a38f;
    5'b10110 : xpb = 1024'h4541d8c6f232d16129dd6a22a3c32860370d989df02dd6cfd49643e63dad6d7dcb9b335c98f73a48c6dbcfa5726ad8d6a83683a9c3bd77dd349d3592cc65c9a6bef949eddcaf7f9a038941ae3a096825bc112b5560c3690166aed94579528afc7ea925ce387dcc66751f537bb37f2d1dc7af848f285cfdb3b539f7b304035123;
    5'b10111 : xpb = 1024'h405fdf7aa2f01e50d115c69a7047ecc99d201f68b7361f19a9fbca32a11247b1b1cd817296bae5b9f732f91e1bd427bff12087d590e0dc925d85d8098d324d8359a3edcdd3199ccc6b9421a31e74356b0afa736998f4bd2f40306825f65ffe4725307df89bc0331edd0c640e7635ad6eb5e7c6458f4684ff8014a046953efeb7;
    5'b11000 : xpb = 1024'h3b7de62e53ad6b40784e23123cccb1330332a6337e3e67637f61507f047721e597ffcf88947e912b278a2296c53d76a93a0a8c015e044147866e7a804dfed15ff44e91adc983b9fed39f019802df02b059e3bb7dd126115d19b1f706736d7191cbb7d622ff0299d744f974a138ec2dbfa42007fbf6300c4b4aef48da267aac4b;
    5'b11001 : xpb = 1024'h369bece2046ab8301f867f8a0951759c69452cfe4546afad54c6d6cb67dbfc197e321d9e92423c9c57e14c0f6ea6c59282f4902d2b27a5fcaf571cf70ecb553c8ef9358dbfedd7313ba9e18ce749cff5a8cd03920957658af33385e6f07ae4dc723f2e4d6245008face68533fba2ae10925849b25d19939715c9f16db7b659df;
    5'b11010 : xpb = 1024'h31b9f395b528051fc6bedc01d5d63a05cf57b3c90c4ef7f72a2c5d17cb40d64d64646bb49005e80d883875881810147bcbde9458f84b0ab1d83fbf6dcf97d91929a3d96db657f463a3b4c181cbb49d3af7b64ba64188b9b8ccb514c76d88582718c68677c587674814d395c6be592e6180908b68c4031ae2e0a49a0148f20773;
    5'b11011 : xpb = 1024'h2cd7fa4965e5520f6df73879a25afe6f356a3a93d3574040ff91e3642ea5b0814a96b9ca8dc9937eb88f9f00c179636514c89884c56e6f67012861e490645cf5c44e7d4dacc211960bbfa176b01f6a80469f93ba79ba0de6a636a3a7ea95cb71bf4ddea228c9ce007cc0a659810faeb26ec8cd1f2aeca22eab7f4294da2db507;
    5'b11100 : xpb = 1024'h27f600fd16a29eff152f94f16edfc2d89b7cc15e9a5f888ad4f769b0920a8ab530c907e08b8d3eefe8e6c8796ae2b24e5db29cb09291d41c2a11045b5130e0d25ef9212da32c2ec873ca816b948a37c59588dbceb1eb62147fb8328867a33ebc65d536cc8c0c34b8e4adb6ec43c62f035d010ed591d6297a7659eb286b69629b;
    5'b11101 : xpb = 1024'h231407b0c75febeebc67f1693b648742018f48296167d0d4aa5ceffcf56f64e916fb55f68950ea61193df1f2144c0137a69ca0dc5fb538d152f9a6d211fd64aef9a3c50d99964bfadbd5616078f5050ae47223e2ea1cb6425939c168e4b0b2070c5c8ef6ef4e9b714c9ac77f067caf544b39508bf8bfb0c6413493bbfca5102f;
    5'b11110 : xpb = 1024'h1e320e64781d38de63a04de107e94bab67a1cef42870191e7fc2764958d43f1cfd2da40c871495d249951b6abdb55020ef86a5082cd89d867be24948d2c9e88b944e68ed9000692d43e041555d5fd250335b6bf7224e0a7032bb504961be2551b2e3e72152910229b487d811c9332fa5397192425fa938120c0f3c4f8de0bdc3;
    5'b11111 : xpb = 1024'h1950151828da85ce0ad8aa58d46e1014cdb455beef7861685527fc95bc391950e35ff22284d8414379ec44e3671e9f0a3870a933f9fc023ba4caebbf93966c682ef90ccd866a865fabeb214a41ca9f958244b40b5a7f5e9e0c3cdf29decb989c596b3f4bb5d368e21c74e8a48be9aff627a9d3f8c692bf5dd6e9e4e31f1c6b57;
    endcase
end

endmodule

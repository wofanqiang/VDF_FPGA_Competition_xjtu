module xpb_5_920
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3d5365c20d6f6fcee914fb53ea3449e6d40e7f295e37f06f728b1c9dfdb174492d111260905abf73e66f7d90ac75922b7bb0ab224dbccf3f4876c1b0ddafdf2f248b1ba99f402d0daf0069b8f8f3332ec47a79e854feb49886ba3b74f13f64f1ede8c172843028f5fc0f68e4e8c60fa4076384e227f5f59f546229c80e16f90;
    5'b00010 : xpb = 1024'h7aa6cb841adedf9dd229f6a7d46893cda81cfe52bc6fe0dee516393bfb62e8925a2224c120b57ee7ccdefb2158eb2456f76156449b799e7e90ed8361bb5fbe5e491637533e805a1b5e00d371f1e6665d88f4f3d0a9fd69310d7476e9e27ec9e3dbd182e5086051ebf81ed1c9d18c1f480ec709c44febeb3ea8c453901c2df20;
    5'b00011 : xpb = 1024'hb7fa3146284e4f6cbb3ef1fbbe9cddb47c2b7d7c1aa7d14e57a155d9f9145cdb87333721b1103e5bb34e78b20560b68273120166e9366dbdd9644512990f9d8d6da152fcddc087290d013d2aead9998c4d6f6db8fefc1dc9942eb25ed3be2ed5c9ba44578c907ae1f42e3aaeba522eec162a8ea677e1e0ddfd267d582a44eb0;
    5'b00100 : xpb = 1024'hf54d970835bdbf3ba453ed4fa8d1279b5039fca578dfc1bdca2c7277f6c5d124b4444982416afdcf99bdf642b1d648adeec2ac8936f33cfd21db06c376bf7cbc922c6ea67d00b436bc01a6e3e3ccccbb11e9e7a153fad2621ae8edd3c4fd93c7b7a305ca10c0a3d7f03da393a3183e901d8e13889fd7d67d5188a720385be40;
    5'b00101 : xpb = 1024'h132a0fcca432d2f0a8d68e8a39305718224487bced717b22d3cb78f15f477456de1555be2d1c5bd43802d73d35e4bdad96a7357ab84b00c3c6a51c874546f5bebb6b78a501c40e1446b02109cdcbfffe9d6646189a8f986faa1a32948b63cf8b9a58bc73c94f0cccdec4d0c788bde4e3424f1986ac7cdcc1ca5ead0e84672dd0;
    5'b00110 : xpb = 1024'h16ff4628c509c9ed9767de3f77d39bb68f856faf8354fa29caf42abb3f228b9b70e666e4362207cb7669cf1640ac16d04e62402cdd26cdb7bb2c88a25321f3b1adb42a5f9bb810e521a027a55d5b333189adedb71fdf83b93285d64bda77c5dab937488af1920f5c3e85c755d74a45dd82c551d4cefc3c1bbfa4cfab05489d60;
    5'b00111 : xpb = 1024'h1ad47c84e5e0c0ea85f92df4b676e054fcc657a219387930c21cdc851efda2e003b7780a3f27b3c2b4d0c6ef4b736ff3061d4adf02029aabafb3f4bd60fcf1a49ffcdc1a35ac13b5fc902e40ecea666475f59555a52f6f02baf17a03298bbc29d815d4a219d511eb9e46bde425d6a6d7c33b8a22f17b9b75b4eaf247862a0cf0;
    5'b01000 : xpb = 1024'h1ea9b2e106b7b7e7748a7da9f51a24f36a073f94af1bf837b9458e4efed8ba2496888930482d5fb9f337bec8563ac915bdd8559126de679fa43b60d86ed7ef9792458dd4cfa01686d78034dc7c799997623d3cf42a7f5a4c435d1dba789fb278f6f460b94218147afe07b472746307d203b1c27113fafacfaa3114e4070b7c80;
    5'b01001 : xpb = 1024'h227ee93d278eaee4631bcd5f33bd6991d748278744ff773eb06e4018deb3d16929599a5651330bb1319eb6a161022238759360434bba349398c2ccf37cb2ed8a848e3f8f69941957b2703b780c08ccca4e84e492afcf4595cbc8c171c7b3a8c815d2ecd06a5b170a5dc8ab00c2ef68cc4427fabf367a5a299f77378087ecec10;
    5'b01010 : xpb = 1024'h26541f994865a5e151ad1d147260ae3044890f79dae2f645a796f1e2be8ee8adbc2aab7c5a38b7a87005ae7a6bc97b5b2d4e6af5709601878d4a390e8a8deb7d76d6f14a03881c288d6042139b97fffd3acc8c31351f30df5434652916c79f1734b178e7929e1999bd89a18f117bc9c6849e330d58f9b98394bd5a1d08ce5ba0;
    5'b01011 : xpb = 1024'h2a2955f5693c9cde403e6cc9b103f2ceb1c9f76c70c6754c9ebfa3ac9e69fff24efbbca2633e639fae6ca6537690d47de50975a79571ce7b81d1a5299868e970691fa3049d7c1ef9685048af2b273330271433cfba6f1c28dca008e065db9566539004febae11c291d4a981d60082ac0c5146b5b7b7918dd8a037cb989afcb30;
    5'b01100 : xpb = 1024'h2dfe8c518a1393db2ecfbc7eefa7376d1f0adf5f06a9f45395e855767e451736e1cccdc86c440f96ecd39e2c81582da09cc48059ba4d9b6f76591144a643e7635b6854bf377021ca43404f4abab66663135bdb6e3fbf0772650bac97b4ef8bb5726e9115e3241eb87d0b8eabae948bbb058aa3a99df878377f499f560a913ac0;
    5'b01101 : xpb = 1024'h31d3c2adaaea8ad81d610c342e4a7c0b8c4bc7519c8d735a8d1107405e202e7b749ddeee7549bb8e2b3a96058c1f86c3547f8b0bdf2968636ae07d5fb41ee5564db10679d164249b1e3055e64a459995ffa3830cc50ef2bbed77504f04038204914d1d2d0b672147dccc8539fd20ecb54600dbf7c077d791748fc1f28b72aa50;
    5'b01110 : xpb = 1024'h35a8f909cbc181d50bf25be96cedc0a9f98caf443270f2618439b90a3dfb45c0076ef0147e4f678569a18dde96e6dfe60c3a95be040535575f67e97ac1f9e3493ff9b8346b58276bf9205c81d9d4ccc8ebeb2aab4a5ede0575e2f40653177853b02ba94433aa23d73c8d7bc84bad4daf86771445e2f736eb69d5e48f0c5419e0;
    5'b01111 : xpb = 1024'h397e2f65ec9878d1fa83ab9eab91054866cd9736c85471687b626ad41dd65d049a40013a8755137ca80885b7a1ae3908c3f5a07028e1024b53ef5595cfd4e13c324269ef054c2a3cd410631d6963fffbd832d249cfaec94efe4e97bda22b6ea2cf0a355b5bed26669c4e72569a39aea9c6ed4c94057696455f1c072b8d358970;
    5'b10000 : xpb = 1024'h3d5365c20d6f6fcee914fb53ea3449e6d40e7f295e37f06f728b1c9dfdb174492d111260905abf73e66f7d90ac75922b7bb0ab224dbccf3f4876c1b0ddafdf2f248b1ba99f402d0daf0069b8f8f3332ec47a79e854feb49886ba3b74f13f64f1ede8c172843028f5fc0f68e4e8c60fa4076384e227f5f59f546229c80e16f900;
    5'b10001 : xpb = 1024'h41289c1e2e4666cbd7a64b0928d78e85414f671bf41b6f7669b3ce67dd8c8b8dbfe2238699606b6b24d67569b73ceb4e336bb5d472989c333cfe2dcbeb8add2216d3cd6439342fde89f0705488826661b0c22186da4e9fe20f25df2c40535b410cc74d89ac732b855bd05f733752709e47d9bd304a7554f949a84c648ef86890;
    5'b10010 : xpb = 1024'h44fdd27a4f1d5dc8c6379abe677ad323ae904f0e89feee7d60dc8031bd67a2d252b334aca2661762633d6d42c2044470eb26c08697746927318599e6f965db15091c7f1ed32832af64e076f0181199949d09c9255f9e8b2b979182e38f6751902ba5d9a0d4b62e14bb91560185ded198884ff57e6cf4b4533eee6f010fd9d820;
    5'b10011 : xpb = 1024'h48d308d66ff454c5b4c8ea73a61e17c21bd137011fe26d84580531fb9d42ba16e58445d2ab6bc359a1a4651bcccb9d93a2e1cb38bc50361b260d06020740d907fb6530d96d1c35803fd07d8ba7a0ccc7895170c3e4ee76751ffd269ade7b47df4a8465b7fcf930a41b524c8fd46b3292c8c62dcc8f7413ad3434919d90bb47b0;
    5'b10100 : xpb = 1024'h4ca83f3290cb4bc2a35a3a28e4c15c6089121ef3b5c5ec8b4f2de3c57d1dd15b785556f8b4716f50e00b5cf4d792f6b65a9cd5eae12c030f1a94721d151bd6faedade294071038511ac08427372ffffa759918626a3e61bea868ca522d8f3e2e6962f1cf253c33337b13431e22f7938d093c661ab1f37307297ab43a119cb740;
    5'b10101 : xpb = 1024'h507d758eb1a242bf91eb89de2364a0fef65306e64ba96b924656958f5cf8e8a00b26681ebd771b481e7254cde25a4fd91257e09d0607d0030f1bde3822f6d4eddff6944ea1043b21f5b08ac2c6bf332d61e0c000ef8e4d0830d46e097ca3347d88417de64d7f35c2dad439ac7183f48749b29e68d472d2611ec0d6d6927e26d0;
    5'b10110 : xpb = 1024'h5452abead27939bc807cd9936207e59d6393eed8e18cea993d7f47593cd3ffe49df77944c67cc73f5cd94ca6ed21a8fbca12eb4f2ae39cf703a34a5330d1d2e0d23f46093af83df2d0a0915e564e66604e28679f74de3851b94011c0cbb72acca72009fd75c238523a95303ac01055818a28d6b6f6f231bb1406f973135f9660;
    5'b10111 : xpb = 1024'h5827e246f35030b96f0e2948a0ab2a3bd0d4d6cb777069a034a7f9231caf172930c88a6acf8273369b40447ff7e9021e81cdf6014fbf69eaf82ab66e3eacd0d3c487f7c3d4ec40c3ab9097f9e5dd99933a700f3dfa2e239b41abb5781acb211bc5fe96149e053ae19a5626c90e9cb67bca9f0f0519719115094d1c0f944105f0;
    5'b11000 : xpb = 1024'h5bfd18a3142727b65d9f78fddf4e6eda3e15bebe0d53e8a72bd0aaecfc8a2e6dc3999b90d8881f2dd9a73c5902b05b41398900b3749b36deecb222894c87cec6b6d0a97e6ee0439486809e95756cccc626b7b6dc7f7e0ee4ca17592f69df176ae4dd222bc6483d70fa171d575d2917760b1547533bf0f06efe933eac15227580;
    5'b11001 : xpb = 1024'h5fd24eff34fe1eb34c30c8b31df1b378ab56a6b0a33767ae22f95cb6dc6545b2566aacb6e18dcb25180e34320d77b463f1440b65997703d2e1398ea45a62ccb9a9195b3908d446656170a53104fbfff912ff5e7b04cdfa2e5282fce6b8f30dba03bbae42ee8b400059d813e5abb578704b8b7fa15e704fc8f3d961489603e510;
    5'b11010 : xpb = 1024'h63a7855b55d515b03ac218685c94f81718978ea3391ae6b51a220e80bc405cf6e93bbddcea93771c56752c0b183f0d86a8ff1617be52d0c6d5c0fabf683dcaac9b620cf3a2c849363c60abcc948b332bff4706198a1de577daeea09e08070409229a3a5a16ce428fb9990a73fa41d96a8c01b7ef80efaf22e91f83e516e554a0;
    5'b11011 : xpb = 1024'h677cbbb776ac0cad2953681d9b383cb585d87695cefe65bc114ac04a9c1b743b7c0ccf02f399231394dc23e4230666a960ba20c9e32e9dbaca4866da7618c89f8daabeae3cbc4c071750b268241a665eeb8eadb80f6dd0c1635a4455571afa584178c6713f11451f195a010248ce3a64cc77f03da36f0e7cde65a68197c6c430;
    5'b11100 : xpb = 1024'h6b51f213978303aa17e4b7d2d9db8153f3195e8864e1e4c3087372147bf68b800edde028fc9ecf0ad3431bbd2dcdbfcc18752b7c080a6aaebecfd2f583f3c6927ff37068d6b04ed7f240b903b3a99991d7d6555694bdbc0aebc5e80ca62ef0a760575288675447ae791af790975a9b5f0cee288bc5ee6dd6d3abc91e18a833c0;
    5'b11101 : xpb = 1024'h6f27286fb859faa706760788187ec5f2605a467afac563c9ff9c23de5bd1a2c4a1aef14f05a47b0211aa1396389518eed030362e2ce637a2b3573f1091cec485723c222370a451a8cd30bf9f4338ccc4c41dfcf51a0da75474318bc3f542e6f67f35de9f8f974a3dd8dbee1ee5e6fc594d6460d9e86dcd30c8f1ebba9989a350;
    5'b11110 : xpb = 1024'h72fc5ecbd930f1a3f507573d57220a90cd9b2e6d90a8e2d0f6c4d5a83bacba09348002750eaa26f950110b6f435c721187eb40e051c20496a7deab2b9fa9c2786484d3de0a985479a820c63ad2c7fff7b065a4939f5d929dfc9d2f7b4456dd459e146ab6b7da4ccd389ce4ad34735d538dda99280aed2c8abe380e571a6b12e0;
    5'b11111 : xpb = 1024'h76d19527fa07e8a0e398a6f295c54f2f3adc1660268c61d7eded87721b87d14dc751139b17afd2f08e7803484e23cb343fa64b92769dd18a9c661746ad84c06b56cd8598a48c574a8310ccd66257332a9cad4c3224ad7de78508d332936ad394bcf2f6cde01d4f5c985ddb3b82ffbe4dce50d1762d6c8be4b37e30f39b4c8270;
    endcase
end

endmodule

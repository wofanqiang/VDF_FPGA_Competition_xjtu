module xpb_5_895
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5b9766e3231227e5cd8e6b60f6a12a4f42d745378555772b24e738906133c788d47c9aac76fb684d497579d696a497436a320a380f353e5ee379d3c6689e39eb8034f546a5a3142fcce95f7c4027ff7eb8f9c5d58289021b5d06291d85dcbbf678d86d2bcffcb6a1b2b6e796ea491b704d41feb05bac9d63d97ae9e3979a55d9;
    5'b00010 : xpb = 1024'h681887084361b02d0175eeadce80d4d1438873e35334ddecbf1b7cb0f64e209a5b0b7e023d0520bf38cb46649eb1dbc7049ec89fbb7ac721654682e9669ff258c1ab5de9bb52b1a8738bc55e7743acc7dee9212788bd726047fc040518ed55ac2a9482def3074b5deade84edcc210b74baa1e7e670ddd976c8658c2a6524547;
    5'b00011 : xpb = 1024'h6218ef53a74842e89da5ca4bd389379c570fcc75ba88c509f0d8f05b7098a9927a2d528c9acbba593d022e3ce08fb4ffda7bf6c20aecead0f9ce3bf4ff0839110c4fab2541583f4a54221bd2279c3a4b36e857e7fb14d9416185e95dd76b91513b81b559bf2d2b579164cfe5c70b2c2798ec1d2ec2ba7afb460142a63dec9b20;
    5'b00100 : xpb = 1024'hd0310e1086c3605a02ebdd5b9d01a9a28710e7c6a669bbd97e36f961ec9c4134b616fc047a0a417e71968cc93d63b78e093d913f76f58e42ca8d05d2cd3fe4b18356bbd376a56350e7178abcee87598fbdd2424f117ae4c08ff8080a31daab58552905bde60e96bbd5bd09db984216e97543cfcce1bbb2ed90cb1854ca48a8e;
    5'b00101 : xpb = 1024'h689a77c42b7e5deb6dbd2936b07144e96b4853b3efbc12e8bccaa8267ffd8b9c1fde0a6cbe9c0c65308ee2a32a7ad2bc4ac5e34c06a497431022a42395723836986a6103dd0d6a64db5ad8280f107517b4d6e9fa73a0b0676605a99e28fa66abfe2afd87ae5da00d7012b834a3cd3cdee4963bad29c85892b2879b68e43ee067;
    5'b00110 : xpb = 1024'h138499518ca2510870461cc096b827e73ca995ba9f99e99c63d527612e2ea61cf11227a06b70f623daa61d32ddc1593550ddc59df327055642fd388bc33dfd70a450219bd31f814f95aa3501b65cb06579cbb63769a385720d7f40c0f4ac801047fbd889cd915e219c09b8ec96463225e2fe5b7b352998c645930a47f2f6cfd5;
    5'b00111 : xpb = 1024'h6f1c0034afb478ee3dd488218d5952367f80daf224ef60c788bc5ff18f626da5c58ec24ce26c5e71241b97097465f078bb0fcfd6025c43b526770c522bdc375c248516e278c2957f6293947df684afe432c57c0cec2c878d6a8569de7a893c06c0d445b59d8e14c34ec0a083808f4d9630405a2b90d6362a1f0df42b8a9125ae;
    5'b01000 : xpb = 1024'h1a0621c210d86c0b405d7bab73a0353450e21cf8d4cd377b2fc6df2c3d93882696c2df808f41482fce32d19927ac76f1c127b227eedeb1c85951a0ba59a7fc96306ad77a6ed4ac6a1ce2f1579dd0eb31f7ba4849e22f5c9811ff0101463b556b0aa520b7bcc1d2d77ab7a13b730842dd2ea879f99c37765db219630a9949151c;
    5'b01001 : xpb = 1024'h759d88a533ea93f10debe70c6a415f8393b962305a22aea654ae17bc9ec74faf6b3f7a2d063cb07d17a84b6fbe510e352b59bc5ffe13f0273ccb7480c2463681b09fccc11477c099e9cc50d3ddf8eab0b0b40e1f64b85eb36f052a1ecc181161837d8de38cbe89792d6e88d25d515e4d7bea78a9f7e413c18b944cee30e36af5;
    5'b01010 : xpb = 1024'h2087aa32950e870e1074da9650884281651aa4370a008559fbb896f74cf86a303c739760b3119a3bc1bf85ff719794ae31719eb1ea965e3a6fa608e8f011fbbbbc858d590a89d784a41badad854525fe75a8da5c5abb33be167ec14197ca2ac5cd4e68e5abf2478d5965898a4fca53947a529878034553f51e9fbbcd3f9b5a63;
    5'b01011 : xpb = 1024'h7c1f1115b820aef3de0345f747296cd0a7f1e96e8f55fc85209fcf87ae2c31b910f0320d2a0d02890b34ffd6083c2bf19ba3a8e9f9cb9c99531fdcaf58b035a73cba829fb02cebb471050d29c56d257d2ea2a031dd4435d97384ea5f1da6e6bc4626d6117beefe2f0c1c71213a136f04c79497285ef1f158f81aa5b0d735b03c;
    5'b01100 : xpb = 1024'h270932a31944a210e08c39812d704fce79532b753f33d338c7aa4ec25c5d4c39e2244f40d6e1ec47b54c3a65bb82b26aa1bb8b3be64e0aac85fa7117867bfae148a04337a63f029f2b546a036cb960caf3976c6ed3470ae41afe8181e95900208ff7b1139b22bc43381371d92c8c644bc5fcb6f66a53318c8b26148fe5ed9faa;
    5'b01101 : xpb = 1024'h82a099863c56c9f6ae1aa4e224117a1dbc2a70acc4894a63ec918752bd9113c2b6a0e9ed4ddd5494fec1b43c522749ae0bed9573f583490b697444ddef1a34ccc8d5387e4be216cef83dc97face16049ac91324455d00cff7804aa9f6f35bc1708d01e3f6b1f72e4eaca597016d57fbc133eb5a6c5ffcef064a0fe737d87f583;
    5'b01110 : xpb = 1024'h2d8abb139d7abd13b0a3986c0a585d1b8d8bb2b374672117939c068d6bc22e4387d50720fab23e53a8d8eecc056dd027120577c5e205b71e9c4ed9461ce5fa06d4baf91641f42db9b28d2659542d9b977185fe814bd2e20a1f7e41c23ae7d57b52a0f9418a5330f916c15a28094e750311a6d574d1610f23f7ac6d528c3fe4f1;
    5'b01111 : xpb = 1024'h892221f6c08ce4f97e3203cd00f9876ad062f7eaf9bc9842b8833f1dccf5f5cc5c51a1cd71ada6a0f24e68a29c12676a7c3781fdf13af57d7fc8ad0c858433f254efee5ce79741e97f7685d594559b162a7fc456ce5be4257c846adfc0c49171cb79666d5a4fe79ac97841bef39790735ee8d4252d0dac87d127573623da3aca;
    5'b10000 : xpb = 1024'h340c438421b0d81680baf756e7406a68a1c439f1a99a6ef65f8dbe587b27104d2d85bf011e82905f9c65a3324f58ede3824f644fddbd6390b2a34174b34ff92c60d5aef4dda958d439c5e2af3ba1d663ef749093c45eb93023fe02028c76aad6154a416f7983a5aef56f4276e61085ba5d50f3f3386eecbb6432c61532922a38;
    5'b10001 : xpb = 1024'h8fa3aa6744c2fffc4e4962b7dde194b7e49b7f292eefe6218474f6e8dc5ad7d6020259ad957df8ace5db1d08e5fd8526ec816e87ecf2a1ef961d153b1bee3317e10aa43b834c6d0406af422b7bc9d5e2a86e566946e7bb4b81042b20125366cc8e22ae9b49805c50a8262a0dd059a12aaa92f2a3941b8a1f3dadaff8ca2c8011;
    5'b10010 : xpb = 1024'h3a8dcbf4a5e6f31950d25641c42877b5b5fcc12fdecdbcd52b7f76238a8bf256d33676e14252e26b8ff2579899440b9ff29950d9d9751002c8f7a9a349b9f851ecf064d3795e83eec0fe9f05231611306d6322a63cea9056287dc242de058030d7f3899d68b41a64d41d2ac5c2d29671a8fb12719f7cca52d0b91ed7d8e46f7f;
    5'b10011 : xpb = 1024'h962532d7c8f91aff1e60c1a2bac9a204f8d40667642334005066aeb3ebbfb9dfa7b3118db94e4ab8d967d16f2fe8a2e35ccb5b11e8aa4e61ac717d69b258323d6d255a1a1f01981e8de7fe81633e10af265ce87bbf7392718583eb6063e23c2750cbf6c938b0d10686d4125cad1bb1e1f63d1121fb2967b6aa3408bb707ec558;
    5'b10100 : xpb = 1024'h410f54652a1d0e1c20e9b52ca1108502ca35486e14010ab3f7712dee99f0d46078e72ec166233477837f0bfee32f295c62e33d63d52cbc74df4c11d1e023f777790b1ab21513af0948375b5b0a8a4bfceb51b4b8b576677c2cfd82832f94558b9a9cd1cb57e48f1ab2cb13149f94a728f4a530f0068aa7ea3d3f779a7f36b4c6;
    5'b10101 : xpb = 1024'h9ca6bb484d2f3601ee78208d97b1af520d0c8da5995681df1c58667efb249be94d63c96ddd1e9cc4ccf485d579d3c09fcd15479be461fad3c2c5e59848c23162f9400ff8bab6c3391520bad74ab24b7ba44b7a8e37ff69978a03aba0b571118213753ef727e145bc6581faab89ddc29941e72fa06237454e16ba617e16d10a9f;
    5'b10110 : xpb = 1024'h4790dcd5ae53291ef10114177df8924fde6dcfac49345892c362e5b9a955b66a1e97e6a189f38683770bc0652d1a4718d32d29edd0e468e6f5a07a00768df69d0525d090b0c8da23cf7017b0f1fe86c9694046cb2e023ea2317d42c381232ae65d4619f9471503d09178fb637c56b7e0404f4f6e6d988581a9c5d05d2588fa0d;
    5'b10111 : xpb = 1024'ha32843b8d1655104be8f7f787499bc9f214514e3ce89cfbde84a1e4a0a897df2f314814e00eeeed0c0813a3bc3bede5c3d5f3425e019a745d91a4dc6df2c3088855ac5d7566bee539c59772d32268648223a0ca0b08b40bd8e836be106ffe6dcd61e87251711ba72442fe2fa669fd3508d914e1ec94522e58340ba40bd234fe6;
    5'b11000 : xpb = 1024'h4e12654632894421c11873025ae09f9cf2a656ea7e67a6718f549d84b8ba9873c4489e81adc3d88f6a9874cb770564d543771677cc9c15590bf4e22f0cf7f5c29140866f4c7e053e56a8d406d972c195e72ed8dda68e15c835fd0303d2b200411fef6227364578867026e3b25918c8978bf96decd4a66319164c291fcbdb3f54;
    5'b11001 : xpb = 1024'ha9a9cc29559b6c078ea6de635181c9ec357d9c2203bd1d9cb43bd61519ee5ffc98c5392e24bf40dcb40deea20da9fc18ada920afdbd153b7ef6eb5f575962fae11757bb5f221196e23923383199ac114a0289eb3291717e393032c21588ebc3798c7cf5306422f2822ddcb494361e407d93b6c9d3053007cefc713036375952d;
    5'b11010 : xpb = 1024'h5493edb6b6bf5f24912fd1ed37c8acea06dede28b39af4505b46554fc81f7a7d69f95661d1942a9b5e252931c0f08291b3c10301c853c1cb22494a5da361f4e81d5b3c4de8333058dde1905cc0e6fc62651d6af01f19ecee3a7cc3442440d59be298aa552575ed3c4ed4cc0135dad94ed7a38c6b3bb440b082d281e2722d849b;
    5'b11011 : xpb = 1024'hb02b5499d9d1870a5ebe3d4e2e69d73949b6236038f06b7b802d8de0295342063e75f10e488f92e8a79aa308579519d51df30d39d789002a05c31e240c002ed39d9031948dd64488aacaefd9010efbe11e1730c5a1a2ef099782ec61aa1d91925b711780f572a3de018bb3982023f4bf24e58b1b9760de145c4d6bc609c7da74;
    5'b11100 : xpb = 1024'h5b1576273af57a27614730d814b0ba371b176566e8ce422f27380d1ad7845c870faa0e41f5647ca751b1dd980adba04e240aef8bc40b6e3d389db28c39cbf40da975f22c83e85b73651a4cb2a85b372ee30bfd0297a5c4143efc838475cfaaf6a541f28314a661f22d82b450129cea06234daae9a2c21e47ef58daa5187fc9e2;
    5'b11101 : xpb = 1024'h5ff97b49c196d4463d02461faf79d34ec78a76d98ac18e2ce428c5585b57707e0de2b75a2396665fbc91827be2226c72a22d1ddb08ddc506b7846f46797b947b55bb2c479fa725e1f69a98c4fa7727ca800c93f8da8991ee6761aa74181c45aef12cd8533da20065979b5080515df4d21b5cab7ae235e7b826449842737b950;
    5'b11110 : xpb = 1024'h6196fe97bf2b952a315e8fc2f198c7842f4feca51e01900df329c4e5e6e93e90b55ac6221934ceb3453e91fe54c6be0a9454dc15bfc31aaf4ef21abad035f3333590a80b1f9d868dec5309088fcf71fb60fa8f1510319b3a437c43c4c75e805167eb3ab103d6d6a80c309c9eef5efabd6ef7c96809cffbdf5bdf3367bed20f29;
    5'b11111 : xpb = 1024'hc812025204f884733e7834cd7dfaa8200b12eabcddf66c19a344420951a5911868ee355c609b871ef55cc8e080d44839a6cbe67ac4588c281ccaf22fe01b86d417668a315af9d78a6a265e2371bad4925ef5b5206347044eaf5dae7931099b5b1bc15b3230a94bc38279d56e1d7f0046d5fe93615313c12eeeaa246cd89fe97;
    endcase
end

endmodule

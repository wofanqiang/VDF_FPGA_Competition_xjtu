/*******************************************************************************
  Copyright 2019 xjtu

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
*******************************************************************************/

module xpb_lut_low
(
    input logic [16:0] flag[3],
    output logic [1023:0] xpb[9]
);
        
        
    always_comb begin
        case(flag[0][5:0])
            6'd0: xpb[0] = 1024'd0;
            6'd1: xpb[0] = 1024'd55702617802106849374131591674088040617099270768494973145298226092755780468191824222693406107749861711676964472413899923079725927973196287937687305623143083444077218855294267938671980409728888398142885343697765922473789832121566108508934540857597787896530607270469240209840717864551083287716666502998629652885;
            6'd2: xpb[0] = 1024'd111405235604213698748263183348176081234198541536989946290596452185511560936383648445386812215499723423353928944827799846159451855946392575875374611246286166888154437710588535877343960819457776796285770687395531844947579664243132217017869081715195575793061214540938480419681435729102166575433333005997259305770;
            6'd3: xpb[0] = 1024'd43041157722195806723595847617449689106599385179749235307762823213290446067266333758065147108591910825587744009784206334660113943078368529257901791853098209398540981996311586478385702037669459473118458422706057921057008646143801552561825052889563914422771918397290662599415625519724616846031309682370294474324;
            6'd4: xpb[0] = 1024'd98743775524302656097727439291537729723698655948244208453061049306046226535458157980758553216341772537264708482198106257739839871051564817195589097476241292842618200851605854417057682447398347871261343766403823843530798478265367661070759593747161702319302525667759902809256343384275700133747976185368924127209;
            6'd5: xpb[0] = 1024'd30379697642284764073060103560811337596099499591003497470227420333825111666340843293436888109433959939498523547154512746240501958183540770578116278083053335353004745137328905018099423665610030548094031501714349919640227460166036996614715564921530040949013229524112084988990533174898150404345952861741959295763;
            6'd6: xpb[0] = 1024'd86082315444391613447191695234899378213198770359498470615525646426580892134532667516130294217183821651175488019568412669320227886156737058515803583706196418797081963992623172956771404075338918946236916845412115842114017292287603105123650105779127828845543836794581325198831251039449233692062619364740588948648;
            6'd7: xpb[0] = 1024'd17718237562373721422524359504172986085599614002257759632692017454359777265415352828808629110276009053409303084524819157820889973288713011898330764313008461307468508278346223557813145293550601623069604580722641918223446274188272440667606076953496167475254540650933507378565440830071683962660596041113624117202;
            6'd8: xpb[0] = 1024'd73420855364480570796655951178261026702698884770752732777990243547115557733607177051502035218025870765086267556938719080900615901261909299836018069936151544751545727133640491496485125703279490021212489924420407840697236106309838549176540617811093955371785147921402747588406158694622767250377262544112253770087;
            6'd9: xpb[0] = 1024'd5056777482462678771988615447534634575099728413512021795156614574894442864489862364180370111118058167320082621895125569401277988393885253218545250542963587261932271419363542097526866921491172698045177659730933916806665088210507884720496588985462294001495851777754929768140348485245217520975239220485288938641;
            6'd10: xpb[0] = 1024'd60759395284569528146120207121622675192198999182006994940454840667650223332681686586873776218867919878997047094309025492481003916367081541156232556166106670706009490274657810036198847331220061096188063003428699839280454920332073993229431129843060081898026459048224169977981066349796300808691905723483918591526;
            6'd11: xpb[0] = 1024'd116462013086676377520251798795710715809298269950501968085753066760406003800873510809567182326617781590674011566722925415560729844340277829093919861789249754150086709129952077974870827740948949494330948347126465761754244752453640101738365670700657869794557066318693410187821784214347384096408572226482548244411;
            6'd12: xpb[0] = 1024'd48097935204658485495584463064984323681699113593261257102919437788184888931756196122245517219709968992907826631679331904061391931472253782476447042396061796660473253415675128575912568959160632171163636082436991837863673734354309437282321641875026208424267770175045592367555974004969834367006548902855583412965;
            6'd13: xpb[0] = 1024'd103800553006765334869716054739072364298798384361756230248217663880940669399948020344938923327459830704584791104093231827141117859445450070414134348019204880104550472270969396514584549368889520569306521426134757760337463566475875545791256182732623996320798377445514832577396691869520917654723215405854213065850;
            6'd14: xpb[0] = 1024'd35436475124747442845048719008345972171199228004515519265384034908719554530830705657617258220552018106818606169049638315641779946577426023796661528626016922614937016556692447115626290587101203246139209161445283836446892548376544881335212153906992334950509081301867014757130881660143367925321192082227248234404;
            6'd15: xpb[0] = 1024'd91139092926854292219180310682434012788298498773010492410682261001475334999022529880310664328301879818495570641463538238721505874550622311734348834249160006059014235411986715054298270996830091644282094505143049758920682380498110989844146694764590122847039688572336254966971599524694451213037858585225877887289;
            6'd16: xpb[0] = 1024'd22775015044836400194512974951707620660699342415769781427848632029254220129905215192988999221394067220729385706419944727222167961682598265116876014855972048569400779697709765655340012215041774321114782240453575835030111362398780325388102665938958461476750392428688437146705789315316901483635835261598913055843;
            6'd17: xpb[0] = 1024'd78477632846943249568644566625795661277798613184264754573146858122010000598097039415682405329143928932406350178833844650301893889655794553054563320479115132013477998553004033594011992624770662719257667584151341757503901194520346433897037206796556249373280999699157677356546507179867984771352501764597542708728;
            6'd18: xpb[0] = 1024'd10113554964925357543977230895069269150199456827024043590313229149788885728979724728360740222236116334640165243790251138802555976787770506437090501085927174523864542838727084195053733842982345396090355319461867833613330176421015769440993177970924588002991703555509859536280696970490435041950478440970577877282;
            6'd19: xpb[0] = 1024'd65816172767032206918108822569157309767298727595519016735611455242544666197171548951054146329985978046317129716204151061882281904760966794374777806709070257967941761694021352133725714252711233794233240663159633756087120008542581877949927718828522375899522310825979099746121414835041518329667144943969207530167;
            6'd20: xpb[0] = 1024'd121518790569139056292240414243245350384397998364013989880909681335300446665363373173747552437735839757994094188618050984962007832734163082312465112332213341412018980549315620072397694662440122192376126006857399678560909840664147986458862259686120163796052918096448339955962132699592601617383811446967837183052;
            6'd21: xpb[0] = 1024'd53154712687121164267573078512518958256798842006773278898076052363079331796246058486425887330828027160227909253574457473462669919866139035694992292939025383922405524835038670673439435880651804869208813742167925754670338822564817322002818230860488502425763621952800522135696322490215051887981788123340872351606;
            6'd22: xpb[0] = 1024'd108857330489228013641704670186606998873898112775268252043374278455835112264437882709119293438577888871904873725988357396542395847839335323632679598562168467366482743690332938612111416290380693267351699085865691677144128654686383430511752771718086290322294229223269762345537040354766135175698454626339502004491;
            6'd23: xpb[0] = 1024'd40493252607210121617037334455880606746298956418027541060540649483613997395320568021797628331670076274138688790944763885043057934971311277015206779168980509876869287976055989213153157508592375944184386821176217753253557636587052766055708742892454628952004933079621944525271230145388585446296431302712537173045;
            6'd24: xpb[0] = 1024'd96195870409316970991168926129968647363398227186522514205838875576369777863512392244491034439419937985815653263358663808122783862944507564952894084792123593320946506831350257151825137918321264342327272164873983675727347468708618874564643283750052416848535540350091184735111948009939668734013097805711166825930;
            6'd25: xpb[0] = 1024'd27831792527299078966501590399242255235799070829281803223005246604148662994395077557169369332512125388049468328315070296623445950076483518335421265398935635831333051117073307752866879136532947019159959900184509751836776450609288210108599254924420755478246244206443366914846137800562119004611074482084201994484;
            6'd26: xpb[0] = 1024'd83534410329405928340633182073330295852898341597776776368303472696904443462586901779862775440261987099726432800728970219703171878049679806273108571022078719275410269972367575691538859546261835417302845243882275674310566282730854318617533795782018543374776851476912607124686855665113202292327740985082831647369;
            6'd27: xpb[0] = 1024'd15170332447388036315965846342603903725299185240536065385469843724683328593469587092541110333354174501960247865685376708203833965181655759655635751628890761785796814258090626292580600764473518094135532979192801750419995264631523654161489766956386882004487555333264789304421045455735652562925717661455866815923;
            6'd28: xpb[0] = 1024'd70872950249494885690097438016691944342398456009031038530768069817439109061661411315234516441104036213637212338099276631283559893154852047593323057252033845229874033113384894231252581174202406492278418322890567672893785096753089762670424307813984669901018162603734029514261763320286735850642384164454496468808;
            6'd29: xpb[0] = 1024'd2508872367476993665430102285965552214799299651790327547934440845217994192544096627912851334196223615871027403055683119784221980286828000975850237858845887740260577399107944832294322392414089169111106058201093749003214078653759098214380278988353008530728866460086211693995953110909186121240360840827531637362;
            6'd30: xpb[0] = 1024'd58211490169583843039561693960053592831898570420285300693232666937973774660735920850606257441946085327547991875469583042863947908260024288913537543481988971184337796254402212770966302802142977567253991401898859671477003910775325206723314819845950796427259473730555451903836670975460269408957027343826161290247;
            6'd31: xpb[0] = 1024'd113914107971690692413693285634141633448997841188780273838530893030729555128927745073299663549695947039224956347883482965943673836233220576851224849105132054628415015109696480709638283211871865965396876745596625593950793742896891315232249360703548584323790081001024692113677388840011352696673693846824790943132;
            6'd32: xpb[0] = 1024'd45550030089672800389025949903415241321398684831539562855697264058508440259810430385977998442788134441458771412839889454444335923365196530233752029711944097138801559395419531310680024430083548642229564480907151670060222724797560650776205331877916922953500784857376874293411578630633802967271670523197826111686;
            6'd33: xpb[0] = 1024'd101252647891779649763157541577503281938497955600034536000995490151264220728002254608671404550537996153135735885253789377524061851338392818171439335335087180582878778250713799249352004839812437040372449824604917592534012556919126759285139872735514710850031392127846114503252296495184886254988337026196455764571;
            6'd34: xpb[0] = 1024'd32888570009761757738490205846776889810898799242793825018161861179043105858884939921349739443630183555369550950210195866024723938470368771553966515941899223093265322536436849850393746058024119717205137559915443668643441538819796094829095843909883049479742095984198296682986486285807336525586313702569490933125;
            6'd35: xpb[0] = 1024'd88591187811868607112621797520864930427998070011288798163460087271798886327076764144043145551380045267046515422624095789104449866443565059491653821565042306537342541391731117789065726467753008115348022903613209591117231370941362203338030384767480837376272703254667536892827204150358419813302980205568120586010;
            6'd36: xpb[0] = 1024'd20227109929850715087954461790138538300398913654048087180626458299577771457959449456721480444472232669280330487580502277605111953575541012874181002171854349047729085677454168390107467685964690792180710638923735667226660352842031538881986355941849176005983407111019719072561393940980870083900956881941155754564;
            6'd37: xpb[0] = 1024'd75929727731957564462086053464226578917498184422543060325924684392333551926151273679414886552222094380957294959994402200684837881548737300811868307794997432491806304532748436328779448095693579190323595982621501589700450184963597647390920896799446963902514014381488959282402111805531953371617623384939785407449;
            6'd38: xpb[0] = 1024'd7565649849939672437418717733500186789899028065302349343091055420112437057033958992093221445314281783191110024950808689185499968680713254194395488401809475002192848818471486929821189313905261867156283717932027665809879166864266982934876867973815302532224718237841141462136301596154403642215600061312820576003;
            6'd39: xpb[0] = 1024'd63268267652046521811550309407588227406998298833797322488389281512868217525225783214786627553064143494868074497364708612265225896653909542132082794024952558446270067673765754868493169723634150265299169061629793588283668998985833091443811408831413090428755325508310381671977019460705486929932266564311450228888;
            6'd40: xpb[0] = 1024'd118970885454153371185681901081676268024097569602292295633687507605623997993417607437480033660814005206545038969778608535344951824627105830069770099648095641890347286529060022807165150133363038663442054405327559510757458831107399199952745949689010878325285932778779621881817737325256570217648933067310079881773;
            6'd41: xpb[0] = 1024'd50606807572135479161014565350949875896498413245051584650853878633402883124300292750158368553906192608778854034735015023845613911759081783452297280254907684400733830814783073408206891351574721340274742140638085586866887813008068535496701920863379216954996636635131804061551927115879020488246909743683115050327;
            6'd42: xpb[0] = 1024'd106309425374242328535146157025037916513597684013546557796152104726158663592492116972851774661656054320455818507148914946925339839732278071389984585878050767844811049670077341346878871761303609738417627484335851509340677645129634644005636461720977004851527243905601044271392644980430103775963576246681744703212;
            6'd43: xpb[0] = 1024'd37945347492224436510478821294311524385998527656305846813318475753937548723374802285530109554748241722689633572105321435426001926864254024772511766484862810355197593955800391947920612979515292415250315219646377585450106627030303979549592432895345343481237947761953226451126834771052554046561552923054779871766;
            6'd44: xpb[0] = 1024'd93647965294331285884610412968399565003097798424800819958616701846693329191566626508223515662498103434366598044519221358505727854837450312710199072108005893799274812811094659886592593389244180813393200563344143507923896459151870088058526973752943131377768555032422466660967552635603637334278219426053409524651;
            6'd45: xpb[0] = 1024'd25283887412313393859943077237673172875498642067560108975783072874472214322449311820901850555590290836600413109475627847006389941969426266092726252714817936309661357096817710487634334607455863490225888298654669584033325441052539423602482944927311470007479258888774648840701742426226087604876196102426444693205;
            6'd46: xpb[0] = 1024'd80986505214420243234074668911761213492597912836055082121081298967227994790641136043595256663340152548277377581889527770086115869942622554030413558337961019753738575952111978426306315017184751888368773642352435506507115273174105532111417485784909257904009866159243889050542460290777170892592862605425074346090;
            6'd47: xpb[0] = 1024'd12622427332402351209407333181034821364998756478814371138247669995006879921523821356273591556432339950511192646845934258586777957074598507412940738944773062264125120237835029027348056235396434565201461377662961582616544255074774867655373456959277596533720570015596071230276650081399621163190839281798109514644;
            6'd48: xpb[0] = 1024'd68325045134509200583538924855122861982098027247309344283545896087762660389715645578966997664182201662188157119259834181666503885047794795350628044567916145708202339093129296966020036645125322963344346721360727505090334087196340976164307997816875384430251177286065311440117367945950704450907505784796739167529;
            6'd49: xpb[0] = 1024'd124027662936616049957670516529210902599197298015804317428844122180518440857907469801660403771932063373865121591673734104746229813020991083288315350191059229152279557948423564904692017054854211361487232065058493427564123919317907084673242538674473172326781784556534551649958085810501787738624172287795368820414;
            6'd50: xpb[0] = 1024'd55663585054598157933003180798484510471598141658563606446010493208297325988790155114338738665024250776098936656630140593246891900152967036670842530797871271662666102234146615505733758273065894038319919800369019503673552901218576420217198509848841510956492488412886733829692275601124238009222148964168403988968;
            6'd51: xpb[0] = 1024'd111366202856705007307134772472572551088697412427058579591308719301053106456981979337032144772774112487775901129044040516326617828126163324608529836421014355106743321089440883444405738682794782436462805144066785426147342733340142528726133050706439298853023095683355974039532993465675321296938815467167033641853;
            6'd52: xpb[0] = 1024'd43002124974687115282467436741846158961098256069817868608475090328831991587864664649710479665866299890009716194000447004827279915258139277991057017027826397617129865375163934045447479901006465113295492879377311502256771715240811864270089021880807637482733799539708156219267183256297771567536792143540068810407;
            6'd53: xpb[0] = 1024'd98704742776793964656599028415934199578197526838312841753773316421587772056056488872403885773616161601686680666414346927907005843231335565928744322650969481061207084230458201984119460310735353511438378223075077424730561547362377972779023562738405425379264406810177396429107901120848854855253458646538698463292;
            6'd54: xpb[0] = 1024'd30340664894776072631931692685207807450598370481072130770939687449366657186939174185082220666708349003920495731370753416407667930363311519311271503257781523571593628516181252585161201528947036188271065958385603500839990529263047308322979533912773764008975110666529578608842090911471305125851435322911733631846;
            6'd55: xpb[0] = 1024'd86043282696882922006063284359295848067697641249567103916237913542122437655130998407775626774458210715597460203784653339487393858336507807248958808880924607015670847371475520523833181938675924586413951302083369423313780361384613416831914074770371551905505717936998818818682808776022388413568101825910363284731;
            6'd56: xpb[0] = 1024'd17679204814865029981395948628569455940098484892326392933404284569901322786013683720453961667550398117831275268741059827988055945468483760631485989487736649526057391657198571124874923156887607263246639037393895499423209343285282752375870045944739890535216421793351000998416998566644838684166078502283398453285;
            6'd57: xpb[0] = 1024'd73381822616971879355527540302657496557197755660821366078702510662657103254205507943147367775300259829508239741154959751067781873441680048569173295110879732970134610512492839063546903566616495661389524381091661421896999175406848860884804586802337678431747029063820241208257716431195921971882745005282028106170;
            6'd58: xpb[0] = 1024'd5017744734953987330860204571931104429598599303580655095868881690435988385088193255825702668392447231742054806111366239568443960573656001951700475717691775480521154798215889664588644784828178338222212116402187498006428157307518196428760557976706017061457732920172423387991906221818372242480721681655063274724;
            6'd59: xpb[0] = 1024'd60720362537060836704991796246019145046697870072075628241167107783191768853280017478519108776142308943419019278525266162648169888546852289889387781340834858924598373653510157603260625194557066736365097460099953420480217989429084304937695098834303804957988340190641663597832624086369455530197388184653692927609;
            6'd60: xpb[0] = 1024'd116422980339167686079123387920107185663797140840570601386465333875947549321471841701212514883892170655095983750939166085727895816520048577827075086963977942368675592508804425541932605604285955134507982803797719342954007821550650413446629639691901592854518947461110903807673341950920538817914054687652322580494;
            6'd61: xpb[0] = 1024'd48058902457149794054456052189380793536197984483329890403631704903726434452354527013890849776984358057329798815895572574228557903652024531209602267570789984879062136794527476142974346822497637811340670539108245419063436803451319748990585610866269931484229651317463085987407531741542989088512031364025357749048;
            6'd62: xpb[0] = 1024'd103761520259256643428587643863468834153297255251824863548929930996482214920546351236584255884734219769006763288309472497308283831625220819147289573193933068323139355649821744081646327232226526209483555882806011341537226635572885857499520151723867719380760258587932326197248249606094072376228697867023987401933;
            6'd63: xpb[0] = 1024'd35397442377238751403920308132742442025698098894584152566096302024261100051429036549262590777826407171240578353265878985808945918757196772529816753800745110833525899935544794682688068450438208886316243618116537417646655617473555193043476122898236058010470962444284508376982439396716522646826674543397022570487;
        endcase
    end

    always_comb begin
        case(flag[0][11:6])
            6'd0: xpb[1] = 1024'd0;
            6'd1: xpb[1] = 1024'd91100060179345600778051899806830482642797369663079125711394528117016880519620860771955996885576268882917542825679778908888671846730393060467504059423888194277603118790839062621360048860167097284459128961814303340120445449595121301552410663755833845907001569714753748586823157261267605934543341046395652223372;
            6'd2: xpb[1] = 1024'd58133424674566460157304872208846532540896312200422567294657201169056865701932582633896922556494863456391936243902064383198279852619565786379847993831445347621515563012106907905089858528816988847608060315241366833876530048969345830139842757828438242547183236015390439143539786448606578851967992266165709962413;
            6'd3: xpb[1] = 1024'd25166789169787319536557844610862582438995254737766008877919874221096850884244304495837848227413458029866329662124349857507887858508738512292191928239002500965428007233374753188819668197466880410756991668668430327632614648343570358727274851901042639187364902316027129700256415635945551769392643485935767701454;
            6'd4: xpb[1] = 1024'd116266849349132920314609744417693065081792624400845134589314402338113731403865165267793845112989726912783872487804128766396559705239131572759695987662890695243031126024213815810179717057633977695216120630482733667753060097938691660279685515656876485094366472030780878287079572897213157703935984532331419924826;
            6'd5: xpb[1] = 1024'd83300213844353779693862716819709114979891566938188576172577075390153716586176887129734770783908321486258265906026414240706167711128304298672039922070447848586943570245481661093909526726283869258365051983909797161509144697312916188867117609729480881734548138331417568843796202084552130621360635752101477663867;
            6'd6: xpb[1] = 1024'd50333578339574639073115689221725164877990509475532017755839748442193701768488608991675696454826916059732659324248699715015775717017477024584383856478005001930856014466749506377639336394933760821513983337336860655265229296687140717454549703802085278374729804632054259400512831271891103538785286971871535402908;
            6'd7: xpb[1] = 1024'd17366942834795498452368661623741214776089452012875459339102421494233686950800330853616622125745510633207052742470985189325383722906649750496727790885562155274768458688017351661369146063583652384662914690763924149021313896061365246041981797874689675014911470932690949957229460459230076456209938191641593141949;
            6'd8: xpb[1] = 1024'd108467003014141099230420561430571697418886821675954585050496949611250567470421191625572619011321779516124595568150764098214055569637042810964231850309450349552371577478856414282729194923750749669122043652578227489141759345656486547594392461630523520921913040647444698544052617720497682390753279238037245365321;
            6'd9: xpb[1] = 1024'd75500367509361958609673533832587747316985764213298026633759622663290552652732913487513544682240374089598988986373049572523663575526215536876575784717007502896284021700124259566459004592400641232270975006005290982897843945030711076181824555703127917562094706948081389100769246907836655308177930457807303104362;
            6'd10: xpb[1] = 1024'd42533732004582817988926506234603797215084706750641468217022295715330537835044635349454470353158968663073382404595335046833271581415388262788919719124564656240196465921392104850188814261050532795419906359432354476653928544404935604769256649775732314202276373248718079657485876095175628225602581677577360843403;
            6'd11: xpb[1] = 1024'd9567096499803677368179478636619847113183649287984909800284968767370523017356357211395396024077563236547775822817620521142879587304560988701263653532121809584108910142659950133918623929700424358568837712859417970410013143779160133356688743848336710842458039549354770214202505282514601143027232897347418582444;
            6'd12: xpb[1] = 1024'd100667156679149278146231378443450329755981018951064035511679496884387403536977217983351392909653832119465318648497399430031551434034954049168767712956010003861712028933499012755278672789867521643027966674673721310530458593374281434909099407604170556749459609264108518801025662543782207077570573943743070805816;
            6'd13: xpb[1] = 1024'd67700521174370137525484350845466379654079961488407477094942169936427388719288939845292318580572426692939712066719684904341159439924126775081111647363567157205624473154766858039008482458517413206176898028100784804286543192748505963496531501676774953389641275564745209357742291731121179994995225163513128544857;
            6'd14: xpb[1] = 1024'd34733885669590996904737323247482429552178904025750918678204842988467373901600661707233244251491021266414105484941970378650767445813299500993455581771124310549536917376034703322738292127167304769325829381527848298042627792122730492083963595749379350029822941865381899914458920918460152912419876383283186283898;
            6'd15: xpb[1] = 1024'd1767250164811856283990295649498479450277846563094360261467516040507359083912383569174169922409615839888498903164255852960375451702472226905799516178681463893449361597302548606468101795817196332474760734954911791798712391496955020671395689821983746670004608166018590471175550105799125829844527603053244022939;
            6'd16: xpb[1] = 1024'd92867310344157457062042195456328962093075216226173485972862044157524239603533244341130166807985884722806041728844034761849047298432865287373303575602569658171052480388141611227828150655984293616933889696769215131919157841092076322223806353577817592577006177880772339057998707367066731764387868649448896246311;
            6'd17: xpb[1] = 1024'd59900674839378316441295167858345011991174158763516927556124717209564224785844966203071092478904479296280435147066320236158655304322038013285647510010126811514964924609409456511557960324634185180082821050196278625675242440466300850811238447650421989217187844181409029614715336554405704681812519869218953985352;
            6'd18: xpb[1] = 1024'd26934039334599175820548140260361061889273101300860369139387390261604209968156688065012018149823073869754828565288605710468263310211210739197991444417683964858877368830677301795287769993284076743231752403623342119431327039840525379398670541723026385857369510482045720171431965741744677599237171088989011724393;
            6'd19: xpb[1] = 1024'd118034099513944776598600040067191544532070470963939494850781918378621090487777548836968015035399342752672371390968384619356935156941603799665495503841572159136480487621516364416647818853451174027690881365437645459551772489435646680951081205478860231764371080196799468758255123003012283533780512135384663947765;
            6'd20: xpb[1] = 1024'd85067464009165635977853012469207594430169413501282936434044591430661075670089270698908940706317937326146764809190670093666543162830776525577839438249129312480392931842784209700377628522101065590839812718864708953307857088809871209538513299551464628404552746497436159314971752190351256451205163355154721686806;
            6'd21: xpb[1] = 1024'd52100828504386495357105984871223644328268356038626378017307264482701060852400992560849866377236531899621158227412955567976151168719949251490183372656686465824305376064052054984107438190750957153988744072291772447063941688184095738125945393624069025044734412798072849871688381377690229368629814574924779425847;
            6'd22: xpb[1] = 1024'd19134192999607354736358957273239694226367298575969819600569937534741046034712714422790792048155126473095551645635241042285759174609121977402527307064243619168217820285319900267837247859400848717137675425718835940820026287558320266713377487696673421684916079098709540428405010565029202286054465794694837164888;
            6'd23: xpb[1] = 1024'd110234253178952955514410857080070176869164668239048945311964465651757926554333575194746788933731395356013094471315019951174431021339515037870031366488131813445820939076158962889197296719567946001596804387533139280940471737153441568265788151452507267591917648813463289015228167826296808220597806841090489388260;
            6'd24: xpb[1] = 1024'd77267617674173814893663829482086226767263610776392386895227138703797911736645297056687714604649989929487487889537305425484039027228687763782375300895688966789733383297426808172927106388217837564745735740960202774696556336527666096853220245525111664232099315114099979571944797013635781138022458060860547127301;
            6'd25: xpb[1] = 1024'd44300982169394674272916801884102276665362553313735828478489811755837896918957018918628640275568584502961881307759590899793647033117860489694719235303246120133645827518694653456656916056867729127894667094387266268452640935901890625440652339597716060872280981414736670128661426200974754055447109280630604866342;
            6'd26: xpb[1] = 1024'd11334346664615533652169774286118326563461495851079270061752484807877882101268740780569565946487179076436274725981876374103255039007033215607063169710803273477558271739962498740386725725517620691043598447814329762208725535276115154028084433670320457512462647715373360685378055388313726972871760500400662605383;
            6'd27: xpb[1] = 1024'd102434406843961134430221674092948809206258865514158395773147012924894762620889601552525562832063447959353817551661655282991926885737426276074567229134691467755161390530801561361746774585684717975502727409628633102329170984871236455580495097426154303419464217430127109272201212649581332907415101546796314828755;
            6'd28: xpb[1] = 1024'd69467771339181993809474646494964859104357808051501837356409685976934747803201323414466488502982042532828210969883940757301534891626599001986911163542248621099073834752069406645476584254334609538651658763055696596085255584245460984167927191498758700059645883730763799828917841836920305824839752766566372567796;
            6'd29: xpb[1] = 1024'd36501135834402853188727618896980909002456750588845278939672359028974732985513045276407414173900637106302604388106226231611142897515771727899255097949805774442986278973337251929206393922984501101800590116482760089841340183619685512755359285571363096699827550031400490385634471024259278742264403986336430306837;
            6'd30: xpb[1] = 1024'd3534500329623712567980591298996958900555693126188720522935032081014718167824767138348339844819231679776997806328511705920750903404944453811599032357362927786898723194605097212936203591634392664949521469909823583597424782993910041342791379643967493340009216332037180942351100211598251659689055206106488045878;
            6'd31: xpb[1] = 1024'd94634560508969313346032491105827441543353062789267846234329560198031598687445627910304336730395500562694540632008290614809422750135337514279103091781251122064501841985444159834296252451801489949408650431724126923717870232589031342895202043399801339247010786046790929529174257472865857594232396252502140269250;
            6'd32: xpb[1] = 1024'd61667925004190172725285463507843491441452005326611287817592233250071583869757349772245262401314095136168934050230576089119030756024510240191447026188808275408414286206712005118026062120451381512557581785151190417473954831963255871482634137472405735887192452347427620085890886660204830511657047472272198008291;
            6'd33: xpb[1] = 1024'd28701289499411032104538435909859541339550947863954729400854906302111569052069071634186188072232689709643327468452861563428638761913682966103790960596365428752326730427979850401755871789101273075706513138578253911230039431337480400070066231545010132527374118648064310642607515847543803429081698692042255747332;
            6'd34: xpb[1] = 1024'd119801349678756632882590335716690023982348317527033855112249434419128449571689932406142184957808958592560870294132640472317310608644076026571295020020253623029929849218818913023115920649268370360165642100392557251350484880932601701622476895300843978434375688362818059229430673108811409363625039738437907970704;
            6'd35: xpb[1] = 1024'd86834714173977492261843308118706073880447260064377296695512107471168434754001654268083110628727553166035263712354925946626918614533248752483638954427810776373842293440086758306845730317918261923314573453819620745106569480306826230209908989373448375074557354663454749786147302296150382281049690958207965709745;
            6'd36: xpb[1] = 1024'd53868078669198351641096280520722123778546202601720738278774780523208419936313376130024036299646147739509657130577211420936526620422421478395982888835367929717754737661354603590575539986568153486463504807246684238862654079681050758797341083446052771714739020964091440342863931483489355198474342177978023448786;
            6'd37: xpb[1] = 1024'd20901443164419211020349252922738173676645145139064179862037453575248405118625097991964961970564742312984050548799496895246134626311594204308326823242925083061667181882622448874305349655218045049612436160673747732618738679055275287384773177518657168354920687264728130899580560670828328115898993397748081187827;
            6'd38: xpb[1] = 1024'd112001503343764811798401152729568656319442514802143305573431981692265285638245958763920958856141011195901593374479275804134806473041987264775830882666813277339270300673461511495665398515385142334071565122488051072739184128650396588937183841274491014261922256979481879486403717932095934050442334444143733411199;
            6'd39: xpb[1] = 1024'd79034867838985671177654125131584706217541457339486747156694654744305270820557680625861884527059605769375986792701561278444414478931159990688174817074370430683182744894729356779395208184035033897220496475915114566495268728024621117524615935347095410902103923280118570043120347119434906967866985663913791150240;
            6'd40: xpb[1] = 1024'd46068232334206530556907097533600756115640399876830188739957327796345256002869402487802810197978200342850380210923846752754022484820332716600518751481927584027095189115997202063125017852684925460369427829342178060251353327398845646112048029419699807542285589580755260599836976306773879885291636883683848889281;
            6'd41: xpb[1] = 1024'd13101596829427389936160069935616806013739342414173630323220000848385241185181124349743735868896794916324773629146132227063630490709505442512862685889484737371007633337265047346854827521334817023518359182769241554007437926773070174699480123492304204182467255881391951156553605494112852802716288103453906628322;
            6'd42: xpb[1] = 1024'd104201657008772990714211969742447288656536712077252756034614528965402121704801985121699732754473063799242316454825911135952302337439898502980366745313372931648610752128104109968214876381501914307977488144583544894127883376368191476251890787248138050089468825596145699743376762755380458737259629149849558851694;
            6'd43: xpb[1] = 1024'd71235021503993850093464942144463338554635654614596197617877202017442106887113706983640658425391658372716709873048196610261910343329071228892710679720930084992523196349371955251944686050151805871126419498010608387883967975742416004839322881320742446729650491896782390300093391942719431654684280369619616590735;
            6'd44: xpb[1] = 1024'd38268385999214709472717914546479388452734597151939639201139875069482092069425428845581584096310252946191103291270482084571518349218243954805054614128487238336435640570639800535674495718801697434275350851437671881640052575116640533426754975393346843369832158197419080856810021130058404572108931589389674329776;
            6'd45: xpb[1] = 1024'd5301750494435568851970886948495438350833539689283080784402548121522077251737150707522509767228847519665496709492767558881126355107416680717398548536044391680348084791907645819404305387451588997424282204864735375396137174490865062014187069465951240010013824498055771413526650317397377489533582809159732068817;
            6'd46: xpb[1] = 1024'd96401810673781169630022786755325920993630909352362206495797076238538957771358011479478506652805116402583039535172546467769798201837809741184902607959932585957951203582746708440764354247618686281883411166679038715516582624085986363566597733221785085917015394212809520000349807578664983424076923855555384292189;
            6'd47: xpb[1] = 1024'd63435175169002029009275759157341970891729851889705648079059749290578942953669733341419432323723710976057432953394831942079406207726982467097246542367489739301863647804014553724494163916268577845032342520106102209272667223460210892154029827294389482557197060513446210557066436766003956341501575075325442031230;
            6'd48: xpb[1] = 1024'd30468539664222888388528731559358020789828794427049089662322422342618928135981455203360357994642305549531826371617117416389014213616155193009590476775046892645776092025282399008223973584918469408181273873533165703028751822834435420741461921366993879197378726814082901113783065953342929258926226295095499770271;
            6'd49: xpb[1] = 1024'd121568599843568489166580631366188503432626164090128215373716950459635808655602315975316354880218574432449369197296896325277686060346548253477094536198935086923379210816121461629584022445085566692640402835347469043149197272429556722293872585122827725104380296528836649700606223214610535193469567341491151993643;
            6'd50: xpb[1] = 1024'd88601964338789348545833603768204553330725106627471656956979623511675793837914037837257280551137169005923762615519181799587294066235720979389438470606492240267291655037389306913313832113735458255789334188774532536905281871803781250881304679195432121744561962829473340257322852401949508110894218561261209732684;
            6'd51: xpb[1] = 1024'd55635328834010207925086576170220603228824049164815098540242296563715779020225759699198206222055763579398156033741467273896902072124893705301782405014049393611204099258657152197043641782385349818938265542201596030661366471178005779468736773268036518384743629130110030814039481589288481028318869781031267471725;
            6'd52: xpb[1] = 1024'd22668693329231067304339548572236653126922991702158540123504969615755764202537481561139131892974358152872549451963752748206510078014066431214126339421606546955116543479924997480773451451035241382087196895628659524417451070552230308056168867340640915024925295430746721370756110776627453945743521000801325210766;
            6'd53: xpb[1] = 1024'd113768753508576668082391448379067135769720361365237665834899497732772644722158342333095128778550627035790092277643531657095181924744459491681630398845494741232719662270764060102133500311202338666546325857442962864537896520147351609608579531096474760931926865145500469957579268037895059880286862047196977434138;
            6'd54: xpb[1] = 1024'd80802118003797527461644420781083185667819303902581107418162170784812629904470064195036054449469221609264485695865817131404789930633632217593974333253051894576632106492031905385863309979852230229695257210870026358293981119521576138196011625169079157572108531446137160514295897225234032797711513266967035173179;
            6'd55: xpb[1] = 1024'd47835482499018386840897393183099235565918246439924549001424843836852615086781786056976980120387816182738879114088102605714397936522804943506318267660609047920544550713299750669593119648502121792844188564297089852050065718895800666783443719241683554212290197746773851071012526412573005715136164486737092912220;
            6'd56: xpb[1] = 1024'd14868846994239246220150365585115285464017188977267990584687516888892600269093507918917905791306410756213272532310388080024005942411977669418662202068166201264456994934567595953322929317152013355993119917724153345806150318270025195370875813314287950852471864047410541627729155599911978632560815706507150651261;
            6'd57: xpb[1] = 1024'd105968907173584846998202265391945768106814558640347116296082045005909480788714368690873902676882679639130815357990166988912677789142370729886166261492054395542060113725406658574682978177319110640452248879538456685926595767865146496923286477070121796759473433762164290214552312861179584567104156752902802874633;
            6'd58: xpb[1] = 1024'd73002271668805706377455237793961818004913501177690557879344718057949465971026090552814828347801274212605208776212452463222285795031543455798510195899611548885972557946674503858412787845969002203601180232965520179682680367239371025510718571142726193399655100062800980771268942048518557484528807972672860613674;
            6'd59: xpb[1] = 1024'd40035636164026565756708210195977867903012443715033999462607391109989451153337812414755754018719868786079602194434737937531893800920716181710854130307168702229885002167942349142142597514618893766750111586392583673438764966613595554098150665215330590039836766363437671327985571235857530401953459192442918352715;
            6'd60: xpb[1] = 1024'd7069000659247425135961182597993917801111386252377441045870064162029436335649534276696679689638463359553995612657023411841501806809888907623198064714725855573797446389210194425872407183268785329899042939819647167194849565987820082685582759287934986680018432664074361884702200423196503319378110412212976091756;
            6'd61: xpb[1] = 1024'd98169060838593025914013082404824400443908755915456566757264592279046316855270395048652676575214732242471538438336802320730173653540281968090702124138614049851400565180049257047232456043435882614358171901633950507315295015582941384237993423043768832587020002378828110471525357684464109253921451458608628315128;
            6'd62: xpb[1] = 1024'd65202425333813885293266054806840450342007698452800008340527265331086302037582116910593602246133326815945931856559087795039781659429454694003046058546171203195313009401317102330962265712085774177507103255061014001071379614957165912825425517116373229227201668679464801028241986871803082171346102678378686054169;
            6'd63: xpb[1] = 1024'd32235789829034744672519027208856500240106640990143449923789938383126287219893838772534527917051921389420325274781373269349389665318627419915389992953728356539225453622584947614692075380735665740656034608488077494827464214331390441412857611188977625867383334980101491584958616059142055088770753898148743793210;
        endcase
    end

    always_comb begin
        case(flag[0][16:12])
            5'd0: xpb[2] = 1024'd0;
            5'd1: xpb[2] = 1024'd123335850008380345450570927015686982882904010653222575635184466500143167739514699544490524802628190272337868100461152178238061512049020480382894052377616550816828572413424010236052124240902763025115163570302380834947909663926511742965268274944811471774384904694855240171781773320409661023314094944544396016582;
            5'd2: xpb[2] = 1024'd122605004332635949502342926626559533021109594180709467142237077935309440141720260178965978390598706235232586793464810921897059183256820626210627979738902060699966470257276803134474009290288320328920129532217521823531458477632126712965557980206393494281949905975593422313457018566890689029509500062463197548833;
            5'd3: xpb[2] = 1024'd121874158656891553554114926237432083159315177708196358649289689370475712543925820813441431978569222198127305486468469665556056854464620772038361907100187570583104368101129596032895894339673877632725095494132662812115007291337741682965847685467975516789514907256331604455132263813371717035704905180381999081084;
            5'd4: xpb[2] = 1024'd121143312981147157605886925848304633297520761235683250156342300805641984946131381447916885566539738161022024179472128409215054525672420917866095834461473080466242265944982388931317779389059434936530061456047803800698556105043356652966137390729557539297079908537069786596807509059852745041900310298300800613335;
            5'd5: xpb[2] = 1024'd120412467305402761657658925459177183435726344763170141663394912240808257348336942082392339154510254123916742872475787152874052196880221063693829761822758590349380163788835181829739664438444992240335027417962944789282104918748971622966427095991139561804644909817807968738482754306333773048095715416219602145586;
            5'd6: xpb[2] = 1024'd119681621629658365709430925070049733573931928290657033170447523675974529750542502716867792742480770086811461565479445896533049868088021209521563689184044100232518061632687974728161549487830549544139993379878085777865653732454586592966716801252721584312209911098546150880157999552814801054291120534138403677837;
            5'd7: xpb[2] = 1024'd118950775953913969761202924680922283712137511818143924677500135111140802152748063351343246330451286049706180258483104640192047539295821355349297616545329610115655959476540767626583434537216106847944959341793226766449202546160201562967006506514303606819774912379284333021833244799295829060486525652057205210088;
            5'd8: xpb[2] = 1024'd118219930278169573812974924291794833850343095345630816184552746546307074554953623985818699918421802012600898951486763383851045210503621501177031543906615119998793857320393560525005319586601664151749925303708367755032751359865816532967296211775885629327339913660022515163508490045776857066681930769976006742339;
            5'd9: xpb[2] = 1024'd117489084602425177864746923902667383988548678873117707691605357981473346957159184620294153506392317975495617644490422127510042881711421647004765471267900629881931755164246353423427204635987221455554891265623508743616300173571431502967585917037467651834904914940760697305183735292257885072877335887894808274590;
            5'd10: xpb[2] = 1024'd116758238926680781916518923513539934126754262400604599198657969416639619359364745254769607094362833938390336337494080871169040552919221792832499398629186139765069653008099146321849089685372778759359857227538649732199848987277046472967875622299049674342469916221498879446858980538738913079072741005813609806841;
            5'd11: xpb[2] = 1024'd116027393250936385968290923124412484264959845928091490705710580851805891761570305889245060682333349901285055030497739614828038224127021938660233325990471649648207550851951939220270974734758336063164823189453790720783397800982661442968165327560631696850034917502237061588534225785219941085268146123732411339092;
            5'd12: xpb[2] = 1024'd115296547575191990020062922735285034403165429455578382212763192286972164163775866523720514270303865864179773723501398358487035895334822084487967253351757159531345448695804732118692859784143893366969789151368931709366946614688276412968455032822213719357599918782975243730209471031700969091463551241651212871343;
            5'd13: xpb[2] = 1024'd114565701899447594071834922346157584541371012983065273719815803722138436565981427158195967858274381827074492416505057102146033566542622230315701180713042669414483346539657525017114744833529450670774755113284072697950495428393891382968744738083795741865164920063713425871884716278181997097658956359570014403594;
            5'd14: xpb[2] = 1024'd113834856223703198123606921957030134679576596510552165226868415157304708968186987792671421446244897789969211109508715845805031237750422376143435108074328179297621244383510317915536629882915007974579721075199213686534044242099506352969034443345377764372729921344451608013559961524663025103854361477488815935845;
            5'd15: xpb[2] = 1024'd113104010547958802175378921567902684817782180038039056733921026592470981370392548427146875034215413752863929802512374589464028908958222521971169035435613689180759142227363110813958514932300565278384687037114354675117593055805121322969324148606959786880294922625189790155235206771144053110049766595407617468096;
            5'd16: xpb[2] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            5'd17: xpb[2] = 1024'd111642319196470010278922920789647785094193347093012839748026249462803526174803669696097782210156445678653367188519692076782024251373822813626636890158184708947034937915068696610802285031071679885994618960944636652284690683216351262969903559130123831895424925186666154438585697264106109122440576831245220532598;
            5'd18: xpb[2] = 1024'd110911473520725614330694920400520335232398930620499731255078860897969798577009230330573235798126961641548085881523350820441021922581622959454370817519470218830172835758921489509224170080457237189799584922859777640868239496921966232970193264391705854402989926467404336580260942510587137128635981949164022064849;
            5'd19: xpb[2] = 1024'd110180627844981218382466920011392885370604514147986622762131472333136070979214790965048689386097477604442804574527009564100019593789423105282104744880755728713310733602774282407646055129842794493604550884774918629451788310627581202970482969653287876910554927748142518721936187757068165134831387067082823597100;
            5'd20: xpb[2] = 1024'd109449782169236822434238919622265435508810097675473514269184083768302343381420351599524142974067993567337523267530668307759017264997223251109838672242041238596448631446627075306067940179228351797409516846690059618035337124333196172970772674914869899418119929028880700863611433003549193141026792185001625129351;
            5'd21: xpb[2] = 1024'd108718936493492426486010919233137985647015681202960405776236695203468615783625912233999596562038509530232241960534327051418014936205023396937572599603326748479586529290479868204489825228613909101214482808605200606618885938038811142971062380176451921925684930309618883005286678250030221147222197302920426661602;
            5'd22: xpb[2] = 1024'd107988090817748030537782918844010535785221264730447297283289306638634888185831472868475050150009025493126960653537985795077012607412823542765306526964612258362724427134332661102911710277999466405019448770520341595202434751744426112971352085438033944433249931590357065146961923496511249153417602420839228193853;
            5'd23: xpb[2] = 1024'd107257245142003634589554918454883085923426848257934188790341918073801160588037033502950503737979541456021679346541644538736010278620623688593040454325897768245862324978185454001333595327385023708824414732435482583785983565450041082971641790699615966940814932871095247288637168742992277159613007538758029726104;
            5'd24: xpb[2] = 1024'd106526399466259238641326918065755636061632431785421080297394529508967432990242594137425957325950057418916398039545303282395007949828423834420774381687183278129000222822038246899755480376770581012629380694350623572369532379155656052971931495961197989448379934151833429430312413989473305165808412656676831258355;
            5'd25: xpb[2] = 1024'd105795553790514842693098917676628186199838015312907971804447140944133705392448154771901410913920573381811116732548962026054005621036223980248508309048468788012138120665891039798177365426156138316434346656265764560953081192861271022972221201222780011955944935432571611571987659235954333172003817774595632790606;
            5'd26: xpb[2] = 1024'd105064708114770446744870917287500736338043598840394863311499752379299977794653715406376864501891089344705835425552620769713003292244024126076242236409754297895276018509743832696599250475541695620239312618180905549536630006566885992972510906484362034463509936713309793713662904482435361178199222892514434322857;
            5'd27: xpb[2] = 1024'd104333862439026050796642916898373286476249182367881754818552363814466250196859276040852318089861605307600554118556279513372000963451824271903976163771039807778413916353596625595021135524927252924044278580096046538120178820272500962972800611745944056971074937994047975855338149728916389184394628010433235855108;
            5'd28: xpb[2] = 1024'd103603016763281654848414916509245836614454765895368646325604975249632522599064836675327771677832121270495272811559938257030998634659624417731710091132325317661551814197449418493443020574312810227849244542011187526703727633978115932973090317007526079478639939274786157997013394975397417190590033128352037387359;
            5'd29: xpb[2] = 1024'd102872171087537258900186916120118386752660349422855537832657586684798795001270397309803225265802637233389991504563597000689996305867424563559444018493610827544689712041302211391864905623698367531654210503926328515287276447683730902973380022269108101986204940555524340138688640221878445196785438246270838919610;
            5'd30: xpb[2] = 1024'd102141325411792862951958915730990936890865932950342429339710198119965067403475957944278678853773153196284710197567255744348993977075224709387177945854896337427827609885155004290286790673083924835459176465841469503870825261389345872973669727530690124493769941836262522280363885468359473202980843364189640451861;
            5'd31: xpb[2] = 1024'd101410479736048467003730915341863487029071516477829320846762809555131339805681518578754132441743669159179428890570914488007991648283024855214911873216181847310965507729007797188708675722469482139264142427756610492454374075094960842973959432792272147001334943117000704422039130714840501209176248482108441984112;
        endcase
    end

    always_comb begin
        case(flag[1][5:0])
            6'd0: xpb[3] = 1024'd0;
            6'd1: xpb[3] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            6'd2: xpb[3] = 1024'd100679634060304071055502914952736037167277100005316212353815420990297612207887079213229586029714185122074147583574573231666989319490825001042645800577467357194103405572860590087130560771855039443069108389671751481037922888800575812974249138053854169508899944397738886563714375961321529215371653600027243516363;
            6'd3: xpb[3] = 1024'd88986103248393735883854908726696839378566436445106476466657203952957970643176049364836843437242440528389646671633113130210952058815627334286388638358035515324309771074505276461880721562023956303948563780314007298374703908090415332978884422239166529629939964889549800830518299905017977314498135486728068032379;
            6'd4: xpb[3] = 1024'd77292572436483400712206902500657641589855772884896740579498986915618329078465019516444100844770695934705145759691653028754914798140429667530131476138603673454516136576149962836630882352192873164828019170956263115711484927380254852983519706424478889750979985381360715097322223848714425413624617373428892548395;
            6'd5: xpb[3] = 1024'd65599041624573065540558896274618443801145109324687004692340769878278687513753989668051358252298951341020644847750192927298877537465232000773874313919171831584722502077794649211381043142361790025707474561598518933048265946670094372988154990609791249872020005873171629364126147792410873512751099260129717064411;
            6'd6: xpb[3] = 1024'd53905510812662730368910890048579246012434445764477268805182552840939045949042959819658615659827206747336143935808732825842840276790034334017617151699739989714928867579439335586131203932530706886586929952240774750385046965959933892992790274795103609993060026364982543630930071736107321611877581146830541580427;
            6'd7: xpb[3] = 1024'd42211980000752395197262883822540048223723782204267532918024335803599404384331929971265873067355462153651643023867272724386803016114836667261359989480308147845135233081084021960881364722699623747466385342883030567721827985249773412997425558980415970114100046856793457897733995679803769711004063033531366096443;
            6'd8: xpb[3] = 1024'd30518449188842060025614877596500850435013118644057797030866118766259762819620900122873130474883717559967142111925812622930765755439639000505102827260876305975341598582728708335631525512868540608345840733525286385058609004539612933002060843165728330235140067348604372164537919623500217810130544920232190612459;
            6'd9: xpb[3] = 1024'd18824918376931724853966871370461652646302455083848061143707901728920121254909870274480387882411972966282641199984352521474728494764441333748845665041444464105547964084373394710381686303037457469225296124167542202395390023829452453006696127351040690356180087840415286431341843567196665909257026806933015128475;
            6'd10: xpb[3] = 1024'd7131387565021389682318865144422454857591791523638325256549684691580479690198840426087645289940228372598140288042892420018691234089243666992588502822012622235754329586018081085131847093206374330104751514809798019732171043119291973011331411536353050477220108332226200698145767510893114008383508693633839644491;
            6'd11: xpb[3] = 1024'd119504552437235795909469786323197689813579555089164273497523322719217733462796949487709973912126158088356788783558925753141717814255266334791491465618911821299651369657233984797512247074892496912294404513839293683433312912630028265980945265404894859865080032238154172995056219528518195124628680406960258644838;
            6'd12: xpb[3] = 1024'd107811021625325460737821780097158492024868891528954537610365105681878091898085919639317231319654413494672287871617465651685680553580068668035234303399479979429857735158878671172262407865061413773173859904481549500770093931919867785985580549590207219986120052729965087261860143472214643223755162293661083160854;
            6'd13: xpb[3] = 1024'd96117490813415125566173773871119294236158227968744801723206888644538450333374889790924488727182668900987786959676005550229643292904871001278977141180048137560064100660523357547012568655230330634053315295123805318106874951209707305990215833775519580107160073221776001528664067415911091322881644180361907676870;
            6'd14: xpb[3] = 1024'd84423960001504790394525767645080096447447564408535065836048671607198808768663859942531746134710924307303286047734545448773606032229673334522719978960616295690270466162168043921762729445399247494932770685766061135443655970499546825994851117960831940228200093713586915795467991359607539422008126067062732192886;
            6'd15: xpb[3] = 1024'd72730429189594455222877761419040898658736900848325329948890454569859167203952830094139003542239179713618785135793085347317568771554475667766462816741184453820476831663812730296512890235568164355812226076408316952780436989789386345999486402146144300349240114205397830062271915303303987521134607953763556708902;
            6'd16: xpb[3] = 1024'd61036898377684120051229755193001700870026237288115594061732237532519525639241800245746260949767435119934284223851625245861531510879278001010205654521752611950683197165457416671263051025737081216691681467050572770117218009079225866004121686331456660470280134697208744329075839247000435620261089840464381224918;
            6'd17: xpb[3] = 1024'd49343367565773784879581748966962503081315573727905858174574020495179884074530770397353518357295690526249783311910165144405494250204080334253948492302320770080889562667102103046013211815905998077571136857692828587453999028369065386008756970516769020591320155189019658595879763190696883719387571727165205740934;
            6'd18: xpb[3] = 1024'd37649836753863449707933742740923305292604910167696122287415803457840242509819740548960775764823945932565282399968705042949456989528882667497691330082888928211095928168746789420763372606074914938450592248335084404790780047658904906013392254702081380712360175680830572862683687134393331818514053613866030256950;
            6'd19: xpb[3] = 1024'd25956305941953114536285736514884107503894246607486386400257586420500600945108710700568033172352201338880781488027244941493419728853685000741434167863457086341302293670391475795513533396243831799330047638977340222127561066948744426018027538887393740833400196172641487129487611078089779917640535500566854772966;
            6'd20: xpb[3] = 1024'd14262775130042779364637730288844909715183583047276650513099369383160959380397680852175290579880456745196280576085784840037382468178487333985177005644025244471508659172036162170263694186412748660209503029619596039464342086238583946022662823072706100954440216664452401396291535021786228016767017387267679288982;
            6'd21: xpb[3] = 1024'd2569244318132444192989724062805711926472919487066914625941152345821317815686651003782547987408712151511779664144324738581345207503289667228919843424593402601715024673680848545013854976581665521088958420261851856801123105528423466027298107258018461075480237156263315663095458965482676115893499273968503804998;
            6'd22: xpb[3] = 1024'd114942409190346850420140645241580946882460683052592862866914790373458571588284760065404876609594641867270428159660358071704371787669312335027822806221492601665612064744896752257394254958267788103278611419291347520502264975039159758996911961126560270463340161062191287960005910983107757232138670987294922805345;
            6'd23: xpb[3] = 1024'd103248878378436515248492639015541749093750019492383126979756573336118930023573730217012134017122897273585927247718897970248334526994114668271565644002060759795818430246541438632144415748436704964158066809933603337839045994328999279001547245311872630584380181554002202226809834926804205331265152873995747321361;
            6'd24: xpb[3] = 1024'd91555347566526180076844632789502551305039355932173391092598356298779288458862700368619391424651152679901426335777437868792297266318917001515308481782628917926024795748186125006894576538605621825037522200575859155175827013618838799006182529497184990705420202045813116493613758870500653430391634760696571837377;
            6'd25: xpb[3] = 1024'd79861816754615844905196626563463353516328692371963655205440139261439646894151670520226648832179408086216925423835977767336260005643719334759051319563197076056231161249830811381644737328774538685916977591218114972512608032908678319010817813682497350826460222537624030760417682814197101529518116647397396353393;
            6'd26: xpb[3] = 1024'd68168285942705509733548620337424155727618028811753919318281922224100005329440640671833906239707663492532424511894517665880222744968521668002794157343765234186437526751475497756394898118943455546796432981860370789849389052198517839015453097867809710947500243029434945027221606757893549628644598534098220869409;
            6'd27: xpb[3] = 1024'd56474755130795174561900614111384957938907365251544183431123705186760363764729610823441163647235918898847923599953057564424185484293324001246536995124333392316643892253120184131145058909112372407675888372502626607186170071488357359020088382053122071068540263521245859294025530701589997727771080420799045385425;
            6'd28: xpb[3] = 1024'd44781224318884839390252607885345760150196701691334447543965488149420722200018580975048421054764174305163422688011597462968148223618126334490279832904901550446850257754764870505895219699281289268555343763144882424522951090778196879024723666238434431189580284013056773560829454645286445826897562307499869901441;
            6'd29: xpb[3] = 1024'd33087693506974504218604601659306562361486038131124711656807271112081080635307551126655678462292429711478921776070137361512110962942928667734022670685469708577056623256409556880645380489450206129434799153787138241859732110068036399029358950423746791310620304504867687827633378588982893926024044194200694417457;
            6'd30: xpb[3] = 1024'd21394162695064169046956595433267364572775374570914975769649054074741439070596521278262935869820685117794420864128677260056073702267731000977765508466037866707262988758054243255395541279619122990314254544429394059196513129357875919033994234609059151431660324996678602094437302532679342025150526080901518933473;
            6'd31: xpb[3] = 1024'd9700631883153833875308589207228166784064711010705239882490837037401797505885491429870193277348940524109919952187217158600036441592533334221508346246606024837469354259698929630145702069788039851193709935071649876533294148647715439038629518794371511552700345488489516361241226476375790124277007967602343449489;
            6'd32: xpb[3] = 1024'd122073796755368240102459510386003401740052474576231188123464475065039051278483600491492521899534870239868568447703250491723063021758556002020411309043505223901366394330914833342526102051474162433383362934101145540234436018158451732008243372662913320940560269394417488658151678494000871240522179680928762449836;
            6'd33: xpb[3] = 1024'd110380265943457904930811504159964203951341811016021452236306258027699409713772570643099779307063125646184067535761790390267025761083358335264154146824073382031572759832559519717276262841643079294262818324743401357571217037448291252012878656848225681061600289886228402924955602437697319339648661567629586965852;
            6'd34: xpb[3] = 1024'd98686735131547569759163497933925006162631147455811716349148040990359768149061540794707036714591381052499566623820330288810988500408160668507896984604641540161779125334204206092026423631811996155142273715385657174907998056738130772017513941033538041182640310378039317191759526381393767438775143454330411481868;
            6'd35: xpb[3] = 1024'd86993204319637234587515491707885808373920483895601980461989823953020126584350510946314294122119636458815065711878870187354951239732963001751639822385209698291985490835848892466776584421980913016021729106027912992244779076027970292022149225218850401303680330869850231458563450325090215537901625341031235997884;
            6'd36: xpb[3] = 1024'd75299673507726899415867485481846610585209820335392244574831606915680485019639481097921551529647891865130564799937410085898913979057765334995382660165777856422191856337493578841526745212149829876901184496670168809581560095317809812026784509404162761424720351361661145725367374268786663637028107227732060513900;
            6'd37: xpb[3] = 1024'd63606142695816564244219479255807412796499156775182508687673389878340843454928451249528808937176147271446063887995949984442876718382567668239125497946346014552398221839138265216276906002318746737780639887312424626918341114607649332031419793589475121545760371853472059992171298212483111736154589114432885029916;
            6'd38: xpb[3] = 1024'd51912611883906229072571473029768215007788493214972772800515172841001201890217421401136066344704402677761562976054489882986839457707370001482868335726914172682604587340782951591027066792487663598660095277954680444255122133897488852036055077774787481666800392345282974258975222156179559835281071001133709545932;
            6'd39: xpb[3] = 1024'd40219081071995893900923466803729017219077829654763036913356955803661560325506391552743323752232658084077062064113029781530802197032172334726611173507482330812810952842427637965777227582656580459539550668596936261591903153187328372040690361960099841787840412837093888525779146099876007934407552887834534061948;
            6'd40: xpb[3] = 1024'd28525550260085558729275460577689819430367166094553301026198738766321918760795361704350581159760913490392561152171569680074764936356974667970354011288050488943017318344072324340527388372825497320419006059239192078928684172477167892045325646145412201908880433328904802792583070043572456033534034774535358577964;
            6'd41: xpb[3] = 1024'd16832019448175223557627454351650621641656502534343565139040521728982277196084331855957838567289168896708060240230109578618727675681777001214096849068618647073223683845717010715277549162994414181298461449881447896265465191767007412049960930330724562029920453820715717059386993987268904132660516661236183093980;
            6'd42: xpb[3] = 1024'd5138488636264888385979448125611423852945838974133829251882304691642635631373302007565095974817424303023559328288649477162690415006579334457839686849186805203430049347361697090027709953163331042177916840523703713602246211056846932054596214516036922150960474312526631326190917930965352231786998547937007609996;
            6'd43: xpb[3] = 1024'd117511653508479294613130369304386658808933602539659777492855942719279889403971411069187424597003354018782207823804682810285716995172602002256742649646086004267327089418577600802408109934849453624367569839553199377303388080567583225024210068384578731538820398218454603623101369948590433348032170261263426610343;
            6'd44: xpb[3] = 1024'd105818122696568959441482363078347461020222938979450041605697725681940247839260381220794682004531609425097706911863222708829679734497404335500485487426654162397533454920222287177158270725018370485247025230195455194640169099857422745028845352569891091659860418710265517889905293892286881447158652147964251126359;
            6'd45: xpb[3] = 1024'd94124591884658624269834356852308263231512275419240305718539508644600606274549351372401939412059864831413205999921762607373642473822206668744228325207222320527739820421866973551908431515187287346126480620837711011976950119147262265033480636755203451780900439202076432156709217835983329546285134034665075642375;
            6'd46: xpb[3] = 1024'd82431061072748289098186350626269065442801611859030569831381291607260964709838321524009196819588120237728705087980302505917605213147009001987971162987790478657946185923511659926658592305356204207005936011479966829313731138437101785038115920940515811901940459693887346423513141779679777645411615921365900158391;
            6'd47: xpb[3] = 1024'd70737530260837953926538344400229867654090948298820833944223074569921323145127291675616454227116375644044204176038842404461567952471811335231714000768358636788152551425156346301408753095525121067885391402122222646650512157726941305042751205125828172022980480185698260690317065723376225744538097808066724674407;
            6'd48: xpb[3] = 1024'd59043999448927618754890338174190669865380284738611098057064857532581681580416261827223711634644631050359703264097382303005530691796613668475456838548926794918358916926801032676158913885694037928764846792764478463987293177016780825047386489311140532144020500677509174957120989667072673843664579694767549190423;
            6'd49: xpb[3] = 1024'd47350468637017283583242331948151472076669621178401362169906640495242040015705231978830969042172886456675202352155922201549493431121416001719199676329494953048565282428445719050909074675862954789644302183406734281324074196306620345052021773496452892265060521169320089223924913610769121942791061581468373706439;
            6'd50: xpb[3] = 1024'd35656937825106948411594325722112274287958957618191626282748423457902398450994202130438226449701141862990701440214462100093456170446218334962942514110063111178771647930090405425659235466031871650523757574048990098660855215596459865056657057681765252386100541661131003490728837554465570041917543468169198222455;
            6'd51: xpb[3] = 1024'd23963407013196613239946319496073076499248294057981890395590206420562756886283172282045483857229397269306200528273001998637418909771020668206685351890631269308978013431735091800409396256200788511403212964691245915997636234886299385061292341867077612507140562152941917757532761498162018141044025354870022738471;
            6'd52: xpb[3] = 1024'd12269876201286278068298313270033878710537630497772154508431989383223115321572142433652741264757652675621699616331541897181381649095823001450428189671199427439184378933379778175159557046369705372282668355333501733334417254176138905065927626052389972628180582644752832024336685441858466240170507241570847254487;
            6'd53: xpb[3] = 1024'd576345389375942896650307043994680921826966937562418621273772345883473756861112585259998672285908081937198704390081795725344388420625334694171027451767585569390744435024464549909717836538622233162123745975757550671198273465978425070562910237702332749220603136563746291140609385554914339296989128271671770503;
            6'd54: xpb[3] = 1024'd112949510261590349123801228222769915877814730503088366862247410373520727529459221646882327294471837797695847199906115128848370968586648002493073990248666784633287784506240368262290117818224744815351776745005253214372340142976714718040176764106244142137080527042491718588051061403179995455542160841598090770850;
            6'd55: xpb[3] = 1024'd101255979449680013952153221996730718089104066942878630975089193336181085964748191798489584702000093204011346287964655027392333707911450335736816828029234942763494150007885054637040278608393661676231232135647509031709121162266554238044812048291556502258120547534302632854854985346876443554668642728298915286866;
            6'd56: xpb[3] = 1024'd89562448637769678780505215770691520300393403382668895087930976298841444400037161950096842109528348610326845376023194925936296447236252668980559665809803100893700515509529741011790439398562578537110687526289764849045902181556393758049447332476868862379160568026113547121658909290572891653795124614999739802882;
            6'd57: xpb[3] = 1024'd77868917825859343608857209544652322511682739822459159200772759261501802835326132101704099517056604016642344464081734824480259186561055002224302503590371259023906881011174427386540600188731495397990142916932020666382683200846233278054082616662181222500200588517924461388462833234269339752921606501700564318898;
            6'd58: xpb[3] = 1024'd66175387013949008437209203318613124722972076262249423313614542224162161270615102253311356924584859422957843552140274723024221925885857335468045341370939417154113246512819113761290760978900412258869598307574276483719464220136072798058717900847493582621240609009735375655266757177965787852048088388401388834914;
            6'd59: xpb[3] = 1024'd54481856202038673265561197092573926934261412702039687426456325186822519705904072404918614332113114829273342640198814621568184665210659668711788179151507575284319612014463800136040921769069329119749053698216532301056245239425912318063353185032805942742280629501546289922070681121662235951174570275102213350930;
            6'd60: xpb[3] = 1024'd42788325390128338093913190866534729145550749141829951539298108149482878141193042556525871739641370235588841728257354520112147404535462001955531016932075733414525977516108486510791082559238245980628509088858788118393026258715751838067988469218118302863320649993357204188874605065358684050301052161803037866946;
            6'd61: xpb[3] = 1024'd31094794578218002922265184640495531356840085581620215652139891112143236576482012708133129147169625641904340816315894418656110143860264335199273854712643891544732343017753172885541243349407162841507964479501043935729807278005591358072623753403430662984360670485168118455678529009055132149427534048503862382962;
            6'd62: xpb[3] = 1024'd19401263766307667750617178414456333568129422021410479764981674074803595011770982859740386554697881048219839904374434317200072883185066668443016692493212049674938708519397859260291404139576079702387419870143299753066588297295430878077259037588743023105400690976979032722482452952751580248554015935204686898978;
            6'd63: xpb[3] = 1024'd7707732954397332578969172188417135779418758461200743877823457037463953447059953011347643962226136454535338992432974215744035622509869001686759530273780207805145074021042545635041564929744996563266875260785555570403369316585270398081894321774055383226440711468789946989286376896448028347680497821905511414994;
        endcase
    end

    always_comb begin
        case(flag[1][11:6])
            6'd0: xpb[4] = 1024'd0;
            6'd1: xpb[4] = 1024'd120080897826611738806120093367192370735406522026726692118797095065101207219658062072969972584412066170293987487949007548867062202675891669485662493070679406869042114092258449347421964911431119145456528259815051234104511186096006691051508175642597192614300635374717919286196828914073109463925669535231930415341;
            6'd2: xpb[4] = 1024'd116095099969098736213441259329570308726114616927717700109462335065225519102006985235924873954166458031144825568440521663155060564510563004416164861125027772804393553614945681357213690631345032569602858911242862621844661521971116609138037781601964935961781367335318780542287129754217585910732649243838266346351;
            6'd3: xpb[4] = 1024'd112109302111585733620762425291948246716822711828708708100127575065349830984355908398879775323920849891995663648932035777443058926345234339346667229179376138739744993137632913367005416351258945993749189562670674009584811857846226527224567387561332679309262099295919641798377430594362062357539628952444602277361;
            6'd4: xpb[4] = 1024'd108123504254072731028083591254326184707530806729699716090792815065474142866704831561834676693675241752846501729423549891731057288179905674277169597233724504675096432660320145376797142071172859417895520214098485397324962193721336445311096993520700422656742831256520503054467731434506538804346608661050938208371;
            6'd5: xpb[4] = 1024'd104137706396559728435404757216704122698238901630690724081458055065598454749053754724789578063429633613697339809915064006019055650014577009207671965288072870610447872183007377386588867791086772842041850865526296785065112529596446363397626599480068166004223563217121364310558032274651015251153588369657274139381;
            6'd6: xpb[4] = 1024'd100151908539046725842725923179082060688946996531681732072123295065722766631402677887744479433184025474548177890406578120307054011849248344138174333342421236545799311705694609396380593511000686266188181516954108172805262865471556281484156205439435909351704295177722225566648333114795491697960568078263610070391;
            6'd7: xpb[4] = 1024'd96166110681533723250047089141459998679655091432672740062788535065847078513751601050699380802938417335399015970898092234595052373683919679068676701396769602481150751228381841406172319230914599690334512168381919560545413201346666199570685811398803652699185027138323086822738633954939968144767547786869946001401;
            6'd8: xpb[4] = 1024'd92180312824020720657368255103837936670363186333663748053453775065971390396100524213654282172692809196249854051389606348883050735518591013999179069451117968416502190751069073415964044950828513114480842819809730948285563537221776117657215417358171396046665759098923948078828934795084444591574527495476281932411;
            6'd9: xpb[4] = 1024'd88194514966507718064689421066215874661071281234654756044119015066095702278449447376609183542447201057100692131881120463171049097353262348929681437505466334351853630273756305425755770670742426538627173471237542336025713873096886035743745023317539139394146491059524809334919235635228921038381507204082617863421;
            6'd10: xpb[4] = 1024'd84208717108994715472010587028593812651779376135645764034784255066220014160798370539564084912201592917951530212372634577459047459187933683860183805559814700287205069796443537435547496390656339962773504122665353723765864208971995953830274629276906882741627223020125670591009536475373397485188486912688953794431;
            6'd11: xpb[4] = 1024'd80222919251481712879331752990971750642487471036636772025449495066344326043147293702518986281955984778802368292864148691747045821022605018790686173614163066222556509319130769445339222110570253386919834774093165111506014544847105871916804235236274626089107954980726531847099837315517873931995466621295289725441;
            6'd12: xpb[4] = 1024'd76237121393968710286652918953349688633195565937627780016114735066468637925496216865473887651710376639653206373355662806035044182857276353721188541668511432157907948841818001455130947830484166811066165425520976499246164880722215790003333841195642369436588686941327393103190138155662350378802446329901625656451;
            6'd13: xpb[4] = 1024'd72251323536455707693974084915727626623903660838618788006779975066592949807845140028428789021464768500504044453847176920323042544691947688651690909722859798093259388364505233464922673550398080235212496076948787886986315216597325708089863447155010112784069418901928254359280438995806826825609426038507961587461;
            6'd14: xpb[4] = 1024'd68265525678942705101295250878105564614611755739609795997445215066717261690194063191383690391219160361354882534338691034611040906526619023582193277777208164028610827887192465474714399270311993659358826728376599274726465552472435626176393053114377856131550150862529115615370739835951303272416405747114297518471;
            6'd15: xpb[4] = 1024'd64279727821429702508616416840483502605319850640600803988110455066841573572542986354338591760973552222205720614830205148899039268361290358512695645831556529963962267409879697484506124990225907083505157379804410662466615888347545544262922659073745599479030882823129976871461040676095779719223385455720633449481;
            6'd16: xpb[4] = 1024'd60293929963916699915937582802861440596027945541591811978775695066965885454891909517293493130727944083056558695321719263187037630195961693443198013885904895899313706932566929494297850710139820507651488031232222050206766224222655462349452265033113342826511614783730838127551341516240256166030365164326969380491;
            6'd17: xpb[4] = 1024'd56308132106403697323258748765239378586736040442582819969440935067090197337240832680248394500482335943907396775813233377475035992030633028373700381940253261834665146455254161504089576430053733931797818682660033437946916560097765380435981870992481086173992346744331699383641642356384732612837344872933305311501;
            6'd18: xpb[4] = 1024'd52322334248890694730579914727617316577444135343573827960106175067214509219589755843203295870236727804758234856304747491763034353865304363304202749994601627770016585977941393513881302149967647355944149334087844825687066895972875298522511476951848829521473078704932560639731943196529209059644324581539641242511;
            6'd19: xpb[4] = 1024'd48336536391377692137901080689995254568152230244564835950771415067338821101938679006158197239991119665609072936796261606051032715699975698234705118048949993705368025500628625523673027869881560780090479985515656213427217231847985216609041082911216572868953810665533421895822244036673685506451304290145977173521;
            6'd20: xpb[4] = 1024'd44350738533864689545222246652373192558860325145555843941436655067463132984287602169113098609745511526459911017287775720339031077534647033165207486103298359640719465023315857533464753589795474204236810636943467601167367567723095134695570688870584316216434542626134283151912544876818161953258283998752313104531;
            6'd21: xpb[4] = 1024'd40364940676351686952543412614751130549568420046546851932101895067587444866636525332067999979499903387310749097779289834627029439369318368095709854157646725576070904546003089543256479309709387628383141288371278988907517903598205052782100294829952059563915274586735144408002845716962638400065263707358649035541;
            6'd22: xpb[4] = 1024'd36379142818838684359864578577129068540276514947537859922767135067711756748985448495022901349254295248161587178270803948915027801203989703026212222211995091511422344068690321553048205029623301052529471939799090376647668239473314970868629900789319802911396006547336005664093146557107114846872243415964984966551;
            6'd23: xpb[4] = 1024'd32393344961325681767185744539507006530984609848528867913432375067836068631334371657977802719008687109012425258762318063203026163038661037956714590266343457446773783591377553562839930749537214476675802591226901764387818575348424888955159506748687546258876738507936866920183447397251591293679223124571320897561;
            6'd24: xpb[4] = 1024'd28407547103812679174506910501884944521692704749519875904097615067960380513683294820932704088763078969863263339253832177491024524873332372887216958320691823382125223114064785572631656469451127900822133242654713152127968911223534807041689112708055289606357470468537728176273748237396067740486202833177656828571;
            6'd25: xpb[4] = 1024'd24421749246299676581828076464262882512400799650510883894762855068084692396032217983887605458517470830714101419745346291779022886708003707817719326375040189317476662636752017582423382189365041324968463894082524539868119247098644725128218718667423032953838202429138589432364049077540544187293182541783992759581;
            6'd26: xpb[4] = 1024'd20435951388786673989149242426640820503108894551501891885428095068209004278381141146842506828271862691564939500236860406067021248542675042748221694429388555252828102159439249592215107909278954749114794545510335927608269582973754643214748324626790776301318934389739450688454349917685020634100162250390328690591;
            6'd27: xpb[4] = 1024'd16450153531273671396470408389018758493816989452492899876093335068333316160730064309797408198026254552415777580728374520355019610377346377678724062483736921188179541682126481602006833629192868173261125196938147315348419918848864561301277930586158519648799666350340311944544650757829497080907141958996664621601;
            6'd28: xpb[4] = 1024'd12464355673760668803791574351396696484525084353483907866758575068457628043078987472752309567780646413266615661219888634643017972212017712609226430538085287123530981204813713611798559349106781597407455848365958703088570254723974479387807536545526262996280398310941173200634951597973973527714121667603000552611;
            6'd29: xpb[4] = 1024'd8478557816247666211112740313774634475233179254474915857423815068581939925427910635707210937535038274117453741711402748931016334046689047539728798592433653058882420727500945621590285069020695021553786499793770090828720590599084397474337142504894006343761130271542034456725252438118449974521101376209336483621;
            6'd30: xpb[4] = 1024'd4492759958734663618433906276152572465941274155465923848089055068706251807776833798662112307289430134968291822202916863219014695881360382470231166646782018994233860250188177631382010788934608445700117151221581478568870926474194315560866748464261749691241862232142895712815553278262926421328081084815672414631;
            6'd31: xpb[4] = 1024'd506962101221661025755072238530510456649369056456931838754295068830563690125756961617013677043821995819129902694430977507013057716031717400733534701130384929585299772875409641173736508848521869846447802649392866309021262349304233647396354423629493038722594192743756968905854118407402868135060793422008345641;
            6'd32: xpb[4] = 1024'd120587859927833399831875165605722881192055891083183623957551390133931770909783819034586986261455888166113117390643438526374075260391923386886396027771809791798627413865133858988595701420279641015302976062464444100413532448445310924698904530066226685653023229567461676255102683032480512332060730328653938760982;
            6'd33: xpb[4] = 1024'd116602062070320397239196331568100819182763985984174631948216630134056082792132742197541887631210280026963955471134952640662073622226594721816898395826158157733978853387821090998387427140193554439449306713892255488153682784320420842785434136025594429000503961528062537511192983872624988778867710037260274691992;
            6'd34: xpb[4] = 1024'd112616264212807394646517497530478757173472080885165639938881870134180394674481665360496789000964671887814793551626466754950071984061266056747400763880506523669330292910508323008179152860107467863595637365320066875893833120195530760871963741984962172347984693488663398767283284712769465225674689745866610623002;
            6'd35: xpb[4] = 1024'd108630466355294392053838663492856695164180175786156647929547110134304706556830588523451690370719063748665631632117980869238070345895937391677903131934854889604681732433195555017970878580021381287741968016747878263633983456070640678958493347944329915695465425449264260023373585552913941672481669454472946554012;
            6'd36: xpb[4] = 1024'd104644668497781389461159829455234633154888270687147655920212350134429018439179511686406591740473455609516469712609494983526068707730608726608405499989203255540033171955882787027762604299935294711888298668175689651374133791945750597045022953903697659042946157409865121279463886393058418119288649163079282485022;
            6'd37: xpb[4] = 1024'd100658870640268386868480995417612571145596365588138663910877590134553330321528434849361493110227847470367307793101009097814067069565280061538907868043551621475384611478570019037554330019849208136034629319603501039114284127820860515131552559863065402390426889370465982535554187233202894566095628871685618416032;
            6'd38: xpb[4] = 1024'd96673072782755384275802161379990509136304460489129671901542830134677642203877358012316394479982239331218145873592523212102065431399951396469410236097899987410736051001257251047346055739763121560180959971031312426854434463695970433218082165822433145737907621331066843791644488073347371012902608580291954347042;
            6'd39: xpb[4] = 1024'd92687274925242381683123327342368447127012555390120679892208070134801954086226281175271295849736631192068983954084037326390063793234622731399912604152248353346087490523944483057137781459677034984327290622459123814594584799571080351304611771781800889085388353291667705047734788913491847459709588288898290278052;
            6'd40: xpb[4] = 1024'd88701477067729379090444493304746385117720650291111687882873310134926265968575204338226197219491023052919822034575551440678062155069294066330414972206596719281438930046631715066929507179590948408473621273886935202334735135446190269391141377741168632432869085252268566303825089753636323906516567997504626209062;
            6'd41: xpb[4] = 1024'd84715679210216376497765659267124323108428745192102695873538550135050577850924127501181098589245414913770660115067065554966060516903965401260917340260945085216790369569318947076721232899504861832619951925314746590074885471321300187477670983700536375780349817212869427559915390593780800353323547706110962140072;
            6'd42: xpb[4] = 1024'd80729881352703373905086825229502261099136840093093703864203790135174889733273050664135999958999806774621498195558579669254058878738636736191419708315293451152141809092006179086512958619418775256766282576742557977815035807196410105564200589659904119127830549173470288816005691433925276800130527414717298071082;
            6'd43: xpb[4] = 1024'd76744083495190371312407991191880199089844934994084711854869030135299201615621973827090901328754198635472336276050093783542057240573308071121922076369641817087493248614693411096304684339332688680912613228170369365555186143071520023650730195619271862475311281134071150072095992274069753246937507123323634002092;
            6'd44: xpb[4] = 1024'd72758285637677368719729157154258137080553029895075719845534270135423513497970896990045802698508590496323174356541607897830055602407979406052424444423990183022844688137380643106096410059246602105058943879598180753295336478946629941737259801578639605822792013094672011328186293114214229693744486831929969933102;
            6'd45: xpb[4] = 1024'd68772487780164366127050323116636075071261124796066727836199510135547825380319820153000704068262982357174012437033122012118053964242650740982926812478338548958196127660067875115888135779160515529205274531025992141035486814821739859823789407538007349170272745055272872584276593954358706140551466540536305864112;
            6'd46: xpb[4] = 1024'd64786689922651363534371489079014013061969219697057735826864750135672137262668743315955605438017374218024850517524636126406052326077322075913429180532686914893547567182755107125679861499074428953351605182453803528775637150696849777910319013497375092517753477015873733840366894794503182587358446249142641795122;
            6'd47: xpb[4] = 1024'd60800892065138360941692655041391951052677314598048743817529990135796449145017666478910506807771766078875688598016150240694050687911993410843931548587035280828899006705442339135471587218988342377497935833881614916515787486571959695996848619456742835865234208976474595096457195634647659034165425957748977726132;
            6'd48: xpb[4] = 1024'd56815094207625358349013821003769889043385409499039751808195230135920761027366589641865408177526157939726526678507664354982049049746664745774433916641383646764250446228129571145263312938902255801644266485309426304255937822447069614083378225416110579212714940937075456352547496474792135480972405666355313657142;
            6'd49: xpb[4] = 1024'd52829296350112355756334986966147827034093504400030759798860470136045072909715512804820309547280549800577364758999178469270047411581336080704936284695732012699601885750816803155055038658816169225790597136737237691996088158322179532169907831375478322560195672897676317608637797314936611927779385374961649588152;
            6'd50: xpb[4] = 1024'd48843498492599353163656152928525765024801599301021767789525710136169384792064435967775210917034941661428202839490692583558045773416007415635438652750080378634953325273504035164846764378730082649936927788165049079736238494197289450256437437334846065907676404858277178864728098155081088374586365083567985519162;
            6'd51: xpb[4] = 1024'd44857700635086350570977318890903703015509694202012775780190950136293696674413359130730112286789333522279040919982206697846044135250678750565941020804428744570304764796191267174638490098643996074083258439592860467476388830072399368342967043294213809255157136818878040120818398995225564821393344792174321450172;
            6'd52: xpb[4] = 1024'd40871902777573347978298484853281641006217789103003783770856190136418008556762282293685013656543725383129879000473720812134042497085350085496443388858777110505656204318878499184430215818557909498229589091020671855216539165947509286429496649253581552602637868779478901376908699835370041268200324500780657381182;
            6'd53: xpb[4] = 1024'd36886104920060345385619650815659578996925884003994791761521430136542320439111205456639915026298117243980717080965234926422040858920021420426945756913125476441007643841565731194221941538471822922375919742448483242956689501822619204516026255212949295950118600740079762632999000675514517715007304209386993312192;
            6'd54: xpb[4] = 1024'd32900307062547342792940816778037516987633978904985799752186670136666632321460128619594816396052509104831555161456749040710039220754692755357448124967473842376359083364252963204013667258385736346522250393876294630696839837697729122602555861172317039297599332700680623889089301515658994161814283917993329243202;
            6'd55: xpb[4] = 1024'd28914509205034340200261982740415454978342073805976807742851910136790944203809051782549717765806900965682393241948263154998037582589364090287950493021822208311710522886940195213805392978299649770668581045304106018436990173572839040689085467131684782645080064661281485145179602355803470608621263626599665174212;
            6'd56: xpb[4] = 1024'd24928711347521337607583148702793392969050168706967815733517150136915256086157974945504619135561292826533231322439777269286035944424035425218452861076170574247061962409627427223597118698213563194814911696731917406177140509447948958775615073091052525992560796621882346401269903195947947055428243335206001105222;
            6'd57: xpb[4] = 1024'd20942913490008335014904314665171330959758263607958823724182390137039567968506898108459520505315684687384069402931291383574034306258706760148955229130518940182413401932314659233388844418127476618961242348159728793917290845323058876862144679050420269340041528582483207657360204036092423502235223043812337036232;
            6'd58: xpb[4] = 1024'd16957115632495332422225480627549268950466358508949831714847630137163879850855821271414421875070076548234907483422805497862032668093378095079457597184867306117764841455001891243180570138041390043107572999587540181657441181198168794948674285009788012687522260543084068913450504876236899949042202752418672967242;
            6'd59: xpb[4] = 1024'd12971317774982329829546646589927206941174453409940839705512870137288191733204744434369323244824468409085745563914319612150031029928049430009959965239215672053116280977689123252972295857955303467253903651015351569397591517073278713035203890969155756035002992503684930169540805716381376395849182461025008898252;
            6'd60: xpb[4] = 1024'd8985519917469327236867812552305144931882548310931847696178110137412503615553667597324224614578860269936583644405833726438029391762720764940462333293564037988467720500376355262764021577869216891400234302443162957137741852948388631121733496928523499382483724464285791425631106556525852842656162169631344829262;
            6'd61: xpb[4] = 1024'd4999722059956324644188978514683082922590643211922855686843350137536815497902590760279125984333252130787421724897347840726027753597392099870964701347912403923819160023063587272555747297783130315546564953870974344877892188823498549208263102887891242729964456424886652681721407396670329289463141878237680760272;
            6'd62: xpb[4] = 1024'd1013924202443322051510144477061020913298738112913863677508590137661127380251513923234027354087643991638259805388861955014026115432063434801467069402260769859170599545750819282347473017697043739692895605298785732618042524698608467294792708847258986077445188385487513937811708236814805736270121586844016691282;
            6'd63: xpb[4] = 1024'd121094822029055060857630237844253391648705260139640555796305685202762334599909575996203999938499710161932247293337869503881088318107955104287129562472940176728212713638009268629769437929128162885149423865113836966722553710794615158346300884489856178691745823760205433224008537150887915200195791122075947106623;
        endcase
    end

    always_comb begin
        case(flag[1][16:12])
            5'd0: xpb[5] = 1024'd0;
            5'd1: xpb[5] = 1024'd117109024171542058264951403806631329639413355040631563786970925202886646482258499159158901308254102022783085373829383618169086679942626439217631930527288542663564153160696500639561163649042076309295754516541648354462704046669725076432830490449223922039226555720806294480098837991032391647002770830682283037633;
            5'd2: xpb[5] = 1024'd110151352658959375131103880208448226534128282955527443445809995340796397627207859408302731401850529736123021340201273801759109519044032543880103736038246044393437631751821783941492088106566946897281311424696056862561047243118553379900682411215218394811633208027495530930091147908136150276886851834738971590935;
            5'd3: xpb[5] = 1024'd103193681146376691997256356610265123428843210870423323104649065478706148772157219657446561495446957449462957306573163985349132358145438648542575541549203546123311110342947067243423012564091817485266868332850465370659390439567381683368534331981212867584039860334184767380083457825239908906770932838795660144237;
            5'd4: xpb[5] = 1024'd96236009633794008863408833012082020323558138785319202763488135616615899917106579906590391589043385162802893272945054168939155197246844753205047347060161047853184588934072350545353937021616688073252425241004873878757733636016209986836386252747207340356446512640874003830075767742343667536655013842852348697539;
            5'd5: xpb[5] = 1024'd89278338121211325729561309413898917218273066700215082422327205754525651062055940155734221682639812876142829239316944352529178036348250857867519152571118549583058067525197633847284861479141558661237982149159282386856076832465038290304238173513201813128853164947563240280068077659447426166539094846909037250841;
            5'd6: xpb[5] = 1024'd82320666608628642595713785815715814112987994615110962081166275892435402207005300404878051776236240589482765205688834536119200875449656962529990958082076051312931546116322917149215785936666429249223539057313690894954420028913866593772090094279196285901259817254252476730060387576551184796423175850965725804143;
            5'd7: xpb[5] = 1024'd75362995096045959461866262217532711007702922530006841740005346030345153351954660654021881869832668302822701172060724719709223714551063067192462763593033553042805024707448200451146710394191299837209095965468099403052763225362694897239942015045190758673666469560941713180052697493654943426307256855022414357445;
            5'd8: xpb[5] = 1024'd68405323583463276328018738619349607902417850444902721398844416168254904496904020903165711963429096016162637138432614903299246553652469171854934569103991054772678503298573483753077634851716170425194652873622507911151106421811523200707793935811185231446073121867630949630045007410758702056191337859079102910747;
            5'd9: xpb[5] = 1024'd61447652070880593194171215021166504797132778359798601057683486306164655641853381152309542057025523729502573104804505086889269392753875276517406374614948556502551981889698767055008559309241041013180209781776916419249449618260351504175645856577179704218479774174320186080037317327862460686075418863135791464049;
            5'd10: xpb[5] = 1024'd54489980558297910060323691422983401691847706274694480716522556444074406786802741401453372150621951442842509071176395270479292231855281381179878180125906058232425460480824050356939483766765911601165766689931324927347792814709179807643497777343174176990886426481009422530029627244966219315959499867192480017351;
            5'd11: xpb[5] = 1024'd47532309045715226926476167824800298586562634189590360375361626581984157931752101650597202244218379156182445037548285454069315070956687485842349985636863559962298939071949333658870408224290782189151323598085733435446136011158008111111349698109168649763293078787698658980021937162069977945843580871249168570653;
            5'd12: xpb[5] = 1024'd40574637533132543792628644226617195481277562104486240034200696719893909076701461899741032337814806869522381003920175637659337910058093590504821791147821061692172417663074616960801332681815652777136880506240141943544479207606836414579201618875163122535699731094387895430014247079173736575727661875305857123955;
            5'd13: xpb[5] = 1024'd33616966020549860658781120628434092375992490019382119693039766857803660221650822148884862431411234582862316970292065821249360749159499695167293596658778563422045896254199900262732257139340523365122437414394550451642822404055664718047053539641157595308106383401077131880006556996277495205611742879362545677257;
            5'd14: xpb[5] = 1024'd26659294507967177524933597030250989270707417934277999351878836995713411366600182398028692525007662296202252936663956004839383588260905799829765402169736065151919374845325183564663181596865393953107994322548958959741165600504493021514905460407152068080513035707766368329998866913381253835495823883419234230559;
            5'd15: xpb[5] = 1024'd19701622995384494391086073432067886165422345849173879010717907133623162511549542647172522618604090009542188903035846188429406427362311904492237207680693566881792853436450466866594106054390264541093551230703367467839508796953321324982757381173146540852919688014455604779991176830485012465379904887475922783861;
            5'd16: xpb[5] = 1024'd12743951482801811257238549833884783060137273764069758669556977271532913656498902896316352712200517722882124869407736372019429266463718009154709013191651068611666332027575750168525030511915135129079108138857775975937851993402149628450609301939141013625326340321144841229983486747588771095263985891532611337163;
            5'd17: xpb[5] = 1024'd5786279970219128123391026235701679954852201678965638328396047409442664801448263145460182805796945436222060835779626555609452105565124113817180818702608570341539810618701033470455954969440005717064665047012184484036195189850977931918461222705135486397732992627834077679975796664692529725148066895589299890465;
            5'd18: xpb[5] = 1024'd122895304141761186388342430042333009594265556719597202115366972612329311283706762304619084114051047459005146209609010173778538785507750553034812749229897113005103963779397534110017118618482082026360419563553832838498899236520703008351291713154359408436959548348640372160074634655724921372150837726271582928098;
            5'd19: xpb[5] = 1024'd115937632629178503254494906444149906488980484634493081774206042750239062428656122553762914207647475172345082175980900357368561624609156657697284554740854614734977442370522817411948043076006952614345976471708241346597242432969531311819143633920353881209366200655329608610066944572828680002034918730328271481400;
            5'd20: xpb[5] = 1024'd108979961116595820120647382845966803383695412549388961433045112888148813573605482802906744301243902885685018142352790540958584463710562762359756360251812116464850920961648100713878967533531823202331533379862649854695585629418359615286995554686348353981772852962018845060059254489932438631918999734384960034702;
            5'd21: xpb[5] = 1024'd102022289604013136986799859247783700278410340464284841091884183026058564718554843052050574394840330599024954108724680724548607302811968867022228165762769618194724399552773384015809891991056693790317090288017058362793928825867187918754847475452342826754179505268708081510051564407036197261803080738441648588004;
            5'd22: xpb[5] = 1024'd95064618091430453852952335649600597173125268379180720750723253163968315863504203301194404488436758312364890075096570908138630141913374971684699971273727119924597878143898667317740816448581564378302647196171466870892272022316016222222699396218337299526586157575397317960043874324139955891687161742498337141306;
            5'd23: xpb[5] = 1024'd88106946578847770719104812051417494067840196294076600409562323301878067008453563550338234582033186025704826041468461091728652981014781076347171776784684621654471356735023950619671740906106434966288204104325875378990615218764844525690551316984331772298992809882086554410036184241243714521571242746555025694608;
            5'd24: xpb[5] = 1024'd81149275066265087585257288453234390962555124208972480068401393439787818153402923799482064675629613739044762007840351275318675820116187181009643582295642123384344835326149233921602665363631305554273761012480283887088958415213672829158403237750326245071399462188775790860028494158347473151455323750611714247910;
            5'd25: xpb[5] = 1024'd74191603553682404451409764855051287857270052123868359727240463577697569298352284048625894769226041452384697974212241458908698659217593285672115387806599625114218313917274517223533589821156176142259317920634692395187301611662501132626255158516320717843806114495465027310020804075451231781339404754668402801212;
            5'd26: xpb[5] = 1024'd67233932041099721317562241256868184751984980038764239386079533715607320443301644297769724862822469165724633940584131642498721498318999390334587193317557126844091792508399800525464514278681046730244874828789100903285644808111329436094107079282315190616212766802154263760013113992554990411223485758725091354514;
            5'd27: xpb[5] = 1024'd60276260528517038183714717658685081646699907953660119044918603853517071588251004546913554956418896879064569906956021826088744337420405494997058998828514628573965271099525083827395438736205917318230431736943509411383988004560157739561959000048309663388619419108843500210005423909658749041107566762781779907816;
            5'd28: xpb[5] = 1024'd53318589015934355049867194060501978541414835868555998703757673991426822733200364796057385050015324592404505873327912009678767176521811599659530804339472130303838749690650367129326363193730787906215988645097917919482331201008986043029810920814304136161026071415532736659997733826762507670991647766838468461118;
            5'd29: xpb[5] = 1024'd46360917503351671916019670462318875436129763783451878362596744129336573878149725045201215143611752305744441839699802193268790015623217704322002609850429632033712228281775650431257287651255658494201545553252326427580674397457814346497662841580298608933432723722221973109990043743866266300875728770895157014420;
            5'd30: xpb[5] = 1024'd39403245990768988782172146864135772330844691698347758021435814267246325023099085294345045237208180019084377806071692376858812854724623808984474415361387133763585706872900933733188212108780529082187102461406734935679017593906642649965514762346293081705839376028911209559982353660970024930759809774951845567722;
            5'd31: xpb[5] = 1024'd32445574478186305648324623265952669225559619613243637680274884405156076168048445543488875330804607732424313772443582560448835693826029913646946220872344635493459185464026217035119136566305399670172659369561143443777360790355470953433366683112287554478246028335600446009974663578073783560643890779008534121024;
        endcase
    end

    always_comb begin
        case(flag[2][5:0])
            6'd0: xpb[6] = 1024'd0;
            6'd1: xpb[6] = 1024'd12743951482801811257238549833884783060137273764069758669556977271532913656498902896316352712200517722882124869407736372019429266463718009154709013191651068611666332027575750168525030511915135129079108138857775975937851993402149628450609301939141013625326340321144841229983486747588771095263985891532611337163;
            6'd2: xpb[6] = 1024'd25487902965603622514477099667769566120274547528139517339113954543065827312997805792632705424401035445764249738815472744038858532927436018309418026383302137223332664055151500337050061023830270258158216277715551951875703986804299256901218603878282027250652680642289682459966973495177542190527971783065222674326;
            6'd3: xpb[6] = 1024'd38231854448405433771715649501654349180411821292209276008670931814598740969496708688949058136601553168646374608223209116058287799391154027464127039574953205834998996082727250505575091535745405387237324416573327927813555980206448885351827905817423040875979020963434523689950460242766313285791957674597834011489;
            6'd4: xpb[6] = 1024'd50975805931207245028954199335539132240549095056279034678227909086131654625995611585265410848802070891528499477630945488077717065854872036618836052766604274446665328110303000674100122047660540516316432555431103903751407973608598513802437207756564054501305361284579364919933946990355084381055943566130445348652;
            6'd5: xpb[6] = 1024'd63719757414009056286192749169423915300686368820348793347784886357664568282494514481581763561002588614410624347038681860097146332318590045773545065958255343058331660137878750842625152559575675645395540694288879879689259967010748142253046509695705068126631701605724206149917433737943855476319929457663056685815;
            6'd6: xpb[6] = 1024'd76463708896810867543431299003308698360823642584418552017341863629197481938993417377898116273203106337292749216446418232116575598782308054928254079149906411669997992165454501011150183071490810774474648833146655855627111960412897770703655811634846081751958041926869047379900920485532626571583915349195668022978;
            6'd7: xpb[6] = 1024'd89207660379612678800669848837193481420960916348488310686898840900730395595492320274214468985403624060174874085854154604136004865246026064082963092341557480281664324193030251179675213583405945903553756972004431831564963953815047399154265113573987095377284382248013888609884407233121397666847901240728279360141;
            6'd8: xpb[6] = 1024'd101951611862414490057908398671078264481098190112558069356455818172263309251991223170530821697604141783056998955261890976155434131709744073237672105533208548893330656220606001348200244095321081032632865110862207807502815947217197027604874415513128109002610722569158729839867893980710168762111887132260890697304;
            6'd9: xpb[6] = 1024'd114695563345216301315146948504963047541235463876627828026012795443796222908490126066847174409804659505939123824669627348174863398173462082392381118724859617504996988248181751516725274607236216161711973249719983783440667940619346656055483717452269122627937062890303571069851380728298939857375873023793502034467;
            6'd10: xpb[6] = 1024'd3372819143893371173586570934033397856674310514961902567437917650352241227679890053148455907347502919378099286619870285615228823795959756991930006900179645182972645706186284347620065927634145569480883780190519913014159083800599511541114449708180686986443499797331354269728339401959077935521169088700518887299;
            6'd11: xpb[6] = 1024'd16116770626695182430825120767918180916811584279031661236994894921885154884178792949464808619548020642260224156027606657634658090259677766146639020091830713794638977733762034516145096439549280698559991919048295888952011077202749139991723751647321700611769840118476195499711826149547849030785154980233130224462;
            6'd12: xpb[6] = 1024'd28860722109496993688063670601802963976948858043101419906551872193418068540677695845781161331748538365142349025435343029654087356723395775301348033283481782406305309761337784684670126951464415827639100057906071864889863070604898768442333053586462714237096180439621036729695312897136620126049140871765741561625;
            6'd13: xpb[6] = 1024'd41604673592298804945302220435687747037086131807171178576108849464950982197176598742097514043949056088024473894843079401673516623187113784456057046475132851017971641788913534853195157463379550956718208196763847840827715064007048396892942355525603727862422520760765877959678799644725391221313126763298352898788;
            6'd14: xpb[6] = 1024'd54348625075100616202540770269572530097223405571240937245665826736483895853675501638413866756149573810906598764250815773692945889650831793610766059666783919629637973816489285021720187975294686085797316335621623816765567057409198025343551657464744741487748861081910719189662286392314162316577112654830964235951;
            6'd15: xpb[6] = 1024'd67092576557902427459779320103457313157360679335310695915222804008016809510174404534730219468350091533788723633658552145712375156114549802765475072858434988241304305844065035190245218487209821214876424474479399792703419050811347653794160959403885755113075201403055560419645773139902933411841098546363575573114;
            6'd16: xpb[6] = 1024'd79836528040704238717017869937342096217497953099380454584779781279549723166673307431046572180550609256670848503066288517731804422578267811920184086050086056852970637871640785358770248999124956343955532613337175768641271044213497282244770261343026768738401541724200401649629259887491704507105084437896186910277;
            6'd17: xpb[6] = 1024'd92580479523506049974256419771226879277635226863450213254336758551082636823172210327362924892751126979552973372474024889751233689041985821074893099241737125464636969899216535527295279511040091473034640752194951744579123037615646910695379563282167782363727882045345242879612746635080475602369070329428798247440;
            6'd18: xpb[6] = 1024'd105324431006307861231494969605111662337772500627519971923893735822615550479671113223679277604951644702435098241881761261770662955505703830229602112433388194076303301926792285695820310022955226602113748891052727720516975031017796539145988865221308795989054222366490084109596233382669246697633056220961409584603;
            6'd19: xpb[6] = 1024'd118068382489109672488733519438996445397909774391589730593450713094148464136170016119995630317152162425317223111289497633790092221969421839384311125625039262687969633954368035864345340534870361731192857029910503696454827024419946167596598167160449809614380562687634925339579720130258017792897042112494020921766;
            6'd20: xpb[6] = 1024'd6745638287786742347173141868066795713348621029923805134875835300704482455359780106296911814695005838756198573239740571230457647591919513983860013800359290365945291412372568695240131855268291138961767560381039826028318167601199023082228899416361373972886999594662708539456678803918155871042338177401037774598;
            6'd21: xpb[6] = 1024'd19489589770588553604411691701951578773485894793993563804432812572237396111858683002613264526895523561638323442647476943249886914055637523138569026992010358977611623439948318863765162367183426268040875699238815801966170161003348651532838201355502387598213339915807549769440165551506926966306324068933649111761;
            6'd22: xpb[6] = 1024'd32233541253390364861650241535836361833623168558063322473989789843770309768357585898929617239096041284520448312055213315269316180519355532293278040183661427589277955467524069032290192879098561397119983838096591777904022154405498279983447503294643401223539680236952390999423652299095698061570309960466260448924;
            6'd23: xpb[6] = 1024'd44977492736192176118888791369721144893760442322133081143546767115303223424856488795245969951296559007402573181462949687288745446983073541447987053375312496200944287495099819200815223391013696526199091976954367753841874147807647908434056805233784414848866020558097232229407139046684469156834295851998871786087;
            6'd24: xpb[6] = 1024'd57721444218993987376127341203605927953897716086202839813103744386836137081355391691562322663497076730284698050870686059308174713446791550602696066566963564812610619522675569369340253902928831655278200115812143729779726141209797536884666107172925428474192360879242073459390625794273240252098281743531483123250;
            6'd25: xpb[6] = 1024'd70465395701795798633365891037490711014034989850272598482660721658369050737854294587878675375697594453166822920278422431327603979910509559757405079758614633424276951550251319537865284414843966784357308254669919705717578134611947165335275409112066442099518701200386914689374112541862011347362267635064094460413;
            6'd26: xpb[6] = 1024'd83209347184597609890604440871375494074172263614342357152217698929901964394353197484195028087898112176048947789686158803347033246374227568912114092950265702035943283577827069706390314926759101913436416393527695681655430128014096793785884711051207455724845041521531755919357599289450782442626253526596705797576;
            6'd27: xpb[6] = 1024'd95953298667399421147842990705260277134309537378412115821774676201434878050852100380511380800098629898931072659093895175366462512837945578066823106141916770647609615605402819874915345438674237042515524532385471657593282121416246422236494012990348469350171381842676597149341086037039553537890239418129317134739;
            6'd28: xpb[6] = 1024'd108697250150201232405081540539145060194446811142481874491331653472967791707351003276827733512299147621813197528501631547385891779301663587221532119333567839259275947632978570043440375950589372171594632671243247633531134114818396050687103314929489482975497722163821438379324572784628324633154225309661928471902;
            6'd29: xpb[6] = 1024'd121441201633003043662320090373029843254584084906551633160888630744500705363849906173144086224499665344695322397909367919405321045765381596376241132525218907870942279660554320211965406462504507300673740810101023609468986108220545679137712616868630496600824062484966279609308059532217095728418211201194539809065;
            6'd30: xpb[6] = 1024'd10118457431680113520759712802100193570022931544885707702313752951056723683039670159445367722042508758134297859859610856845686471387879270975790020700538935548917937118558853042860197782902436708442651340571559739042477251401798534623343349124542060959330499391994062809185018205877233806563507266101556661897;
            6'd31: xpb[6] = 1024'd22862408914481924777998262635984976630160205308955466371870730222589637339538573055761720434243026481016422729267347228865115737851597280130499033892190004160584269146134603211385228294817571837521759479429335714980329244803948163073952651063683074584656839713138904039168504953466004901827493157634167999060;
            6'd32: xpb[6] = 1024'd35606360397283736035236812469869759690297479073025225041427707494122550996037475952078073146443544203898547598675083600884545004315315289285208047083841072772250601173710353379910258806732706966600867618287111690918181238206097791524561953002824088209983180034283745269151991701054775997091479049166779336223;
            6'd33: xpb[6] = 1024'd48350311880085547292475362303754542750434752837094983710984684765655464652536378848394425858644061926780672468082819972903974270779033298439917060275492141383916933201286103548435289318647842095679975757144887666856033231608247419975171254941965101835309520355428586499135478448643547092355464940699390673386;
            6'd34: xpb[6] = 1024'd61094263362887358549713912137639325810572026601164742380541662037188378309035281744710778570844579649662797337490556344923403537242751307594626073467143209995583265228861853716960319830562977224759083896002663642793885225010397048425780556881106115460635860676573427729118965196232318187619450832232002010549;
            6'd35: xpb[6] = 1024'd73838214845689169806952461971524108870709300365234501050098639308721291965534184641027131283045097372544922206898292716942832803706469316749335086658794278607249597256437603885485350342478112353838192034860439618731737218412546676876389858820247129085962200997718268959102451943821089282883436723764613347712;
            6'd36: xpb[6] = 1024'd86582166328490981064191011805408891930846574129304259719655616580254205622033087537343483995245615095427047076306029088962262070170187325904044099850445347218915929284013354054010380854393247482917300173718215594669589211814696305326999160759388142711288541318863110189085938691409860378147422615297224684875;
            6'd37: xpb[6] = 1024'd99326117811292792321429561639293674990983847893374018389212593851787119278531990433659836707446132818309171945713765460981691336633905335058753113042096415830582261311589104222535411366308382611996408312575991570607441205216845933777608462698529156336614881640007951419069425438998631473411408506829836022038;
            6'd38: xpb[6] = 1024'd112070069294094603578668111473178458051121121657443777058769571123320032935030893329976189419646650541191296815121501833001120603097623344213462126233747484442248593339164854391060441878223517741075516451433767546545293198618995562228217764637670169961941221961152792649052912186587402568675394398362447359201;
            6'd39: xpb[6] = 1024'd747325092771673437107733902248808366559968295777851600194693329876051254220657316277470917189493954630272277071744770441486028720121018813011014409067512120224250797169387221955233198621447148844426981904303676118784341800248417713848496893581734320447658868180575848929870860247540646820690463269464212033;
            6'd40: xpb[6] = 1024'd13491276575573484694346283736133591426697242059847610269751670601408964910719560212593823629390011677512397146479481142460915295183839027967720027600718580731890582824745137390480263710536582277923535120762079652056636335202398046164457798832722747945773999189325417078913357607836311742084676354802075549196;
            6'd41: xpb[6] = 1024'd26235228058375295951584833570018374486834515823917368939308647872941878567218463108910176341590529400394522015887217514480344561647557037122429040792369649343556914852320887559005294222451717407002643259619855627994488328604547674615067100771863761571100339510470258308896844355425082837348662246334686886359;
            6'd42: xpb[6] = 1024'd38979179541177107208823383403903157546971789587987127608865625144474792223717366005226529053791047123276646885294953886499773828111275046277138053984020717955223246879896637727530324734366852536081751398477631603932340322006697303065676402711004775196426679831615099538880331103013853932612648137867298223522;
            6'd43: xpb[6] = 1024'd51723131023978918466061933237787940607109063352056886278422602416007705880216268901542881765991564846158771754702690258519203094574993055431847067175671786566889578907472387896055355246281987665160859537335407579870192315408846931516285704650145788821753020152759940768863817850602625027876634029399909560685;
            6'd44: xpb[6] = 1024'd64467082506780729723300483071672723667246337116126644947979579687540619536715171797859234478192082569040896624110426630538632361038711064586556080367322855178555910935048138064580385758197122794239967676193183555808044308810996559966895006589286802447079360473904781998847304598191396123140619920932520897848;
            6'd45: xpb[6] = 1024'd77211033989582540980539032905557506727383610880196403617536556959073533193214074694175587190392600291923021493518163002558061627502429073741265093558973923790222242962623888233105416270112257923319075815050959531745896302213146188417504308528427816072405700795049623228830791345780167218404605812465132235011;
            6'd46: xpb[6] = 1024'd89954985472384352237777582739442289787520884644266162287093534230606446849712977590491939902593118014805146362925899374577490893966147082895974106750624992401888574990199638401630446782027393052398183953908735507683748295615295816868113610467568829697732041116194464458814278093368938313668591703997743572174;
            6'd47: xpb[6] = 1024'd102698936955186163495016132573327072847658158408335920956650511502139360506211880486808292614793635737687271232333635746596920160429865092050683119942276061013554907017775388570155477293942528181477292092766511483621600289017445445318722912406709843323058381437339305688797764840957709408932577595530354909337;
            6'd48: xpb[6] = 1024'd115442888437987974752254682407211855907795432172405679626207488773672274162710783383124645326994153460569396101741372118616349426893583101205392133133927129625221239045351138738680507805857663310556400231624287459559452282419595073769332214345850856948384721758484146918781251588546480504196563487062966246500;
            6'd49: xpb[6] = 1024'd4120144236665044610694304836282206223234278810739754167632610980228292481900547369425926824536996874008371563691615056056714852516080775804941021309247157303196896503355671569575299126255592718325310762094823589132943425600847929254962946601762421306891158665511930118658210262206618582341859551969983099332;
            6'd50: xpb[6] = 1024'd16864095719466855867932854670166989283371552574809512837189588251761206138399450265742279536737514596890496433099351428076144118979798784959650034500898225914863228530931421738100329638170727847404418900952599565070795419002997557705572248540903434932217498986656771348641697009795389677605845443502594436495;
            6'd51: xpb[6] = 1024'd29608047202268667125171404504051772343508826338879271506746565523294119794898353162058632248938032319772621302507087800095573385443516794114359047692549294526529560558507171906625360150085862976483527039810375541008647412405147186156181550480044448557543839307801612578625183757384160772869831335035205773658;
            6'd52: xpb[6] = 1024'd42351998685070478382409954337936555403646100102949030176303542794827033451397256058374984961138550042654746171914824172115002651907234803269068060884200363138195892586082922075150390662000998105562635178668151516946499405807296814606790852419185462182870179628946453808608670504972931868133817226567817110821;
            6'd53: xpb[6] = 1024'd55095950167872289639648504171821338463783373867018788845860520066359947107896158954691337673339067765536871041322560544134431918370952812423777074075851431749862224613658672243675421173916133234641743317525927492884351399209446443057400154358326475808196519950091295038592157252561702963397803118100428447984;
            6'd54: xpb[6] = 1024'd67839901650674100896887054005706121523920647631088547515417497337892860764395061851007690385539585488418995910730296916153861184834670821578486087267502500361528556641234422412200451685831268363720851456383703468822203392611596071508009456297467489433522860271236136268575644000150474058661789009633039785147;
            6'd55: xpb[6] = 1024'd80583853133475912154125603839590904584057921395158306184974474609425774420893964747324043097740103211301120780138033288173290451298388830733195100459153568973194888668810172580725482197746403492799959595241479444760055386013745699958618758236608503058849200592380977498559130747739245153925774901165651122310;
            6'd56: xpb[6] = 1024'd93327804616277723411364153673475687644195195159228064854531451880958688077392867643640395809940620934183245649545769660192719717762106839887904113650804637584861220696385922749250512709661538621879067734099255420697907379415895328409228060175749516684175540913525818728542617495328016249189760792698262459473;
            6'd57: xpb[6] = 1024'd106071756099079534668602703507360470704332468923297823524088429152491601733891770539956748522141138657065370518953506032212148984225824849042613126842455706196527552723961672917775543221576673750958175872957031396635759372818044956859837362114890530309501881234670659958526104242916787344453746684230873796636;
            6'd58: xpb[6] = 1024'd118815707581881345925841253341245253764469742687367582193645406424024515390390673436273101234341656379947495388361242404231578250689542858197322140034106774808193884751537423086300573733491808880037284011814807372573611366220194585310446664054031543934828221555815501188509590990505558439717732575763485133799;
            6'd59: xpb[6] = 1024'd7492963380558415784280875770315604079908589325701656735070528630580533709580437422574382731884499793386470850311485341671943676312040532796871028209426802486169542209541955917195365053889738287806194542285343502147102509401447440796077396309943108293334658462843284388386549664165696517863028640670501986631;
            6'd60: xpb[6] = 1024'd20236914863360227041519425604200387140045863089771415404627505902113447366079340318890735444085017516268595719719221713691372942775758541951580041401077871097835874237117706085720395565804873416885302681143119478084954502803597069246686698249084121918660998783988125618370036411754467613127014532203113323794;
            6'd61: xpb[6] = 1024'd32980866346162038298757975438085170200183136853841174074184483173646361022578243215207088156285535239150720589126958085710802209239476551106289054592728939709502206264693456254245426077720008545964410820000895454022806496205746697697296000188225135543987339105132966848353523159343238708391000423735724660957;
            6'd62: xpb[6] = 1024'd45724817828963849555996525271969953260320410617910932743741460445179274679077146111523440868486052962032845458534694457730231475703194560260998067784380008321168538292269206422770456589635143675043518958858671429960658489607896326147905302127366149169313679426277808078337009906932009803654986315268335998120;
            6'd63: xpb[6] = 1024'd58468769311765660813235075105854736320457684381980691413298437716712188335576049007839793580686570684914970327942430829749660742166912569415707080976031076932834870319844956591295487101550278804122627097716447405898510483010045954598514604066507162794640019747422649308320496654520780898918972206800947335283;
        endcase
    end

    always_comb begin
        case(flag[2][11:6])
            6'd0: xpb[7] = 1024'd0;
            6'd1: xpb[7] = 1024'd71212720794567472070473624939739519380594958146050450082855414988245101992074951904156146292887088407797095197350167201769090008630630578570416094167682145544501202347420706759820517613465413933201735236574223381836362476412195583049123906005648176419966360068567490538303983402109551994182958098333558672446;
            6'd2: xpb[7] = 1024'd18358745905010202742148322474664606016491489166365216037578974911513308646840764898297221371116502506151040987242840968959116176420040822585672063319033250155311730125270196182010796035413622145093272864761206917308364102603494393133269242328066903573112816723017923046501438730290470971247226370041522860561;
            6'd3: xpb[7] = 1024'd89571466699577674812621947414404125397086447312415666120434389899758410638915716802453367664003590913948136184593008170728206185050671401156088157486715395699812932472690902941831313648879036078295008101335430299144726579015689976182393148333715079993079176791585413584805422132400022965430184468375081533007;
            6'd4: xpb[7] = 1024'd36717491810020405484296644949329212032982978332730432075157949823026617293681529796594442742233005012302081974485681937918232352840081645171344126638066500310623460250540392364021592070827244290186545729522413834616728205206988786266538484656133807146225633446035846093002877460580941942494452740083045721122;
            6'd5: xpb[7] = 1024'd107930212604587877554770269889068731413577936478780882158013364811271719285756481700750589035120093420099177171835849139687322361470712223741760220805748645855124662597961099123842109684292658223388280966096637216453090681619184369315662390661781983566191993514603336631306860862690493936677410838416604393568;
            6'd6: xpb[7] = 1024'd55076237715030608226444967423993818049474467499095648112736924734539925940522294694891664113349507518453122961728522906877348529260122467757016189957099750465935190375810588546032388106240866435279818594283620751925092307810483179399807726984200710719338450169053769139504316190871412913741679110124568581683;
            6'd7: xpb[7] = 1024'd2222262825473338898119664958918904685370998519410414067460484657808132595288107689032739191578921616807068751621196674067374697049532711772272159108450855076745718153660077968222666528189074647171356222470604287397093934001781989483953063306619437872484906823504201647701771519052331890805947381832532769798;
            6'd8: xpb[7] = 1024'd73434983620040810968593289898658424065965956665460864150315899646053234587363059593188885484466010024604163948971363875836464705680163290342688253276133000621246920501080784728043184141654488580373091459044827669233456410413977572533076969312267614292451266892071692186005754921161883884988905480166091442244;
            6'd9: xpb[7] = 1024'd20581008730483541640267987433583510701862487685775630105039459569321441242128872587329960562695424122958109738864037643026490873469573534357944222427484105232057448278930274150233462563602696792264629087231811204705458036605276382617222305634686341445597723546522124694203210249342802862053173751874055630359;
            6'd10: xpb[7] = 1024'd91793729525051013710741612373323030082457445831826080187894874557566543234203824491486106855582512530755204936214204844795580882100204112928360316595166250776558650626350980910053980177068110725466364323806034586541820513017471965666346211640334517865564083615089615232507193651452354856236131850207614302805;
            6'd11: xpb[7] = 1024'd38939754635493744382416309908248116718353976852140846142618434480834749888969637485627181933811926629109150726106878611985607049889614356943616285746517355387369178404200470332244258599016318937357901951993018122013822139208770775750491547962753245018710540269540047740704648979633273833300400121915578490920;
            6'd12: xpb[7] = 1024'd110152475430061216452889934847987636098948934998191296225473849469079851881044589389783328226699015036906245923457045813754697058520244935514032379914199500931870380751621177092064776212481732870559637188567241503850184615620966358799615453968401421438676900338107538279008632381742825827483358220249137163366;
            6'd13: xpb[7] = 1024'd57298500540503947124564632382912722734845466018506062180197409392348058535810402383924403304928429135260191713349719580944723226309655179529288349065550605542680908529470666514255054634429941082451174816754225039322186241812265168883760790290820148591823356992557970787206087709923744804547626491957101351481;
            6'd14: xpb[7] = 1024'd4444525650946677796239329917837809370741997038820828134920969315616265190576215378065478383157843233614137503242393348134749394099065423544544318216901710153491436307320155936445333056378149294342712444941208574794187868003563978967906126613238875744969813647008403295403543038104663781611894763665065539596;
            6'd15: xpb[7] = 1024'd75657246445514149866712954857577328751336955184871278217776384303861367182651167282221624676044931641411232700592560549903839402729696002114960412384583855697992638654740862696265850669843563227544447681515431956630550344415759562017030032618887052164936173715575893833707526440214215775794852861998624212042;
            6'd16: xpb[7] = 1024'd22803271555956880538387652392502415387233486205186044172499944227129573837416980276362699754274345739765178490485234317093865570519106246130216381535934960308803166432590352118456129091791771439435985309702415492102551970607058372101175368941305779318082630370026326341904981768395134752859121133706588400157;
            6'd17: xpb[7] = 1024'd94015992350524352608861277332241934767828444351236494255355359215374675829491932180518846047161434147562273687835401518862955579149736824700632475703617105853304368780011058878276646705257185372637720546276638873938914447019253955150299274946953955738048990438593816880208965170504686747042079232040147072603;
            6'd18: xpb[7] = 1024'd41162017460967083280535974867167021403724975371551260210078919138642882484257745174659921125390848245916219477728075286052981746939147068715888444854968210464114896557860548300466925127205393584529258174463622409410916073210552765234444611269372682891195447093044249388406420498685605724106347503748111260718;
            6'd19: xpb[7] = 1024'd112374738255534555351009599806906540784319933517601710292934334126887984476332697078816067418277936653713314675078242487822071755569777647286304539022650356008616098905281255060287442740670807517730993411037845791247278549622748348283568517275020859311161807161611739926710403900795157718289305602081669933164;
            6'd20: xpb[7] = 1024'd59520763365977286022684297341831627420216464537916476247657894050156191131098510072957142496507350752067260464970916255012097923359187891301560508174001460619426626683130744482477721162619015729622531039224829326719280175814047158367713853597439586464308263816062172434907859228976076695353573873789634121279;
            6'd21: xpb[7] = 1024'd6666788476420016694358994876756714056112995558231242202381453973424397785864323067098217574736764850421206254863590022202124091148598135316816477325352565230237154460980233904667999584567223941514068667411812862191281802005345968451859189919858313617454720470512604943105314557156995672417842145497598309394;
            6'd22: xpb[7] = 1024'd77879509270987488764832619816496233436707953704281692285236868961669499777939274971254363867623853258218301452213757223971214099779228713887232571493034710774738356808400940664488517198032637874715803903986036244027644278417541551500983095925506490037421080539080095481409297959266547666600800243831156981840;
            6'd23: xpb[7] = 1024'd25025534381430219436507317351421320072604484724596458239960428884937706432705087965395438945853267356572247242106430991161240267568638957902488540644385815385548884586250430086678795619980846086607341532173019779499645904608840361585128432247925217190567537193530527989606753287447466643665068515539121169955;
            6'd24: xpb[7] = 1024'd96238255175997691506980942291160839453199442870646908322815843873182808424780039869551585238740355764369342439456598192930330276199269536472904634812067960930050086933671136846499313233446260019809076768747243161336008381021035944634252338253573393610533897262098018527910736689557018637848026613872679842401;
            6'd25: xpb[7] = 1024'd43384280286440422178655639826085926089095973890961674277539403796451015079545852863692660316969769862723288229349271960120356443988679780488160603963419065540860614711520626268689591655394468231700614396934226696808010007212334754718397674575992120763680353916548451036108192017737937614912294885580644030516;
            6'd26: xpb[7] = 1024'd114597001081007894249129264765825445469690932037012124360394818784696117071620804767848806609856858270520383426699439161889446452619310359058576698131101211085361817058941333028510109268859882164902349633508450078644372483624530337767521580581640297183646713985115941574412175419847489609095252983914202702962;
            6'd27: xpb[7] = 1024'd61743026191450624920803962300750532105587463057326890315118378707964323726386617761989881688086272368874329216592112929079472620408720603073832667282452315696172344836790822450700387690808090376793887261695433614116374109815829147851666916904059024336793170639566374082609630748028408586159521255622166891077;
            6'd28: xpb[7] = 1024'd8889051301893355592478659835675618741483994077641656269841938631232530381152430756130956766315686467228275006484786696269498788198130847089088636433803420306982872614640311872890666112756298588685424889882417149588375736007127957935812253226477751489939627294016806590807086076209327563223789527330131079192;
            6'd29: xpb[7] = 1024'd80101772096460827662952284775415138122078952223692106352697353619477632373227382660287103059202774875025370203834953898038588796828761425659504730601485565851484074962061018632711183726221712521887160126456640531424738212419323540984936159232125927909905987362584297129111069478318879557406747625663689751638;
            6'd30: xpb[7] = 1024'd27247797206903558334626982310340224757975483244006872307420913542745839027993195654428178137432188973379315993727627665228614964618171669674760699752836670462294602739910508054901462148169920733778697754643624066896739838610622351069081495554544655063052444017034729637308524806499798534471015897371653939753;
            6'd31: xpb[7] = 1024'd98460518001471030405100607250079744138570441390057322390276328530990941020068147558584324430319277381176411191077794866997704973248802248245176793920518816006795805087331214814721979761635334666980432991217847448733102315022817934118205401560192831483018804085602220175612508208609350528653973995705212612199;
            6'd32: xpb[7] = 1024'd45606543111913761076775304785004830774466972410372088344999888454259147674833960552725399508548691479530356980970468634187731141038212492260432763071869920617606332865180704236912258183583542878871970619404830984205103941214116744202350737882611558636165260740052652683809963536790269505718242267413176800314;
            6'd33: xpb[7] = 1024'd116819263906481233147248929724744350155061930556422538427855303442504249666908912456881545801435779887327452178320635835956821149668843070830848857239552066162107535212601410996732775797048956812073705855979054366041466417626312327251474643888259735056131620808620143222113946938899821499901200365746735472760;
            6'd34: xpb[7] = 1024'd63965289016923963818923627259669436790958461576737304382578863365772456321674725451022620879665193985681397968213309603146847317458253314846104826390903170772918062990450900418923054218997165023965243484166037901513468043817611137335619980210678462209278077463070575730311402267080740476965468637454699660875;
            6'd35: xpb[7] = 1024'd11111314127366694490598324794594523426854992597052070337302423289040662976440538445163695957894608084035343758105983370336873485247663558861360795542254275383728590768300389841113332640945373235856781112353021436985469670008909947419765316533097189362424534117521008238508857595261659454029736909162663848990;
            6'd36: xpb[7] = 1024'd82324034921934166561071949734334042807449950743102520420157838277285764968515490349319842250781696491832438955456150572105963493878294137431776889709936420928229793115721096600933850254410787169058516348927244818821832146421105530468889222538745365782390894186088498776812840997371211448212695007496222521436;
            6'd37: xpb[7] = 1024'd29470060032376897232746647269259129443346481763417286374881398200553971623281303343460917329011110590186384745348824339295989661667704381447032858861287525539040320893570586023124128676358995380950053977114228354293833772612404340553034558861164092935537350840538931285010296325552130425276963279204186709551;
            6'd38: xpb[7] = 1024'd100682780826944369303220272208998648823941439909467736457736813188799073615356255247617063621898198997983479942698991541065079670298334960017448953028969671083541523240991292782944646289824409314151789213688451736130196249024599923602158464866812269355503710909106421823314279727661682419459921377537745381997;
            6'd39: xpb[7] = 1024'd47828805937387099974894969743923735459837970929782502412460373112067280270122068241758138700127613096337425732591665308255105838087745204032704922180320775694352051018840782205134924711772617526043326841875435271602197875215898733686303801189230996508650167563556854331511735055842601396524189649245709570112;
            6'd40: xpb[7] = 1024'd119041526731954572045368594683663254840432929075832952495315788100312382262197020145914284993014701504134520929941832510024195846718375782603121016348002921238853253366261488964955442325238031459245062078449658653438560351628094316735427707194879172928616527632124344869815718457952153390707147747579268242558;
            6'd41: xpb[7] = 1024'd66187551842397302717043292218588341476329460096147718450039348023580588916962833140055360071244115602488466719834506277214222014507786026618376985499354025849663781144110978387145720747186239671136599706636642188910561977819393126819573043517297900081762984286574777378013173786133072367771416019287232430673;
            6'd42: xpb[7] = 1024'd13333576952840033388717989753513428112225991116462484404762907946848795571728646134196435149473529700842412509727180044404248182297196270633632954650705130460474308921960467809335999169134447883028137334823625724382563604010691936903718379839716627234909440941025209886210629114313991344835684290995196618788;
            6'd43: xpb[7] = 1024'd84546297747407505459191614693252947492820949262512934487618322935093897563803598038352581442360618108639507707077347246173338190927826849204049048818387276004975511269381174569156516782599861816229872571397849106218926080422887519952842285845364803654875801009592700424514612516423543339018642389328755291234;
            6'd44: xpb[7] = 1024'd31692322857850236130866312228178034128717480282827700442341882858362104218569411032493656520590032206993453496970021013363364358717237093219305017969738380615786039047230663991346795204548070028121410199584832641690927706614186330036987622167783530808022257664043132932712067844604462316082910661036719479349;
            6'd45: xpb[7] = 1024'd102905043652417708201339937167917553509312438428878150525197297846607206210644362936649802813477120614790548694320188215132454367347867671789721112137420526160287241394651370751167312818013483961323145436159056023527290183026381913086111528173431707227988617732610623471016051246714014310265868759370278151795;
            6'd46: xpb[7] = 1024'd50051068762860438873014634702842640145208969449192916479920857769875412865410175930790877891706534713144494484212861982322480535137277915804977081288771630771097769172500860173357591239961692173214683064346039558999291809217680723170256864495850434381135074387061055979213506574894933287330137031078242339910;
            6'd47: xpb[7] = 1024'd121263789557427910943488259642582159525803927595243366562776272758120514857485127834947024184593623120941589681563029184091570543767908494375393175456453776315598971519921566933178108853427106106416418300920262940835654285629876306219380770501498610801101434455628546517517489977004485281513095129411801012356;
            6'd48: xpb[7] = 1024'd68409814667870641615162957177507246161700458615558132517499832681388721512250940829088099262823037219295535471455702951281596711557318738390649144607804880926409499297771056355368387275375314318307955929107246476307655911821175116303526106823917337954247891110078979025714945305185404258577363401119765200471;
            6'd49: xpb[7] = 1024'd15555839778313372286837654712432332797596989635872898472223392604656928167016753823229174341052451317649481261348376718471622879346728982405905113759155985537220027075620545777558665697323522530199493557294230011779657538012473926387671443146336065107394347764529411533912400633366323235641631672827729388586;
            6'd50: xpb[7] = 1024'd86768560572880844357311279652171852178191947781923348555078807592902030159091705727385320633939539725446576458698543920240712887977359560976321207926838131081721229423041252537379183310788936463401228793868453393616020014424669509436795349151984241527360707833096902072216384035475875229824589771161288061032;
            6'd51: xpb[7] = 1024'd33914585683323575028985977187096938814088478802238114509802367516170236813857518721526395712168953823800522248591217687430739055766769804991577177078189235692531757200890741959569461732737144675292766422055436929088021640615968319520940685474402968680507164487547334580413839363656794206888858042869252249147;
            6'd52: xpb[7] = 1024'd105127306477891047099459602126836458194683436948288564592657782504415338805932470625682542005056042231597617445941384889199829064397400383561993271245871381237032959548311448719389979346202558608494501658629660310924384117028163902570064591480051145100473524556114825118717822765766346201071816141202810921593;
            6'd53: xpb[7] = 1024'd52273331588333777771134299661761544830579967968603330547381342427683545460698283619823617083285456329951563235834058656389855232186810627577249240397222485847843487326160938141580257768150766820386039286816643846396385743219462712654209927802469872253619981210565257626915278093947265178136084412910775109708;
            6'd54: xpb[7] = 1024'd123486052382901249841607924601501064211174926114653780630236757415928647452773235523979763376172544737748658433184225858158945240817441206147665334564904631392344689673581644901400775381616180753587774523390867228232748219631658295703333833808118048673586341279132748165219261496056817172319042511244333782154;
            6'd55: xpb[7] = 1024'd70632077493343980513282622136426150847071457134968546584960317339196854107539048518120838454401958836102604223076899625348971408606851450162921303716255736003155217451431134323591053803564388965479312151577850763704749845822957105787479170130536775826732797933583180673416716824237736149383310782952297970269;
            6'd56: xpb[7] = 1024'd17778102603786711184957319671351237482967988155283312539683877262465060762304861512261913532631372934456550012969573392538997576396261694178177272867606840613965745229280623745781332225512597177370849779764834299176751472014255915871624506452955502979879254588033613181614172152418655126447579054660262158384;
            6'd57: xpb[7] = 1024'd88990823398354183255430944611090756863562946301333762622539292250710162754379813416418059825518461342253645210319740594308087585026892272748593367035288986158466947576701330505601849838978011110572585016339057681013113948426451498920748412458603679399845614656601103719918155554528207120630537152993820830830;
            6'd58: xpb[7] = 1024'd36136848508796913927105642146015843499459477321648528577262852173978369409145626410559134903747875440607591000212414361498113752816302516763849336186640090769277475354550819927792128260926219322464122644526041216485115574617750309004893748781022406552992071311051536228115610882709126097694805424701785018945;
            6'd59: xpb[7] = 1024'd107349569303364385997579267085755362880054435467698978660118267162223471401220578314715281196634963848404686197562581563267203761446933095334265430354322236313778677701971526687612645874391633255665857881100264598321478051029945892054017654786670582972958431379619026766419594284818678091877763523035343691391;
            6'd60: xpb[7] = 1024'd54495594413807116669253964620680449515950966488013744614841827085491678055986391308856356274864377946758631987455255330457229929236343339349521399505673340924589205479821016109802924296339841467557395509287248133793479677221244702138162991109089310126104888034069459274617049612999597068942031794743307879506;
            6'd61: xpb[7] = 1024'd1641619524249847340928662155605536151847497508328510569565387008759884710752204302997431353093792045112577777347929097647256097025753583364777368657024445535399733257670505531993202718288049679448933137474231669265481303412543512222308327431508037279251344688519891782814504941180516046006300066451272067621;
            6'd62: xpb[7] = 1024'd72854340318817319411402287095345055532442455654378960652420801997004986702827156207153577645980880452909672974698096299416346105656384161935193462824706591079900935605091212291813720331753463612650668374048455051101843779824739095271432233437156213699217704757087382321118488343290068040189258164784830740067;
            6'd63: xpb[7] = 1024'd20000365429260050083076984630270142168338986674693726607144361920273193357592969201294652724210294551263618764590770066606372273445794405950449431976057695690711463382940701714003998753701671824542206002235438586573845406016037905355577569759574940852364161411537814829315943671470987017253526436492794928182;
        endcase
    end

    always_comb begin
        case(flag[2][16:12])
            5'd0: xpb[8] = 1024'd0;
            5'd1: xpb[8] = 1024'd91213086223827522153550609570009661548933944820744176689999776908518295349667921105450799017097382959060713961940937268375462282076424984520865526143739841235212665730361408473824516367167085757743941238809661968410207882428233488404701475765223117272330521480105305367619927073580539011436484534826353600628;
            5'd2: xpb[8] = 1024'd58359476763530302908302291735204890353169462515752669251867698752059695362026703300886526819537091608678278516424381102171860723311629634486570927271148641536734656891151599610018793542816965794177684869232084090456054914635570203844424381847216785277841139546093552705133326073232445005754279243027112716925;
            5'd3: xpb[8] = 1024'd25505867303233083663053973900400119157404980210761161813735620595601095374385485496322254621976800258295843070907824935968259164546834284452276328398557441838256648051941790746213070718466845830611428499654506212501901946842906919284147287929210453283351757612081800042646725072884351000072073951227871833222;
            5'd4: xpb[8] = 1024'd116718953527060605816604583470409780706338925031505338503735397504119390724053406601773053639074183217356557032848762204343721446623259268973141854542297283073469313782303199220037587085633931588355369738464168180912109829271140407688848763694433570555682279092187105410266652146464890011508558486054225433850;
            5'd5: xpb[8] = 1024'd83865344066763386571356265635605009510574442726513831065603319347660790736412188797208781441513891866974121587332206038140119887858463918938847255669706083374991304943093390356231864261283811624789113368886590302957956861478477123128571669776427238561192897158175352747780051146116796005826353194254984550147;
            5'd6: xpb[8] = 1024'd51011734606466167326107947800800238314809960421522323627471241191202190748770970992644509243953600516591686141815649871936518329093668568904552656797114883676513296103883581492426141436933691661222856999309012425003803893685813838568294575858420906566703515224163600085293450145768702000144147902455743666444;
            5'd7: xpb[8] = 1024'd18158125146168948080859629965995467119045478116530816189339163034743590761129753188080237046393309166209250696299093705732916770328873218870258057924523683978035287264673772628620418612583571697656600629731434547049650925893150554008017481940414574572214133290151847422806849145420607994461942610656502782741;
            5'd8: xpb[8] = 1024'd109371211369996470234410239536005128667979422937274992879338939943261886110797674293531036063490692125269964658240030974108379052405298203391123584068263525213247952995035181102444934979750657455400541868541096515459858808321384042412718957705637691844544654770257152790426776219001147005898427145482856383369;
            5'd9: xpb[8] = 1024'd76517601909699250989161921701200357472214940632283485441206861786803286123156456488966763865930400774887529212723474807904777493640502853356828985195672325514769944155825372238639212155400537491834285498963518637505705840528720757852441863787631359850055272836245400127940175218653053000216221853683615499666;
            5'd10: xpb[8] = 1024'd43663992449402031743913603866395586276450458327291978003074783630344686135515238684402491668370109424505093767206918641701175934875707503322534386323081125816291935316615563374833489331050417528268029129385940759551552872736057473292164769869625027855565890902233647465453574218304958994534016561884374615963;
            5'd11: xpb[8] = 1024'd10810382989104812498665286031590815080685976022300470564942705473886086147874020879838219470809818074122658321690362475497574376110912153288239787450489926117813926477405754511027766506700297564701772759808362881597399904943394188731887675951618695861076508968221894802966973217956864988851811270085133732260;
            5'd12: xpb[8] = 1024'd102023469212932334652215895601600476629619920843044647254942482382404381497541941985289018487907201033183372283631299743873036658187337137809105313594229767353026592207767162984852282873867383322445713998618024850007607787371627677136589151716841813133407030448327200170586900291537404000288295804911487332888;
            5'd13: xpb[8] = 1024'd69169859752635115406967577766795705433855438538053139816810404225945781509900724180724746290346909682800936838114743577669435099422541787774810714721638567654548583368557354121046560049517263358879457629040446972053454819578964392576312057798835481138917648514315447508100299291189309994606090513112246449185;
            5'd14: xpb[8] = 1024'd36316250292337896161719259931990934238090956233061632378678326069487181522259506376160474092786618332418501392598187411465833540657746437740516115849047367956070574529347545257240837225167143395313201259462869094099301851786301108016034963880829149144428266580303694845613698290841215988923885221313005565482;
            5'd15: xpb[8] = 1024'd3462640832040676916470942097186163042326473928070124940546247913028581534618288571596201895226326982036065947081631245262231981892951087706221516976456168257592565690137736393435114400817023431746944889885291216145148883993637823455757869962822817149938884646291942183127097290493121983241679929513764681779;
            5'd16: xpb[8] = 1024'd94675727055868199070021551667195824591260418748814301630546024821546876884286209677047000912323709941096779909022568513637694263969376072227087043120196009492805231420499144867259630767984109189490886128694953184555356766421871311860459345728045934422269406126397247550747024364073660994678164464340118282407;
            5'd17: xpb[8] = 1024'd61822117595570979824773233832391053395495936443822794192413946665088276896644991872482728714763418590714344463506012347434092705204580722192792444247604809794327222581289336003453907943633989225924629759117375306601203798629208027300182251810039602427780024192385494888260423363725566988995959172540877398704;
            5'd18: xpb[8] = 1024'd28968508135273760579524915997586282199731454138831286754281868508629676909003774067918456517203127240331909017989456181230491146439785372158497845375013610095849213742079527139648185119283869262358373389539797428647050830836544742739905157892033270433290642258373742225773822363377472983313753880741636515001;
            5'd19: xpb[8] = 1024'd120181594359101282733075525567595943748665398959575463444281645417147972258671695173369255534300510199392622979930393449605953428516210356679363371518753451331061879472440935613472701486450955020102314628349459397057258713264778231144606633657256387705621163738479047593393749436958011994750238415567990115629;
            5'd20: xpb[8] = 1024'd87327984898804063487827207732791172552900916654583956006149567260689372271030477368804983336740218849010187534413837283402351869751415006645068772646162251632583870633231126749666978662100835056536058258771881519103105745472114946584329539739250055711131781804467294930907148436609917989068033123768749231926;
            5'd21: xpb[8] = 1024'd54474375438506844242578889897986401357136434349592448568017489104230772283389259564240711139179927498627752088897281117198750310986619656610774173773571051934105861794021317885861255837750715092969801889194303641148952777679451662024052445821243723716642399870455542268420547436261823983385827831969508348223;
            5'd22: xpb[8] = 1024'd21620765978209624997330572063181630161371952044600941129885410947772172295748041759676438941619636148245316643380724950995148752221824306576479574900979852235627852954811509022055533013400595129403545519616725763194799809886788377463775351903237391722153017936443789605933946435913729977703622540170267464520;
            5'd23: xpb[8] = 1024'd112833852202037147150881181633191291710305896865345117819885187856290467645415962865127237958717019107306030605321662219370611034298249291097345101044719693470840518685172917495880049380567680887147486758426387731605007692315021865868476827668460508994483539416549094973553873509494268989140107074996621065148;
            5'd24: xpb[8] = 1024'd79980242741739927905632863798386520514541414560353610381753109699831867657774745060562965761156727756923595159805106053167009475533453941063050502172128493772362509845963108632074326556217560923581230388848809853650854724522358581308199733750454176999994157482537342311067272509146174983457901783197380181445;
            5'd25: xpb[8] = 1024'd47126633281442708660384545963581749318776932255362102943621031543373267670133527255998693563596436406541159714288549886963407916768658591028755903299537294073884501006753299768268603731867440960014974019271231975696701756729695296747922639832447845005504775548525589648580671508798080977775696491398139297742;
            5'd26: xpb[8] = 1024'd14273023821145489415136228128776978123012449950370595505488953386914667682492309451434421366036145056158724268771993720759806358003863240994461304426946094375406492167543490904462880907517320996448717649693654097742548788937032012187645545914441513011015393614513836986094070508449986972093491199598898414039;
            5'd27: xpb[8] = 1024'd105486110044973011568686837698786639671946394771114772195488730295432963032160230556885220383133528015219438230712930989135268640080288225515326830570685935610619157897904899378287397274684406754192658888503316066152756671365265500592347021679664630283345915094619142353713997582030525983529975734425252014667;
            5'd28: xpb[8] = 1024'd72632500584675792323438519863981868476181912466123264757356652138974363044519012752320948185573236664837002785196374822931667081315492875481032231698094735912141149058695090514481674450334286790626402518925738188198603703572602216032069927761658298288856533160607389691227396581682431977847770442626011130964;
            5'd29: xpb[8] = 1024'd39778891124378573078190202029177097280417430161131757319224573982515763056877794947756675988012945314454567339679818656728065522550697525446737632825503536213663140219485281650675951625984166827060146149348160310244450735779938931471792833843651966294367151226595637028740795581334337972165565150826770247261;
            5'd30: xpb[8] = 1024'd6925281664081353832941884194372326084652947856140249881092495826057163069236577143192403790452653964072131894163262490524463963785902175412443033952912336515185131380275472786870228801634046863493889779770582432290297767987275646911515739925645634299877769292583884366254194580986243966483359859027529363558;
            5'd31: xpb[8] = 1024'd98138367887908875986492493764381987633586892676884426571092272734575458418904498248643202807550036923132845856104199758899926245862327159933308560096652177750397797110636881260694745168801132621237831018580244400700505650415509135316217215690868751572208290772689189733874121654566782977919844393853882964186;
        endcase
    end



endmodule



module xpb_lut_high
(
    input logic [16:0] flag[66],
    output logic [1023:0] xpb[198]
);
        
        
    always_comb begin
        case(flag[0][5:0])
            6'd0: xpb[0] = 1024'd0;
            6'd1: xpb[0] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            6'd2: xpb[0] = 1024'd100679634060304071055502914952736037167277100005316212353815420990297612207887079213229586029714185122074147583574573231666989319490825001042645800577467357194103405572860590087130560771855039443069108389671751481037922888800575812974249138053854169508899944397738886563714375961321529215371653600027243516363;
            6'd3: xpb[0] = 1024'd88986103248393735883854908726696839378566436445106476466657203952957970643176049364836843437242440528389646671633113130210952058815627334286388638358035515324309771074505276461880721562023956303948563780314007298374703908090415332978884422239166529629939964889549800830518299905017977314498135486728068032379;
            6'd4: xpb[0] = 1024'd77292572436483400712206902500657641589855772884896740579498986915618329078465019516444100844770695934705145759691653028754914798140429667530131476138603673454516136576149962836630882352192873164828019170956263115711484927380254852983519706424478889750979985381360715097322223848714425413624617373428892548395;
            6'd5: xpb[0] = 1024'd65599041624573065540558896274618443801145109324687004692340769878278687513753989668051358252298951341020644847750192927298877537465232000773874313919171831584722502077794649211381043142361790025707474561598518933048265946670094372988154990609791249872020005873171629364126147792410873512751099260129717064411;
            6'd6: xpb[0] = 1024'd53905510812662730368910890048579246012434445764477268805182552840939045949042959819658615659827206747336143935808732825842840276790034334017617151699739989714928867579439335586131203932530706886586929952240774750385046965959933892992790274795103609993060026364982543630930071736107321611877581146830541580427;
            6'd7: xpb[0] = 1024'd42211980000752395197262883822540048223723782204267532918024335803599404384331929971265873067355462153651643023867272724386803016114836667261359989480308147845135233081084021960881364722699623747466385342883030567721827985249773412997425558980415970114100046856793457897733995679803769711004063033531366096443;
            6'd8: xpb[0] = 1024'd30518449188842060025614877596500850435013118644057797030866118766259762819620900122873130474883717559967142111925812622930765755439639000505102827260876305975341598582728708335631525512868540608345840733525286385058609004539612933002060843165728330235140067348604372164537919623500217810130544920232190612459;
            6'd9: xpb[0] = 1024'd18824918376931724853966871370461652646302455083848061143707901728920121254909870274480387882411972966282641199984352521474728494764441333748845665041444464105547964084373394710381686303037457469225296124167542202395390023829452453006696127351040690356180087840415286431341843567196665909257026806933015128475;
            6'd10: xpb[0] = 1024'd7131387565021389682318865144422454857591791523638325256549684691580479690198840426087645289940228372598140288042892420018691234089243666992588502822012622235754329586018081085131847093206374330104751514809798019732171043119291973011331411536353050477220108332226200698145767510893114008383508693633839644491;
            6'd11: xpb[0] = 1024'd119504552437235795909469786323197689813579555089164273497523322719217733462796949487709973912126158088356788783558925753141717814255266334791491465618911821299651369657233984797512247074892496912294404513839293683433312912630028265980945265404894859865080032238154172995056219528518195124628680406960258644838;
            6'd12: xpb[0] = 1024'd107811021625325460737821780097158492024868891528954537610365105681878091898085919639317231319654413494672287871617465651685680553580068668035234303399479979429857735158878671172262407865061413773173859904481549500770093931919867785985580549590207219986120052729965087261860143472214643223755162293661083160854;
            6'd13: xpb[0] = 1024'd96117490813415125566173773871119294236158227968744801723206888644538450333374889790924488727182668900987786959676005550229643292904871001278977141180048137560064100660523357547012568655230330634053315295123805318106874951209707305990215833775519580107160073221776001528664067415911091322881644180361907676870;
            6'd14: xpb[0] = 1024'd84423960001504790394525767645080096447447564408535065836048671607198808768663859942531746134710924307303286047734545448773606032229673334522719978960616295690270466162168043921762729445399247494932770685766061135443655970499546825994851117960831940228200093713586915795467991359607539422008126067062732192886;
            6'd15: xpb[0] = 1024'd72730429189594455222877761419040898658736900848325329948890454569859167203952830094139003542239179713618785135793085347317568771554475667766462816741184453820476831663812730296512890235568164355812226076408316952780436989789386345999486402146144300349240114205397830062271915303303987521134607953763556708902;
            6'd16: xpb[0] = 1024'd61036898377684120051229755193001700870026237288115594061732237532519525639241800245746260949767435119934284223851625245861531510879278001010205654521752611950683197165457416671263051025737081216691681467050572770117218009079225866004121686331456660470280134697208744329075839247000435620261089840464381224918;
            6'd17: xpb[0] = 1024'd49343367565773784879581748966962503081315573727905858174574020495179884074530770397353518357295690526249783311910165144405494250204080334253948492302320770080889562667102103046013211815905998077571136857692828587453999028369065386008756970516769020591320155189019658595879763190696883719387571727165205740934;
            6'd18: xpb[0] = 1024'd37649836753863449707933742740923305292604910167696122287415803457840242509819740548960775764823945932565282399968705042949456989528882667497691330082888928211095928168746789420763372606074914938450592248335084404790780047658904906013392254702081380712360175680830572862683687134393331818514053613866030256950;
            6'd19: xpb[0] = 1024'd25956305941953114536285736514884107503894246607486386400257586420500600945108710700568033172352201338880781488027244941493419728853685000741434167863457086341302293670391475795513533396243831799330047638977340222127561066948744426018027538887393740833400196172641487129487611078089779917640535500566854772966;
            6'd20: xpb[0] = 1024'd14262775130042779364637730288844909715183583047276650513099369383160959380397680852175290579880456745196280576085784840037382468178487333985177005644025244471508659172036162170263694186412748660209503029619596039464342086238583946022662823072706100954440216664452401396291535021786228016767017387267679288982;
            6'd21: xpb[0] = 1024'd2569244318132444192989724062805711926472919487066914625941152345821317815686651003782547987408712151511779664144324738581345207503289667228919843424593402601715024673680848545013854976581665521088958420261851856801123105528423466027298107258018461075480237156263315663095458965482676115893499273968503804998;
            6'd22: xpb[0] = 1024'd114942409190346850420140645241580946882460683052592862866914790373458571588284760065404876609594641867270428159660358071704371787669312335027822806221492601665612064744896752257394254958267788103278611419291347520502264975039159758996911961126560270463340161062191287960005910983107757232138670987294922805345;
            6'd23: xpb[0] = 1024'd103248878378436515248492639015541749093750019492383126979756573336118930023573730217012134017122897273585927247718897970248334526994114668271565644002060759795818430246541438632144415748436704964158066809933603337839045994328999279001547245311872630584380181554002202226809834926804205331265152873995747321361;
            6'd24: xpb[0] = 1024'd91555347566526180076844632789502551305039355932173391092598356298779288458862700368619391424651152679901426335777437868792297266318917001515308481782628917926024795748186125006894576538605621825037522200575859155175827013618838799006182529497184990705420202045813116493613758870500653430391634760696571837377;
            6'd25: xpb[0] = 1024'd79861816754615844905196626563463353516328692371963655205440139261439646894151670520226648832179408086216925423835977767336260005643719334759051319563197076056231161249830811381644737328774538685916977591218114972512608032908678319010817813682497350826460222537624030760417682814197101529518116647397396353393;
            6'd26: xpb[0] = 1024'd68168285942705509733548620337424155727618028811753919318281922224100005329440640671833906239707663492532424511894517665880222744968521668002794157343765234186437526751475497756394898118943455546796432981860370789849389052198517839015453097867809710947500243029434945027221606757893549628644598534098220869409;
            6'd27: xpb[0] = 1024'd56474755130795174561900614111384957938907365251544183431123705186760363764729610823441163647235918898847923599953057564424185484293324001246536995124333392316643892253120184131145058909112372407675888372502626607186170071488357359020088382053122071068540263521245859294025530701589997727771080420799045385425;
            6'd28: xpb[0] = 1024'd44781224318884839390252607885345760150196701691334447543965488149420722200018580975048421054764174305163422688011597462968148223618126334490279832904901550446850257754764870505895219699281289268555343763144882424522951090778196879024723666238434431189580284013056773560829454645286445826897562307499869901441;
            6'd29: xpb[0] = 1024'd33087693506974504218604601659306562361486038131124711656807271112081080635307551126655678462292429711478921776070137361512110962942928667734022670685469708577056623256409556880645380489450206129434799153787138241859732110068036399029358950423746791310620304504867687827633378588982893926024044194200694417457;
            6'd30: xpb[0] = 1024'd21394162695064169046956595433267364572775374570914975769649054074741439070596521278262935869820685117794420864128677260056073702267731000977765508466037866707262988758054243255395541279619122990314254544429394059196513129357875919033994234609059151431660324996678602094437302532679342025150526080901518933473;
            6'd31: xpb[0] = 1024'd9700631883153833875308589207228166784064711010705239882490837037401797505885491429870193277348940524109919952187217158600036441592533334221508346246606024837469354259698929630145702069788039851193709935071649876533294148647715439038629518794371511552700345488489516361241226476375790124277007967602343449489;
            6'd32: xpb[0] = 1024'd122073796755368240102459510386003401740052474576231188123464475065039051278483600491492521899534870239868568447703250491723063021758556002020411309043505223901366394330914833342526102051474162433383362934101145540234436018158451732008243372662913320940560269394417488658151678494000871240522179680928762449836;
            6'd33: xpb[0] = 1024'd110380265943457904930811504159964203951341811016021452236306258027699409713772570643099779307063125646184067535761790390267025761083358335264154146824073382031572759832559519717276262841643079294262818324743401357571217037448291252012878656848225681061600289886228402924955602437697319339648661567629586965852;
            6'd34: xpb[0] = 1024'd98686735131547569759163497933925006162631147455811716349148040990359768149061540794707036714591381052499566623820330288810988500408160668507896984604641540161779125334204206092026423631811996155142273715385657174907998056738130772017513941033538041182640310378039317191759526381393767438775143454330411481868;
            6'd35: xpb[0] = 1024'd86993204319637234587515491707885808373920483895601980461989823953020126584350510946314294122119636458815065711878870187354951239732963001751639822385209698291985490835848892466776584421980913016021729106027912992244779076027970292022149225218850401303680330869850231458563450325090215537901625341031235997884;
            6'd36: xpb[0] = 1024'd75299673507726899415867485481846610585209820335392244574831606915680485019639481097921551529647891865130564799937410085898913979057765334995382660165777856422191856337493578841526745212149829876901184496670168809581560095317809812026784509404162761424720351361661145725367374268786663637028107227732060513900;
            6'd37: xpb[0] = 1024'd63606142695816564244219479255807412796499156775182508687673389878340843454928451249528808937176147271446063887995949984442876718382567668239125497946346014552398221839138265216276906002318746737780639887312424626918341114607649332031419793589475121545760371853472059992171298212483111736154589114432885029916;
            6'd38: xpb[0] = 1024'd51912611883906229072571473029768215007788493214972772800515172841001201890217421401136066344704402677761562976054489882986839457707370001482868335726914172682604587340782951591027066792487663598660095277954680444255122133897488852036055077774787481666800392345282974258975222156179559835281071001133709545932;
            6'd39: xpb[0] = 1024'd40219081071995893900923466803729017219077829654763036913356955803661560325506391552743323752232658084077062064113029781530802197032172334726611173507482330812810952842427637965777227582656580459539550668596936261591903153187328372040690361960099841787840412837093888525779146099876007934407552887834534061948;
            6'd40: xpb[0] = 1024'd28525550260085558729275460577689819430367166094553301026198738766321918760795361704350581159760913490392561152171569680074764936356974667970354011288050488943017318344072324340527388372825497320419006059239192078928684172477167892045325646145412201908880433328904802792583070043572456033534034774535358577964;
            6'd41: xpb[0] = 1024'd16832019448175223557627454351650621641656502534343565139040521728982277196084331855957838567289168896708060240230109578618727675681777001214096849068618647073223683845717010715277549162994414181298461449881447896265465191767007412049960930330724562029920453820715717059386993987268904132660516661236183093980;
            6'd42: xpb[0] = 1024'd5138488636264888385979448125611423852945838974133829251882304691642635631373302007565095974817424303023559328288649477162690415006579334457839686849186805203430049347361697090027709953163331042177916840523703713602246211056846932054596214516036922150960474312526631326190917930965352231786998547937007609996;
            6'd43: xpb[0] = 1024'd117511653508479294613130369304386658808933602539659777492855942719279889403971411069187424597003354018782207823804682810285716995172602002256742649646086004267327089418577600802408109934849453624367569839553199377303388080567583225024210068384578731538820398218454603623101369948590433348032170261263426610343;
            6'd44: xpb[0] = 1024'd105818122696568959441482363078347461020222938979450041605697725681940247839260381220794682004531609425097706911863222708829679734497404335500485487426654162397533454920222287177158270725018370485247025230195455194640169099857422745028845352569891091659860418710265517889905293892286881447158652147964251126359;
            6'd45: xpb[0] = 1024'd94124591884658624269834356852308263231512275419240305718539508644600606274549351372401939412059864831413205999921762607373642473822206668744228325207222320527739820421866973551908431515187287346126480620837711011976950119147262265033480636755203451780900439202076432156709217835983329546285134034665075642375;
            6'd46: xpb[0] = 1024'd82431061072748289098186350626269065442801611859030569831381291607260964709838321524009196819588120237728705087980302505917605213147009001987971162987790478657946185923511659926658592305356204207005936011479966829313731138437101785038115920940515811901940459693887346423513141779679777645411615921365900158391;
            6'd47: xpb[0] = 1024'd70737530260837953926538344400229867654090948298820833944223074569921323145127291675616454227116375644044204176038842404461567952471811335231714000768358636788152551425156346301408753095525121067885391402122222646650512157726941305042751205125828172022980480185698260690317065723376225744538097808066724674407;
            6'd48: xpb[0] = 1024'd59043999448927618754890338174190669865380284738611098057064857532581681580416261827223711634644631050359703264097382303005530691796613668475456838548926794918358916926801032676158913885694037928764846792764478463987293177016780825047386489311140532144020500677509174957120989667072673843664579694767549190423;
            6'd49: xpb[0] = 1024'd47350468637017283583242331948151472076669621178401362169906640495242040015705231978830969042172886456675202352155922201549493431121416001719199676329494953048565282428445719050909074675862954789644302183406734281324074196306620345052021773496452892265060521169320089223924913610769121942791061581468373706439;
            6'd50: xpb[0] = 1024'd35656937825106948411594325722112274287958957618191626282748423457902398450994202130438226449701141862990701440214462100093456170446218334962942514110063111178771647930090405425659235466031871650523757574048990098660855215596459865056657057681765252386100541661131003490728837554465570041917543468169198222455;
            6'd51: xpb[0] = 1024'd23963407013196613239946319496073076499248294057981890395590206420562756886283172282045483857229397269306200528273001998637418909771020668206685351890631269308978013431735091800409396256200788511403212964691245915997636234886299385061292341867077612507140562152941917757532761498162018141044025354870022738471;
            6'd52: xpb[0] = 1024'd12269876201286278068298313270033878710537630497772154508431989383223115321572142433652741264757652675621699616331541897181381649095823001450428189671199427439184378933379778175159557046369705372282668355333501733334417254176138905065927626052389972628180582644752832024336685441858466240170507241570847254487;
            6'd53: xpb[0] = 1024'd576345389375942896650307043994680921826966937562418621273772345883473756861112585259998672285908081937198704390081795725344388420625334694171027451767585569390744435024464549909717836538622233162123745975757550671198273465978425070562910237702332749220603136563746291140609385554914339296989128271671770503;
            6'd54: xpb[0] = 1024'd112949510261590349123801228222769915877814730503088366862247410373520727529459221646882327294471837797695847199906115128848370968586648002493073990248666784633287784506240368262290117818224744815351776745005253214372340142976714718040176764106244142137080527042491718588051061403179995455542160841598090770850;
            6'd55: xpb[0] = 1024'd101255979449680013952153221996730718089104066942878630975089193336181085964748191798489584702000093204011346287964655027392333707911450335736816828029234942763494150007885054637040278608393661676231232135647509031709121162266554238044812048291556502258120547534302632854854985346876443554668642728298915286866;
            6'd56: xpb[0] = 1024'd89562448637769678780505215770691520300393403382668895087930976298841444400037161950096842109528348610326845376023194925936296447236252668980559665809803100893700515509529741011790439398562578537110687526289764849045902181556393758049447332476868862379160568026113547121658909290572891653795124614999739802882;
            6'd57: xpb[0] = 1024'd77868917825859343608857209544652322511682739822459159200772759261501802835326132101704099517056604016642344464081734824480259186561055002224302503590371259023906881011174427386540600188731495397990142916932020666382683200846233278054082616662181222500200588517924461388462833234269339752921606501700564318898;
            6'd58: xpb[0] = 1024'd66175387013949008437209203318613124722972076262249423313614542224162161270615102253311356924584859422957843552140274723024221925885857335468045341370939417154113246512819113761290760978900412258869598307574276483719464220136072798058717900847493582621240609009735375655266757177965787852048088388401388834914;
            6'd59: xpb[0] = 1024'd54481856202038673265561197092573926934261412702039687426456325186822519705904072404918614332113114829273342640198814621568184665210659668711788179151507575284319612014463800136040921769069329119749053698216532301056245239425912318063353185032805942742280629501546289922070681121662235951174570275102213350930;
            6'd60: xpb[0] = 1024'd42788325390128338093913190866534729145550749141829951539298108149482878141193042556525871739641370235588841728257354520112147404535462001955531016932075733414525977516108486510791082559238245980628509088858788118393026258715751838067988469218118302863320649993357204188874605065358684050301052161803037866946;
            6'd61: xpb[0] = 1024'd31094794578218002922265184640495531356840085581620215652139891112143236576482012708133129147169625641904340816315894418656110143860264335199273854712643891544732343017753172885541243349407162841507964479501043935729807278005591358072623753403430662984360670485168118455678529009055132149427534048503862382962;
            6'd62: xpb[0] = 1024'd19401263766307667750617178414456333568129422021410479764981674074803595011770982859740386554697881048219839904374434317200072883185066668443016692493212049674938708519397859260291404139576079702387419870143299753066588297295430878077259037588743023105400690976979032722482452952751580248554015935204686898978;
            6'd63: xpb[0] = 1024'd7707732954397332578969172188417135779418758461200743877823457037463953447059953011347643962226136454535338992432974215744035622509869001686759530273780207805145074021042545635041564929744996563266875260785555570403369316585270398081894321774055383226440711468789946989286376896448028347680497821905511414994;
        endcase
    end

    always_comb begin
        case(flag[0][11:6])
            6'd0: xpb[1] = 1024'd0;
            6'd1: xpb[1] = 1024'd120080897826611738806120093367192370735406522026726692118797095065101207219658062072969972584412066170293987487949007548867062202675891669485662493070679406869042114092258449347421964911431119145456528259815051234104511186096006691051508175642597192614300635374717919286196828914073109463925669535231930415341;
            6'd2: xpb[1] = 1024'd116095099969098736213441259329570308726114616927717700109462335065225519102006985235924873954166458031144825568440521663155060564510563004416164861125027772804393553614945681357213690631345032569602858911242862621844661521971116609138037781601964935961781367335318780542287129754217585910732649243838266346351;
            6'd3: xpb[1] = 1024'd112109302111585733620762425291948246716822711828708708100127575065349830984355908398879775323920849891995663648932035777443058926345234339346667229179376138739744993137632913367005416351258945993749189562670674009584811857846226527224567387561332679309262099295919641798377430594362062357539628952444602277361;
            6'd4: xpb[1] = 1024'd108123504254072731028083591254326184707530806729699716090792815065474142866704831561834676693675241752846501729423549891731057288179905674277169597233724504675096432660320145376797142071172859417895520214098485397324962193721336445311096993520700422656742831256520503054467731434506538804346608661050938208371;
            6'd5: xpb[1] = 1024'd104137706396559728435404757216704122698238901630690724081458055065598454749053754724789578063429633613697339809915064006019055650014577009207671965288072870610447872183007377386588867791086772842041850865526296785065112529596446363397626599480068166004223563217121364310558032274651015251153588369657274139381;
            6'd6: xpb[1] = 1024'd100151908539046725842725923179082060688946996531681732072123295065722766631402677887744479433184025474548177890406578120307054011849248344138174333342421236545799311705694609396380593511000686266188181516954108172805262865471556281484156205439435909351704295177722225566648333114795491697960568078263610070391;
            6'd7: xpb[1] = 1024'd96166110681533723250047089141459998679655091432672740062788535065847078513751601050699380802938417335399015970898092234595052373683919679068676701396769602481150751228381841406172319230914599690334512168381919560545413201346666199570685811398803652699185027138323086822738633954939968144767547786869946001401;
            6'd8: xpb[1] = 1024'd92180312824020720657368255103837936670363186333663748053453775065971390396100524213654282172692809196249854051389606348883050735518591013999179069451117968416502190751069073415964044950828513114480842819809730948285563537221776117657215417358171396046665759098923948078828934795084444591574527495476281932411;
            6'd9: xpb[1] = 1024'd88194514966507718064689421066215874661071281234654756044119015066095702278449447376609183542447201057100692131881120463171049097353262348929681437505466334351853630273756305425755770670742426538627173471237542336025713873096886035743745023317539139394146491059524809334919235635228921038381507204082617863421;
            6'd10: xpb[1] = 1024'd84208717108994715472010587028593812651779376135645764034784255066220014160798370539564084912201592917951530212372634577459047459187933683860183805559814700287205069796443537435547496390656339962773504122665353723765864208971995953830274629276906882741627223020125670591009536475373397485188486912688953794431;
            6'd11: xpb[1] = 1024'd80222919251481712879331752990971750642487471036636772025449495066344326043147293702518986281955984778802368292864148691747045821022605018790686173614163066222556509319130769445339222110570253386919834774093165111506014544847105871916804235236274626089107954980726531847099837315517873931995466621295289725441;
            6'd12: xpb[1] = 1024'd76237121393968710286652918953349688633195565937627780016114735066468637925496216865473887651710376639653206373355662806035044182857276353721188541668511432157907948841818001455130947830484166811066165425520976499246164880722215790003333841195642369436588686941327393103190138155662350378802446329901625656451;
            6'd13: xpb[1] = 1024'd72251323536455707693974084915727626623903660838618788006779975066592949807845140028428789021464768500504044453847176920323042544691947688651690909722859798093259388364505233464922673550398080235212496076948787886986315216597325708089863447155010112784069418901928254359280438995806826825609426038507961587461;
            6'd14: xpb[1] = 1024'd68265525678942705101295250878105564614611755739609795997445215066717261690194063191383690391219160361354882534338691034611040906526619023582193277777208164028610827887192465474714399270311993659358826728376599274726465552472435626176393053114377856131550150862529115615370739835951303272416405747114297518471;
            6'd15: xpb[1] = 1024'd64279727821429702508616416840483502605319850640600803988110455066841573572542986354338591760973552222205720614830205148899039268361290358512695645831556529963962267409879697484506124990225907083505157379804410662466615888347545544262922659073745599479030882823129976871461040676095779719223385455720633449481;
            6'd16: xpb[1] = 1024'd60293929963916699915937582802861440596027945541591811978775695066965885454891909517293493130727944083056558695321719263187037630195961693443198013885904895899313706932566929494297850710139820507651488031232222050206766224222655462349452265033113342826511614783730838127551341516240256166030365164326969380491;
            6'd17: xpb[1] = 1024'd56308132106403697323258748765239378586736040442582819969440935067090197337240832680248394500482335943907396775813233377475035992030633028373700381940253261834665146455254161504089576430053733931797818682660033437946916560097765380435981870992481086173992346744331699383641642356384732612837344872933305311501;
            6'd18: xpb[1] = 1024'd52322334248890694730579914727617316577444135343573827960106175067214509219589755843203295870236727804758234856304747491763034353865304363304202749994601627770016585977941393513881302149967647355944149334087844825687066895972875298522511476951848829521473078704932560639731943196529209059644324581539641242511;
            6'd19: xpb[1] = 1024'd48336536391377692137901080689995254568152230244564835950771415067338821101938679006158197239991119665609072936796261606051032715699975698234705118048949993705368025500628625523673027869881560780090479985515656213427217231847985216609041082911216572868953810665533421895822244036673685506451304290145977173521;
            6'd20: xpb[1] = 1024'd44350738533864689545222246652373192558860325145555843941436655067463132984287602169113098609745511526459911017287775720339031077534647033165207486103298359640719465023315857533464753589795474204236810636943467601167367567723095134695570688870584316216434542626134283151912544876818161953258283998752313104531;
            6'd21: xpb[1] = 1024'd40364940676351686952543412614751130549568420046546851932101895067587444866636525332067999979499903387310749097779289834627029439369318368095709854157646725576070904546003089543256479309709387628383141288371278988907517903598205052782100294829952059563915274586735144408002845716962638400065263707358649035541;
            6'd22: xpb[1] = 1024'd36379142818838684359864578577129068540276514947537859922767135067711756748985448495022901349254295248161587178270803948915027801203989703026212222211995091511422344068690321553048205029623301052529471939799090376647668239473314970868629900789319802911396006547336005664093146557107114846872243415964984966551;
            6'd23: xpb[1] = 1024'd32393344961325681767185744539507006530984609848528867913432375067836068631334371657977802719008687109012425258762318063203026163038661037956714590266343457446773783591377553562839930749537214476675802591226901764387818575348424888955159506748687546258876738507936866920183447397251591293679223124571320897561;
            6'd24: xpb[1] = 1024'd28407547103812679174506910501884944521692704749519875904097615067960380513683294820932704088763078969863263339253832177491024524873332372887216958320691823382125223114064785572631656469451127900822133242654713152127968911223534807041689112708055289606357470468537728176273748237396067740486202833177656828571;
            6'd25: xpb[1] = 1024'd24421749246299676581828076464262882512400799650510883894762855068084692396032217983887605458517470830714101419745346291779022886708003707817719326375040189317476662636752017582423382189365041324968463894082524539868119247098644725128218718667423032953838202429138589432364049077540544187293182541783992759581;
            6'd26: xpb[1] = 1024'd20435951388786673989149242426640820503108894551501891885428095068209004278381141146842506828271862691564939500236860406067021248542675042748221694429388555252828102159439249592215107909278954749114794545510335927608269582973754643214748324626790776301318934389739450688454349917685020634100162250390328690591;
            6'd27: xpb[1] = 1024'd16450153531273671396470408389018758493816989452492899876093335068333316160730064309797408198026254552415777580728374520355019610377346377678724062483736921188179541682126481602006833629192868173261125196938147315348419918848864561301277930586158519648799666350340311944544650757829497080907141958996664621601;
            6'd28: xpb[1] = 1024'd12464355673760668803791574351396696484525084353483907866758575068457628043078987472752309567780646413266615661219888634643017972212017712609226430538085287123530981204813713611798559349106781597407455848365958703088570254723974479387807536545526262996280398310941173200634951597973973527714121667603000552611;
            6'd29: xpb[1] = 1024'd8478557816247666211112740313774634475233179254474915857423815068581939925427910635707210937535038274117453741711402748931016334046689047539728798592433653058882420727500945621590285069020695021553786499793770090828720590599084397474337142504894006343761130271542034456725252438118449974521101376209336483621;
            6'd30: xpb[1] = 1024'd4492759958734663618433906276152572465941274155465923848089055068706251807776833798662112307289430134968291822202916863219014695881360382470231166646782018994233860250188177631382010788934608445700117151221581478568870926474194315560866748464261749691241862232142895712815553278262926421328081084815672414631;
            6'd31: xpb[1] = 1024'd506962101221661025755072238530510456649369056456931838754295068830563690125756961617013677043821995819129902694430977507013057716031717400733534701130384929585299772875409641173736508848521869846447802649392866309021262349304233647396354423629493038722594192743756968905854118407402868135060793422008345641;
            6'd32: xpb[1] = 1024'd120587859927833399831875165605722881192055891083183623957551390133931770909783819034586986261455888166113117390643438526374075260391923386886396027771809791798627413865133858988595701420279641015302976062464444100413532448445310924698904530066226685653023229567461676255102683032480512332060730328653938760982;
            6'd33: xpb[1] = 1024'd116602062070320397239196331568100819182763985984174631948216630134056082792132742197541887631210280026963955471134952640662073622226594721816898395826158157733978853387821090998387427140193554439449306713892255488153682784320420842785434136025594429000503961528062537511192983872624988778867710037260274691992;
            6'd34: xpb[1] = 1024'd112616264212807394646517497530478757173472080885165639938881870134180394674481665360496789000964671887814793551626466754950071984061266056747400763880506523669330292910508323008179152860107467863595637365320066875893833120195530760871963741984962172347984693488663398767283284712769465225674689745866610623002;
            6'd35: xpb[1] = 1024'd108630466355294392053838663492856695164180175786156647929547110134304706556830588523451690370719063748665631632117980869238070345895937391677903131934854889604681732433195555017970878580021381287741968016747878263633983456070640678958493347944329915695465425449264260023373585552913941672481669454472946554012;
            6'd36: xpb[1] = 1024'd104644668497781389461159829455234633154888270687147655920212350134429018439179511686406591740473455609516469712609494983526068707730608726608405499989203255540033171955882787027762604299935294711888298668175689651374133791945750597045022953903697659042946157409865121279463886393058418119288649163079282485022;
            6'd37: xpb[1] = 1024'd100658870640268386868480995417612571145596365588138663910877590134553330321528434849361493110227847470367307793101009097814067069565280061538907868043551621475384611478570019037554330019849208136034629319603501039114284127820860515131552559863065402390426889370465982535554187233202894566095628871685618416032;
            6'd38: xpb[1] = 1024'd96673072782755384275802161379990509136304460489129671901542830134677642203877358012316394479982239331218145873592523212102065431399951396469410236097899987410736051001257251047346055739763121560180959971031312426854434463695970433218082165822433145737907621331066843791644488073347371012902608580291954347042;
            6'd39: xpb[1] = 1024'd92687274925242381683123327342368447127012555390120679892208070134801954086226281175271295849736631192068983954084037326390063793234622731399912604152248353346087490523944483057137781459677034984327290622459123814594584799571080351304611771781800889085388353291667705047734788913491847459709588288898290278052;
            6'd40: xpb[1] = 1024'd88701477067729379090444493304746385117720650291111687882873310134926265968575204338226197219491023052919822034575551440678062155069294066330414972206596719281438930046631715066929507179590948408473621273886935202334735135446190269391141377741168632432869085252268566303825089753636323906516567997504626209062;
            6'd41: xpb[1] = 1024'd84715679210216376497765659267124323108428745192102695873538550135050577850924127501181098589245414913770660115067065554966060516903965401260917340260945085216790369569318947076721232899504861832619951925314746590074885471321300187477670983700536375780349817212869427559915390593780800353323547706110962140072;
            6'd42: xpb[1] = 1024'd80729881352703373905086825229502261099136840093093703864203790135174889733273050664135999958999806774621498195558579669254058878738636736191419708315293451152141809092006179086512958619418775256766282576742557977815035807196410105564200589659904119127830549173470288816005691433925276800130527414717298071082;
            6'd43: xpb[1] = 1024'd76744083495190371312407991191880199089844934994084711854869030135299201615621973827090901328754198635472336276050093783542057240573308071121922076369641817087493248614693411096304684339332688680912613228170369365555186143071520023650730195619271862475311281134071150072095992274069753246937507123323634002092;
            6'd44: xpb[1] = 1024'd72758285637677368719729157154258137080553029895075719845534270135423513497970896990045802698508590496323174356541607897830055602407979406052424444423990183022844688137380643106096410059246602105058943879598180753295336478946629941737259801578639605822792013094672011328186293114214229693744486831929969933102;
            6'd45: xpb[1] = 1024'd68772487780164366127050323116636075071261124796066727836199510135547825380319820153000704068262982357174012437033122012118053964242650740982926812478338548958196127660067875115888135779160515529205274531025992141035486814821739859823789407538007349170272745055272872584276593954358706140551466540536305864112;
            6'd46: xpb[1] = 1024'd64786689922651363534371489079014013061969219697057735826864750135672137262668743315955605438017374218024850517524636126406052326077322075913429180532686914893547567182755107125679861499074428953351605182453803528775637150696849777910319013497375092517753477015873733840366894794503182587358446249142641795122;
            6'd47: xpb[1] = 1024'd60800892065138360941692655041391951052677314598048743817529990135796449145017666478910506807771766078875688598016150240694050687911993410843931548587035280828899006705442339135471587218988342377497935833881614916515787486571959695996848619456742835865234208976474595096457195634647659034165425957748977726132;
            6'd48: xpb[1] = 1024'd56815094207625358349013821003769889043385409499039751808195230135920761027366589641865408177526157939726526678507664354982049049746664745774433916641383646764250446228129571145263312938902255801644266485309426304255937822447069614083378225416110579212714940937075456352547496474792135480972405666355313657142;
            6'd49: xpb[1] = 1024'd52829296350112355756334986966147827034093504400030759798860470136045072909715512804820309547280549800577364758999178469270047411581336080704936284695732012699601885750816803155055038658816169225790597136737237691996088158322179532169907831375478322560195672897676317608637797314936611927779385374961649588152;
            6'd50: xpb[1] = 1024'd48843498492599353163656152928525765024801599301021767789525710136169384792064435967775210917034941661428202839490692583558045773416007415635438652750080378634953325273504035164846764378730082649936927788165049079736238494197289450256437437334846065907676404858277178864728098155081088374586365083567985519162;
            6'd51: xpb[1] = 1024'd44857700635086350570977318890903703015509694202012775780190950136293696674413359130730112286789333522279040919982206697846044135250678750565941020804428744570304764796191267174638490098643996074083258439592860467476388830072399368342967043294213809255157136818878040120818398995225564821393344792174321450172;
            6'd52: xpb[1] = 1024'd40871902777573347978298484853281641006217789103003783770856190136418008556762282293685013656543725383129879000473720812134042497085350085496443388858777110505656204318878499184430215818557909498229589091020671855216539165947509286429496649253581552602637868779478901376908699835370041268200324500780657381182;
            6'd53: xpb[1] = 1024'd36886104920060345385619650815659578996925884003994791761521430136542320439111205456639915026298117243980717080965234926422040858920021420426945756913125476441007643841565731194221941538471822922375919742448483242956689501822619204516026255212949295950118600740079762632999000675514517715007304209386993312192;
            6'd54: xpb[1] = 1024'd32900307062547342792940816778037516987633978904985799752186670136666632321460128619594816396052509104831555161456749040710039220754692755357448124967473842376359083364252963204013667258385736346522250393876294630696839837697729122602555861172317039297599332700680623889089301515658994161814283917993329243202;
            6'd55: xpb[1] = 1024'd28914509205034340200261982740415454978342073805976807742851910136790944203809051782549717765806900965682393241948263154998037582589364090287950493021822208311710522886940195213805392978299649770668581045304106018436990173572839040689085467131684782645080064661281485145179602355803470608621263626599665174212;
            6'd56: xpb[1] = 1024'd24928711347521337607583148702793392969050168706967815733517150136915256086157974945504619135561292826533231322439777269286035944424035425218452861076170574247061962409627427223597118698213563194814911696731917406177140509447948958775615073091052525992560796621882346401269903195947947055428243335206001105222;
            6'd57: xpb[1] = 1024'd20942913490008335014904314665171330959758263607958823724182390137039567968506898108459520505315684687384069402931291383574034306258706760148955229130518940182413401932314659233388844418127476618961242348159728793917290845323058876862144679050420269340041528582483207657360204036092423502235223043812337036232;
            6'd58: xpb[1] = 1024'd16957115632495332422225480627549268950466358508949831714847630137163879850855821271414421875070076548234907483422805497862032668093378095079457597184867306117764841455001891243180570138041390043107572999587540181657441181198168794948674285009788012687522260543084068913450504876236899949042202752418672967242;
            6'd59: xpb[1] = 1024'd12971317774982329829546646589927206941174453409940839705512870137288191733204744434369323244824468409085745563914319612150031029928049430009959965239215672053116280977689123252972295857955303467253903651015351569397591517073278713035203890969155756035002992503684930169540805716381376395849182461025008898252;
            6'd60: xpb[1] = 1024'd8985519917469327236867812552305144931882548310931847696178110137412503615553667597324224614578860269936583644405833726438029391762720764940462333293564037988467720500376355262764021577869216891400234302443162957137741852948388631121733496928523499382483724464285791425631106556525852842656162169631344829262;
            6'd61: xpb[1] = 1024'd4999722059956324644188978514683082922590643211922855686843350137536815497902590760279125984333252130787421724897347840726027753597392099870964701347912403923819160023063587272555747297783130315546564953870974344877892188823498549208263102887891242729964456424886652681721407396670329289463141878237680760272;
            6'd62: xpb[1] = 1024'd1013924202443322051510144477061020913298738112913863677508590137661127380251513923234027354087643991638259805388861955014026115432063434801467069402260769859170599545750819282347473017697043739692895605298785732618042524698608467294792708847258986077445188385487513937811708236814805736270121586844016691282;
            6'd63: xpb[1] = 1024'd121094822029055060857630237844253391648705260139640555796305685202762334599909575996203999938499710161932247293337869503881088318107955104287129562472940176728212713638009268629769437929128162885149423865113836966722553710794615158346300884489856178691745823760205433224008537150887915200195791122075947106623;
        endcase
    end

    always_comb begin
        case(flag[0][16:12])
            5'd0: xpb[2] = 1024'd0;
            5'd1: xpb[2] = 1024'd117109024171542058264951403806631329639413355040631563786970925202886646482258499159158901308254102022783085373829383618169086679942626439217631930527288542663564153160696500639561163649042076309295754516541648354462704046669725076432830490449223922039226555720806294480098837991032391647002770830682283037633;
            5'd2: xpb[2] = 1024'd110151352658959375131103880208448226534128282955527443445809995340796397627207859408302731401850529736123021340201273801759109519044032543880103736038246044393437631751821783941492088106566946897281311424696056862561047243118553379900682411215218394811633208027495530930091147908136150276886851834738971590935;
            5'd3: xpb[2] = 1024'd103193681146376691997256356610265123428843210870423323104649065478706148772157219657446561495446957449462957306573163985349132358145438648542575541549203546123311110342947067243423012564091817485266868332850465370659390439567381683368534331981212867584039860334184767380083457825239908906770932838795660144237;
            5'd4: xpb[2] = 1024'd96236009633794008863408833012082020323558138785319202763488135616615899917106579906590391589043385162802893272945054168939155197246844753205047347060161047853184588934072350545353937021616688073252425241004873878757733636016209986836386252747207340356446512640874003830075767742343667536655013842852348697539;
            5'd5: xpb[2] = 1024'd89278338121211325729561309413898917218273066700215082422327205754525651062055940155734221682639812876142829239316944352529178036348250857867519152571118549583058067525197633847284861479141558661237982149159282386856076832465038290304238173513201813128853164947563240280068077659447426166539094846909037250841;
            5'd6: xpb[2] = 1024'd82320666608628642595713785815715814112987994615110962081166275892435402207005300404878051776236240589482765205688834536119200875449656962529990958082076051312931546116322917149215785936666429249223539057313690894954420028913866593772090094279196285901259817254252476730060387576551184796423175850965725804143;
            5'd7: xpb[2] = 1024'd75362995096045959461866262217532711007702922530006841740005346030345153351954660654021881869832668302822701172060724719709223714551063067192462763593033553042805024707448200451146710394191299837209095965468099403052763225362694897239942015045190758673666469560941713180052697493654943426307256855022414357445;
            5'd8: xpb[2] = 1024'd68405323583463276328018738619349607902417850444902721398844416168254904496904020903165711963429096016162637138432614903299246553652469171854934569103991054772678503298573483753077634851716170425194652873622507911151106421811523200707793935811185231446073121867630949630045007410758702056191337859079102910747;
            5'd9: xpb[2] = 1024'd61447652070880593194171215021166504797132778359798601057683486306164655641853381152309542057025523729502573104804505086889269392753875276517406374614948556502551981889698767055008559309241041013180209781776916419249449618260351504175645856577179704218479774174320186080037317327862460686075418863135791464049;
            5'd10: xpb[2] = 1024'd54489980558297910060323691422983401691847706274694480716522556444074406786802741401453372150621951442842509071176395270479292231855281381179878180125906058232425460480824050356939483766765911601165766689931324927347792814709179807643497777343174176990886426481009422530029627244966219315959499867192480017351;
            5'd11: xpb[2] = 1024'd47532309045715226926476167824800298586562634189590360375361626581984157931752101650597202244218379156182445037548285454069315070956687485842349985636863559962298939071949333658870408224290782189151323598085733435446136011158008111111349698109168649763293078787698658980021937162069977945843580871249168570653;
            5'd12: xpb[2] = 1024'd40574637533132543792628644226617195481277562104486240034200696719893909076701461899741032337814806869522381003920175637659337910058093590504821791147821061692172417663074616960801332681815652777136880506240141943544479207606836414579201618875163122535699731094387895430014247079173736575727661875305857123955;
            5'd13: xpb[2] = 1024'd33616966020549860658781120628434092375992490019382119693039766857803660221650822148884862431411234582862316970292065821249360749159499695167293596658778563422045896254199900262732257139340523365122437414394550451642822404055664718047053539641157595308106383401077131880006556996277495205611742879362545677257;
            5'd14: xpb[2] = 1024'd26659294507967177524933597030250989270707417934277999351878836995713411366600182398028692525007662296202252936663956004839383588260905799829765402169736065151919374845325183564663181596865393953107994322548958959741165600504493021514905460407152068080513035707766368329998866913381253835495823883419234230559;
            5'd15: xpb[2] = 1024'd19701622995384494391086073432067886165422345849173879010717907133623162511549542647172522618604090009542188903035846188429406427362311904492237207680693566881792853436450466866594106054390264541093551230703367467839508796953321324982757381173146540852919688014455604779991176830485012465379904887475922783861;
            5'd16: xpb[2] = 1024'd12743951482801811257238549833884783060137273764069758669556977271532913656498902896316352712200517722882124869407736372019429266463718009154709013191651068611666332027575750168525030511915135129079108138857775975937851993402149628450609301939141013625326340321144841229983486747588771095263985891532611337163;
            5'd17: xpb[2] = 1024'd5786279970219128123391026235701679954852201678965638328396047409442664801448263145460182805796945436222060835779626555609452105565124113817180818702608570341539810618701033470455954969440005717064665047012184484036195189850977931918461222705135486397732992627834077679975796664692529725148066895589299890465;
            5'd18: xpb[2] = 1024'd122895304141761186388342430042333009594265556719597202115366972612329311283706762304619084114051047459005146209609010173778538785507750553034812749229897113005103963779397534110017118618482082026360419563553832838498899236520703008351291713154359408436959548348640372160074634655724921372150837726271582928098;
            5'd19: xpb[2] = 1024'd115937632629178503254494906444149906488980484634493081774206042750239062428656122553762914207647475172345082175980900357368561624609156657697284554740854614734977442370522817411948043076006952614345976471708241346597242432969531311819143633920353881209366200655329608610066944572828680002034918730328271481400;
            5'd20: xpb[2] = 1024'd108979961116595820120647382845966803383695412549388961433045112888148813573605482802906744301243902885685018142352790540958584463710562762359756360251812116464850920961648100713878967533531823202331533379862649854695585629418359615286995554686348353981772852962018845060059254489932438631918999734384960034702;
            5'd21: xpb[2] = 1024'd102022289604013136986799859247783700278410340464284841091884183026058564718554843052050574394840330599024954108724680724548607302811968867022228165762769618194724399552773384015809891991056693790317090288017058362793928825867187918754847475452342826754179505268708081510051564407036197261803080738441648588004;
            5'd22: xpb[2] = 1024'd95064618091430453852952335649600597173125268379180720750723253163968315863504203301194404488436758312364890075096570908138630141913374971684699971273727119924597878143898667317740816448581564378302647196171466870892272022316016222222699396218337299526586157575397317960043874324139955891687161742498337141306;
            5'd23: xpb[2] = 1024'd88106946578847770719104812051417494067840196294076600409562323301878067008453563550338234582033186025704826041468461091728652981014781076347171776784684621654471356735023950619671740906106434966288204104325875378990615218764844525690551316984331772298992809882086554410036184241243714521571242746555025694608;
            5'd24: xpb[2] = 1024'd81149275066265087585257288453234390962555124208972480068401393439787818153402923799482064675629613739044762007840351275318675820116187181009643582295642123384344835326149233921602665363631305554273761012480283887088958415213672829158403237750326245071399462188775790860028494158347473151455323750611714247910;
            5'd25: xpb[2] = 1024'd74191603553682404451409764855051287857270052123868359727240463577697569298352284048625894769226041452384697974212241458908698659217593285672115387806599625114218313917274517223533589821156176142259317920634692395187301611662501132626255158516320717843806114495465027310020804075451231781339404754668402801212;
            5'd26: xpb[2] = 1024'd67233932041099721317562241256868184751984980038764239386079533715607320443301644297769724862822469165724633940584131642498721498318999390334587193317557126844091792508399800525464514278681046730244874828789100903285644808111329436094107079282315190616212766802154263760013113992554990411223485758725091354514;
            5'd27: xpb[2] = 1024'd60276260528517038183714717658685081646699907953660119044918603853517071588251004546913554956418896879064569906956021826088744337420405494997058998828514628573965271099525083827395438736205917318230431736943509411383988004560157739561959000048309663388619419108843500210005423909658749041107566762781779907816;
            5'd28: xpb[2] = 1024'd53318589015934355049867194060501978541414835868555998703757673991426822733200364796057385050015324592404505873327912009678767176521811599659530804339472130303838749690650367129326363193730787906215988645097917919482331201008986043029810920814304136161026071415532736659997733826762507670991647766838468461118;
            5'd29: xpb[2] = 1024'd46360917503351671916019670462318875436129763783451878362596744129336573878149725045201215143611752305744441839699802193268790015623217704322002609850429632033712228281775650431257287651255658494201545553252326427580674397457814346497662841580298608933432723722221973109990043743866266300875728770895157014420;
            5'd30: xpb[2] = 1024'd39403245990768988782172146864135772330844691698347758021435814267246325023099085294345045237208180019084377806071692376858812854724623808984474415361387133763585706872900933733188212108780529082187102461406734935679017593906642649965514762346293081705839376028911209559982353660970024930759809774951845567722;
            5'd31: xpb[2] = 1024'd32445574478186305648324623265952669225559619613243637680274884405156076168048445543488875330804607732424313772443582560448835693826029913646946220872344635493459185464026217035119136566305399670172659369561143443777360790355470953433366683112287554478246028335600446009974663578073783560643890779008534121024;
        endcase
    end

    always_comb begin
        case(flag[1][5:0])
            6'd0: xpb[3] = 1024'd0;
            6'd1: xpb[3] = 1024'd12743951482801811257238549833884783060137273764069758669556977271532913656498902896316352712200517722882124869407736372019429266463718009154709013191651068611666332027575750168525030511915135129079108138857775975937851993402149628450609301939141013625326340321144841229983486747588771095263985891532611337163;
            6'd2: xpb[3] = 1024'd25487902965603622514477099667769566120274547528139517339113954543065827312997805792632705424401035445764249738815472744038858532927436018309418026383302137223332664055151500337050061023830270258158216277715551951875703986804299256901218603878282027250652680642289682459966973495177542190527971783065222674326;
            6'd3: xpb[3] = 1024'd38231854448405433771715649501654349180411821292209276008670931814598740969496708688949058136601553168646374608223209116058287799391154027464127039574953205834998996082727250505575091535745405387237324416573327927813555980206448885351827905817423040875979020963434523689950460242766313285791957674597834011489;
            6'd4: xpb[3] = 1024'd50975805931207245028954199335539132240549095056279034678227909086131654625995611585265410848802070891528499477630945488077717065854872036618836052766604274446665328110303000674100122047660540516316432555431103903751407973608598513802437207756564054501305361284579364919933946990355084381055943566130445348652;
            6'd5: xpb[3] = 1024'd63719757414009056286192749169423915300686368820348793347784886357664568282494514481581763561002588614410624347038681860097146332318590045773545065958255343058331660137878750842625152559575675645395540694288879879689259967010748142253046509695705068126631701605724206149917433737943855476319929457663056685815;
            6'd6: xpb[3] = 1024'd76463708896810867543431299003308698360823642584418552017341863629197481938993417377898116273203106337292749216446418232116575598782308054928254079149906411669997992165454501011150183071490810774474648833146655855627111960412897770703655811634846081751958041926869047379900920485532626571583915349195668022978;
            6'd7: xpb[3] = 1024'd89207660379612678800669848837193481420960916348488310686898840900730395595492320274214468985403624060174874085854154604136004865246026064082963092341557480281664324193030251179675213583405945903553756972004431831564963953815047399154265113573987095377284382248013888609884407233121397666847901240728279360141;
            6'd8: xpb[3] = 1024'd101951611862414490057908398671078264481098190112558069356455818172263309251991223170530821697604141783056998955261890976155434131709744073237672105533208548893330656220606001348200244095321081032632865110862207807502815947217197027604874415513128109002610722569158729839867893980710168762111887132260890697304;
            6'd9: xpb[3] = 1024'd114695563345216301315146948504963047541235463876627828026012795443796222908490126066847174409804659505939123824669627348174863398173462082392381118724859617504996988248181751516725274607236216161711973249719983783440667940619346656055483717452269122627937062890303571069851380728298939857375873023793502034467;
            6'd10: xpb[3] = 1024'd3372819143893371173586570934033397856674310514961902567437917650352241227679890053148455907347502919378099286619870285615228823795959756991930006900179645182972645706186284347620065927634145569480883780190519913014159083800599511541114449708180686986443499797331354269728339401959077935521169088700518887299;
            6'd11: xpb[3] = 1024'd16116770626695182430825120767918180916811584279031661236994894921885154884178792949464808619548020642260224156027606657634658090259677766146639020091830713794638977733762034516145096439549280698559991919048295888952011077202749139991723751647321700611769840118476195499711826149547849030785154980233130224462;
            6'd12: xpb[3] = 1024'd28860722109496993688063670601802963976948858043101419906551872193418068540677695845781161331748538365142349025435343029654087356723395775301348033283481782406305309761337784684670126951464415827639100057906071864889863070604898768442333053586462714237096180439621036729695312897136620126049140871765741561625;
            6'd13: xpb[3] = 1024'd41604673592298804945302220435687747037086131807171178576108849464950982197176598742097514043949056088024473894843079401673516623187113784456057046475132851017971641788913534853195157463379550956718208196763847840827715064007048396892942355525603727862422520760765877959678799644725391221313126763298352898788;
            6'd14: xpb[3] = 1024'd54348625075100616202540770269572530097223405571240937245665826736483895853675501638413866756149573810906598764250815773692945889650831793610766059666783919629637973816489285021720187975294686085797316335621623816765567057409198025343551657464744741487748861081910719189662286392314162316577112654830964235951;
            6'd15: xpb[3] = 1024'd67092576557902427459779320103457313157360679335310695915222804008016809510174404534730219468350091533788723633658552145712375156114549802765475072858434988241304305844065035190245218487209821214876424474479399792703419050811347653794160959403885755113075201403055560419645773139902933411841098546363575573114;
            6'd16: xpb[3] = 1024'd79836528040704238717017869937342096217497953099380454584779781279549723166673307431046572180550609256670848503066288517731804422578267811920184086050086056852970637871640785358770248999124956343955532613337175768641271044213497282244770261343026768738401541724200401649629259887491704507105084437896186910277;
            6'd17: xpb[3] = 1024'd92580479523506049974256419771226879277635226863450213254336758551082636823172210327362924892751126979552973372474024889751233689041985821074893099241737125464636969899216535527295279511040091473034640752194951744579123037615646910695379563282167782363727882045345242879612746635080475602369070329428798247440;
            6'd18: xpb[3] = 1024'd105324431006307861231494969605111662337772500627519971923893735822615550479671113223679277604951644702435098241881761261770662955505703830229602112433388194076303301926792285695820310022955226602113748891052727720516975031017796539145988865221308795989054222366490084109596233382669246697633056220961409584603;
            6'd19: xpb[3] = 1024'd118068382489109672488733519438996445397909774391589730593450713094148464136170016119995630317152162425317223111289497633790092221969421839384311125625039262687969633954368035864345340534870361731192857029910503696454827024419946167596598167160449809614380562687634925339579720130258017792897042112494020921766;
            6'd20: xpb[3] = 1024'd6745638287786742347173141868066795713348621029923805134875835300704482455359780106296911814695005838756198573239740571230457647591919513983860013800359290365945291412372568695240131855268291138961767560381039826028318167601199023082228899416361373972886999594662708539456678803918155871042338177401037774598;
            6'd21: xpb[3] = 1024'd19489589770588553604411691701951578773485894793993563804432812572237396111858683002613264526895523561638323442647476943249886914055637523138569026992010358977611623439948318863765162367183426268040875699238815801966170161003348651532838201355502387598213339915807549769440165551506926966306324068933649111761;
            6'd22: xpb[3] = 1024'd32233541253390364861650241535836361833623168558063322473989789843770309768357585898929617239096041284520448312055213315269316180519355532293278040183661427589277955467524069032290192879098561397119983838096591777904022154405498279983447503294643401223539680236952390999423652299095698061570309960466260448924;
            6'd23: xpb[3] = 1024'd44977492736192176118888791369721144893760442322133081143546767115303223424856488795245969951296559007402573181462949687288745446983073541447987053375312496200944287495099819200815223391013696526199091976954367753841874147807647908434056805233784414848866020558097232229407139046684469156834295851998871786087;
            6'd24: xpb[3] = 1024'd57721444218993987376127341203605927953897716086202839813103744386836137081355391691562322663497076730284698050870686059308174713446791550602696066566963564812610619522675569369340253902928831655278200115812143729779726141209797536884666107172925428474192360879242073459390625794273240252098281743531483123250;
            6'd25: xpb[3] = 1024'd70465395701795798633365891037490711014034989850272598482660721658369050737854294587878675375697594453166822920278422431327603979910509559757405079758614633424276951550251319537865284414843966784357308254669919705717578134611947165335275409112066442099518701200386914689374112541862011347362267635064094460413;
            6'd26: xpb[3] = 1024'd83209347184597609890604440871375494074172263614342357152217698929901964394353197484195028087898112176048947789686158803347033246374227568912114092950265702035943283577827069706390314926759101913436416393527695681655430128014096793785884711051207455724845041521531755919357599289450782442626253526596705797576;
            6'd27: xpb[3] = 1024'd95953298667399421147842990705260277134309537378412115821774676201434878050852100380511380800098629898931072659093895175366462512837945578066823106141916770647609615605402819874915345438674237042515524532385471657593282121416246422236494012990348469350171381842676597149341086037039553537890239418129317134739;
            6'd28: xpb[3] = 1024'd108697250150201232405081540539145060194446811142481874491331653472967791707351003276827733512299147621813197528501631547385891779301663587221532119333567839259275947632978570043440375950589372171594632671243247633531134114818396050687103314929489482975497722163821438379324572784628324633154225309661928471902;
            6'd29: xpb[3] = 1024'd121441201633003043662320090373029843254584084906551633160888630744500705363849906173144086224499665344695322397909367919405321045765381596376241132525218907870942279660554320211965406462504507300673740810101023609468986108220545679137712616868630496600824062484966279609308059532217095728418211201194539809065;
            6'd30: xpb[3] = 1024'd10118457431680113520759712802100193570022931544885707702313752951056723683039670159445367722042508758134297859859610856845686471387879270975790020700538935548917937118558853042860197782902436708442651340571559739042477251401798534623343349124542060959330499391994062809185018205877233806563507266101556661897;
            6'd31: xpb[3] = 1024'd22862408914481924777998262635984976630160205308955466371870730222589637339538573055761720434243026481016422729267347228865115737851597280130499033892190004160584269146134603211385228294817571837521759479429335714980329244803948163073952651063683074584656839713138904039168504953466004901827493157634167999060;
            6'd32: xpb[3] = 1024'd35606360397283736035236812469869759690297479073025225041427707494122550996037475952078073146443544203898547598675083600884545004315315289285208047083841072772250601173710353379910258806732706966600867618287111690918181238206097791524561953002824088209983180034283745269151991701054775997091479049166779336223;
            6'd33: xpb[3] = 1024'd48350311880085547292475362303754542750434752837094983710984684765655464652536378848394425858644061926780672468082819972903974270779033298439917060275492141383916933201286103548435289318647842095679975757144887666856033231608247419975171254941965101835309520355428586499135478448643547092355464940699390673386;
            6'd34: xpb[3] = 1024'd61094263362887358549713912137639325810572026601164742380541662037188378309035281744710778570844579649662797337490556344923403537242751307594626073467143209995583265228861853716960319830562977224759083896002663642793885225010397048425780556881106115460635860676573427729118965196232318187619450832232002010549;
            6'd35: xpb[3] = 1024'd73838214845689169806952461971524108870709300365234501050098639308721291965534184641027131283045097372544922206898292716942832803706469316749335086658794278607249597256437603885485350342478112353838192034860439618731737218412546676876389858820247129085962200997718268959102451943821089282883436723764613347712;
            6'd36: xpb[3] = 1024'd86582166328490981064191011805408891930846574129304259719655616580254205622033087537343483995245615095427047076306029088962262070170187325904044099850445347218915929284013354054010380854393247482917300173718215594669589211814696305326999160759388142711288541318863110189085938691409860378147422615297224684875;
            6'd37: xpb[3] = 1024'd99326117811292792321429561639293674990983847893374018389212593851787119278531990433659836707446132818309171945713765460981691336633905335058753113042096415830582261311589104222535411366308382611996408312575991570607441205216845933777608462698529156336614881640007951419069425438998631473411408506829836022038;
            6'd38: xpb[3] = 1024'd112070069294094603578668111473178458051121121657443777058769571123320032935030893329976189419646650541191296815121501833001120603097623344213462126233747484442248593339164854391060441878223517741075516451433767546545293198618995562228217764637670169961941221961152792649052912186587402568675394398362447359201;
            6'd39: xpb[3] = 1024'd747325092771673437107733902248808366559968295777851600194693329876051254220657316277470917189493954630272277071744770441486028720121018813011014409067512120224250797169387221955233198621447148844426981904303676118784341800248417713848496893581734320447658868180575848929870860247540646820690463269464212033;
            6'd40: xpb[3] = 1024'd13491276575573484694346283736133591426697242059847610269751670601408964910719560212593823629390011677512397146479481142460915295183839027967720027600718580731890582824745137390480263710536582277923535120762079652056636335202398046164457798832722747945773999189325417078913357607836311742084676354802075549196;
            6'd41: xpb[3] = 1024'd26235228058375295951584833570018374486834515823917368939308647872941878567218463108910176341590529400394522015887217514480344561647557037122429040792369649343556914852320887559005294222451717407002643259619855627994488328604547674615067100771863761571100339510470258308896844355425082837348662246334686886359;
            6'd42: xpb[3] = 1024'd38979179541177107208823383403903157546971789587987127608865625144474792223717366005226529053791047123276646885294953886499773828111275046277138053984020717955223246879896637727530324734366852536081751398477631603932340322006697303065676402711004775196426679831615099538880331103013853932612648137867298223522;
            6'd43: xpb[3] = 1024'd51723131023978918466061933237787940607109063352056886278422602416007705880216268901542881765991564846158771754702690258519203094574993055431847067175671786566889578907472387896055355246281987665160859537335407579870192315408846931516285704650145788821753020152759940768863817850602625027876634029399909560685;
            6'd44: xpb[3] = 1024'd64467082506780729723300483071672723667246337116126644947979579687540619536715171797859234478192082569040896624110426630538632361038711064586556080367322855178555910935048138064580385758197122794239967676193183555808044308810996559966895006589286802447079360473904781998847304598191396123140619920932520897848;
            6'd45: xpb[3] = 1024'd77211033989582540980539032905557506727383610880196403617536556959073533193214074694175587190392600291923021493518163002558061627502429073741265093558973923790222242962623888233105416270112257923319075815050959531745896302213146188417504308528427816072405700795049623228830791345780167218404605812465132235011;
            6'd46: xpb[3] = 1024'd89954985472384352237777582739442289787520884644266162287093534230606446849712977590491939902593118014805146362925899374577490893966147082895974106750624992401888574990199638401630446782027393052398183953908735507683748295615295816868113610467568829697732041116194464458814278093368938313668591703997743572174;
            6'd47: xpb[3] = 1024'd102698936955186163495016132573327072847658158408335920956650511502139360506211880486808292614793635737687271232333635746596920160429865092050683119942276061013554907017775388570155477293942528181477292092766511483621600289017445445318722912406709843323058381437339305688797764840957709408932577595530354909337;
            6'd48: xpb[3] = 1024'd115442888437987974752254682407211855907795432172405679626207488773672274162710783383124645326994153460569396101741372118616349426893583101205392133133927129625221239045351138738680507805857663310556400231624287459559452282419595073769332214345850856948384721758484146918781251588546480504196563487062966246500;
            6'd49: xpb[3] = 1024'd4120144236665044610694304836282206223234278810739754167632610980228292481900547369425926824536996874008371563691615056056714852516080775804941021309247157303196896503355671569575299126255592718325310762094823589132943425600847929254962946601762421306891158665511930118658210262206618582341859551969983099332;
            6'd50: xpb[3] = 1024'd16864095719466855867932854670166989283371552574809512837189588251761206138399450265742279536737514596890496433099351428076144118979798784959650034500898225914863228530931421738100329638170727847404418900952599565070795419002997557705572248540903434932217498986656771348641697009795389677605845443502594436495;
            6'd51: xpb[3] = 1024'd29608047202268667125171404504051772343508826338879271506746565523294119794898353162058632248938032319772621302507087800095573385443516794114359047692549294526529560558507171906625360150085862976483527039810375541008647412405147186156181550480044448557543839307801612578625183757384160772869831335035205773658;
            6'd52: xpb[3] = 1024'd42351998685070478382409954337936555403646100102949030176303542794827033451397256058374984961138550042654746171914824172115002651907234803269068060884200363138195892586082922075150390662000998105562635178668151516946499405807296814606790852419185462182870179628946453808608670504972931868133817226567817110821;
            6'd53: xpb[3] = 1024'd55095950167872289639648504171821338463783373867018788845860520066359947107896158954691337673339067765536871041322560544134431918370952812423777074075851431749862224613658672243675421173916133234641743317525927492884351399209446443057400154358326475808196519950091295038592157252561702963397803118100428447984;
            6'd54: xpb[3] = 1024'd67839901650674100896887054005706121523920647631088547515417497337892860764395061851007690385539585488418995910730296916153861184834670821578486087267502500361528556641234422412200451685831268363720851456383703468822203392611596071508009456297467489433522860271236136268575644000150474058661789009633039785147;
            6'd55: xpb[3] = 1024'd80583853133475912154125603839590904584057921395158306184974474609425774420893964747324043097740103211301120780138033288173290451298388830733195100459153568973194888668810172580725482197746403492799959595241479444760055386013745699958618758236608503058849200592380977498559130747739245153925774901165651122310;
            6'd56: xpb[3] = 1024'd93327804616277723411364153673475687644195195159228064854531451880958688077392867643640395809940620934183245649545769660192719717762106839887904113650804637584861220696385922749250512709661538621879067734099255420697907379415895328409228060175749516684175540913525818728542617495328016249189760792698262459473;
            6'd57: xpb[3] = 1024'd106071756099079534668602703507360470704332468923297823524088429152491601733891770539956748522141138657065370518953506032212148984225824849042613126842455706196527552723961672917775543221576673750958175872957031396635759372818044956859837362114890530309501881234670659958526104242916787344453746684230873796636;
            6'd58: xpb[3] = 1024'd118815707581881345925841253341245253764469742687367582193645406424024515390390673436273101234341656379947495388361242404231578250689542858197322140034106774808193884751537423086300573733491808880037284011814807372573611366220194585310446664054031543934828221555815501188509590990505558439717732575763485133799;
            6'd59: xpb[3] = 1024'd7492963380558415784280875770315604079908589325701656735070528630580533709580437422574382731884499793386470850311485341671943676312040532796871028209426802486169542209541955917195365053889738287806194542285343502147102509401447440796077396309943108293334658462843284388386549664165696517863028640670501986631;
            6'd60: xpb[3] = 1024'd20236914863360227041519425604200387140045863089771415404627505902113447366079340318890735444085017516268595719719221713691372942775758541951580041401077871097835874237117706085720395565804873416885302681143119478084954502803597069246686698249084121918660998783988125618370036411754467613127014532203113323794;
            6'd61: xpb[3] = 1024'd32980866346162038298757975438085170200183136853841174074184483173646361022578243215207088156285535239150720589126958085710802209239476551106289054592728939709502206264693456254245426077720008545964410820000895454022806496205746697697296000188225135543987339105132966848353523159343238708391000423735724660957;
            6'd62: xpb[3] = 1024'd45724817828963849555996525271969953260320410617910932743741460445179274679077146111523440868486052962032845458534694457730231475703194560260998067784380008321168538292269206422770456589635143675043518958858671429960658489607896326147905302127366149169313679426277808078337009906932009803654986315268335998120;
            6'd63: xpb[3] = 1024'd58468769311765660813235075105854736320457684381980691413298437716712188335576049007839793580686570684914970327942430829749660742166912569415707080976031076932834870319844956591295487101550278804122627097716447405898510483010045954598514604066507162794640019747422649308320496654520780898918972206800947335283;
        endcase
    end

    always_comb begin
        case(flag[1][11:6])
            6'd0: xpb[4] = 1024'd0;
            6'd1: xpb[4] = 1024'd71212720794567472070473624939739519380594958146050450082855414988245101992074951904156146292887088407797095197350167201769090008630630578570416094167682145544501202347420706759820517613465413933201735236574223381836362476412195583049123906005648176419966360068567490538303983402109551994182958098333558672446;
            6'd2: xpb[4] = 1024'd18358745905010202742148322474664606016491489166365216037578974911513308646840764898297221371116502506151040987242840968959116176420040822585672063319033250155311730125270196182010796035413622145093272864761206917308364102603494393133269242328066903573112816723017923046501438730290470971247226370041522860561;
            6'd3: xpb[4] = 1024'd89571466699577674812621947414404125397086447312415666120434389899758410638915716802453367664003590913948136184593008170728206185050671401156088157486715395699812932472690902941831313648879036078295008101335430299144726579015689976182393148333715079993079176791585413584805422132400022965430184468375081533007;
            6'd4: xpb[4] = 1024'd36717491810020405484296644949329212032982978332730432075157949823026617293681529796594442742233005012302081974485681937918232352840081645171344126638066500310623460250540392364021592070827244290186545729522413834616728205206988786266538484656133807146225633446035846093002877460580941942494452740083045721122;
            6'd5: xpb[4] = 1024'd107930212604587877554770269889068731413577936478780882158013364811271719285756481700750589035120093420099177171835849139687322361470712223741760220805748645855124662597961099123842109684292658223388280966096637216453090681619184369315662390661781983566191993514603336631306860862690493936677410838416604393568;
            6'd6: xpb[4] = 1024'd55076237715030608226444967423993818049474467499095648112736924734539925940522294694891664113349507518453122961728522906877348529260122467757016189957099750465935190375810588546032388106240866435279818594283620751925092307810483179399807726984200710719338450169053769139504316190871412913741679110124568581683;
            6'd7: xpb[4] = 1024'd2222262825473338898119664958918904685370998519410414067460484657808132595288107689032739191578921616807068751621196674067374697049532711772272159108450855076745718153660077968222666528189074647171356222470604287397093934001781989483953063306619437872484906823504201647701771519052331890805947381832532769798;
            6'd8: xpb[4] = 1024'd73434983620040810968593289898658424065965956665460864150315899646053234587363059593188885484466010024604163948971363875836464705680163290342688253276133000621246920501080784728043184141654488580373091459044827669233456410413977572533076969312267614292451266892071692186005754921161883884988905480166091442244;
            6'd9: xpb[4] = 1024'd20581008730483541640267987433583510701862487685775630105039459569321441242128872587329960562695424122958109738864037643026490873469573534357944222427484105232057448278930274150233462563602696792264629087231811204705458036605276382617222305634686341445597723546522124694203210249342802862053173751874055630359;
            6'd10: xpb[4] = 1024'd91793729525051013710741612373323030082457445831826080187894874557566543234203824491486106855582512530755204936214204844795580882100204112928360316595166250776558650626350980910053980177068110725466364323806034586541820513017471965666346211640334517865564083615089615232507193651452354856236131850207614302805;
            6'd11: xpb[4] = 1024'd38939754635493744382416309908248116718353976852140846142618434480834749888969637485627181933811926629109150726106878611985607049889614356943616285746517355387369178404200470332244258599016318937357901951993018122013822139208770775750491547962753245018710540269540047740704648979633273833300400121915578490920;
            6'd12: xpb[4] = 1024'd110152475430061216452889934847987636098948934998191296225473849469079851881044589389783328226699015036906245923457045813754697058520244935514032379914199500931870380751621177092064776212481732870559637188567241503850184615620966358799615453968401421438676900338107538279008632381742825827483358220249137163366;
            6'd13: xpb[4] = 1024'd57298500540503947124564632382912722734845466018506062180197409392348058535810402383924403304928429135260191713349719580944723226309655179529288349065550605542680908529470666514255054634429941082451174816754225039322186241812265168883760790290820148591823356992557970787206087709923744804547626491957101351481;
            6'd14: xpb[4] = 1024'd4444525650946677796239329917837809370741997038820828134920969315616265190576215378065478383157843233614137503242393348134749394099065423544544318216901710153491436307320155936445333056378149294342712444941208574794187868003563978967906126613238875744969813647008403295403543038104663781611894763665065539596;
            6'd15: xpb[4] = 1024'd75657246445514149866712954857577328751336955184871278217776384303861367182651167282221624676044931641411232700592560549903839402729696002114960412384583855697992638654740862696265850669843563227544447681515431956630550344415759562017030032618887052164936173715575893833707526440214215775794852861998624212042;
            6'd16: xpb[4] = 1024'd22803271555956880538387652392502415387233486205186044172499944227129573837416980276362699754274345739765178490485234317093865570519106246130216381535934960308803166432590352118456129091791771439435985309702415492102551970607058372101175368941305779318082630370026326341904981768395134752859121133706588400157;
            6'd17: xpb[4] = 1024'd94015992350524352608861277332241934767828444351236494255355359215374675829491932180518846047161434147562273687835401518862955579149736824700632475703617105853304368780011058878276646705257185372637720546276638873938914447019253955150299274946953955738048990438593816880208965170504686747042079232040147072603;
            6'd18: xpb[4] = 1024'd41162017460967083280535974867167021403724975371551260210078919138642882484257745174659921125390848245916219477728075286052981746939147068715888444854968210464114896557860548300466925127205393584529258174463622409410916073210552765234444611269372682891195447093044249388406420498685605724106347503748111260718;
            6'd19: xpb[4] = 1024'd112374738255534555351009599806906540784319933517601710292934334126887984476332697078816067418277936653713314675078242487822071755569777647286304539022650356008616098905281255060287442740670807517730993411037845791247278549622748348283568517275020859311161807161611739926710403900795157718289305602081669933164;
            6'd20: xpb[4] = 1024'd59520763365977286022684297341831627420216464537916476247657894050156191131098510072957142496507350752067260464970916255012097923359187891301560508174001460619426626683130744482477721162619015729622531039224829326719280175814047158367713853597439586464308263816062172434907859228976076695353573873789634121279;
            6'd21: xpb[4] = 1024'd6666788476420016694358994876756714056112995558231242202381453973424397785864323067098217574736764850421206254863590022202124091148598135316816477325352565230237154460980233904667999584567223941514068667411812862191281802005345968451859189919858313617454720470512604943105314557156995672417842145497598309394;
            6'd22: xpb[4] = 1024'd77879509270987488764832619816496233436707953704281692285236868961669499777939274971254363867623853258218301452213757223971214099779228713887232571493034710774738356808400940664488517198032637874715803903986036244027644278417541551500983095925506490037421080539080095481409297959266547666600800243831156981840;
            6'd23: xpb[4] = 1024'd25025534381430219436507317351421320072604484724596458239960428884937706432705087965395438945853267356572247242106430991161240267568638957902488540644385815385548884586250430086678795619980846086607341532173019779499645904608840361585128432247925217190567537193530527989606753287447466643665068515539121169955;
            6'd24: xpb[4] = 1024'd96238255175997691506980942291160839453199442870646908322815843873182808424780039869551585238740355764369342439456598192930330276199269536472904634812067960930050086933671136846499313233446260019809076768747243161336008381021035944634252338253573393610533897262098018527910736689557018637848026613872679842401;
            6'd25: xpb[4] = 1024'd43384280286440422178655639826085926089095973890961674277539403796451015079545852863692660316969769862723288229349271960120356443988679780488160603963419065540860614711520626268689591655394468231700614396934226696808010007212334754718397674575992120763680353916548451036108192017737937614912294885580644030516;
            6'd26: xpb[4] = 1024'd114597001081007894249129264765825445469690932037012124360394818784696117071620804767848806609856858270520383426699439161889446452619310359058576698131101211085361817058941333028510109268859882164902349633508450078644372483624530337767521580581640297183646713985115941574412175419847489609095252983914202702962;
            6'd27: xpb[4] = 1024'd61743026191450624920803962300750532105587463057326890315118378707964323726386617761989881688086272368874329216592112929079472620408720603073832667282452315696172344836790822450700387690808090376793887261695433614116374109815829147851666916904059024336793170639566374082609630748028408586159521255622166891077;
            6'd28: xpb[4] = 1024'd8889051301893355592478659835675618741483994077641656269841938631232530381152430756130956766315686467228275006484786696269498788198130847089088636433803420306982872614640311872890666112756298588685424889882417149588375736007127957935812253226477751489939627294016806590807086076209327563223789527330131079192;
            6'd29: xpb[4] = 1024'd80101772096460827662952284775415138122078952223692106352697353619477632373227382660287103059202774875025370203834953898038588796828761425659504730601485565851484074962061018632711183726221712521887160126456640531424738212419323540984936159232125927909905987362584297129111069478318879557406747625663689751638;
            6'd30: xpb[4] = 1024'd27247797206903558334626982310340224757975483244006872307420913542745839027993195654428178137432188973379315993727627665228614964618171669674760699752836670462294602739910508054901462148169920733778697754643624066896739838610622351069081495554544655063052444017034729637308524806499798534471015897371653939753;
            6'd31: xpb[4] = 1024'd98460518001471030405100607250079744138570441390057322390276328530990941020068147558584324430319277381176411191077794866997704973248802248245176793920518816006795805087331214814721979761635334666980432991217847448733102315022817934118205401560192831483018804085602220175612508208609350528653973995705212612199;
            6'd32: xpb[4] = 1024'd45606543111913761076775304785004830774466972410372088344999888454259147674833960552725399508548691479530356980970468634187731141038212492260432763071869920617606332865180704236912258183583542878871970619404830984205103941214116744202350737882611558636165260740052652683809963536790269505718242267413176800314;
            6'd33: xpb[4] = 1024'd116819263906481233147248929724744350155061930556422538427855303442504249666908912456881545801435779887327452178320635835956821149668843070830848857239552066162107535212601410996732775797048956812073705855979054366041466417626312327251474643888259735056131620808620143222113946938899821499901200365746735472760;
            6'd34: xpb[4] = 1024'd63965289016923963818923627259669436790958461576737304382578863365772456321674725451022620879665193985681397968213309603146847317458253314846104826390903170772918062990450900418923054218997165023965243484166037901513468043817611137335619980210678462209278077463070575730311402267080740476965468637454699660875;
            6'd35: xpb[4] = 1024'd11111314127366694490598324794594523426854992597052070337302423289040662976440538445163695957894608084035343758105983370336873485247663558861360795542254275383728590768300389841113332640945373235856781112353021436985469670008909947419765316533097189362424534117521008238508857595261659454029736909162663848990;
            6'd36: xpb[4] = 1024'd82324034921934166561071949734334042807449950743102520420157838277285764968515490349319842250781696491832438955456150572105963493878294137431776889709936420928229793115721096600933850254410787169058516348927244818821832146421105530468889222538745365782390894186088498776812840997371211448212695007496222521436;
            6'd37: xpb[4] = 1024'd29470060032376897232746647269259129443346481763417286374881398200553971623281303343460917329011110590186384745348824339295989661667704381447032858861287525539040320893570586023124128676358995380950053977114228354293833772612404340553034558861164092935537350840538931285010296325552130425276963279204186709551;
            6'd38: xpb[4] = 1024'd100682780826944369303220272208998648823941439909467736457736813188799073615356255247617063621898198997983479942698991541065079670298334960017448953028969671083541523240991292782944646289824409314151789213688451736130196249024599923602158464866812269355503710909106421823314279727661682419459921377537745381997;
            6'd39: xpb[4] = 1024'd47828805937387099974894969743923735459837970929782502412460373112067280270122068241758138700127613096337425732591665308255105838087745204032704922180320775694352051018840782205134924711772617526043326841875435271602197875215898733686303801189230996508650167563556854331511735055842601396524189649245709570112;
            6'd40: xpb[4] = 1024'd119041526731954572045368594683663254840432929075832952495315788100312382262197020145914284993014701504134520929941832510024195846718375782603121016348002921238853253366261488964955442325238031459245062078449658653438560351628094316735427707194879172928616527632124344869815718457952153390707147747579268242558;
            6'd41: xpb[4] = 1024'd66187551842397302717043292218588341476329460096147718450039348023580588916962833140055360071244115602488466719834506277214222014507786026618376985499354025849663781144110978387145720747186239671136599706636642188910561977819393126819573043517297900081762984286574777378013173786133072367771416019287232430673;
            6'd42: xpb[4] = 1024'd13333576952840033388717989753513428112225991116462484404762907946848795571728646134196435149473529700842412509727180044404248182297196270633632954650705130460474308921960467809335999169134447883028137334823625724382563604010691936903718379839716627234909440941025209886210629114313991344835684290995196618788;
            6'd43: xpb[4] = 1024'd84546297747407505459191614693252947492820949262512934487618322935093897563803598038352581442360618108639507707077347246173338190927826849204049048818387276004975511269381174569156516782599861816229872571397849106218926080422887519952842285845364803654875801009592700424514612516423543339018642389328755291234;
            6'd44: xpb[4] = 1024'd31692322857850236130866312228178034128717480282827700442341882858362104218569411032493656520590032206993453496970021013363364358717237093219305017969738380615786039047230663991346795204548070028121410199584832641690927706614186330036987622167783530808022257664043132932712067844604462316082910661036719479349;
            6'd45: xpb[4] = 1024'd102905043652417708201339937167917553509312438428878150525197297846607206210644362936649802813477120614790548694320188215132454367347867671789721112137420526160287241394651370751167312818013483961323145436159056023527290183026381913086111528173431707227988617732610623471016051246714014310265868759370278151795;
            6'd46: xpb[4] = 1024'd50051068762860438873014634702842640145208969449192916479920857769875412865410175930790877891706534713144494484212861982322480535137277915804977081288771630771097769172500860173357591239961692173214683064346039558999291809217680723170256864495850434381135074387061055979213506574894933287330137031078242339910;
            6'd47: xpb[4] = 1024'd121263789557427910943488259642582159525803927595243366562776272758120514857485127834947024184593623120941589681563029184091570543767908494375393175456453776315598971519921566933178108853427106106416418300920262940835654285629876306219380770501498610801101434455628546517517489977004485281513095129411801012356;
            6'd48: xpb[4] = 1024'd68409814667870641615162957177507246161700458615558132517499832681388721512250940829088099262823037219295535471455702951281596711557318738390649144607804880926409499297771056355368387275375314318307955929107246476307655911821175116303526106823917337954247891110078979025714945305185404258577363401119765200471;
            6'd49: xpb[4] = 1024'd15555839778313372286837654712432332797596989635872898472223392604656928167016753823229174341052451317649481261348376718471622879346728982405905113759155985537220027075620545777558665697323522530199493557294230011779657538012473926387671443146336065107394347764529411533912400633366323235641631672827729388586;
            6'd50: xpb[4] = 1024'd86768560572880844357311279652171852178191947781923348555078807592902030159091705727385320633939539725446576458698543920240712887977359560976321207926838131081721229423041252537379183310788936463401228793868453393616020014424669509436795349151984241527360707833096902072216384035475875229824589771161288061032;
            6'd51: xpb[4] = 1024'd33914585683323575028985977187096938814088478802238114509802367516170236813857518721526395712168953823800522248591217687430739055766769804991577177078189235692531757200890741959569461732737144675292766422055436929088021640615968319520940685474402968680507164487547334580413839363656794206888858042869252249147;
            6'd52: xpb[4] = 1024'd105127306477891047099459602126836458194683436948288564592657782504415338805932470625682542005056042231597617445941384889199829064397400383561993271245871381237032959548311448719389979346202558608494501658629660310924384117028163902570064591480051145100473524556114825118717822765766346201071816141202810921593;
            6'd53: xpb[4] = 1024'd52273331588333777771134299661761544830579967968603330547381342427683545460698283619823617083285456329951563235834058656389855232186810627577249240397222485847843487326160938141580257768150766820386039286816643846396385743219462712654209927802469872253619981210565257626915278093947265178136084412910775109708;
            6'd54: xpb[4] = 1024'd123486052382901249841607924601501064211174926114653780630236757415928647452773235523979763376172544737748658433184225858158945240817441206147665334564904631392344689673581644901400775381616180753587774523390867228232748219631658295703333833808118048673586341279132748165219261496056817172319042511244333782154;
            6'd55: xpb[4] = 1024'd70632077493343980513282622136426150847071457134968546584960317339196854107539048518120838454401958836102604223076899625348971408606851450162921303716255736003155217451431134323591053803564388965479312151577850763704749845822957105787479170130536775826732797933583180673416716824237736149383310782952297970269;
            6'd56: xpb[4] = 1024'd17778102603786711184957319671351237482967988155283312539683877262465060762304861512261913532631372934456550012969573392538997576396261694178177272867606840613965745229280623745781332225512597177370849779764834299176751472014255915871624506452955502979879254588033613181614172152418655126447579054660262158384;
            6'd57: xpb[4] = 1024'd88990823398354183255430944611090756863562946301333762622539292250710162754379813416418059825518461342253645210319740594308087585026892272748593367035288986158466947576701330505601849838978011110572585016339057681013113948426451498920748412458603679399845614656601103719918155554528207120630537152993820830830;
            6'd58: xpb[4] = 1024'd36136848508796913927105642146015843499459477321648528577262852173978369409145626410559134903747875440607591000212414361498113752816302516763849336186640090769277475354550819927792128260926219322464122644526041216485115574617750309004893748781022406552992071311051536228115610882709126097694805424701785018945;
            6'd59: xpb[4] = 1024'd107349569303364385997579267085755362880054435467698978660118267162223471401220578314715281196634963848404686197562581563267203761446933095334265430354322236313778677701971526687612645874391633255665857881100264598321478051029945892054017654786670582972958431379619026766419594284818678091877763523035343691391;
            6'd60: xpb[4] = 1024'd54495594413807116669253964620680449515950966488013744614841827085491678055986391308856356274864377946758631987455255330457229929236343339349521399505673340924589205479821016109802924296339841467557395509287248133793479677221244702138162991109089310126104888034069459274617049612999597068942031794743307879506;
            6'd61: xpb[4] = 1024'd1641619524249847340928662155605536151847497508328510569565387008759884710752204302997431353093792045112577777347929097647256097025753583364777368657024445535399733257670505531993202718288049679448933137474231669265481303412543512222308327431508037279251344688519891782814504941180516046006300066451272067621;
            6'd62: xpb[4] = 1024'd72854340318817319411402287095345055532442455654378960652420801997004986702827156207153577645980880452909672974698096299416346105656384161935193462824706591079900935605091212291813720331753463612650668374048455051101843779824739095271432233437156213699217704757087382321118488343290068040189258164784830740067;
            6'd63: xpb[4] = 1024'd20000365429260050083076984630270142168338986674693726607144361920273193357592969201294652724210294551263618764590770066606372273445794405950449431976057695690711463382940701714003998753701671824542206002235438586573845406016037905355577569759574940852364161411537814829315943671470987017253526436492794928182;
        endcase
    end

    always_comb begin
        case(flag[1][16:12])
            5'd0: xpb[5] = 1024'd0;
            5'd1: xpb[5] = 1024'd91213086223827522153550609570009661548933944820744176689999776908518295349667921105450799017097382959060713961940937268375462282076424984520865526143739841235212665730361408473824516367167085757743941238809661968410207882428233488404701475765223117272330521480105305367619927073580539011436484534826353600628;
            5'd2: xpb[5] = 1024'd58359476763530302908302291735204890353169462515752669251867698752059695362026703300886526819537091608678278516424381102171860723311629634486570927271148641536734656891151599610018793542816965794177684869232084090456054914635570203844424381847216785277841139546093552705133326073232445005754279243027112716925;
            5'd3: xpb[5] = 1024'd25505867303233083663053973900400119157404980210761161813735620595601095374385485496322254621976800258295843070907824935968259164546834284452276328398557441838256648051941790746213070718466845830611428499654506212501901946842906919284147287929210453283351757612081800042646725072884351000072073951227871833222;
            5'd4: xpb[5] = 1024'd116718953527060605816604583470409780706338925031505338503735397504119390724053406601773053639074183217356557032848762204343721446623259268973141854542297283073469313782303199220037587085633931588355369738464168180912109829271140407688848763694433570555682279092187105410266652146464890011508558486054225433850;
            5'd5: xpb[5] = 1024'd83865344066763386571356265635605009510574442726513831065603319347660790736412188797208781441513891866974121587332206038140119887858463918938847255669706083374991304943093390356231864261283811624789113368886590302957956861478477123128571669776427238561192897158175352747780051146116796005826353194254984550147;
            5'd6: xpb[5] = 1024'd51011734606466167326107947800800238314809960421522323627471241191202190748770970992644509243953600516591686141815649871936518329093668568904552656797114883676513296103883581492426141436933691661222856999309012425003803893685813838568294575858420906566703515224163600085293450145768702000144147902455743666444;
            5'd7: xpb[5] = 1024'd18158125146168948080859629965995467119045478116530816189339163034743590761129753188080237046393309166209250696299093705732916770328873218870258057924523683978035287264673772628620418612583571697656600629731434547049650925893150554008017481940414574572214133290151847422806849145420607994461942610656502782741;
            5'd8: xpb[5] = 1024'd109371211369996470234410239536005128667979422937274992879338939943261886110797674293531036063490692125269964658240030974108379052405298203391123584068263525213247952995035181102444934979750657455400541868541096515459858808321384042412718957705637691844544654770257152790426776219001147005898427145482856383369;
            5'd9: xpb[5] = 1024'd76517601909699250989161921701200357472214940632283485441206861786803286123156456488966763865930400774887529212723474807904777493640502853356828985195672325514769944155825372238639212155400537491834285498963518637505705840528720757852441863787631359850055272836245400127940175218653053000216221853683615499666;
            5'd10: xpb[5] = 1024'd43663992449402031743913603866395586276450458327291978003074783630344686135515238684402491668370109424505093767206918641701175934875707503322534386323081125816291935316615563374833489331050417528268029129385940759551552872736057473292164769869625027855565890902233647465453574218304958994534016561884374615963;
            5'd11: xpb[5] = 1024'd10810382989104812498665286031590815080685976022300470564942705473886086147874020879838219470809818074122658321690362475497574376110912153288239787450489926117813926477405754511027766506700297564701772759808362881597399904943394188731887675951618695861076508968221894802966973217956864988851811270085133732260;
            5'd12: xpb[5] = 1024'd102023469212932334652215895601600476629619920843044647254942482382404381497541941985289018487907201033183372283631299743873036658187337137809105313594229767353026592207767162984852282873867383322445713998618024850007607787371627677136589151716841813133407030448327200170586900291537404000288295804911487332888;
            5'd13: xpb[5] = 1024'd69169859752635115406967577766795705433855438538053139816810404225945781509900724180724746290346909682800936838114743577669435099422541787774810714721638567654548583368557354121046560049517263358879457629040446972053454819578964392576312057798835481138917648514315447508100299291189309994606090513112246449185;
            5'd14: xpb[5] = 1024'd36316250292337896161719259931990934238090956233061632378678326069487181522259506376160474092786618332418501392598187411465833540657746437740516115849047367956070574529347545257240837225167143395313201259462869094099301851786301108016034963880829149144428266580303694845613698290841215988923885221313005565482;
            5'd15: xpb[5] = 1024'd3462640832040676916470942097186163042326473928070124940546247913028581534618288571596201895226326982036065947081631245262231981892951087706221516976456168257592565690137736393435114400817023431746944889885291216145148883993637823455757869962822817149938884646291942183127097290493121983241679929513764681779;
            5'd16: xpb[5] = 1024'd94675727055868199070021551667195824591260418748814301630546024821546876884286209677047000912323709941096779909022568513637694263969376072227087043120196009492805231420499144867259630767984109189490886128694953184555356766421871311860459345728045934422269406126397247550747024364073660994678164464340118282407;
            5'd17: xpb[5] = 1024'd61822117595570979824773233832391053395495936443822794192413946665088276896644991872482728714763418590714344463506012347434092705204580722192792444247604809794327222581289336003453907943633989225924629759117375306601203798629208027300182251810039602427780024192385494888260423363725566988995959172540877398704;
            5'd18: xpb[5] = 1024'd28968508135273760579524915997586282199731454138831286754281868508629676909003774067918456517203127240331909017989456181230491146439785372158497845375013610095849213742079527139648185119283869262358373389539797428647050830836544742739905157892033270433290642258373742225773822363377472983313753880741636515001;
            5'd19: xpb[5] = 1024'd120181594359101282733075525567595943748665398959575463444281645417147972258671695173369255534300510199392622979930393449605953428516210356679363371518753451331061879472440935613472701486450955020102314628349459397057258713264778231144606633657256387705621163738479047593393749436958011994750238415567990115629;
            5'd20: xpb[5] = 1024'd87327984898804063487827207732791172552900916654583956006149567260689372271030477368804983336740218849010187534413837283402351869751415006645068772646162251632583870633231126749666978662100835056536058258771881519103105745472114946584329539739250055711131781804467294930907148436609917989068033123768749231926;
            5'd21: xpb[5] = 1024'd54474375438506844242578889897986401357136434349592448568017489104230772283389259564240711139179927498627752088897281117198750310986619656610774173773571051934105861794021317885861255837750715092969801889194303641148952777679451662024052445821243723716642399870455542268420547436261823983385827831969508348223;
            5'd22: xpb[5] = 1024'd21620765978209624997330572063181630161371952044600941129885410947772172295748041759676438941619636148245316643380724950995148752221824306576479574900979852235627852954811509022055533013400595129403545519616725763194799809886788377463775351903237391722153017936443789605933946435913729977703622540170267464520;
            5'd23: xpb[5] = 1024'd112833852202037147150881181633191291710305896865345117819885187856290467645415962865127237958717019107306030605321662219370611034298249291097345101044719693470840518685172917495880049380567680887147486758426387731605007692315021865868476827668460508994483539416549094973553873509494268989140107074996621065148;
            5'd24: xpb[5] = 1024'd79980242741739927905632863798386520514541414560353610381753109699831867657774745060562965761156727756923595159805106053167009475533453941063050502172128493772362509845963108632074326556217560923581230388848809853650854724522358581308199733750454176999994157482537342311067272509146174983457901783197380181445;
            5'd25: xpb[5] = 1024'd47126633281442708660384545963581749318776932255362102943621031543373267670133527255998693563596436406541159714288549886963407916768658591028755903299537294073884501006753299768268603731867440960014974019271231975696701756729695296747922639832447845005504775548525589648580671508798080977775696491398139297742;
            5'd26: xpb[5] = 1024'd14273023821145489415136228128776978123012449950370595505488953386914667682492309451434421366036145056158724268771993720759806358003863240994461304426946094375406492167543490904462880907517320996448717649693654097742548788937032012187645545914441513011015393614513836986094070508449986972093491199598898414039;
            5'd27: xpb[5] = 1024'd105486110044973011568686837698786639671946394771114772195488730295432963032160230556885220383133528015219438230712930989135268640080288225515326830570685935610619157897904899378287397274684406754192658888503316066152756671365265500592347021679664630283345915094619142353713997582030525983529975734425252014667;
            5'd28: xpb[5] = 1024'd72632500584675792323438519863981868476181912466123264757356652138974363044519012752320948185573236664837002785196374822931667081315492875481032231698094735912141149058695090514481674450334286790626402518925738188198603703572602216032069927761658298288856533160607389691227396581682431977847770442626011130964;
            5'd29: xpb[5] = 1024'd39778891124378573078190202029177097280417430161131757319224573982515763056877794947756675988012945314454567339679818656728065522550697525446737632825503536213663140219485281650675951625984166827060146149348160310244450735779938931471792833843651966294367151226595637028740795581334337972165565150826770247261;
            5'd30: xpb[5] = 1024'd6925281664081353832941884194372326084652947856140249881092495826057163069236577143192403790452653964072131894163262490524463963785902175412443033952912336515185131380275472786870228801634046863493889779770582432290297767987275646911515739925645634299877769292583884366254194580986243966483359859027529363558;
            5'd31: xpb[5] = 1024'd98138367887908875986492493764381987633586892676884426571092272734575458418904498248643202807550036923132845856104199758899926245862327159933308560096652177750397797110636881260694745168801132621237831018580244400700505650415509135316217215690868751572208290772689189733874121654566782977919844393853882964186;
        endcase
    end

    always_comb begin
        case(flag[2][5:0])
            6'd0: xpb[6] = 1024'd0;
            6'd1: xpb[6] = 1024'd94675727055868199070021551667195824591260418748814301630546024821546876884286209677047000912323709941096779909022568513637694263969376072227087043120196009492805231420499144867259630767984109189490886128694953184555356766421871311860459345728045934422269406126397247550747024364073660994678164464340118282407;
            6'd2: xpb[6] = 1024'd65284758427611656741244175929577216437822410371892919132960194578116858431263280444078930609989745572750410410587643592696324687097531809899013961224060978051919788271427072396889022344451012657671574649002666522746352682622845850755940121772862419577718908838677437071387520654218688972237639102054642080483;
            6'd3: xpb[6] = 1024'd35893789799355114412466800191958608284384401994971536635374364334686839978240351211110860307655781204404040912152718671754955110225687547570940879327925946611034345122354999926518413920917916125852263169310379860937348598823820389651420897817678904733168411550957626592028016944363716949797113739769165878559;
            6'd4: xpb[6] = 1024'd6502821171098572083689424454340000130946393618050154137788534091256821525217421978142790005321816836057671413717793750813585533353843285242867797431790915170148901973282927456147805497384819594032951689618093199128344515024794928546901673862495389888617914263237816112668513234508744927356588377483689676635;
            6'd5: xpb[6] = 1024'd101178548226966771153710976121535824722206812366864455768334558912803698409503631655189790917645526777154451322740362264451279797323219357469954840551986924662954133393782072323407436265368928783523837818313046383683701281446666240407361019590541324310887320389635063663415537598582405922034752841823807959042;
            6'd6: xpb[6] = 1024'd71787579598710228824933600383917216568768803989943073270748728669373679956480702422221720615311562408808081824305437343509910220451375095141881758655851893222068690244709999853036827841835832251704526338620759721874697197647640779302841795635357809466336823101915253184056033888727433899594227479538331757118;
            6'd7: xpb[6] = 1024'd42396610970453686496156224646298608415330795613021690773162898425943661503457773189253650312977598040461712325870512422568540643579530832813808676759716861781183247095637927382666219418302735719885214858928473060065693113848615318198322571680174294621786325814195442704696530178872461877153702117252855555194;
            6'd8: xpb[6] = 1024'd13005642342197144167378848908680000261892787236100308275577068182513643050434843956285580010643633672115342827435587501627171066707686570485735594863581830340297803946565854912295610994769639188065903379236186398256689030049589857093803347724990779777235828526475632225337026469017489854713176754967379353270;
            6'd9: xpb[6] = 1024'd107681369398065343237400400575875824853153205984914609906123093004060519934721053633332580922967343613212122736458156015264865330677062642712822637983777839833103035367064999779555241762753748377556789507931139582812045796471461168954262693453036714199505234652872879776084050833091150849391341219307497635677;
            6'd10: xpb[6] = 1024'd78290400769808800908623024838257216699715197607993227408537262760630501481698124400364510620633379244865753238023231094323495753805218380384749556087642808392217592217992927309184633339220651845737478028238852921003041712672435707849743469497853199354954737365153069296724547123236178826950815857022021433753;
            6'd11: xpb[6] = 1024'd48899432141552258579845649100638608546277189231071844910951432517200483028675195167396440318299414876519383739588306173382126176933374118056676474191507776951332149068920854838814024915687555313918166548546566259194037628873410246745224245542669684510404240077433258817365043413381206804510290494736545231829;
            6'd12: xpb[6] = 1024'd19508463513295716251068273363020000392839180854150462413365602273770464575652265934428370015965450508173014241153381252440756600061529855728603392295372745510446705919848782368443416492154458782098855068854279597385033545074384785640705021587486169665853742789713448338005539703526234782069765132451069029905;
            6'd13: xpb[6] = 1024'd114184190569163915321089825030215824984099599602964764043911627095317341459938475611475370928289160449269794150175949766078450864030905927955690435415568755003251937340347927235703047260138567971589741197549232781940390311496256097501164367315532104088123148916110695888752564067599895776747929596791187312312;
            6'd14: xpb[6] = 1024'd84793221940907372992312449292597216830661591226043381546325796851887323006915546378507300625955196080923424651741024845137081287159061665627617353519433723562366494191275854765332438836605471439770429717856946120131386227697230636396645143360348589243572651628390885409393060357744923754307404234505711110388;
            6'd15: xpb[6] = 1024'd55402253312650830663535073554978608677223582849121999048739966608457304553892617145539230323621231712577055153306099924195711710287217403299544271623298692121481051042203782294961830413072374907951118238164659458322382143898205175292125919405165074399022154340671074930033556647889951731866878872220234908464;
            6'd16: xpb[6] = 1024'd26011284684394288334757697817360000523785574472200616551154136365027286100869687912571160021287267344230685654871175003254342133415373140971471189727163660680595607893131709824591221989539278376131806758472372796513378060099179714187606695449981559554471657052951264450674052938034979709426353509934758706540;
            6'd17: xpb[6] = 1024'd120687011740262487404779249484555825115045993221014918181700161186574162985155897589618160933610977285327465563893743516892036397384749213198558232847359670173400839313630854691850852757523387565622692887167325981068734826521051026048066041178027493976741063179348512001421077302108640704104517974274876988947;
            6'd18: xpb[6] = 1024'd91296043112005945076001873746937216961607984844093535684114330943144144532132968356650090631277012916981096065458818595950666820512904950870485150951224638732515396164558782221480244333990291033803381407475039319259730742722025564943546817222843979132190565891628701522061573592253668681663992611989400787023;
            6'd19: xpb[6] = 1024'd61905074483749402747224498009318608808169976467172153186528500699714126079110039123682020328943048548634726567023893675009297243641060688542412069055089607291629953015486709751109635910457194501984069927782752657450726658923000103839027593267660464287640068603908891042702069882398696659223467249703924585099;
            6'd20: xpb[6] = 1024'd32514105855492860418447122271700000654731968090250770688942670456284107626087109890713950026609084180288357068588968754067927666769216426214338987158954575850744509866414637280739027486924097970164758448090465995641722575123974642734508369312476949443089571316189080563342566172543724636782941887418448383175;
            6'd21: xpb[6] = 1024'd3123137227236318089669746534081392501293959713329388191356840212854089173064180657745879724275119811941987570154043833126558089897372163886265905262819544409859066717342564810368419063391001438345446968398179333832718491324949181629989145357293434598539074028469270083983062462688752614342416525132972181251;
            6'd22: xpb[6] = 1024'd97798864283104517159691298201277217092554378462143689821902865034400966057350390334792880636598829753038767479176612346764252353866748236113352948383015553902664298137841709677628049831375110627836333097093132518388075257746820493490448491085339369020808480154866517634730086826762413609020580989473090463658;
            6'd23: xpb[6] = 1024'd68407895654847974830913922463658608939116370085222307324317034790970947604327461101824810334264865384692397980741687425822882776994903973785279866486880522461778854988769637207257441407842014096017021617400845856579071173947795032385929267130155854176257982867146707155370583116907441586580055627187614261734;
            6'd24: xpb[6] = 1024'd39016927026591432502136546726040000785678361708300924826731204547540929151304531868856740031930901016346028482306762504881513200123059711457206784590745491020893411839697564736886832984308917564197710137708559194770067090148769571281410043174972339331707485579426896676011079407052469564139530264902138059810;
            6'd25: xpb[6] = 1024'd9625958398334890173359170988421392632240353331379542329145374304110910698281602635888669729596936647999658983871837583940143623251215449129133702694610459580007968690625492266516224560775821032378398658016272532961063006349744110176890819219788824487156988291707086196651575697197497541699004902616661857886;
            6'd26: xpb[6] = 1024'd104301685454203089243380722655617217223500772080193843959691399125657787582567812312935670641920646589096438892894406097577837887220591521356220745814806469072813200111124637133775855328759930221869284786711225717516419772771615422037350164947834758909426394418104333747398600061271158536377169366956780140293;
            6'd27: xpb[6] = 1024'd74910716825946546914603346917998609070062763703272461462105568882227769129544883079967600339586682220750069394459481176636468310348747259028147663918671437631927756962052564663405246905226833690049973307018939055707415688972589960932830940992651244064875897130384523268039096351416186513936644004671303938369;
            6'd28: xpb[6] = 1024'd45519748197690004585825971180380000916624755326351078964519738638797750676521953846999530037252717852403699896024556255695098733476902996700074582022536406191042313812980492193034638481693737158230661827326652393898411605173564499828311717037467729220325399842664712788679592641561214491496118642385827736445;
            6'd29: xpb[6] = 1024'd16128779569433462257048595442761392763186746949429696466933908395367732223499024614031459734918753484057330397589631334753729156605058734372001500126401374750156870663908419722664030058160640626411350347634365732089407521374539038723792493082284214375774902554944902309320088931706242469055593280100351534521;
            6'd30: xpb[6] = 1024'd110804506625301661327070147109957217354447165698243998097479933216914609107785234291078460647242463425154110306612199848391423420574434806599088543246597384242962102084407564589923660826144749815902236476329318916644764287796410350584251838810330148798044308681342149860067113295779903463733757744440469816928;
            6'd31: xpb[6] = 1024'd81413537997045118998292771372338609201009157321322615599894102973484590654762305058110390344908499056807740808177274927450053843702590544271015461350462352802076658935335492119553052402611653284082924996637032254835760203997384889479732614855146633953493811393622339380707609585924931441293232382154993615004;
            6'd32: xpb[6] = 1024'd52022569368788576669515395634720001047571148944401233102308272730054572201739375825142320042574534688461371309742350006508684266830746281942942379454327321361191215786263419649182443979078556752263613516944745593026756120198359428375213390899963119108943314105902528901348105876069959418852707019869517413080;
            6'd33: xpb[6] = 1024'd22631600740532034340738019897101392894133140567479850604722442486624553748716446592174249740240570320115001811307425085567314689958902019614869297558192289920305772637191347178811835555545460220444302037252458931217752036399333967270694166944779604264392816818182718421988602166214987396412181657584041211156;
            6'd34: xpb[6] = 1024'd117307327796400233410759571564297217485393559316294152235268467308171430633002656269221250652564280261211781720329993599205008953928278091841956340678388299413111004057690492046071466323529569409935188165947412115773108802821205279131153512672825538686662222944579965972735626530288648391090346121924159493563;
            6'd35: xpb[6] = 1024'd87916359168143691081982195826678609331955550939372769737682637064741412179979727036253180350230315892865412221895068678263639377056433829513883258782253267972225560908618419575700857899996472878115876686255125453964104719022179818026634288717642023842111725656860155493376122820433676368649820759638683291639;
            6'd36: xpb[6] = 1024'd58525390539887148753204820089060001178517542562451387240096806821311393726956797803285110047896351524519042723460143757322269800184589567185810176886118236531340117759546347105330249476463376346296565206562838792155100635223154356922115064762458508997561228369140345014016619110578704346209295397353207089715;
            6'd37: xpb[6] = 1024'd29134421911630606424427444351441393025079534185530004742510976577881375273933868570317039745562387156172673225025218836380900223312745304857737094989983205090454674610474274634959641052930279814477253726870552130346096551424128895817595840807274994153010731081420534534657115400723732323768770035067730887791;
            6'd38: xpb[6] = 1024'd123810148967498805494448996018637217616339952934344306373057001399428252158220078247364040657886097097269453134047787350018594487282121377084824138110179214583259906030973419502219271820914389003968139855565505314901453317846000207678055186535320928575280137207817782085404139764797393318446934499407849170198;
            6'd39: xpb[6] = 1024'd94419180339242263165671620281018609462901944557422923875471171155998233705197149014395970355552132728923083635612862429077224910410277114756751056214044183142374462881901347031848663397381292472148828375873218653092449234046974746573535962580137413730729639920097971606044636054942421296006409137122372968274;
            6'd40: xpb[6] = 1024'd65028211710985720836894244543400001309463936180501541377885340912568215252174219781427900053218168360576714137177937508135855333538432852428677974317909151701489019732829274561478054973848195940329516896180931991283445150247949285469016738624953898886179142632378161126685132345087449273565883774836896766350;
            6'd41: xpb[6] = 1024'd35637243082729178508116868805781393156025927803580158880299510669138196799151290548459829750884203992230344638743012587194485756666588590100604892421774120260603576583757202091107446550315099408510205416488645329474441066448923824364497514669770384041628645344658350647325628635232477251125358412551420564426;
            6'd42: xpb[6] = 1024'd6246274454472636179339493068162785002587919426658776382713680425708178346128361315491759448550239623883975140308087666253116179794744327772531810525639088819718133434685129620736838126782002876690893936796358667665436982649898363259978290714586869197078148056938540167966124925377505228684833050265944362502;
            6'd43: xpb[6] = 1024'd100922001510340835249361044735358609593848338175473078013259705247255055230414570992538760360873949564980755049330656179890810443764120399999618853645835098312523364855184274487996468894766112066181780065491311852220793749071769675120437636442632803619347554183335787718713149289451166223362997514606062644909;
            6'd44: xpb[6] = 1024'd71531032882084292920583668997740001440410329798551695515673875003825036777391641759570690058539985196634385550895731258949440866892276137671545771749700066871637921706112202017625860471233015534362468585799025190411789665272744214015918412487449288774797056895615977239353645579596194200922472152320586442985;
            6'd45: xpb[6] = 1024'd42140064253827750591806293260121393286972321421630313018088044760395018324368712526602619756206020828288016052460806338008071290020431875343472689853565035430752478557040129547255252047699919002543157106106738528602785581473718752911399188532265773930246559607896166759994141869741222178481946790035110241061;
            6'd46: xpb[6] = 1024'd12749095625571208263028917522502785133534313044708930520502214516964999871345783293634549453872056459941646554025881417066701713148587613015399607957430003989867035407968057076884643624166822470723845626414451866793781497674693291806879964577082259085696062320176356280634638159886250156041421427749634039137;
            6'd47: xpb[6] = 1024'd107424822681439407333050469189698609724794731793523232151048239338511876755631992970681550366195766401038426463048449930704395977117963685242486651077626013482672266828467201944144274392150931660214731755109405051349138264096564603667339310305128193507965468446573603831381662523959911150719585892089752321544;
            6'd48: xpb[6] = 1024'd78033854053182865004273093452080001571356723416601849653462409095081858302609063737713480063861802032692056964613525009763026400246119422914413569181490982041786823679395129473773665968617835128395420275417118389540134180297539142562820086349944678663414971158853793352022158814104939128279060529804276119620;
            6'd49: xpb[6] = 1024'd48642885424926322675495717714461393417918715039680467155876578851651839849586134504745409761527837664345687466178600088821656823374275160586340487285355950600901380530323057003403057545084738596576108795724831727731130096498513681458300862394761163818864473871133982872662655104249967105838535167518799917696;
            6'd50: xpb[6] = 1024'd19251916796669780346718341976842785264480706662759084658290748608221821396563205271777339459193873295999317967743675167880287246502430898258267405389220919160015937381250984533032449121551642064756797316032545065922126012699488220353781638439577648974313976583414172393303151394394995083398009805233323715772;
            6'd51: xpb[6] = 1024'd113927643852537979416739893644038609855741125411573386288836773429768698280849414948824340371517583237096097876766243681517981510471806970485354448509416928652821168801750129400292079889535751254247683444727498250477482779121359532214240984167623583396583382709811419944050175758468656078076174269573441998179;
            6'd52: xpb[6] = 1024'd84536675224281437087962517906420001702303117034652003791250943186338679827826485715856270069183618868749728378331318760576611933599962708157281366613281897211935725652678056929921471466002654722428371965035211588668478695322334071109721760212440068552032885422091609464690672048613684055635648907287965796255;
            6'd53: xpb[6] = 1024'd55145706596024894759185142168801393548865108657730621293665112942908661374803556482888199766849654500403358879896393839635242356728118445829208284717146865771050282503605984459550863042469558190609060485342924926859474611523308610005202536257256553707482388134371798985331168338758712033195123545002489594331;
            6'd54: xpb[6] = 1024'd25754737967768352430407766431182785395427100280809238796079282699478642921780627249920129464515690132056989381461468918693872779856274183501135202821011834330164839354533911989180254618936461658789749005650638265050470527724283148900683312302073038862931890846651988505971664628903740010754598182717013392407;
            6'd55: xpb[6] = 1024'd120430465023636551500429318098378609986687519029623540426625307521025519806066836926967130376839400073153769290484037432331567043825650255728222245941207843822970070775033056856439885386920570848280635134345591449605827294146154460761142658030118973285201296973049236056718688992977401005432762647057131674814;
            6'd56: xpb[6] = 1024'd91039496395380009171651942360760001833249510652702157929039477277595501353043907693999060074505435704807399792049112511390197466953805993400149164045072812382084627625960984386069276963387474316461323654653304787796823210347128999656623434074935458440650799685329425577359185283122428982992237284771655472890;
            6'd57: xpb[6] = 1024'd61648527767123466842874566623141393679811502275780775431453647034165482900020978461030989772171471336461030293614187590448827890081961731072076082148937780941199184476888911915698668539854377784642012174961018125987819126548103538552104210119751943596100302397609615097999681573267456960551711922486179270966;
            6'd58: xpb[6] = 1024'd32257559138866924514097190885522785526373493898859392933867816790735464446998049228062919469837506968114660795179262669507458313210117468744003000252802749500313741327816839445328060116321281252822700695268731464178815042749078077447584986164568428751549805109889804618640177863412484938111186560200703069042;
            6'd59: xpb[6] = 1024'd2866590510610382185319815147904177372935485521938010436281986547305445993975119995094849167503542599768291296744337748566088736338273206415929918356667718059428298178744766974957451692788184721003389215576444802369810958950052616343065762209384913906999307822169994139280674153557512915670661197915226867118;
            6'd60: xpb[6] = 1024'd97542317566478581255341366815100001964195904270752312066828011368852322878261329672141850079827252540865071205766906262203783000307649278643016961476863727552233529599243911842217082460772293910494275344271397986925167725371923928203525107937430848329268713948567241690027698517631173910348825662255345149525;
            6'd61: xpb[6] = 1024'd68151348938222038926563991077481393810757895893830929569242181125422304425238400439173779777493288172518701707331981341262413423435805016314943879580728696111348086450171839371846474037239197378674963864579111325116163641572898467099005883982247333484718216660847431210668194807776201887908300299969868947601;
            6'd62: xpb[6] = 1024'd38760380309965496597786615339862785657319887516909547071656350881992285972215471206205709475159323804172332208897056420321043846563960753986870797684593664670462643301099766901475865613706100846855652384886824663307159557773873005994486660027063818640167719373127620731308691097921229865467774937684392745677;
            6'd63: xpb[6] = 1024'd9369411681708954269009239602244177503881879139988164574070520638562267519192541973237639172825359435825962710462131499379674269692116491658797715788458633229577200152027694431105257190173004315036340905194538001498155473974847544889967436071880303795617222085407810251949187388066257843027249575398916543753;
        endcase
    end

    always_comb begin
        case(flag[2][11:6])
            6'd0: xpb[7] = 1024'd0;
            6'd1: xpb[7] = 1024'd104045138737577153339030791269440002095142297888802466204616545460109144403478751650284640085149069376922742619484700013017368533661492563885884758908654642722382431572526839298364887958157113504527227033889491186053512240396718856750426781799926238217886628211805057802696211752139918837705414039739034826160;
            6'd2: xpb[7] = 1024'd84023581791029565279262655134065571445586168651869248281101235855241393469648364390554208955640464444402335831511906591455673226481764793216609392800978244511074188575482461259099536724797021287744256459391742525742663630572540940535874993916623027168953353009493057575285895430351204658292138252852475167989;
            6'd3: xpb[7] = 1024'd64002024844481977219494518998691140796030039414936030357585926250373642535817977130823777826131859511881929043539113169893977919302037022547334026693301846299765945578438083219834185491436929070961285884893993865431815020748363024321323206033319816120020077807181057347875579108562490478878862465965915509818;
            6'd4: xpb[7] = 1024'd43980467897934389159726382863316710146473910178002812434070616645505891601987589871093346696623254579361522255566319748332282612122309251878058660585625448088457702581393705180568834258076836854178315310396245205120966410924185108106771418150016605071086802604869057120465262786773776299465586679079355851647;
            6'd5: xpb[7] = 1024'd23958910951386801099958246727942279496917780941069594510555307040638140668157202611362915567114649646841115467593526326770587304942581481208783294477949049877149459584349327141303483024716744637395344735898496544810117801100007191892219630266713394022153527402557056893054946464985062120052310892192796193476;
            6'd6: xpb[7] = 1024'd3937354004839213040190110592567848847361651704136376587039997435770389734326815351632484437606044714320708679620732905208891997762853710539507928370272651665841216587304949102038131791356652420612374161400747884499269191275829275677667842383410182973220252200245056665644630143196347940639035105306236535305;
            6'd7: xpb[7] = 1024'd107982492742416366379220901862007850942503949592938842791656542895879534137805567001917124522755114091243451299105432918226260531424346274425392687278927294388223648159831788400403019749513765925139601195290239070552781431672548132428094624183336421191106880412050114468340841895336266778344449145045271361465;
            6'd8: xpb[7] = 1024'd87960935795868778319452765726633420292947820356005624868141233291011783203975179742186693393246509158723044511132639496664565224244618503756117321171250896176915405162787410361137668516153673708356630620792490410241932821848370216213542836300033210142173605209738114240930525573547552598931173358158711703294;
            6'd9: xpb[7] = 1024'd67939378849321190259684629591258989643391691119072406944625923686144032270144792482456262263737904226202637723159846075102869917064890733086841955063574497965607162165743032321872317282793581491573660046294741749931084212024192299998991048416729999093240330007426114013520209251758838419517897571272152045123;
            6'd10: xpb[7] = 1024'd47917821902773602199916493455884558993835561882139189021110614081276281336314405222725831134229299293682230935187052653541174609885162962417566588955898099754298919168698654282606966049433489274790689471796993089620235602200014383784439260533426788044307054805114113786109892929970124240104621784385592386952;
            6'd11: xpb[7] = 1024'd27896264956226014140148357320510128344279432645205971097595304476408530402484017962995400004720694361161824147214259231979479302705435191748291222848221701542990676171654276243341614816073397058007718897299244429309386992375836467569887472650123576995373779602802113558699576608181410060691345997499032728781;
            6'd12: xpb[7] = 1024'd7874708009678426080380221185135697694723303408272753174079994871540779468653630703264968875212089428641417359241465810417783995525707421079015856740545303331682433174609898204076263582713304841224748322801495768998538382551658551355335684766820365946440504400490113331289260286392695881278070210612473070610;
            6'd13: xpb[7] = 1024'd111919846747255579419411012454575699789865601297075219378696540331649923872132382353549608960361158805564159978726165823435152529187199984964900615649199946054064864747136737502441151540870418345751975356690986955052050622948377408105762466566746604164327132612295171133985472038532614718983484250351507896770;
            6'd14: xpb[7] = 1024'd91898289800707991359642876319201269140309472060142001455181230726782172938301995093819177830852553873043753190753372401873457222007472214295625249541523547842756621750092359463175800307510326128969004782193238294741202013124199491891210678683443393115393857409983170906575155716743900539570208463464948238599;
            6'd15: xpb[7] = 1024'd71876732854160403299874740183826838490753342823208783531665921121914422004471607834088746701343948940523346402780578980311761914827744443626349883433847149631448378753047981423910449074150233912186034207695489634430353403300021575676658890800140182066460582207671170679164839394955186360156932676578388580428;
            6'd16: xpb[7] = 1024'd51855175907612815240106604048452407841197213586275565608150611517046671070641220574358315571835344008002939614807785558750066607648016672957074517326170751420140135756003603384645097840790141695403063633197740974119504793475843659462107102916836971017527307005359170451754523073166472180743656889691828922257;
            6'd17: xpb[7] = 1024'd31833618961065227180338467913077977191641084349342347684635301912178920136810833314627884442326739075482532826834992137188371300468288902287799151218494353208831892758959225345379746607430049478620093058699992313808656183651665743247555315033533759968594031803047170224344206751377758001330381102805269264086;
            6'd18: xpb[7] = 1024'd11812062014517639120570331777703546542084955112409129761119992307311169202980446054897453312818134142962126038862198715626675993288561131618523785110817954997523649761914847306114395374069957261837122484202243653497807573827487827033003527150230548919660756600735169996933890429589043821917105315918709605915;
            6'd19: xpb[7] = 1024'd115857200752094792459601123047143548637227253001211595965736537767420313606459197705182093397967203519884868658346898728644044526950053695504408544019472597719906081334441686604479283332227070766364349518091734839551319814224206683783430308950156787137547384812540227799630102181728962659622519355657744432075;
            6'd20: xpb[7] = 1024'd95835643805547204399832986911769117987671123764278378042221228162552562672628810445451662268458598587364461870374105307082349219770325924835133177911796199508597838337397308565213932098866978549581378943593986179240471204400028767568878521066853576088614109610228227572219785859940248480209243568771184773904;
            6'd21: xpb[7] = 1024'd75814086858999616340064850776394687338114994527345160118705918557684811738798423185721231138949993654844055082401311885520653912590598154165857811804119801297289595340352930525948580865506886332798408369096237518929622594575850851354326733183550365039680834407916227344809469538151534300795967781884625115733;
            6'd22: xpb[7] = 1024'd55792529912452028280296714641020256688558865290411942195190608952817060804968035925990800009441388722323648294428518463958958605410870383496582445696443403085981352343308552486683229632146794116015437794598488858618773984751672935139774945300247153990747559205604227117399153216362820121382691994998065457562;
            6'd23: xpb[7] = 1024'd35770972965904440220528578505645826039002736053478724271675299347949309871137648666260368879932783789803241506455725042397263298231142612827307079588767004874673109346264174447417878398786701899232467220100740198307925374927495018925223157416943942941814284003292226889988836894574105941969416208111505799391;
            6'd24: xpb[7] = 1024'd15749416019356852160760442370271395389446606816545506348159989743081558937307261406529937750424178857282834718482931620835567991051414842158031713481090606663364866349219796408152527165426609682449496645602991537997076765103317102710671369533640731892881008800980226662578520572785391762556140421224946141220;
            6'd25: xpb[7] = 1024'd119794554756934005499791233639711397484588904705347972552776535203190703340786013056814577835573248234205577337967631633852936524712907406043916472389745249385747297921746635706517415123583723186976723679492482724050589005500035959461098151333566970110767637012785284465274732324925310600261554460963980967380;
            6'd26: xpb[7] = 1024'd99772997810386417440023097504336966835032775468414754629261225598322952406955625797084146706064643301685170549994838212291241217533179635374641106282068851174439054924702257667252063890223630970193753104994734063739740395675858043246546363450263759061834361810473284237864416003136596420848278674077421309209;
            6'd27: xpb[7] = 1024'd79751440863838829380254961368962536185476646231481536705745915993455201473125238537353715576556038369164763762022044790729545910353451864705365740174392452963130811927657879627986712656863538753410782530496985403428891785851680127031994575566960548012901086608161284010454099681347882241435002887190861651038;
            6'd28: xpb[7] = 1024'd59729883917291241320486825233588105535920516994548318782230606388587450539294851277623284447047433436644356974049251369167850603173724094036090374066716054751822568930613501588721361423503446536627811955999236743118043176027502210817442787683657336963967811405849283783043783359559168062021727100304301992867;
            6'd29: xpb[7] = 1024'd39708326970743653260718689098213674886364387757615100858715296783719699605464464017892853317538828504123950186076457947606155295993996323366815007959039656540514325933569123549456010190143354319844841381501488082807194566203324294602890999800354125915034536203537283555633467037770453882608451313417742334696;
            6'd30: xpb[7] = 1024'd19686770024196065200950552962839244236808258520681882935199987178851948671634076758162422188030223571603543398103664526044459988814268552697539641851363258329206082936524745510190658956783262103061870807003739422496345956379146378388339211917050914866101261001225283328223150715981739703195175526531182676525;
            6'd31: xpb[7] = 1024'd123731908761773218539981344232279246331950556409484349139816532638961093075112828408447062273179292948526286017588364539061828522475761116583424400760017901051588514509051584808555546914940375607589097840893230608549858196775865235138765993716977153083987889213030341130919362468121658540900589566270217502685;
            6'd32: xpb[7] = 1024'd103710351815225630480213208096904815682394427172551131216301223034093342141282441148716631143670688016005879229615571117500133215296033345914149034652341502840280271512007206769290195681580283390806127266395481948239009586951687318924214205833673942035054614010718340903509046146332944361487313779383657844514;
            6'd33: xpb[7] = 1024'd83688794868678042420445071961530385032838297935617913292785913429225591207452053888986200014162083083485472441642777695938437908116305575244873668544665104628972028514962828730024844448220191174023156691897733287928160977127509402709662417950370730986121338808406340676098729824544230182074037992497098186343;
            6'd34: xpb[7] = 1024'd63667237922130454360676935826155954383282168698684695369270603824357840273621666629255768884653478150965065653669984274376742600936577804575598302436988706417663785517918450690759493214860098957240186117399984627617312367303331486495110630067067519937188063606094340448688413502755516002660762205610538528172;
            6'd35: xpb[7] = 1024'd43645680975582866300908799690781523733726039461751477445755294219490089339791279369525337755144873218444658865697190852815047293756850033906322936329312308206355542520874072651494141981500006740457215542902235967306463757479153570280558842183764308888254788403782340221278097180966801823247486418723978870001;
            6'd36: xpb[7] = 1024'd23624124029035278241140663555407093084169910224818259522239984614622338405960892109794906625636268285924252077724397431253351986577122263237047570221635909995047299523829694612228790748139914523674244968404487306995615147654975654066007054300461097839321513201470339993867780859178087643834210631837419211830;
            6'd37: xpb[7] = 1024'd3602567082487690181372527420032662434613780987885041598724675009754587472130504850064475496127663353403845289751604009691656679397394492567772204113959511783739056526785316572963439514779822306891274393906738646684766537830797737851455266417157886790388237999158339766457464537389373464420934844950859553659;
            6'd38: xpb[7] = 1024'd107647705820064843520403318689472664529756078876687507803341220469863731875609256500349115581276732730326587909236304022709025213058887056453656963022614154506121488099312155871328327472936935811418501427796229832738278778227516594601882048217084125008274866210963397569153676289529292302126348884689894379819;
            6'd39: xpb[7] = 1024'd87626148873517255460635182554098233880199949639754289879825910864995980941778869240618684451768127797806181121263510601147329905879159285784381596914937756294813245102267777832062976239576843594635530853298481172427430168403338678387330260333780913959341591008651397341743359967740578122713073097803334721648;
            6'd40: xpb[7] = 1024'd67604591926969667400867046418723803230643820402821071956310601260128230007948481980888253322259522865285774333290717179585634598699431515115106230807261358083505002105223399792797625006216751377852560278800732512116581558579160762172778472450477702910408315806339397114333043645951863943299797310916775063477;
            6'd41: xpb[7] = 1024'd47583034980422079341098910283349372581087691165887854032795291655260479074118094721157822192750917932765367545317923758023939291519703744445830864699584959872196759108179021753532273772856659161069589704302983851805732948754982845958226684567174491861475040604027396886922727324163149763886521524030215405306;
            6'd42: xpb[7] = 1024'd27561478033874491281330774147974941931531561928954636109279982050392728140287707461427391063242313000244960757345130336462243984339975973776555498591908561660888516111134643714266922539496566944286619129805235191494884338930804929743674896683871280812541765401715396659512411002374435584473245737143655747135;
            6'd43: xpb[7] = 1024'd7539921087326903221562638012600511281975432692021418185764672445524977206457320201696959933733708067724553969372336914900548677160248203107280132484232163449580273114090265675001571306136474727503648555307486531184035729106627013529123108800568069763608490199403396432102094680585721405059969950257096088964;
            6'd44: xpb[7] = 1024'd111585059824904056560593429282040513377117730580823884390381217905634121609936071851981600018882777444647296588857036927917917210821740766993164891392886806171962704686617104973366459264293588232030875589196977717237547969503345870279549890600494307981495118411208454234798306432725640242765383989996130915124;
            6'd45: xpb[7] = 1024'd91563502878356468500825293146666082727561601343890666466865908300766370676105684592251168889374172512126889800884243506356221903642012996323889525285210407960654461689572726934101108030933496015247905014699229056926699359679167954064998102717191096932561843208896454007387990110936926063352108203109571256953;
            6'd46: xpb[7] = 1024'd71541945931808880441057157011291652078005472106957448543350598695898619742275297332520737759865567579606483012911450084794526596462285225654614159177534009749346218692528348894835756797573403798464934440201480396615850749854990037850446314833887885883628568006584453779977673789148211883938832416223011598782;
            6'd47: xpb[7] = 1024'd51520388985261292381289020875917221428449342870024230619835289091030868808444910072790306630356962647086076224938656663232831289282557454985338793069857611538037975695483970855570405564213311581681963865703731736305002140030812121635894526950584674834695292804272453552567357467359497704525556629336451940611;
            6'd48: xpb[7] = 1024'd31498832038713704321520884740542790778893213633091012696319979486163117874614522813059875500848357714565669436965863241671135982102829684316063426962181213326729732698439592816305054330853219364898993291205983075994153530206634205421342739067281463785762017601960453325157041145570783525112280842449892282440;
            6'd49: xpb[7] = 1024'd11477275092166116261752748605168360129337084396157794772804669881295366940784135553329444371339752782045262648993069820109440674923101913646788060854504815115421489701395214777039703097493127148116022716708234415683304920382456289206790951183978252736828742399648453097746724823782069345699005055563332624269;
            6'd50: xpb[7] = 1024'd115522413829743269600783539874608362224479382284960260977421215341404511344262887203614084456488822158968005268477769833126809208584594477532672819763159457837803921273922054075404591055650240652643249750597725601736817160779175145957217732983904490954715370611453510900442936575921988183404419095302367450429;
            6'd51: xpb[7] = 1024'd95500856883195681541015403739233931574923253048027043053905905736536760410432499943883653326980217226447598480504976411565113901404866706863397453655483059626495678276877676036139239822290148435860279176099976941425968550954997229742665945100601279905782095409141510673032620254133274003991143308415807792258;
            6'd52: xpb[7] = 1024'd75479299936648093481247267603859500925367123811093825130390596131669009476602112684153222197471612293927191692532182990003418594225138936194122087547806661415187435279833297996873888588930056219077308601602228281115119941130819313528114157217298068856848820206829510445622303932344559824577867521529248134087;
            6'd53: xpb[7] = 1024'd55457742990100505421479131468485070275810994574160607206875286526801258542771725424422791067963007361406784904559389568441723287045411165524846721440130263203879192282788919957608537355569964002294338027104479620804271331306641397313562369333994857807915545004517510218211987610555845645164591734642688475916;
            6'd54: xpb[7] = 1024'd35436186043552917361710995333110639626254865337227389283359976921933507608941338164692359938454402428886378116586596146880027979865683394855571355332453864992570949285744541918343186122209871785511367452606730960493422721482463481099010581450691646758982269802205509990801671288767131465751315947756128817745;
            6'd55: xpb[7] = 1024'd15414629097005329301942859197736208976698736100294171359844667317065756675110950904961928808945797496365971328613802725318332672685955624186295989224777466781262706288700163879077834888849779568728396878108982300182574111658285564884458793567388435710048994599893509763391354966978417286338040160869569159574;
            6'd56: xpb[7] = 1024'd119459767834582482640973650467176211071841033989096637564461212777174901078589702555246568894094866873288713948098502738335701206347448188072180748133432109503645137861227003177442722847006893073255623911998473486236086352055004421634885575367314673927935622811698567566087566719118336124043454200608603985734;
            6'd57: xpb[7] = 1024'd99438210888034894581205514331801780422284904752163419640945903172307150144759315295516137764586261940768307160125709316774005899167720417402905382025755711292336894864182625138177371613646800856472653337500724825925237742230826505420333787484011462879002347609386567338677250397329621944630178413722044327563;
            6'd58: xpb[7] = 1024'd79416653941487306521437378196427349772728775515230201717430593567439399210928928035785706635077657008247900372152915895212310591987992646733630015918079313081028651867138247098912020380286708639689682763002976165614389132406648589205781999600708251830069072407074567111266934075540907765216902626835484669392;
            6'd59: xpb[7] = 1024'd59395096994939718461669242061052919123172646278296983793915283962571648277098540776055275505569052075727493584180122473650615284808264876064354649810402914869720408870093869059646669146926616422906712188505227505303540522582470672991230211717405040781135797204762566883856617753752193585803626839948925011221;
            6'd60: xpb[7] = 1024'd39373540048392130401901105925678488473616517041363765870399974357703897343268153516324844376060447143207086796207329052088919977628537105395079283702726516658412165873049491020381317913566524206123741614007478844992691912758292756776678423834101829732202522002450566656446301431963479406390351053062365353050;
            6'd61: xpb[7] = 1024'd19351983101844542342132969790304057824060387804430547946884664752836146409437766256594413246551842210686680008234535630527224670448809334725803917595050118447103922876005112981115966680206431989340771039509730184681843302934114840562126635950798618683269246800138566429035985110174765226977075266175805694879;
            6'd62: xpb[7] = 1024'd123397121839421695681163761059744059919202685693233014151501210212945290812916517906879053331700911587609422627719235643544593204110301898611688676503704761169486354448531952279480854638363545493867998073399221370735355543330833697312553417750724856901155875011943624231732196862314684064682489305914840521039;
            6'd63: xpb[7] = 1024'd103375564892874107621395624924369629269646556456299796227985900608077539879086130647148622202192306655089015839746442221982897896930574127942413310396028362958178111451487574240215503405003453277085027498901472710424506933506655781098001629867421645852222599809631624004321880540525969885269213519028280862868;
        endcase
    end

    always_comb begin
        case(flag[2][16:12])
            5'd0: xpb[8] = 1024'd0;
            5'd1: xpb[8] = 1024'd83354007946326519561627488788995198620090427219366578304470591003209788945255743387418191072683701722568609051773648800421202589750846357273137944288351964746869868454443196200950152171643361060302056924403724050113658323682477864883449841984118434803289324607319623776911564218737255705855937732141721204697;
            5'd2: xpb[8] = 1024'd42641320208528297724456050173175964495482427312997472480809326941442682553202347864821310930709729135694068696089804166263341338660472379991115763560372888560049062339315175064270065151769516399293916240420208253862955797144058956801921114285007420339758745800522189523716600363545878394593185637657847925063;
            5'd3: xpb[8] = 1024'd1928632470730075887284611557356730370874427406628366657148062879675576161148952342224430788735756548819528340405959532105480087570098402709093582832393812373228256224187153927589978131895671738285775556436692457612253270605640048720392386585896405876228166993724755270521636508354501083330433543173974645429;
            5'd4: xpb[8] = 1024'd85282640417056595448912100346351928990964854625994944961618653882885365106404695729642621861419458271388137392179608332526682677320944759982231527120745777120098124678630350128540130303539032798587832480840416507725911594288117913603842228570014840679517491601044379047433200727091756789186371275315695850126;
            5'd5: xpb[8] = 1024'd44569952679258373611740661730532694866356854719625839137957389821118258714351300207045741719445485684513597036495763698368821426230570782700209346392766700933277318563502328991860043283665188137579691796856900711475209067749699005522313500870903826215986912794246944794238236871900379477923619180831822570492;
            5'd6: xpb[8] = 1024'd3857264941460151774569223114713460741748854813256733314296125759351152322297904684448861577471513097639056680811919064210960175140196805418187165664787624746456512448374307855179956263791343476571551112873384915224506541211280097440784773171792811752456333987449510541043273016709002166660867086347949290858;
            5'd7: xpb[8] = 1024'd87211272887786671336196711903708659361839282032623311618766716762560941267553648071867052650155214820207665732585567864632162764891043162691325109953139589493326380902817504056130108435434704536873608037277108965338164864893757962324234615155911246555745658594769134317954837235446257872516804818489670495555;
            5'd8: xpb[8] = 1024'd46498585149988449499025273287889425237231282126254205795105452700793834875500252549270172508181242233333125376901723230474301513800669185409302929225160513306505574787689482919450021415560859875865467353293593169087462338355339054242705887456800232092215079787971700064759873380254880561254052724005797215921;
            5'd9: xpb[8] = 1024'd5785897412190227661853834672070191112623282219885099971444188639026728483446857026673292366207269646458585021217878596316440262710295208127280748497181437119684768672561461782769934395687015214857326669310077372836759811816920146161177159757689217628684500981174265811564909525063503249991300629521923936287;
            5'd10: xpb[8] = 1024'd89139905358516747223481323461065389732713709439251678275914779642236517428702600414091483438890971369027194072991527396737642852461141565400418692785533401866554637127004657983720086567330376275159383593713801422950418135499398011044627001741807652431973825588493889588476473743800758955847238361663645140984;
            5'd11: xpb[8] = 1024'd48427217620718525386309884845246155608105709532882572452253515580469411036649204891494603296916998782152653717307682762579781601370767588118396512057554325679733831011876636847039999547456531614151242909730285626699715608960979102963098274042696637968443246781696455335281509888609381644584486267179771861350;
            5'd12: xpb[8] = 1024'd7714529882920303549138446229426921483497709626513466628592251518702304644595809368897723154943026195278113361623838128421920350280393610836374331329575249492913024896748615710359912527582686953143102225746769830449013082422560194881569546343585623504912667974899021082086546033418004333321734172695898581716;
            5'd13: xpb[8] = 1024'd91068537829246823110765935018422120103588136845880044933062842521912093589851552756315914227626727917846722413397486928843122940031239968109512275617927214239782893351191811911310064699226048013445159150150493880562671406105038059765019388327704058308201992582218644858998110252155260039177671904837619786413;
            5'd14: xpb[8] = 1024'd50355850091448601273594496402602885978980136939510939109401578460144987197798157233719034085652755330972182057713642294685261688940865990827490094889948138052962087236063790774629977679352203352437018466166978084311968879566619151683490660628593043844671413775421210605803146396963882727914919810353746506779;
            5'd15: xpb[8] = 1024'd9643162353650379436423057786783651854372137033141833285740314398377880805744761711122153943678782744097641702029797660527400437850492013545467914161969061866141281120935769637949890659478358691428877782183462288061266353028200243601961932929482029381140834968623776352608182541772505416652167715869873227145;
            5'd16: xpb[8] = 1024'd92997170299976898998050546575778850474462564252508411590210905401587669751000505098540345016362484466666250753803446460948603027601338370818605858450321026613011149575378965838900042831121719751730934706587186338174924676710678108485411774913600464184430159575943400129519746760509761122508105448011594431842;
            5'd17: xpb[8] = 1024'd52284482562178677160879107959959616349854564346139305766549641339820563358947109575943464874388511879791710398119601826790741776510964393536583677722341950426190343460250944702219955811247875090722794022603670541924222150172259200403883047214489449720899580769145965876324782905318383811245353353527721152208;
            5'd18: xpb[8] = 1024'd11571794824380455323707669344140382225246564439770199942888377278053456966893714053346584732414539292917170042435757192632880525420590416254561496994362874239369537345122923565539868791374030429714653338620154745673519623633840292322354319515378435257369001962348531623129819050127006499982601259043847872574;
            5'd19: xpb[8] = 1024'd94925802770706974885335158133135580845336991659136778247358968281263245912149457440764775805098241015485779094209405993054083115171436773527699441282714838986239405799566119766490020963017391490016710263023878795787177947316318157205804161499496870060658326569668155400041383268864262205838538991185569077271;
            5'd20: xpb[8] = 1024'd54213115032908753048163719517316346720728991752767672423697704219496139520096061918167895663124268428611238738525561358896221864081062796245677260554735762799418599684438098629809933943143546829008569579040362999536475420777899249124275433800385855597127747762870721146846419413672884894575786896701695797637;
            5'd21: xpb[8] = 1024'd13500427295110531210992280901497112596120991846398566600036440157729033128042666395571015521150295841736698382841716724738360612990688818963655079826756686612597793569310077493129846923269702168000428895056847203285772894239480341042746706101274841133597168956073286893651455558481507583313034802217822518003;
            5'd22: xpb[8] = 1024'd96854435241437050772619769690492311216211419065765144904507031160938822073298409782989206593833997564305307434615365525159563202741535176236793024115108651359467662023753273694079999094913063228302485819460571253399431217921958205926196548085393275936886493563392910670563019777218763289168972534359543722700;
            5'd23: xpb[8] = 1024'd56141747503638828935448331074673077091603419159396039080845767099171715681245014260392326451860024977430767078931520891001701951651161198954770843387129575172646855908625252557399912075039218567294345135477055457148728691383539297844667820386282261473355914756595476417368055922027385977906220439875670443066;
            5'd24: xpb[8] = 1024'd15429059765840607098276892458853842966995419253026933257184503037404609289191618737795446309886052390556226723247676256843840700560787221672748662659150498985826049793497231420719825055165373906286204451493539660898026164845120389763139092687171247009825335949798042164173092066836008666643468345391797163432;
            5'd25: xpb[8] = 1024'd98783067712167126659904381247849041587085846472393511561655094040614398234447362125213637382569754113124835775021325057265043290311633578945886606947502463732695918247940427621669977226808734966588261375897263711011684488527598254646588934671289681813114660557117665941084656285573264372499406077533518368129;
            5'd26: xpb[8] = 1024'd58070379974368904822732942632029807462477846566024405737993829978847291842393966602616757240595781526250295419337480423107182039221259601663864426219523387545875112132812406484989890206934890305580120691913747914760981961989179346565060206972178667349584081750320231687889692430381887061236653983049645088495;
            5'd27: xpb[8] = 1024'd17357692236570682985561504016210573337869846659655299914332565917080185450340571080019877098621808939375755063653635788949320788130885624381842245491544311359054306017684385348309803187061045644571980007930232118510279435450760438483531479273067652886053502943522797434694728575190509749973901888565771808861;
            5'd28: xpb[8] = 1024'd100711700182897202547188992805205771957960273879021878218803156920289974395596314467438068171305510661944364115427284589370523377881731981654980189779896276105924174472127581549259955358704406704874036932333956168623937759133238303366981321257186087689342827550842421211606292793927765455829839620707493013558;
            5'd29: xpb[8] = 1024'd59999012445098980710017554189386537833352273972652772395141892858522868003542918944841188029331538075069823759743439955212662126791358004372958009051917199919103368356999560412579868338830562043865896248350440372373235232594819395285452593558075073225812248744044986958411328938736388144567087526223619733924;
            5'd30: xpb[8] = 1024'd19286324707300758872846115573567303708744274066283666571480628796755761611489523422244307887357565488195283404059595321054800875700984027090935828323938123732282562241871539275899781318956717382857755564366924576122532706056400487203923865858964058762281669937247552705216365083545010833304335431739746454290;
            5'd31: xpb[8] = 1024'd102640332653627278434473604362562502328834701285650244875951219799965550556745266809662498960041267210763892455833244121476003465451830384364073772612290088479152430696314735476849933490600078443159812488770648626236191029738878352087373707843082493565570994544567176482127929302282266539160273163881467658987;
        endcase
    end

    always_comb begin
        case(flag[3][5:0])
            6'd0: xpb[9] = 1024'd0;
            6'd1: xpb[9] = 1024'd92997170299976898998050546575778850474462564252508411590210905401587669751000505098540345016362484466666250753803446460948603027601338370818605858450321026613011149575378965838900042831121719751730934706587186338174924676710678108485411774913600464184430159575943400129519746760509761122508105448011594431842;
            6'd2: xpb[9] = 1024'd61927644915829056597302165746743268204226701379281139052289955738198444164691871287065618818067294623889352100149399487318142214361456407082051591884311012292331624581186714340169846470726233782151671804787132829985488503200459444005844980143971479102040415737769742228932965447090889227897521069397594379353;
            6'd3: xpb[9] = 1024'd30858119531681214196553784917707685933990838506053866514369006074809218578383237475590892619772104781112453446495352513687681401121574443345497325318300997971652099586994462841439650110330747812572408902987079321796052329690240779526278185374342494019650671899596084328346184133672017333286936690783594326864;
            6'd4: xpb[9] = 1024'd123855289831658113194604331493486536408453402758562278104579911476396888329383742574131237636134589247778704200298798974636284428722912814164103183768622024584663249162373428680339692941452467564303343609574265659970977006400918888011689960287942958204080831475539484457865930894181778455795042138795188758706;
            6'd5: xpb[9] = 1024'd92785764447510270793855950664450954138217539885335005566658961813007662743075108762656511437839399405001805546644752001005823615483030850427548917202612010263983724168181177181609496581056981594724080707774212151781540832890700223532123165518313973121691087637365826557279149580762906561184457760181188706217;
            6'd6: xpb[9] = 1024'd61716239063362428393107569835415371867981677012107733028738012149618437156766474951181785239544209562224906892990705027375362802243148886690994650636601995943304199173988925682879300220661495625144817805974158643592104659380481559052556370748684988039301343799192168656692368267344034666573873381567188653728;
            6'd7: xpb[9] = 1024'd30646713679214585992359189006379789597745814138880460490817062486229211570457841139707059041249019719448008239336658053744901989003266922954440384070591981622624674179796674184149103860266009655565554904174105135402668485870262894572989575979056002956911599961018510756105586953925162771963289002953188601239;
            6'd8: xpb[9] = 1024'd123643883979191484990409735582158640072208378391388872081027967887816881321458346238247404057611504186114258993140104514693505016604605293773046242520913008235635823755175640023049146691387729407296489610761291473577593162580941003058401350892656467141341759536961910885625333714434923894471394450964783033081;
            6'd9: xpb[9] = 1024'd92574358595043642589661354753123057801972515518161599543107018224427655735149712426772677859316314343337360339486057541063044203364723330036491975954902993914956298760983388524318950330992243437717226708961237965388156989070722338578834556123027482058952015698788252985038552401016051999860810072350782980592;
            6'd10: xpb[9] = 1024'd61504833210895800188912973924087475531736652644934327005186068561038430148841078615297951661021124500560461685832010567432583390124841366299937709388892979594276773766791137025588753970596757468137963807161184457198720815560503674099267761353398496976562271860614595084451771087597180105250225693736782928103;
            6'd11: xpb[9] = 1024'd30435307826747957788164593095051893261500789771707054467265118897649204562532444803823225462725934657783563032177963593802122576884959402563383442822882965273597248772598885526858557610201271498558700905361130949009284642050285009619700966583769511894172528022440937183864989774178308210639641315122782875614;
            6'd12: xpb[9] = 1024'd123432478126724856786215139670830743735963354024215466057476024299236874313532949902363570479088419124449813785981410054750725604486297773381989301273203991886608398347977851365758600441322991250289635611948317287184209318760963118105112741497369976078602687598384337313384736534688069333147746763134377307456;
            6'd13: xpb[9] = 1024'd92362952742577014385466758841795161465727491150988193519555074635847648727224316090888844280793229281672915132327363081120264791246415809645435034707193977565928873353785599867028404080927505280710372710148263778994773145250744453625545946727740990996212943760210679412797955221269197438537162384520377254967;
            6'd14: xpb[9] = 1024'd61293427358429171984718378012759579195491628277760920981634124972458423140915682279414118082498039438896016478673316107489803978006533845908880768141183963245249348359593348368298207720532019311131109808348210270805336971740525789145979151958112005913823199922037021512211173907850325543926578005906377202478;
            6'd15: xpb[9] = 1024'd30223901974281329583969997183723996925255765404533648443713175309069197554607048467939391884202849596119117825019269133859343164766651882172326501575173948924569823365401096869568011360136533341551846906548156762615900798230307124666412357188483020831433456083863363611624392594431453649315993627292377149989;
            6'd16: xpb[9] = 1024'd123221072274258228582020543759502847399718329657042060033924080710656867305607553566479736900565334062785368578822715594807946192367990252990932360025494975537580972940780062708468054191258253093282781613135343100790825474940985233151824132102083485015863615659806763741144139354941214771824099075303971581831;
            6'd17: xpb[9] = 1024'd92151546890110386181272162930467265129482466783814787496003131047267641719298919755005010702270144220008469925168668621177485379128108289254378093459484961216901447946587811209737857830862767123703518711335289592601389301430766568672257337332454499933473871821633105840557358041522342877213514696689971529342;
            6'd18: xpb[9] = 1024'd61082021505962543780523782101431682859246603910587514958082181383878416132990285943530284503974954377231571271514621647547024565888226325517823826893474946896221922952395559711007661470467281154124255809535236084411953127920547904192690542562825514851084127983459447939970576728103470982602930318075971476853;
            6'd19: xpb[9] = 1024'd30012496121814701379775401272396100589010741037360242420161231720489190546681652132055558305679764534454672617860574673916563752648344361781269560327464932575542397958203308212277465110071795184544992907735182576222516954410329239713123747793196529768694384145285790039383795414684599087992345939461971424364;
            6'd20: xpb[9] = 1024'd123009666421791600377825947848174951063473305289868654010372137122076860297682157230595903322042249001120923371664021134865166780249682732599875418777785959188553547533582274051177507941193514936275927614322368914397441631121007348198535522706796993953124543721229190168903542175194360210500451387473565856206;
            6'd21: xpb[9] = 1024'd91940141037643757977077567019139368793237442416641381472451187458687634711373523419121177123747059158344024718009974161234705967009800768863321152211775944867874022539390022552447311580798028966696664712522315406208005457610788683718968727937168008870734799883055532268316760861775488315889867008859565803717;
            6'd22: xpb[9] = 1024'd60870615653495915576329186190103786523001579543414108934530237795298409125064889607646450925451869315567126064355927187604245153769918805126766885645765930547194497545197771053717115220402542997117401810722261898018569284100570019239401933167539023788345056044881874367729979548356616421279282630245565751228;
            6'd23: xpb[9] = 1024'd29801090269348073175580805361068204252765716670186836396609288131909183538756255796171724727156679472790227410701880213973784340530036841390212619079755916226514972551005519554986918860007057027538138908922208389829133110590351354759835138397910038705955312206708216467143198234937744526668698251631565698739;
            6'd24: xpb[9] = 1024'd122798260569324972173631351936847054727228280922695247986820193533496853289756760894712069743519163939456478164505326674922387368131375212208818477530076942839526122126384485393886961691128776779269073615509394728004057787301029463245246913311510502890385471782651616596662944995447505649176803699643160130581;
            6'd25: xpb[9] = 1024'd91728735185177129772882971107811472456992418049467975448899243870107627703448127083237343545223974096679579510851279701291926554891493248472264210964066928518846597132192233895156765330733290809689810713709341219814621613790810798765680118541881517807995727944477958696076163682028633754566219321029160078092;
            6'd26: xpb[9] = 1024'd60659209801029287372134590278775890186756555176240702910978294206718402117139493271762617346928784253902680857197232727661465741651611284735709944398056914198167072137999982396426568970337804840110547811909287711625185440280592134286113323772252532725605984106304300795489382368609761859955634942415160025603;
            6'd27: xpb[9] = 1024'd29589684416881444971386209449740307916520692303013430373057344543329176530830859460287891148633594411125782203543185754031004928411729320999155677832046899877487547143807730897696372609942318870531284910109234203435749266770373469806546529002623547643216240268130642894902601055190889965345050563801159973114;
            6'd28: xpb[9] = 1024'd122586854716858343969436756025519158390983256555521841963268249944916846281831364558828236164996078877792032957346632214979607956013067691817761536282367926490498696719186696736596415441064038622262219616696420541610673943481051578291958303916224011827646399844074043024422347815700651087853156011812754404956;
            6'd29: xpb[9] = 1024'd91517329332710501568688375196483576120747393682294569425347300281527620695522730747353509966700889035015134303692585241349147142773185728081207269716357912169819171724994445237866219080668552652682956714896367033421237769970832913812391509146595026745256656005900385123835566502281779193242571633198754352467;
            6'd30: xpb[9] = 1024'd60447803948562659167939994367447993850511530809067296887426350618138395109214096935878783768405699192238235650038538267718686329533303764344653003150347897849139646730802193739136022720273066683103693813096313525231801596460614249332824714376966041662866912167726727223248785188862907298631987254584754299978;
            6'd31: xpb[9] = 1024'd29378278564414816767191613538412411580275667935840024349505400954749169522905463124404057570110509349461336996384491294088225516293421800608098736584337883528460121736609942240405826359877580713524430911296260017042365422950395584853257919607337056580477168329553069322662003875444035404021402875970754247489;
            6'd32: xpb[9] = 1024'd122375448864391715765242160114191262054738232188348435939716306356336839273905968222944402586472993816127587750187937755036828543894760171426704595034658910141471271311988908079305869190999300465255365617883446355217290099661073693338669694520937520764907327905496469452181750635953796526529508323982348679331;
            6'd33: xpb[9] = 1024'd91305923480243873364493779285155679784502369315121163401795356692947613687597334411469676388177803973350689096533890781406367730654878207690150328468648895820791746317796656580575672830603814495676102716083392847027853926150855028859102899751308535682517584067322811551594969322534924631918923945368348626842;
            6'd34: xpb[9] = 1024'd60236398096096030963745398456120097514266506441893890863874407029558388101288700599994950189882614130573790442879843807775906917414996243953596061902638881500112221323604405081845476470208328526096839814283339338838417752640636364379536104981679550600127840229149153651008188009116052737308339566754348574353;
            6'd35: xpb[9] = 1024'd29166872711948188562997017627084515244030643568666618325953457366169162514980066788520223991587424287796891789225796834145446104175114280217041795336628867179432696329412153583115280109812842556517576912483285830648981579130417699899969310212050565517738096390975495750421406695697180842697755188140348521864;
            6'd36: xpb[9] = 1024'd122164043011925087561047564202863365718493207821175029916164362767756832265980571887060569007949908754463142543029243295094049131776452651035647653786949893792443845904791119422015322940934562308248511619070472168823906255841095808385381085125651029702168255966918895879941153456206941965205860636151942953706;
            6'd37: xpb[9] = 1024'd91094517627777245160299183373827783448257344947947757378243413104367606679671938075585842809654718911686243889375196321463588318536570687299093387220939879471764320910598867923285126580539076338669248717270418660634470082330877143905814290356022044619778512128745237979354372142788070070595276257537942901217;
            6'd38: xpb[9] = 1024'd60024992243629402759550802544792201178021482074720484840322463440978381093363304264111116611359529068909345235721149347833127505296688723562539120654929865151084795916406616424554930220143590369089985815470365152445033908820658479426247495586393059537388768290571580078767590829369198175984691878923942848728;
            6'd39: xpb[9] = 1024'd28955466859481560358802421715756618907785619201493212302401513777589155507054670452636390413064339226132446582067102374202666692056806759825984854088919850830405270922214364925824733859748104399510722913670311644255597735310439814946680700816764074454999024452397922178180809515950326281374107500309942796239;
            6'd40: xpb[9] = 1024'd121952637159458459356852968291535469382248183454001623892612419179176825258055175551176735429426823692798697335870548835151269719658145130644590712539240877443416420497593330764724776690869824151241657620257497982430522412021117923432092475730364538639429184028341322307700556276460087403882212948321537228081;
            6'd41: xpb[9] = 1024'd90883111775310616956104587462499887112012320580774351354691469515787599671746541739702009231131633850021798682216501861520808906418263166908036445973230863122736895503401079265994580330474338181662394718457444474241086238510899258952525680960735553557039440190167664407113774963041215509271628569707537175592;
            6'd42: xpb[9] = 1024'd59813586391162774555356206633464304841776457707547078816770519852398374085437907928227283032836444007244900028562454887890348093178381203171482179407220848802057370509208827767264383970078852212083131816657390966051650065000680594472958886191106568474649696351994006506526993649622343614661044191093537123103;
            6'd43: xpb[9] = 1024'd28744061007014932154607825804428722571540594834319806278849570189009148499129274116752556834541254164468001374908407914259887279938499239434927912841210834481377845515016576268534187609683366242503868914857337457862213891490461929993392091421477583392259952513820348605940212336203471720050459812479537070614;
            6'd44: xpb[9] = 1024'd121741231306991831152658372380207573046003159086828217869060475590596818250129779215292901850903738631134252128711854375208490307539837610253533771291531861094388995090395542107434230440805085994234803621444523796037138568201140038478803866335078047576690112089763748735459959096713232842558565260491131502456;
            6'd45: xpb[9] = 1024'd90671705922843988751909991551171990775767296213600945331139525927207592663821145403818175652608548788357353475057807401578029494299955646516979504725521846773709470096203290608704034080409600024655540719644470287847702394690921373999237071565449062494300368251590090834873177783294360947947980881877131449967;
            6'd46: xpb[9] = 1024'd59602180538696146351161610722136408505531433340373672793218576263818367077512511592343449454313358945580454821403760427947568681060073682780425238159511832453029945102011039109973837720014114055076277817844416779658266221180702709519670276795820077411910624413416432934286396469875489053337396503263131397478;
            6'd47: xpb[9] = 1024'd28532655154548303950413229893100826235295570467146400255297626600429141491203877780868723256018169102803556167749713454317107867820191719043870971593501818132350420107818787611243641359618628085497014916044363271468830047670484045040103482026191092329520880575242775033699615156456617158726812124649131344989;
            6'd48: xpb[9] = 1024'd121529825454525202948463776468879676709758134719654811845508532002016811242204382879409068272380653569469806921553159915265710895421530089862476830043822844745361569683197753450143684190740347837227949622631549609643754724381162153525515256939791556513951040151186175163219361916966378281234917572660725776831;
            6'd49: xpb[9] = 1024'd90460300070377360547715395639844094439522271846427539307587582338627585655895749067934342074085463726692908267899112941635250082181648126125922563477812830424682044689005501951413487830344861867648686720831496101454318550870943489045948462170162571431561296313012517262632580603547506386624333194046725724342;
            6'd50: xpb[9] = 1024'd59390774686229518146967014810808512169286408973200266769666632675238360069587115256459615875790273883916009614245065968004789268941766162389368296911802816104002519694813250452683291469949375898069423819031442593264882377360724824566381667400533586349171552474838859362045799290128634492013748815432725671853;
            6'd51: xpb[9] = 1024'd28321249302081675746218633981772929899050546099972994231745683011849134483278481444984889677495084041139110960591018994374328455701884198652814030345792801783322994700620998953953095109553889928490160917231389085075446203850506160086814872630904601266781808636665201461459017976709762597403164436818725619364;
            6'd52: xpb[9] = 1024'd121318419602058574744269180557551780373513110352481405821956588413436804234278986543525234693857568507805361714394465455322931483303222569471419888796113828396334144275999964792853137940675609680221095623818575423250370880561184268572226647544505065451211968212608601590978764737219523719911269884830320051206;
            6'd53: xpb[9] = 1024'd90248894217910732343520799728516198103277247479254133284035638750047578647970352732050508495562378665028463060740418481692470670063340605734865622230103814075654619281807713294122941580280123710641832722018521915060934707050965604092659852774876080368822224374434943690391983423800651825300685506216319998717;
            6'd54: xpb[9] = 1024'd59179368833762889942772418899480615833041384606026860746114689086658353061661718920575782297267188822251564407086371508062009856823458641998311355664093799754975094287615461795392745219884637741062569820218468406871498533540746939613093058005247095286432480536261285789805202110381779930690101127602319946228;
            6'd55: xpb[9] = 1024'd28109843449615047542024038070445033562805521732799588208193739423269127475353085109101056098971998979474665753432324534431549043583576678261757089098083785434295569293423210296662548859489151771483306918418414898682062360030528275133526263235618110204042736698087627889218420796962908036079516748988319893739;
            6'd56: xpb[9] = 1024'd121107013749591946540074584646223884037268085985307999798404644824856797226353590207641401115334483446140916507235770995380152071184915049080362947548404812047306718868802176135562591690610871523214241625005601236856987036741206383618938038149218574388472896274031028018738167557472669158587622196999914325581;
            6'd57: xpb[9] = 1024'd90037488365444104139326203817188301767032223112080727260483695161467571640044956396166674917039293603364017853581724021749691257945033085343808680982394797726627193874609924636832395330215385553634978723205547728667550863230987719139371243379589589306083152435857370118151386244053797263977037818385914273092;
            6'd58: xpb[9] = 1024'd58967962981296261738577822988152719496796360238853454722562745498078346053736322584691948718744103760587119199927677048119230444705151121607254414416384783405947668880417673138102198969819899584055715821405494220478114689720769054659804448609960604223693408597683712217564604930634925369366453439771914220603;
            6'd59: xpb[9] = 1024'd27898437597148419337829442159117137226560497365626182184641795834689120467427688773217222520448913917810220546273630074488769631465269157870700147850374769085268143886225421639372002609424413614476452919605440712288678516210550390180237653840331619141303664759510054316977823617216053474755869061157914168114;
            6'd60: xpb[9] = 1024'd120895607897125318335879988734895987701023061618134593774852701236276790218428193871757567536811398384476471300077076535437372659066607528689306006300695795698279293461604387478272045440546133366207387626192627050463603192921228498665649428753932083325733824335453454446497570377725814597263974509169508599956;
            6'd61: xpb[9] = 1024'd89826082512977475935131607905860405430787198744907321236931751572887564632119560060282841338516208541699572646423029561806911845826725564952751739734685781377599768467412135979541849080150647396628124724392573542274167019411009834186082633984303098243344080497279796545910789064306942702653390130555508547467;
            6'd62: xpb[9] = 1024'd58756557128829633534383227076824823160551335871680048699010801909498339045810926248808115140221018698922673992768982588176451032586843601216197473168675767056920243473219884480811652719755161427048861822592520034084730845900791169706515839214674113160954336659106138645324007750888070808042805751941508494978;
            6'd63: xpb[9] = 1024'd27687031744681791133634846247789240890315472998452776161089852246109113459502292437333388941925828856145775339114935614545990219346961637479643206602665752736240718479027632982081456359359675457469598920792466525895294672390572505226949044445045128078564592820932480744737226437469198913432221373327508442489;
        endcase
    end

    always_comb begin
        case(flag[3][11:6])
            6'd0: xpb[10] = 1024'd0;
            6'd1: xpb[10] = 1024'd120684202044658690131685392823568091364778037250961187751300757647696783210502797535873733958288313322812026092918382075494593246948300008298249065052986779349251868054406598820981499190481395209200533627379652864070219349101250613712360819358645592262994752396875880874256973197978960035940326821339102874331;
            6'd2: xpb[10] = 1024'd117301708405192638864571858242321749984857647376186691374469660230416671083696456161732396701918952336180902778379270716410122653055379682041338005089642517764813061539241980304332759189445584697090869646372065881776077847981604454459743069034061735259169601379634703718407418322029287054761963816052611264331;
            6'd3: xpb[10] = 1024'd113919214765726587597458323661075408604937257501412194997638562813136558956890114787591059445549591349549779463840159357325652059162459355784426945126298256180374255024077361787684019188409774184981205665364478899481936346861958295207125318709477878255344450362393526562557863446079614073583600810766119654331;
            6'd4: xpb[10] = 1024'd110536721126260536330344789079829067225016867626637698620807465395856446830083773413449722189180230362918656149301047998241181465269539029527515885162953994595935448508912743271035279187373963672871541684356891917187794845742312135954507568384894021251519299345152349406708308570129941092405237805479628044331;
            6'd5: xpb[10] = 1024'd107154227486794485063231254498582725845096477751863202243976367978576334703277432039308384932810869376287532834761936639156710871376618703270604825199609733011496641993748124754386539186338153160761877703349304934893653344622665976701889818060310164247694148327911172250858753694180268111226874800193136434331;
            6'd6: xpb[10] = 1024'd103771733847328433796117719917336384465176087877088705867145270561296222576471090665167047676441508389656409520222825280072240277483698377013693765236265471427057835478583506237737799185302342648652213722341717952599511843503019817449272067735726307243868997310669995095009198818230595130048511794906644824331;
            6'd7: xpb[10] = 1024'd100389240207862382529004185336090043085255698002314209490314173144016110449664749291025710420072147403025286205683713920987769683590778050756782705272921209842619028963418887721089059184266532136542549741334130970305370342383373658196654317411142450240043846293428817939159643942280922148870148789620153214331;
            6'd8: xpb[10] = 1024'd97006746568396331261890650754843701705335308127539713113483075726735998322858407916884373163702786416394162891144602561903299089697857724499871645309576948258180222448254269204440319183230721624432885760326543988011228841263727498944036567086558593236218695276187640783310089066331249167691785784333661604331;
            6'd9: xpb[10] = 1024'd93624252928930279994777116173597360325414918252765216736651978309455886196052066542743035907333425429763039576605491202818828495804937398242960585346232686673741415933089650687791579182194911112323221779318957005717087340144081339691418816761974736232393544258946463627460534190381576186513422779047169994331;
            6'd10: xpb[10] = 1024'd90241759289464228727663581592351018945494528377990720359820880892175774069245725168601698650964064443131916262066379843734357901912017071986049525382888425089302609417925032171142839181159100600213557798311370023422945839024435180438801066437390879228568393241705286471610979314431903205335059773760678384331;
            6'd11: xpb[10] = 1024'd86859265649998177460550047011104677565574138503216223982989783474895661942439383794460361394594703456500792947527268484649887308019096745729138465419544163504863802902760413654494099180123290088103893817303783041128804337904789021186183316112807022224743242224464109315761424438482230224156696768474186774331;
            6'd12: xpb[10] = 1024'd83476772010532126193436512429858336185653748628441727606158686057615549815633042420319024138225342469869669632988157125565416714126176419472227405456199901920424996387595795137845359179087479575994229836296196058834662836785142861933565565788223165220918091207222932159911869562532557242978333763187695164331;
            6'd13: xpb[10] = 1024'd80094278371066074926322977848611994805733358753667231229327588640335437688826701046177686881855981483238546318449045766480946120233256093215316345492855640335986189872431176621196619178051669063884565855288609076540521335665496702680947815463639308217092940189981755004062314686582884261799970757901203554331;
            6'd14: xpb[10] = 1024'd76711784731600023659209443267365653425812968878892734852496491223055325562020359672036349625486620496607423003909934407396475526340335766958405285529511378751547383357266558104547879177015858551774901874281022094246379834545850543428330065139055451213267789172740577848212759810633211280621607752614711944331;
            6'd15: xpb[10] = 1024'd73329291092133972392095908686119312045892579004118238475665393805775213435214018297895012369117259509976299689370823048312004932447415440701494225566167117167108576842101939587899139175980048039665237893273435111952238333426204384175712314814471594209442638155499400692363204934683538299443244747328220334331;
            6'd16: xpb[10] = 1024'd69946797452667921124982374104872970665972189129343742098834296388495101308407676923753675112747898523345176374831711689227534338554495114444583165602822855582669770326937321071250399174944237527555573912265848129658096832306558224923094564489887737205617487138258223536513650058733865318264881742041728724331;
            6'd17: xpb[10] = 1024'd66564303813201869857868839523626629286051799254569245722003198971214989181601335549612337856378537536714053060292600330143063744661574788187672105639478593998230963811772702554601659173908427015445909931258261147363955331186912065670476814165303880201792336121017046380664095182784192337086518736755237114331;
            6'd18: xpb[10] = 1024'd63181810173735818590755304942380287906131409379794749345172101553934877054794994175471000600009176550082929745753488971058593150768654461930761045676134332413792157296608084037952919172872616503336245950250674165069813830067265906417859063840720023197967185103775869224814540306834519355908155731468745504331;
            6'd19: xpb[10] = 1024'd59799316534269767323641770361133946526211019505020252968341004136654764927988652801329663343639815563451806431214377611974122556875734135673849985712790070829353350781443465521304179171836805991226581969243087182775672328947619747165241313516136166194142034086534692068964985430884846374729792726182253894331;
            6'd20: xpb[10] = 1024'd56416822894803716056528235779887605146290629630245756591509906719374652801182311427188326087270454576820683116675266252889651962982813809416938925749445809244914544266278847004655439170800995479116917988235500200481530827827973587912623563191552309190316883069293514913115430554935173393551429720895762284331;
            6'd21: xpb[10] = 1024'd53034329255337664789414701198641263766370239755471260214678809302094540674375970053046988830901093590189559802136154893805181369089893483160027865786101547660475737751114228488006699169765184967007254007227913218187389326708327428660005812866968452186491732052052337757265875678985500412373066715609270674331;
            6'd22: xpb[10] = 1024'd49651835615871613522301166617394922386449849880696763837847711884814428547569628678905651574531732603558436487597043534720710775196973156903116805822757286076036931235949609971357959168729374454897590026220326235893247825588681269407388062542384595182666581034811160601416320803035827431194703710322779064331;
            6'd23: xpb[10] = 1024'd46269341976405562255187632036148581006529460005922267461016614467534316420763287304764314318162371616927313173057932175636240181304052830646205745859413024491598124720784991454709219167693563942787926045212739253599106324469035110154770312217800738178841430017569983445566765927086154450016340705036287454331;
            6'd24: xpb[10] = 1024'd42886848336939510988074097454902239626609070131147771084185517050254204293956945930622977061793010630296189858518820816551769587411132504389294685896068762907159318205620372938060479166657753430678262064205152271304964823349388950902152561893216881175016279000328806289717211051136481468837977699749795844331;
            6'd25: xpb[10] = 1024'd39504354697473459720960562873655898246688680256373274707354419632974092167150604556481639805423649643665066543979709457467298993518212178132383625932724501322720511690455754421411739165621942918568598083197565289010823322229742791649534811568633024171191127983087629133867656175186808487659614694463304234331;
            6'd26: xpb[10] = 1024'd36121861058007408453847028292409556866768290381598778330523322215693980040344263182340302549054288657033943229440598098382828399625291851875472565969380239738281705175291135904762999164586132406458934102189978306716681821110096632396917061244049167167365976965846451978018101299237135506481251689176812624331;
            6'd27: xpb[10] = 1024'd32739367418541357186733493711163215486847900506824281953692224798413867913537921808198965292684927670402819914901486739298357805732371525618561506006035978153842898660126517388114259163550321894349270121182391324422540319990450473144299310919465310163540825948605274822168546423287462525302888683890321014331;
            6'd28: xpb[10] = 1024'd29356873779075305919619959129916874106927510632049785576861127381133755786731580434057628036315566683771696600362375380213887211839451199361650446042691716569404092144961898871465519162514511382239606140174804342128398818870804313891681560594881453159715674931364097666318991547337789544124525678603829404331;
            6'd29: xpb[10] = 1024'd25974380139609254652506424548670532727007120757275289200030029963853643659925239059916290779946205697140573285823264021129416617946530873104739386079347454984965285629797280354816779161478700870129942159167217359834257317751158154639063810270297596155890523914122920510469436671388116562946162673317337794331;
            6'd30: xpb[10] = 1024'd22591886500143203385392889967424191347086730882500792823198932546573531533118897685774953523576844710509449971284152662044946024053610546847828326116003193400526479114632661838168039160442890358020278178159630377540115816631511995386446059945713739152065372896881743354619881795438443581767799668030846184331;
            6'd31: xpb[10] = 1024'd19209392860677152118279355386177849967166341007726296446367835129293419406312556311633616267207483723878326656745041302960475430160690220590917266152658931816087672599468043321519299159407079845910614197152043395245974315511865836133828309621129882148240221879640566198770326919488770600589436662744354574331;
            6'd32: xpb[10] = 1024'd15826899221211100851165820804931508587245951132951800069536737712013307279506214937492279010838122737247203342205929943876004836267769894334006206189314670231648866084303424804870559158371269333800950216144456412951832814392219676881210559296546025144415070862399389042920772043539097619411073657457862964331;
            6'd33: xpb[10] = 1024'd12444405581745049584052286223685167207325561258177303692705640294733195152699873563350941754468761750616080027666818584791534242374849568077095146225970408647210059569138806288221819157335458821691286235136869430657691313272573517628592808971962168140589919845158211887071217167589424638232710652171371354331;
            6'd34: xpb[10] = 1024'd9061911942278998316938751642438825827405171383402807315874542877453083025893532189209604498099400763984956713127707225707063648481929241820184086262626147062771253053974187771573079156299648309581622254129282448363549812152927358375975058647378311136764768827917034731221662291639751657054347646884879744331;
            6'd35: xpb[10] = 1024'd5679418302812947049825217061192484447484781508628310939043445460172970899087190815068267241730039777353833398588595866622593054589008915563273026299281885478332446538809569254924339155263837797471958273121695466069408311033281199123357308322794454132939617810675857575372107415690078675875984641598388134331;
            6'd36: xpb[10] = 1024'd2296924663346895782711682479946143067564391633853814562212348042892858772280849440926929985360678790722710084049484507538122460696088589306361966335937623893893640023644950738275599154228027285362294292114108483775266809913635039870739557998210597129114466793434680419522552539740405694697621636311896524331;
            6'd37: xpb[10] = 1024'd122981126708005585914397075303514234432342428884815002313513105690589641982783646976800663943648992113534736176967866583032715707644388597604611031388924403243145508078051549559257098344709422494562827919493761347845486159014885653583100377356856189392109219190310561293779525737719365730637948457650999398662;
            6'd38: xpb[10] = 1024'd119598633068539534647283540722267893052422039010040505936682008273309529855977305602659326687279631126903612862428755223948245113751468271347699971425580141658706701562886931042608358343673611982453163938486174365551344657895239494330482627032272332388284068173069384137929970861769692749459585452364507788662;
            6'd39: xpb[10] = 1024'd116216139429073483380170006141021551672501649135266009559850910856029417729170964228517989430910270140272489547889643864863774519858547945090788911462235880074267895047722312525959618342637801470343499957478587383257203156775593335077864876707688475384458917155828206982080415985820019768281222447078016178662;
            6'd40: xpb[10] = 1024'd112833645789607432113056471559775210292581259260491513183019813438749305602364622854376652174540909153641366233350532505779303925965627618833877851498891618489829088532557694009310878341601990958233835976471000400963061655655947175825247126383104618380633766138587029826230861109870346787102859441791524568662;
            6'd41: xpb[10] = 1024'd109451152150141380845942936978528868912660869385717016806188716021469193475558281480235314918171548167010242918811421146694833332072707292576966791535547356905390282017393075492662138340566180446124171995463413418668920154536301016572629376058520761376808615121345852670381306233920673805924496436505032958662;
            6'd42: xpb[10] = 1024'd106068658510675329578829402397282527532740479510942520429357618604189081348751940106093977661802187180379119604272309787610362738179786966320055731572203095320951475502228456976013398339530369934014508014455826436374778653416654857320011625733936904372983464104104675514531751357971000824746133431218541348662;
            6'd43: xpb[10] = 1024'd102686164871209278311715867816036186152820089636168024052526521186908969221945598731952640405432826193747996289733198428525892144286866640063144671608858833736512668987063838459364658338494559421904844033448239454080637152297008698067393875409353047369158313086863498358682196482021327843567770425932049738662;
            6'd44: xpb[10] = 1024'd99303671231743227044602333234789844772899699761393527675695423769628857095139257357811303149063465207116872975194087069441421550393946313806233611645514572152073862471899219942715918337458748909795180052440652471786495651177362538814776125084769190365333162069622321202832641606071654862389407420645558128662;
            6'd45: xpb[10] = 1024'd95921177592277175777488798653543503392979309886619031298864326352348744968332915983669965892694104220485749660654975710356950956501025987549322551682170310567635055956734601426067178336422938397685516071433065489492354150057716379562158374760185333361508011052381144046983086730121981881211044415359066518662;
            6'd46: xpb[10] = 1024'd92538683952811124510375264072297162013058920011844534922033228935068632841526574609528628636324743233854626346115864351272480362608105661292411491718826048983196249441569982909418438335387127885575852090425478507198212648938070220309540624435601476357682860035139966891133531854172308900032681410072574908662;
            6'd47: xpb[10] = 1024'd89156190313345073243261729491050820633138530137070038545202131517788520714720233235387291379955382247223503031576752992188009768715185335035500431755481787398757442926405364392769698334351317373466188109417891524904071147818424061056922874111017619353857709017898789735283976978222635918854318404786083298662;
            6'd48: xpb[10] = 1024'd85773696673879021976148194909804479253218140262295542168371034100508408587913891861245954123586021260592379717037641633103539174822265008778589371792137525814318636411240745876120958333315506861356524128410304542609929646698777901804305123786433762350032558000657612579434422102272962937675955399499591688662;
            6'd49: xpb[10] = 1024'd82391203034412970709034660328558137873297750387521045791539936683228296461107550487104616867216660273961256402498530274019068580929344682521678311828793264229879829896076127359472218332279696349246860147402717560315788145579131742551687373461849905346207406983416435423584867226323289956497592394213100078662;
            6'd50: xpb[10] = 1024'd79008709394946919441921125747311796493377360512746549414708839265948184334301209112963279610847299287330133087959418914934597987036424356264767251865449002645441023380911508842823478331243885837137196166395130578021646644459485583299069623137266048342382255966175258267735312350373616975319229388926608468662;
            6'd51: xpb[10] = 1024'd75626215755480868174807591166065455113456970637972053037877741848668072207494867738821942354477938300699009773420307555850127393143504030007856191902104741061002216865746890326174738330208075325027532185387543595727505143339839424046451872812682191338557104948934081111885757474423943994140866383640116858662;
            6'd52: xpb[10] = 1024'd72243722116014816907694056584819113733536580763197556661046644431387960080688526364680605098108577314067886458881196196765656799250583703750945131938760479476563410350582271809525998329172264812917868204379956613433363642220193264793834122488098334334731953931692903956036202598474271012962503378353625248662;
            6'd53: xpb[10] = 1024'd68861228476548765640580522003572772353616190888423060284215547014107847953882184990539267841739216327436763144342084837681186205357663377494034071975416217892124603835417653292877258328136454300808204223372369631139222141100547105541216372163514477330906802914451726800186647722524598031784140373067133638662;
            6'd54: xpb[10] = 1024'd65478734837082714373466987422326430973695801013648563907384449596827735827075843616397930585369855340805639829802973478596715611464743051237123012012071956307685797320253034776228518327100643788698540242364782648845080639980900946288598621838930620327081651897210549644337092846574925050605777367780642028662;
            6'd55: xpb[10] = 1024'd62096241197616663106353452841080089593775411138874067530553352179547623700269502242256593329000494354174516515263862119512245017571822724980211952048727694723246990805088416259579778326064833276588876261357195666550939138861254787035980871514346763323256500879969372488487537970625252069427414362494150418662;
            6'd56: xpb[10] = 1024'd58713747558150611839239918259833748213855021264099571153722254762267511573463160868115256072631133367543393200724750760427774423678902398723300892085383433138808184289923797742931038325029022764479212280349608684256797637741608627783363121189762906319431349862728195332637983094675579088249051357207658808662;
            6'd57: xpb[10] = 1024'd55331253918684560572126383678587406833934631389325074776891157344987399446656819493973918816261772380912269886185639401343303829785982072466389832122039171554369377774759179226282298323993212252369548299342021701962656136621962468530745370865179049315606198845487018176788428218725906107070688351921167198662;
            6'd58: xpb[10] = 1024'd51948760279218509305012849097341065454014241514550578400060059927707287319850478119832581559892411394281146571646528042258833235893061746209478772158694909969930571259594560709633558322957401740259884318334434719668514635502316309278127620540595192311781047828245841020938873342776233125892325346634675588662;
            6'd59: xpb[10] = 1024'd48566266639752458037899314516094724074093851639776082023228962510427175193044136745691244303523050407650023257107416683174362642000141419952567712195350648385491764744429942192984818321921591228150220337326847737374373134382670150025509870216011335307955896811004663865089318466826560144713962341348183978662;
            6'd60: xpb[10] = 1024'd45183773000286406770785779934848382694173461765001585646397865093147063066237795371549907047153689421018899942568305324089892048107221093695656652232006386801052958229265323676336078320885780716040556356319260755080231633263023990772892119891427478304130745793763486709239763590876887163535599336061692368662;
            6'd61: xpb[10] = 1024'd41801279360820355503672245353602041314253071890227089269566767675866950939431453997408569790784328434387776628029193965005421454214300767438745592268662125216614151714100705159687338319849970203930892375311673772786090132143377831520274369566843621300305594776522309553390208714927214182357236330775200758662;
            6'd62: xpb[10] = 1024'd38418785721354304236558710772355699934332682015452592892735670258586838812625112623267232534414967447756653313490082605920950860321380441181834532305317863632175345198936086643038598318814159691821228394304086790491948631023731672267656619242259764296480443759281132397540653838977541201178873325488709148662;
            6'd63: xpb[10] = 1024'd35036292081888252969445176191109358554412292140678096515904572841306726685818771249125895278045606461125529998950971246836480266428460114924923472341973602047736538683771468126389858317778349179711564413296499808197807129904085513015038868917675907292655292742039955241691098963027868220000510320202217538662;
        endcase
    end

    always_comb begin
        case(flag[3][16:12])
            5'd0: xpb[11] = 1024'd0;
            5'd1: xpb[11] = 1024'd31653798442422201702331641609863017174491902265903600139073475424026614559012429874984558021676245474494406684411859887752009672535539788668012412378629340463297732168606849609741118316742538667601900432288912825903665628784439353762421118593092050288830141724798778085841544087078195238822147314915725928662;
            5'd2: xpb[11] = 1024'd63307596884844403404663283219726034348983804531807200278146950848053229118024859749969116043352490948988813368823719775504019345071079577336024824757258680926595464337213699219482236633485077335203800864577825651807331257568878707524842237186184100577660283449597556171683088174156390477644294629831451857324;
            5'd3: xpb[11] = 1024'd94961395327266605106994924829589051523475706797710800417220426272079843677037289624953674065028736423483220053235579663256029017606619366004037237135888021389893196505820548829223354950227616002805701296866738477710996886353318061287263355779276150866490425174396334257524632261234585716466441944747177785986;
            5'd4: xpb[11] = 1024'd2548498085564065410527639034637635953269181937878716428162046631129562898740580589923160872047307588534477330189946116428974849300938820116889524498186320919500254104856181101334234075452948949097404120768411457250301664916860642084705904689138751888500663485078054313259648274384147938169899433037309230317;
            5'd5: xpb[11] = 1024'd34202296527986267112859280644500653127761084203782316567235522055156177457753010464907718893723553063028884014601806004180984521836478608784901936876815661382797986273463030711075352392195487616699304553057324283153967293701299995847127023282230802177330805209876832399101192361462343176992046747953035158979;
            5'd6: xpb[11] = 1024'd65856094970408468815190922254363670302252986469685916706308997479182792016765440339892276915399798537523290699013665891932994194372018397452914349255445001846095718442069880320816470708938026284301204985346237109057632922485739349609548141875322852466160946934675610484942736448540538415814194062868761087641;
            5'd7: xpb[11] = 1024'd97509893412830670517522563864226687476744888735589516845382472903209406575777870214876834937076044012017697383425525779685003866907558186120926761634074342309393450610676729930557589025680564951903105417635149934961298551270178703371969260468414902754991088659474388570784280535618733654636341377784487016303;
            5'd8: xpb[11] = 1024'd5096996171128130821055278069275271906538363875757432856324093262259125797481161179846321744094615177068954660379892232857949698601877640233779048996372641839000508209712362202668468150905897898194808241536822914500603329833721284169411809378277503777001326970156108626519296548768295876339798866074618460634;
            5'd9: xpb[11] = 1024'd36750794613550332523386919679138289081030266141661032995397568686285740356493591054830879765770860651563361344791752120609959371137417428901791461375001982302298240378319211812409586467648436565796708673825735740404268958618160637931832927971369554065831468694954886712360840635846491115161946180990344389296;
            5'd10: xpb[11] = 1024'd68404593055972534225718561289001306255522168407564633134471044110312354915506020929815437787447106126057768029203612008361969043672957217569803873753631322765595972546926061422150704784390975233398609106114648566307934587402599991694254046564461604354661610419753664798202384722924686353984093495906070317958;
            5'd11: xpb[11] = 1024'd100058391498394735928050202898864323430014070673468233273544519534338969474518450804799995809123351600552174713615471896113978716208497006237816286132260663228893704715532911031891823101133513901000509538403561392211600216187039345456675165157553654643491752144552442884043928810002881592806240810821796246620;
            5'd12: xpb[11] = 1024'd7645494256692196231582917103912907859807545813636149284486139893388688696221741769769482616141922765603431990569838349286924547902816460350668573494558962758500762314568543304002702226358846847292212362305234371750904994750581926254117714067416255665501990455234162939778944823152443814509698299111927690951;
            5'd13: xpb[11] = 1024'd39299292699114397933914558713775925034299448079539749423559615317415303255234171644754040637818168240097838674981698237038934220438356249018680985873188303221798494483175392913743820543101385514894112794594147197654570623535021280016538832660508305954332132180032941025620488910230639053331845614027653619613;
            5'd14: xpb[11] = 1024'd70953091141536599636246200323638942208791350345443349562633090741441917814246601519738598659494413714592245359393558124790943892973896037686693398251817643685096226651782242523484938859843924182496013226883060023558236252319460633778959951253600356243162273904831719111462032997308834292153992928943379548275;
            5'd15: xpb[11] = 1024'd102606889583958801338577841933501959383283252611346949701706566165468532373259031394723156681170659189086652043805418012542953565509435826354705810630446984148393958820389092133226057176586462850097913659171972849461901881103899987541381069846692406531992415629630497197303577084387029530976140243859105476937;
            5'd16: xpb[11] = 1024'd10193992342256261642110556138550543813076727751514865712648186524518251594962322359692643488189230354137909320759784465715899397203755280467558097992745283678001016419424724405336936301811795796389616483073645829001206659667442568338823618756555007554002653940312217253038593097536591752679597732149236921268;
            5'd17: xpb[11] = 1024'd41847790784678463344442197748413560987568630017418465851721661948544866153974752234677201509865475828632316005171644353467909069739295069135570510371374624141298748588031574015078054618554334463991516915362558654904872288451881922101244737349647057842832795665110995338880137184614786991501745047064962849930;
            5'd18: xpb[11] = 1024'd73501589227100665046773839358276578162060532283322065990795137372571480712987182109661759531541721303126722689583504241219918742274834857803582922750003964604596480756638423624819172935296873131593417347651471480808537917236321275863665855942739108131662937389909773424721681271692982230323892361980688778592;
            5'd19: xpb[11] = 1024'd105155387669522866749105480968139595336552434549225666129868612796598095271999611984646317553217966777621129373995364128971928414810374646471595335128633305067894212925245273234560291252039411799195317779940384306712203546020760629626086974535831158420493079114708551510563225358771177469146039676896414707254;
            5'd20: xpb[11] = 1024'd12742490427820327052638195173188179766345909689393582140810233155647814493702902949615804360236537942672386650949730582144874246504694100584447622490931604597501270524280905506671170377264744745487020603842057286251508324584303210423529523445693759442503317425390271566298241371920739690849497165186546151585;
            5'd21: xpb[11] = 1024'd44396288870242528754969836783051196940837811955297182279883708579674429052715332824600362381912783417166793335361590469896883919040233889252460034869560945060799002692887755116412288694007283413088921036130970112155173953368742564185950642038785809731333459150189049652139785458998934929671644480102272080247;
            5'd22: xpb[11] = 1024'd76050087312664730457301478392914214115329714221200782418957184003701043611727762699584920403589028891661200019773450357648893591575773677920472447248190285524096734861494604726153407010749822080690821468419882938058839582153181917948371760631877860020163600874987827737981329546077130168493791795017998008909;
            5'd23: xpb[11] = 1024'd107703885755086932159633120002777231289821616487104382558030659427727658170740192574569478425265274366155606704185310245400903264111313466588484859626819625987394467030101454335894525327492360748292721900708795763962505210937621271710792879224969910308993742599786605823822873633155325407315939109933723937571;
            5'd24: xpb[11] = 1024'd15290988513384392463165834207825815719615091627272298568972279786777377392443483539538965232283845531206863981139676698573849095805632920701337146989117925517001524629137086608005404452717693694584424724610468743501809989501163852508235428134832511331003980910468325879557889646304887629019396598223855381902;
            5'd25: xpb[11] = 1024'd46944786955806594165497475817688832894106993893175898708045755210803991951455913414523523253960091005701270665551536586325858768341172709369349559367747265980299256797743936217746522769460232362186325156899381569405475618285603206270656546727924561619834122635267103965399433733383082867841543913139581310564;
            5'd26: xpb[11] = 1024'd78598585398228795867829117427551850068598896159079498847119230634830606510468343289508081275636336480195677349963396474077868440876712498037361971746376606443596988966350785827487641086202771029788225589188294395309141247070042560033077665321016611908664264360065882051240977820461278106663691228055307239226;
            5'd27: xpb[11] = 1024'd110252383840650997570160759037414867243090798424983098986192706058857221069480773164492639297312581954690084034375256361829878113412252286705374384125005946906894721134957635437228759402945309697390126021477207221212806875854481913795498783914108662197494406084864660137082521907539473345485838542971033167888;
            5'd28: xpb[11] = 1024'd17839486598948457873693473242463451672884273565151014997134326417906940291184064129462126104331153119741341311329622815002823945106571740818226671487304246436501778733993267709339638528170642643681828845378880200752111654418024494592941332823971263219504644395546380192817537920689035567189296031261164612219;
            5'd29: xpb[11] = 1024'd49493285041370659576025114852326468847376175831054615136207801841933554850196494004446684126007398594235747995741482702754833617642111529486239083865933586899799510902600117319080756844913181311283729277667793026655777283202463848355362451417063313508334786120345158278659082007767230806011443346176890540881;
            5'd30: xpb[11] = 1024'd81147083483792861278356756462189486021868078096958215275281277265960169409208923879431242147683644068730154680153342590506843290177651318154251496244562927363097243071206966928821875161655719978885629709956705852559442911986903202117783570010155363797164927845143936364500626094845426044833590661092616469543;
            5'd31: xpb[11] = 1024'd112800881926215062980688398072052503196359980362861815414354752689986783968221353754415800169359889543224561364565202478258852962713191106822263908623192267826394975239813816538562993478398258646487530142245618678463108540771342555880204688603247414085995069569942714450342170181923621283655737976008342398205;
        endcase
    end

    always_comb begin
        case(flag[4][5:0])
            6'd0: xpb[12] = 1024'd0;
            6'd1: xpb[12] = 1024'd10193992342256261642110556138550543813076727751514865712648186524518251594962322359692643488189230354137909320759784465715899397203755280467558097992745283678001016419424724405336936301811795796389616483073645829001206659667442568338823618756555007554002653940312217253038593097536591752679597732149236921268;
            6'd2: xpb[12] = 1024'd20387984684512523284221112277101087626153455503029731425296373049036503189924644719385286976378460708275818641519568931431798794407510560935116195985490567356002032838849448810673872603623591592779232966147291658002413319334885136677647237513110015108005307880624434506077186195073183505359195464298473842536;
            6'd3: xpb[12] = 1024'd30581977026768784926331668415651631439230183254544597137944559573554754784886967079077930464567691062413727962279353397147698191611265841402674293978235851034003049258274173216010808905435387389168849449220937487003619979002327705016470856269665022662007961820936651759115779292609775258038793196447710763804;
            6'd4: xpb[12] = 1024'd40775969369025046568442224554202175252306911006059462850592746098073006379849289438770573952756921416551637283039137862863597588815021121870232391970981134712004065677698897621347745207247183185558465932294583316004826638669770273355294475026220030216010615761248869012154372390146367010718390928596947685072;
            6'd5: xpb[12] = 1024'd50969961711281308210552780692752719065383638757574328563240932622591257974811611798463217440946151770689546603798922328579496986018776402337790489963726418390005082097123622026684681509058978981948082415368229145006033298337212841694118093782775037770013269701561086265192965487682958763397988660746184606340;
            6'd6: xpb[12] = 1024'd61163954053537569852663336831303262878460366509089194275889119147109509569773934158155860929135382124827455924558706794295396383222531682805348587956471702068006098516548346432021617810870774778337698898441874974007239958004655410032941712539330045324015923641873303518231558585219550516077586392895421527608;
            6'd7: xpb[12] = 1024'd71357946395793831494773892969853806691537094260604059988537305671627761164736256517848504417324612478965365245318491260011295780426286963272906685949216985746007114935973070837358554112682570574727315381515520803008446617672097978371765331295885052878018577582185520771270151682756142268757184125044658448876;
            6'd8: xpb[12] = 1024'd81551938738050093136884449108404350504613822012118925701185492196146012759698578877541147905513842833103274566078275725727195177630042243740464783941962269424008131355397795242695490414494366371116931864589166632009653277339540546710588950052440060432021231522497738024308744780292734021436781857193895370144;
            6'd9: xpb[12] = 1024'd91745931080306354778995005246954894317690549763633791413833678720664264354660901237233791393703073187241183886838060191443094574833797524208022881934707553102009147774822519648032426716306162167506548347662812461010859937006983115049412568808995067986023885462809955277347337877829325774116379589343132291412;
            6'd10: xpb[12] = 1024'd101939923422562616421105561385505438130767277515148657126481865245182515949623223596926434881892303541379093207597844657158993972037552804675580979927452836780010164194247244053369363018117957963896164830736458290012066596674425683388236187565550075540026539403122172530385930975365917526795977321492369212680;
            6'd11: xpb[12] = 1024'd112133915764818878063216117524055981943844005266663522839130051769700767544585545956619078370081533895517002528357629122874893369241308085143139077920198120458011180613671968458706299319929753760285781313810104119013273256341868251727059806322105083094029193343434389783424524072902509279475575053641606133948;
            6'd12: xpb[12] = 1024'd122327908107075139705326673662606525756920733018178388551778238294219019139547868316311721858270764249654911849117413588590792766445063365610697175912943404136012197033096692864043235621741549556675397796883749948014479916009310820065883425078660090648031847283746607036463117170439101032155172785790843055216;
            6'd13: xpb[12] = 1024'd8455204765206659948638302396342636825299033643957570136294569753760375397201051765989294131802320294349671762419704619727628322807598311523095148889357646880322538882950199931749932732036139631754816671570155930651325725455856615439728474151985648935214597809941766259395182194047059767716080691314485492153;
            6'd14: xpb[12] = 1024'd18649197107462921590748858534893180638375761395472435848942756278278626992163374125681937619991550648487581083179489085443527720011353591990653246882102930558323555302374924337086869033847935428144433154643801759652532385123299183778552092908540656489217251750253983512433775291583651520395678423463722413421;
            6'd15: xpb[12] = 1024'd28843189449719183232859414673443724451452489146987301561590942802796878587125696485374581108180781002625490403939273551159427117215108872458211344874848214236324571721799648742423805335659731224534049637717447588653739044790741752117375711665095664043219905690566200765472368389120243273075276155612959334689;
            6'd16: xpb[12] = 1024'd39037181791975444874969970811994268264529216898502167274239129327315130182088018845067224596370011356763399724699058016875326514418864152925769442867593497914325588141224373147760741637471527020923666120791093417654945704458184320456199330421650671597222559630878418018510961486656835025754873887762196255957;
            6'd17: xpb[12] = 1024'd49231174134231706517080526950544812077605944650017032986887315851833381777050341204759868084559241710901309045458842482591225911622619433393327540860338781592326604560649097553097677939283322817313282603864739246656152364125626888795022949178205679151225213571190635271549554584193426778434471619911433177225;
            6'd18: xpb[12] = 1024'd59425166476487968159191083089095355890682672401531898699535502376351633372012663564452511572748472065039218366218626948307125308826374713860885638853084065270327620980073821958434614241095118613702899086938385075657359023793069457133846567934760686705227867511502852524588147681730018531114069352060670098493;
            6'd19: xpb[12] = 1024'd69619158818744229801301639227645899703759400153046764412183688900869884966974985924145155060937702419177127686978411414023024706030129994328443736845829348948328637399498546363771550542906914410092515570012030904658565683460512025472670186691315694259230521451815069777626740779266610283793667084209907019761;
            6'd20: xpb[12] = 1024'd79813151161000491443412195366196443516836127904561630124831875425388136561937308283837798549126932773315037007738195879738924103233885274796001834838574632626329653818923270769108486844718710206482132053085676733659772343127954593811493805447870701813233175392127287030665333876803202036473264816359143941029;
            6'd21: xpb[12] = 1024'd90007143503256753085522751504746987329912855656076495837480061949906388156899630643530442037316163127452946328497980345454823500437640555263559932831319916304330670238347995174445423146530506002871748536159322562660979002795397162150317424204425709367235829332439504283703926974339793789152862548508380862297;
            6'd22: xpb[12] = 1024'd100201135845513014727633307643297531142989583407591361550128248474424639751861953003223085525505393481590855649257764811170722897641395835731118030824065199982331686657772719579782359448342301799261365019232968391662185662462839730489141042960980716921238483272751721536742520071876385541832460280657617783565;
            6'd23: xpb[12] = 1024'd110395128187769276369743863781848074956066311159106227262776434998942891346824275362915729013694623835728764970017549276886622294845151116198676128816810483660332703077197443985119295750154097595650981502306614220663392322130282298827964661717535724475241137213063938789781113169412977294512058012806854704833;
            6'd24: xpb[12] = 1024'd120589120530025538011854419920398618769143038910621092975424621523461142941786597722608372501883854189866674290777333742602521692048906396666234226809555767338333719496622168390456232051965893392040597985380260049664598981797724867166788280474090732029243791153376156042819706266949569047191655744956091626101;
            6'd25: xpb[12] = 1024'd6716417188157058255166048654134729837521339536400274559940952983002499199439781172285944775415410234561434204079624773739357248411441342578632199785970010082644061346475675458162929162260483467120016860066666032301444791244270662540633329547416290316426541679571315265751771290557527782752563650479734063038;
            6'd26: xpb[12] = 1024'd16910409530413319897276604792685273650598067287915140272589139507520750794402103531978588263604640588699343524839409239455256645615196623046190297778715293760645077765900399863499865464072279263509633343140311861302651450911713230879456948303971297870429195619883532518790364388094119535432161382628970984306;
            6'd27: xpb[12] = 1024'd27104401872669581539387160931235817463674795039430005985237326032039002389364425891671231751793870942837252845599193705171156042818951903513748395771460577438646094185325124268836801765884075059899249826213957690303858110579155799218280567060526305424431849560195749771828957485630711288111759114778207905574;
            6'd28: xpb[12] = 1024'd37298394214925843181497717069786361276751522790944871697885512556557253984326748251363875239983101296975162166358978170887055440022707183981306493764205861116647110604749848674173738067695870856288866309287603519305064770246598367557104185817081312978434503500507967024867550583167303040791356846927444826842;
            6'd29: xpb[12] = 1024'd47492386557182104823608273208336905089828250542459737410533699081075505579289070611056518728172331651113071487118762636602954837226462464448864591756951144794648127024174573079510674369507666652678482792361249348306271429914040935895927804573636320532437157440820184277906143680703894793470954579076681748110;
            6'd30: xpb[12] = 1024'd57686378899438366465718829346887448902904978293974603123181885605593757174251392970749162216361562005250980807878547102318854234430217744916422689749696428472649143443599297484847610671319462449068099275434895177307478089581483504234751423330191328086439811381132401530944736778240486546150552311225918669378;
            6'd31: xpb[12] = 1024'd67880371241694628107829385485437992715981706045489468835830072130112008769213715330441805704550792359388890128638331568034753631633973025383980787742441712150650159863024021890184546973131258245457715758508541006308684749248926072573575042086746335640442465321444618783983329875777078298830150043375155590646;
            6'd32: xpb[12] = 1024'd78074363583950889749939941623988536529058433797004334548478258654630260364176037690134449192740022713526799449398116033750653028837728305851538885735186995828651176282448746295521483274943054041847332241582186835309891408916368640912398660843301343194445119261756836037021922973313670051509747775524392511914;
            6'd33: xpb[12] = 1024'd88268355926207151392050497762539080342135161548519200261126445179148511959138360049827092680929253067664708770157900499466552426041483586319096983727932279506652192701873470700858419576754849838236948724655832664311098068583811209251222279599856350748447773202069053290060516070850261804189345507673629433182;
            6'd34: xpb[12] = 1024'd98462348268463413034161053901089624155211889300034065973774631703666763554100682409519736169118483421802618090917684965182451823245238866786655081720677563184653209121298195106195355878566645634626565207729478493312304728251253777590045898356411358302450427142381270543099109168386853556868943239822866354450;
            6'd35: xpb[12] = 1024'd108656340610719674676271610039640167968288617051548931686422818228185015149063004769212379657307713775940527411677469430898351220448994147254213179713422846862654225540722919511532292180378441431016181690803124322313511387918696345928869517112966365856453081082693487796137702265923445309548540971972103275718;
            6'd36: xpb[12] = 1024'd118850332952975936318382166178190711781365344803063797399071004752703266744025327128905023145496944130078436732437253896614250617652749427721771277706168130540655241960147643916869228482190237227405798173876770151314718047586138914267693135869521373410455735023005705049176295363460037062228138704121340196986;
            6'd37: xpb[12] = 1024'd4977629611107456561693794911926822849743645428842978983587336212244623001678510578582595419028500174773196645739544927751086174015284373634169250682582373284965583810001150984575925592484827302485217048563176133951563857032684709641538184942846931697638485549200864272108360387067995797789046609644982633923;
            6'd38: xpb[12] = 1024'd15171621953363718203804351050477366662820373180357844696235522736762874596640832938275238907217730528911105966499329393466985571219039654101727348675327656962966600229425875389912861894296623098874833531636821962952770516700127277980361803699401939251641139489513081525146953484604587550468644341794219555191;
            6'd39: xpb[12] = 1024'd25365614295619979845914907189027910475897100931872710408883709261281126191603155297967882395406960883049015287259113859182884968422794934569285446668072940640967616648850599795249798196108418895264450014710467791953977176367569846319185422455956946805643793429825298778185546582141179303148242073943456476459;
            6'd40: xpb[12] = 1024'd35559606637876241488025463327578454288973828683387576121531895785799377786565477657660525883596191237186924608018898324898784365626550215036843544660818224318968633068275324200586734497920214691654066497784113620955183836035012414658009041212511954359646447370137516031224139679677771055827839806092693397727;
            6'd41: xpb[12] = 1024'd45753598980132503130136019466128998102050556434902441834180082310317629381527800017353169371785421591324833928778682790614683762830305495504401642653563507996969649487700048605923670799732010488043682980857759449956390495702454982996832659969066961913649101310449733284262732777214362808507437538241930318995;
            6'd42: xpb[12] = 1024'd55947591322388764772246575604679541915127284186417307546828268834835880976490122377045812859974651945462743249538467256330583160034060775971959740646308791674970665907124773011260607101543806284433299463931405278957597155369897551335656278725621969467651755250761950537301325874750954561187035270391167240263;
            6'd43: xpb[12] = 1024'd66141583664645026414357131743230085728204011937932173259476455359354132571452444736738456348163882299600652570298251722046482557237816056439517838639054075352971682326549497416597543403355602080822915947005051107958803815037340119674479897482176977021654409191074167790339918972287546313866633002540404161531;
            6'd44: xpb[12] = 1024'd76335576006901288056467687881780629541280739689447038972124641883872384166414767096431099836353112653738561891058036187762381954441571336907075936631799359030972698745974221821934479705167397877212532430078696936960010474704782688013303516238731984575657063131386385043378512069824138066546230734689641082799;
            6'd45: xpb[12] = 1024'd86529568349157549698578244020331173354357467440961904684772828408390635761377089456123743324542343007876471211817820653478281351645326617374634034624544642708973715165398946227271416006979193673602148913152342765961217134372225256352127134995286992129659717071698602296417105167360729819225828466838878004067;
            6'd46: xpb[12] = 1024'd96723560691413811340688800158881717167434195192476770397421014932908887356339411815816386812731573362014380532577605119194180748849081897842192132617289926386974731584823670632608352308790989469991765396225988594962423794039667824690950753751841999683662371012010819549455698264897321571905426198988114925335;
            6'd47: xpb[12] = 1024'd106917553033670072982799356297432260980510922943991636110069201457427138951301734175509030300920803716152289853337389584910080146052837178309750230610035210064975748004248395037945288610602785266381381879299634423963630453707110393029774372508397007237665024952323036802494291362433913324585023931137351846603;
            6'd48: xpb[12] = 1024'd117111545375926334624909912435982804793587650695506501822717387981945390546264056535201673789110034070290199174097174050625979543256592458777308328602780493742976764423673119443282224912414581062770998362373280252964837113374552961368597991264952014791667678892635254055532884459970505077264621663286588767871;
            6'd49: xpb[12] = 1024'd3238842034057854868221541169718915861965951321285683407233719441486746803917239984879246062641590114984959087399465081762815099619127404689706301579194736487287106273526626510988922022709171137850417237059686235601682922821098756742443040338277573078850429418830413278464949483578463812825529568810231204808;
            6'd50: xpb[12] = 1024'd13432834376314116510332097308269459675042679072800549119881905966004998398879562344571889550830820469122868408159249547478714496822882685157264399571940020165288122692951350916325858324520966934240033720133332064602889582488541325081266659094832580632853083359142630531503542581115055565505127300959468126076;
            6'd51: xpb[12] = 1024'd23626826718570378152442653446820003488119406824315414832530092490523249993841884704264533039020050823260777728919034013194613894026637965624822497564685303843289139112376075321662794626332762730629650203206977893604096242155983893420090277851387588186855737299454847784542135678651647318184725033108705047344;
            6'd52: xpb[12] = 1024'd33820819060826639794553209585370547301196134575830280545178279015041501588804207063957176527209281177398687049678818478910513291230393246092380595557430587521290155531800799726999730928144558527019266686280623722605302901823426461758913896607942595740858391239767065037580728776188239070864322765257941968612;
            6'd53: xpb[12] = 1024'd44014811403082901436663765723921091114272862327345146257826465539559753183766529423649820015398511531536596370438602944626412688434148526559938693550175871199291171951225524132336667229956354323408883169354269551606509561490869030097737515364497603294861045180079282290619321873724830823543920497407178889880;
            6'd54: xpb[12] = 1024'd54208803745339163078774321862471634927349590078860011970474652064078004778728851783342463503587741885674505691198387410342312085637903807027496791542921154877292188370650248537673603531768150119798499652427915380607716221158311598436561134121052610848863699120391499543657914971261422576223518229556415811148;
            6'd55: xpb[12] = 1024'd64402796087595424720884878001022178740426317830374877683122838588596256373691174143035106991776972239812415011958171876058211482841659087495054889535666438555293204790074972943010539833579945916188116135501561209608922880825754166775384752877607618402866353060703716796696508068798014328903115961705652732416;
            6'd56: xpb[12] = 1024'd74596788429851686362995434139572722553503045581889743395771025113114507968653496502727750479966202593950324332717956341774110880045414367962612987528411722233294221209499697348347476135391741712577732618575207038610129540493196735114208371634162625956869007001015934049735101166334606081582713693854889653684;
            6'd57: xpb[12] = 1024'd84790780772107948005105990278123266366579773333404609108419211637632759563615818862420393968155432948088233653477740807490010277249169648430171085521157005911295237628924421753684412437203537508967349101648852867611336200160639303453031990390717633510871660941328151302773694263871197834262311426004126574952;
            6'd58: xpb[12] = 1024'd94984773114364209647216546416673810179656501084919474821067398162151011158578141222113037456344663302226142974237525273205909674452924928897729183513902289589296254048349146159021348739015333305356965584722498696612542859828081871791855609147272641064874314881640368555812287361407789586941909158153363496220;
            6'd59: xpb[12] = 1024'd105178765456620471289327102555224353992733228836434340533715584686669262753540463581805680944533893656364052294997309738921809071656680209365287281506647573267297270467773870564358285040827129101746582067796144525613749519495524440130679227903827648618876968821952585808850880458944381339621506890302600417488;
            6'd60: xpb[12] = 1024'd115372757798876732931437658693774897805809956587949206246363771211187514348502785941498324432723124010501961615757094204637708468860435489832845379499392856945298286887198594969695221342638924898136198550869790354614956179162967008469502846660382656172879622762264803061889473556480973092301104622451837338756;
            6'd61: xpb[12] = 1024'd1500054457008253174749287427511008874188257213728387830880102670728870606155969391175896706254680055196721529059385235774544025222970435745243352475807099689608628737052102037401918452933514973215617425556196337251801988609512803843347895733708214460062373288459962284821538580088931827862012527975479775693;
            6'd62: xpb[12] = 1024'd11694046799264514816859843566061552687264984965243253543528289195247122201118291750868540194443910409334630849819169701490443422426725716212801450468552383367609645156476826442738854754745310769605233908629842166253008648276955372182171514490263222014065027228772179537860131677625523580541610260124716696961;
            6'd63: xpb[12] = 1024'd21888039141520776458970399704612096500341712716758119256176475719765373796080614110561183682633140763472540170578954167206342819630480996680359548461297667045610661575901550848075791056557106565994850391703487995254215307944397940520995133246818229568067681169084396790898724775162115333221207992273953618229;
        endcase
    end

    always_comb begin
        case(flag[4][11:6])
            6'd0: xpb[13] = 1024'd0;
            6'd1: xpb[13] = 1024'd32082031483777038101080955843162640313418440468272984968824662244283625391042936470253827170822371117610449491338738632922242216834236277147917646454042950723611677995326275253412727358368902362384466874777133824255421967611840508859818752003373237122070335109396614043937317872698707085900805724423190539497;
            6'd2: xpb[13] = 1024'd64164062967554076202161911686325280626836880936545969937649324488567250782085872940507654341644742235220898982677477265844484433668472554295835292908085901447223355990652550506825454716737804724768933749554267648510843935223681017719637504006746474244140670218793228087874635745397414171801611448846381078994;
            6'd3: xpb[13] = 1024'd96246094451331114303242867529487920940255321404818954906473986732850876173128809410761481512467113352831348474016215898766726650502708831443752939362128852170835033985978825760238182075106707087153400624331401472766265902835521526579456256010119711366211005328189842131811953618096121257702417173269571618491;
            6'd4: xpb[13] = 1024'd4261430250983411005524895967836128508975334747356255747166793912157606226862606971000237468631810160998648557897461097109905026495724774036510460799840761960756037411733883676020670241958403728227669890721295450657327020226465262474296438330263499221461437023469398145642743416866195326484533071067167673657;
            6'd5: xpb[13] = 1024'd36343461734760449106605851810998768822393775215629240715991456156441231617905543441254064639454181278609098049236199730032147243329961051184428107253883712684367715407060158929433397600327306090612136765498429274912748987838305771334115190333636736343531772132866012189580061289564902412385338795490358213154;
            6'd6: xpb[13] = 1024'd68425493218537487207686807654161409135812215683902225684816118400724857008948479911507891810276552396219547540574938362954389460164197328332345753707926663407979393402386434182846124958696208452996603640275563099168170955450146280193933942337009973465602107242262626233517379162263609498286144519913548752651;
            6'd7: xpb[13] = 1024'd100507524702314525308767763497324049449230656152175210653640780645008482399991416381761718981098923513829997031913676995876631676998433605480263400161969614131591071397712709436258852317065110815381070515052696923423592923061986789053752694340383210587672442351659240277454697034962316584186950244336739292148;
            6'd8: xpb[13] = 1024'd8522860501966822011049791935672257017950669494712511494333587824315212453725213942000474937263620321997297115794922194219810052991449548073020921599681523921512074823467767352041340483916807456455339781442590901314654040452930524948592876660526998442922874046938796291285486833732390652969066142134335347314;
            6'd9: xpb[13] = 1024'd40604891985743860112130747778834897331369109962985496463158250068598837844768150412254302108085991439607746607133660827142052269825685825220938568053724474645123752818794042605454067842285709818839806656219724725570076008064771033808411628663900235564993209156335410335222804706431097738869871866557525886811;
            6'd10: xpb[13] = 1024'd72686923469520898213211703621997537644787550431258481431982912312882463235811086882508129278908362557218196098472399460064294486659922102368856214507767425368735430814120317858866795200654612181224273530996858549825497975676611542668230380667273472687063544265732024379160122579129804824770677590980716426308;
            6'd11: xpb[13] = 1024'd104768954953297936314292659465160177958205990899531466400807574557166088626854023352761956449730733674828645589811138092986536703494158379516773860961810376092347108809446593112279522559023514543608740405773992374080919943288452051528049132670646709809133879375128638423097440451828511910671483315403906965805;
            6'd12: xpb[13] = 1024'd12784290752950233016574687903508385526926004242068767241500381736472818680587820913000712405895430482995945673692383291329715079487174322109531382399522285882268112235201651028062010725875211184683009672163886351971981060679395787422889314990790497664384311070408194436928230250598585979453599213201503020971;
            6'd13: xpb[13] = 1024'd44866322236727271117655643746671025840344444710341752210325043980756444071630757383254539576717801600606395165031121924251957296321410599257449028853565236605879790230527926281474738084244113547067476546941020176227403028291236296282708066994163734786454646179804808480865548123297293065354404937624693560468;
            6'd14: xpb[13] = 1024'd76948353720504309218736599589833666153762885178614737179149706225040069462673693853508366747540172718216844656369860557174199513155646876405366675307608187329491468225854201534887465442613015909451943421718154000482824995903076805142526818997536971908524981289201422524802865995996000151255210662047884099965;
            6'd15: xpb[13] = 1024'd109030385204281347319817555432996306467181325646887722147974368469323694853716630323762193918362543835827294147708599190096441729989883153553284321761651138053103146221180476788300192800981918271836410296495287824738246963514917314002345571000910209030595316398598036568740183868694707237156016386471074639462;
            6'd16: xpb[13] = 1024'd17045721003933644022099583871344514035901338989425022988667175648630424907450427884000949874527240643994594231589844388439620105982899096146041843199363047843024149646935534704082680967833614912910679562885181802629308080905861049897185753321053996885845748093877592582570973667464781305938132284268670694628;
            6'd17: xpb[13] = 1024'd49127752487710682123180539714507154349319779457698007957491837892914050298493364354254777045349611761605043722928583021361862322817135373293959489653405998566635827642261809957495408326202517275295146437662315626884730048517701558757004505324427234007916083203274206626508291540163488391838938008691861234125;
            6'd18: xpb[13] = 1024'd81209783971487720224261495557669794662738219925970992926316500137197675689536300824508604216171982879215493214267321654284104539651371650441877136107448949290247505637588085210908135684571419637679613312439449451140152016129542067616823257327800471129986418312670820670445609412862195477739743733115051773622;
            6'd19: xpb[13] = 1024'd113291815455264758325342451400832434976156660394243977895141162381481301080579237294762431386994353996825942705606060287206346756485607927589794782561491900013859183632914360464320863042940322000064080187216583275395573983741382576476642009331173708252056753422067434714382927285560902563640549457538242313119;
            6'd20: xpb[13] = 1024'd21307151254917055027624479839180642544876673736781278735833969560788031134313034855001187343159050804993242789487305485549525132478623870182552303999203809803780187058669418380103351209792018641138349453606477253286635101132326312371482191651317496107307185117346990728213717084330976632422665355335838368285;
            6'd21: xpb[13] = 1024'd53389182738694093128705435682343282858295114205054263704658631805071656525355971325255014513981421922603692280826044118471767349312860147330469950453246760527391865053995693633516078568160921003522816328383611077542057068744166821231300943654690733229377520226743604772151034957029683718323471079759028907782;
            6'd22: xpb[13] = 1024'd85471214222471131229786391525505923171713554673327248673483294049355281916398907795508841684803793040214141772164782751394009566147096424478387596907289711251003543049321968886928805926529823365907283203160744901797479036356007330091119695658063970351447855336140218816088352829728390804224276804182219447279;
            6'd23: xpb[13] = 1024'd117553245706248169330867347368668563485131995141600233642307956293638907307441844265762668855626164157824591263503521384316251782981332701626305243361332661974615221044648244140341533284898725728291750077937878726052901003967847838950938447661437207473518190445536832860025670702427097890125082528605409986776;
            6'd24: xpb[13] = 1024'd25568581505900466033149375807016771053852008484137534483000763472945637361175641826001424811790860965991891347384766582659430158974348644219062764799044571764536224470403302056124021451750422369366019344327772703943962121358791574845778629981580995328768622140816388873856460501197171958907198426403006041942;
            6'd25: xpb[13] = 1024'd57650612989677504134230331650179411367270448952410519451825425717229262752218578296255251982613232083602340838723505215581672375808584921366980411253087522488147902465729577309536748810119324731750486219104906528199384088970632083705597381984954232450838957250213002917793778373895879044808004150826196581439;
            6'd26: xpb[13] = 1024'd89732644473454542235311287493342051680688889420683504420650087961512888143261514766509079153435603201212790330062243848503914592642821198514898057707130473211759580461055852562949476168488227094134953093882040352454806056582472592565416133988327469572909292359609616961731096246594586130708809875249387120936;
            6'd27: xpb[13] = 1024'd121814675957231580336392243336504691994107329888956489389474750205796513534304451236762906324257974318823239821400982481426156809477057475662815704161173423935371258456382127816362203526857129456519419968659174176710228024194313101425234885991700706694979627469006231005668414119293293216609615599672577660433;
            6'd28: xpb[13] = 1024'd29830011756883877038674271774852899562827343231493790230167557385103243588038248797001662280422671126990539905282227679769335185470073418255573225598885333725292261882137185732144691693708826097593689235049068154601289141585256837320075068311844494550230059164285787019499203918063367285391731497470173715599;
            6'd29: xpb[13] = 1024'd61912043240660915139755227618015539876245783699766775198992219629386868979081185267255489451245042244600989396620966312691577402304309695403490872052928284448903939877463460985557419052077728459978156109826201978856711109197097346179893820315217731672300394273682401063436521790762074371292537221893364255096;
            6'd30: xpb[13] = 1024'd93994074724437953240836183461178180189664224168039760167816881873670494370124121737509316622067413362211438887959704945613819619138545972551408518506971235172515617872789736238970146410446630822362622984603335803112133076808937855039712572318590968794370729383079015107373839663460781457193342946316554794593;
            6'd31: xpb[13] = 1024'd2009410524090249943118211899526387758384237510577061008509689052977224423857919297748072578232110170378738971840950143956997995131561915144166039944683144962436621298544794154752634577298327463436892250993229781003194194199881590934552754638734756649621161078358571121204629462230855525975458844114150849759;
            6'd32: xpb[13] = 1024'd34091442007867288044199167742689028071802677978850045977334351297260849814900855768001899749054481287989188463179688776879240211965798192292083686398726095686048299293871069408165361935667229825821359125770363605258616161811722099794371506642107993771691496187755185165141947334929562611876264568537341389256;
            6'd33: xpb[13] = 1024'd66173473491644326145280123585851668385221118447123030946159013541544475205943792238255726919876852405599637954518427409801482428800034469440001332852769046409659977289197344661578089294036132188205826000547497429514038129423562608654190258645481230893761831297151799209079265207628269697777070292960531928753;
            6'd34: xpb[13] = 1024'd98255504975421364246361079429014308698639558915396015914983675785828100596986728708509554090699223523210087445857166042723724645634270746587918979306811997133271655284523619914990816652405034550590292875324631253769460097035403117514009010648854468015832166406548413253016583080326976783677876017383722468250;
            6'd35: xpb[13] = 1024'd6270840775073660948643107867362516267359572257933316755676482965134830650720526268748310046863920331377387529738411241066903021627286689180676500744523906923192658710278677830773304819256731191664562141714525231660521214426346853408849192968998255871082598101827969266847372879097050852459991915181318523416;
            6'd36: xpb[13] = 1024'd38352872258850699049724063710525156580778012726206301724501145209418456041763462739002137217686291448987837021077149873989145238461522966328594147198566857646804336705604953084186032177625633554049029016491659055915943182038187362268667944972371492993152933211224583310784690751795757938360797639604509062913;
            6'd37: xpb[13] = 1024'd70434903742627737150805019553687796894196453194479286693325807453702081432806399209255964388508662566598286512415888506911387455295759243476511793652609808370416014700931228337598759535994535916433495891268792880171365149650027871128486696975744730115223268320621197354722008624494465024261603364027699602410;
            6'd38: xpb[13] = 1024'd102516935226404775251885975396850437207614893662752271662150469697985706823849335679509791559331033684208736003754627139833629672129995520624429440106652759094027692696257503591011486894363438278817962766045926704426787117261868379988305448979117967237293603430017811398659326497193172110162409088450890141907;
            6'd39: xpb[13] = 1024'd10532271026057071954168003835198644776334907005289572502843276877292436877583133239748547515495730492376036087635872338176808048123011463217186961544364668883948696122012561506793975061215134919892232032435820682317848234652812115883145631299261755092544035125297367412490116295963246178944524986248486197073;
            6'd40: xpb[13] = 1024'd42614302509834110055248959678361285089753347473562557471667939121576062268626069710002374686318101609986485578974610971099050264957247740365104607998407619607560374117338836760206702419584037282276698907212954506573270202264652624742964383302634992214614370234693981456427434168661953264845330710671676736570;
            6'd41: xpb[13] = 1024'd74696333993611148156329915521523925403171787941835542440492601365859687659669006180256201857140472727596935070313349604021292481791484017513022254452450570331172052112665112013619429777952939644661165781990088330828692169876493133602783135306008229336684705344090595500364752041360660350746136435094867276067;
            6'd42: xpb[13] = 1024'd106778365477388186257410871364686565716590228410108527409317263610143313050711942650510029027962843845207384561652088236943534698625720294660939900906493521054783730107991387267032157136321842007045632656767222155084114137488333642462601887309381466458755040453487209544302069914059367436646942159518057815564;
            6'd43: xpb[13] = 1024'd14793701277040482959692899803034773285310241752645828250010070789450043104445740210748784984127540653374684645533333435286713074618736237253697422344205430844704733533746445182814645303173538648119901923157116132975175254879277378357442069629525254314005472148766765558132859712829441505429058057315653870730;
            6'd44: xpb[13] = 1024'd46875732760817521060773855646197413598728682220918813218834733033733668495488676681002612154949911770985134136872072068208955291452972514401615068798248381568316411529072720436227372661542441010504368797934249957230597222491117887217260821632898491436075807258163379602070177585528148591329863781738844410227;
            6'd45: xpb[13] = 1024'd78957764244594559161854811489360053912147122689191798187659395278017293886531613151256439325772282888595583628210810701131197508287208791549532715252291332291928089524398995689640100019911343372888835672711383781486019190102958396077079573636271728558146142367559993646007495458226855677230669506162034949724;
            6'd46: xpb[13] = 1024'd111039795728371597262935767332522694225565563157464783156484057522300919277574549621510266496594654006206033119549549334053439725121445068697450361706334283015539767519725270943052827378280245735273302547488517605741441157714798904936898325639644965680216477476956607689944813330925562763131475230585225489221;
            6'd47: xpb[13] = 1024'd19055131528023893965217795770870901794285576500002083997176864701607649331308347181749022452759350814373333203430794532396618101114461011290207883144046192805460770945480328858835315545131942376347571813878411583632502275105742640831738507959788753535466909172236163703775603129695636831913591128382821544387;
            6'd48: xpb[13] = 1024'd51137163011800932066298751614033542107704016968275068966001526945891274722351283652002849623581721931983782694769533165318860317948697288438125529598089143529072448940806604112248042903500844738732038688655545407887924242717583149691557259963161990657537244281632777747712921002394343917814396852806012083884;
            6'd49: xpb[13] = 1024'd83219194495577970167379707457196182421122457436548053934826189190174900113394220122256676794404093049594232186108271798241102534782933565586043176052132094252684126936132879365660770261869747101116505563432679232143346210329423658551376011966535227779607579391029391791650238875093051003715202577229202623381;
            6'd50: xpb[13] = 1024'd115301225979355008268460663300358822734540897904821038903650851434458525504437156592510503965226464167204681677447010431163344751617169842733960822506175044976295804931459154619073497620238649463500972438209813056398768177941264167411194763969908464901677914500426005835587556747791758089616008301652393162878;
            6'd51: xpb[13] = 1024'd23316561779007304970742691738707030303260911247358339744343658613765255558170954152749259921391160975371981761328255629506523127610185785326718343943886954766216808357214212534855985787090346104575241704599707034289829295332207903306034946290052252756928346195705561849418346546561832158398124199449989218044;
            6'd52: xpb[13] = 1024'd55398593262784343071823647581869670616679351715631324713168320858048880949213890623003087092213532092982431252666994262428765344444422062474635990397929905489828486352540487788268713145459248466959708579376840858545251262944048412165853698293425489878998681305102175893355664419260539244298929923873179757541;
            6'd53: xpb[13] = 1024'd87480624746561381172904603425032310930097792183904309681992983102332506340256827093256914263035903210592880744005732895351007561278658339622553636851972856213440164347866763041681440503828150829344175454153974682800673230555888921025672450296798727001069016414498789937292982291959246330199735648296370297038;
            6'd54: xpb[13] = 1024'd119562656230338419273985559268194951243516232652177294650817645346616131731299763563510741433858274328203330235344471528273249778112894616770471283306015806937051842343193038295094167862197053191728642328931108507056095198167729429885491202300171964123139351523895403981230300164657953416100541372719560836535;
            6'd55: xpb[13] = 1024'd27577992029990715976267587706543158812236245994714595491510452525922861785033561123749497390022971136370630319225716726616428154105910559363228804743727716726972845768948096210876656029048749832802911595321002484947156315558673165780331384620315751978389783219174959995061089963428027484882657270517156891701;
            6'd56: xpb[13] = 1024'd59660023513767754077348543549705799125654686462987580460335114770206487176076497594003324560845342253981079810564455359538670370940146836511146451197770667450584523764274371464289383387417652195187378470098136309202578283170513674640150136623688989100460118328571574038998407836126734570783462994940347431198;
            6'd57: xpb[13] = 1024'd91742054997544792178429499392868439439073126931260565429159777014490112567119434064257151731667713371591529301903193992460912587774383113659064097651813618174196201759600646717702110745786554557571845344875270133458000250782354183499968888627062226222530453437968188082935725708825441656684268719363537970695;
            6'd58: xpb[13] = 1024'd123824086481321830279510455236031079752491567399533550397984439258773737958162370534510978902490084489201978793241932625383154804608619390806981744105856568897807879754926921971114838104155456919956312219652403957713422218394194692359787640630435463344600788547364802126873043581524148742585074443786728510192;
            6'd59: xpb[13] = 1024'd31839422280974126981792483674379287321211580742070851238677246438080468011896168094749734858654781297369278877123177823726333180601635333399739265543568478687728883180681979886897326271007153561030581486042297935604483335785138428254627822950579251199851220242644358140703833380294222811367190341584324565358;
            6'd60: xpb[13] = 1024'd63921453764751165082873439517541927634630021210343836207501908682364093402939104565003562029477152414979728368461916456648575397435871610547656911997611429411340561176008255140310053629376055923415048360819431759859905303396978937114446574953952488321921555352040972184641151252992929897267996066007515104855;
            6'd61: xpb[13] = 1024'd96003485248528203183954395360704567948048461678616821176326570926647718793982041035257389200299523532590177859800655089570817614270107887695574558451654380134952239171334530393722780987744958285799515235596565584115327271008819445974265326957325725443991890461437586228578469125691636983168801790430705644352;
            6'd62: xpb[13] = 1024'd4018821048180499886236423799052775516768475021154122017019378105954448847715838595496145156464220340757477943681900287913995990263123830288332079889366289924873242597089588309505269154596654926873784501986459562006388388399763181869105509277469513299242322156717142242409258924461711051950917688228301699518;
            6'd63: xpb[13] = 1024'd36100852531957537987317379642215415830186915489427106985844040350238074238758775065749972327286591458367927435020638920836238207097360107436249726343409240648484920592415863562917996512965557289258251376763593386261810356011603690728924261280842750421312657266113756286346576797160418137851723412651492239015;
        endcase
    end

    always_comb begin
        case(flag[4][16:12])
            5'd0: xpb[14] = 1024'd0;
            5'd1: xpb[14] = 1024'd68182884015734576088398335485378056143605355957700091954668702594521699629801711536003799498108962575978376926359377553758480423931596384584167372797452191372096598587742138816330723871334459651642718251540727210517232323623444199588743013284215987543382992375510370330283894669859125223752529137074682778512;
            5'd2: xpb[14] = 1024'd12299072347344410777997743565941679542512284789664499781205550124066503922294284161992527781560250842513604445261261672937897007021972434613174620578573341810502522605913060295031208551151713581975238894694214574670103797025991626212507456885202525819946081336903682630461261265789617430386368447523771072693;
            5'd3: xpb[14] = 1024'd80481956363078986866396079051319735686117640747364591735874252718588203552095995697996327279669213418491981371620639226696377430953568819197341993376025533182599121193655199111361932422486173233617957146234941785187336120649435825801250470169418513363329073712414052960745155935648742654138897584598453851205;
            5'd4: xpb[14] = 1024'd24598144694688821555995487131883359085024569579328999562411100248133007844588568323985055563120501685027208890522523345875794014043944869226349241157146683621005045211826120590062417102303427163950477789388429149340207594051983252425014913770405051639892162673807365260922522531579234860772736895047542145386;
            5'd5: xpb[14] = 1024'd92781028710423397644393822617261415228629925537029091517079802842654707474390279859988855061229464261005585816881900899634274437975541253810516613954598874993101643799568259406393140973637886815593196040929156359857439917675427452013757927054621039183275155049317735591206417201438360084525266032122224923898;
            5'd6: xpb[14] = 1024'd36897217042033232333993230697825038627536854368993499343616650372199511766882852485977583344680752527540813335783785018813691021065917303839523861735720025431507567817739180885093625653455140745925716684082643724010311391077974878637522370655607577459838244010711047891383783797368852291159105342571313218079;
            5'd7: xpb[14] = 1024'd105080101057767808422391566183203094771142210326693591298285352966721211396684564021981382842789715103519190262143162572572171444997513688423691234533172216803604166405481319701424349524789600397568434935623370934527543714701419078226265383939823565003221236386221418221667678467227977514911634479645995996591;
            5'd8: xpb[14] = 1024'd49196289389377643111990974263766718170049139158657999124822200496266015689177136647970111126241003370054417781045046691751588028087889738452698482314293367242010090423652241180124834204606854327900955578776858298680415188103966504850029827540810103279784325347614730521845045063158469721545473790095084290772;
            5'd9: xpb[14] = 1024'd117379173405112219200389309749144774313654495116358091079490903090787715318978848183973910624349965946032794707404424245510068452019486123036865855111745558614106689011394379996455558075941313979543673830317585509197647511727410704438772840825026090823167317723125100852128939733017594945298002927169767069284;
            5'd10: xpb[14] = 1024'd61495361736722053889988717829708397712561423948322498906027750620332519611471420809962638907801254212568022226306308364689485035109862173065873102892866709052512613029565301475156042755758567909876194473471072873350518985129958131062537284426012629099730406684518413152306306328948087151931842237618855363465;
            5'd11: xpb[14] = 1024'd5611550068331888579588125910272021111468352780286906732564598149877323903963993435951367191252542479103249745208192483868901618200238223094880350673987859490918537047736222953856527435575821840208715116624560237503390458532505557686301728026999167376293495645911725452483672924878579358565681548067943657646;
            5'd12: xpb[14] = 1024'd73794434084066464667986461395650077255073708737986998687233300744399023533765704971955166689361505055081626671567570037627382042131834607679047723471440050863015135635478361770187251306910281491851433368165287448020622782155949757275044741311215154919676488021422095782767567594737704582318210685142626436158;
            5'd13: xpb[14] = 1024'd17910622415676299357585869476213700653980637569951406513770148273943827826258277597943894972812793321616854190469454156806798625222210657708054971252561201301421059653649283248887735986727535422183954011318774812173494255558497183898809184912201693196239576982815408082944934190668196788952049995591714730339;
            5'd14: xpb[14] = 1024'd86093506431410875445984204961591756797585993527651498468438850868465527456059989133947694470921755897595231116828831710565279049153807042292222344050013392673517658241391422065218459858061995073826672262859502022690726579181941383487552198196417680739622569358325778413228828860527322012704579132666397508851;
            5'd15: xpb[14] = 1024'd30209694763020710135583613042155380196492922359615906294975698398010331748552561759936422754373044164130458635730715829744695632244183092321229591831134543111923582259562343543918944537879249004159192906012989386843598052584488810111316641797404219016185658319719090713406195456457814219338418443115485803032;
            5'd16: xpb[14] = 1024'd98392578778755286223981948527533436340098278317315998249644400992532031378354273295940222252482006740108835562090093383503176056175779476905396964628586734484020180847304482360249668409213708655801911157553716597360830376207933009700059655081620206559568650695229461043690090126316939443090947580190168581544;
            5'd17: xpb[14] = 1024'd42508767110365120913581356608097059739005207149280406076181248522076835670846845921928950535933295006644063080991977502682592639266155526934404212409707884922426104865475403838950153089030962586134431800707203961513701849610480436323824098682606744836131739656622773343867456722247431649724786890639256875725;
            5'd18: xpb[14] = 1024'd110691651126099697001979692093475115882610563106980498030849951116598535300648557457932750034042257582622440007351355056441073063197751911518571585207160076294522703453217542655280876960365422237777150052247931172030934173233924635912567111966822732379514732032133143674151351392106556873477316027713939654237;
            5'd19: xpb[14] = 1024'd54807839457709531691579100174038739281517491938944905857386798646143339593141130083921478317493545849157667526253239175620489646288127961547578832988281226732928627471388464133981361640182676168109670695401418536183805646636472062536331555567809270656077820993526455974328717988037049080111155338163027948418;
            5'd20: xpb[14] = 1024'd122990723473444107779977435659416795425122847896644997812055501240665039222942841619925277815602508425136044452612616729378970070219724346131746205785733418105025226059130602950312085511517135819752388946942145746701037970259916262125074568852025258199460813369036826304612612657896174303863684475237710726930;
            5'd21: xpb[14] = 1024'd67106911805053942469576843739980418824029776728609405638592348770209843515435414245914006099053796691671271971514500848558386653310100396160753453566854568543431150077301524429012570191334389750084909590095633110853909443662463688748839012453011796476023902330430138604789979253826666510497523785686799021111;
            5'd22: xpb[14] = 1024'd11223100136663777159176251820544042222936705560573813465129196299754647807927986871902734382505084958206499490416384967737803236400476446189760701347975718981837074095472445907713054871151643680417430233249120475006780917065011115372603456053998334752586991291823450904967345849757158717131363096135887315292;
            5'd23: xpb[14] = 1024'd79405984152398353247574587305922098366542061518273905419797898894276347437729698407906533880614047534184876416775762521496283660332072830773928074145427910353933672683214584724043778742486103332060148484789847685524013240688455314961346469338214322295969983667333821235251240519616283940883892233210570093804;
            5'd24: xpb[14] = 1024'd23522172484008187937173995386485721765448990350238313246334746423821151730222271033895262164065335800720103935677646640675700243422448880802935321926549060792339596701385506202744263422303357262392669127943335049676884714091002741585110912939200860572533072628727133535428607115546776147517731543659658387985;
            5'd25: xpb[14] = 1024'd91705056499742764025572330871863777909054346307938405201003449018342851360023982569899061662174298376698480862037024194434180667354045265387102694724001252164436195289127645019074987293637816914035387379484062260194117037714446941173853926223416848115916065004237503865712501785405901371270260680734341166497;
            5'd26: xpb[14] = 1024'd35821244831352598715171738952427401307961275139902813027540296547887655652516555195887789945625586643233708380938908313613597250444421315416109942505122402602842119307298566497775471973455070844367908022637549624346988511116994367797618369824403386392479153965630816165889868381336393577904099991183429460678;
            5'd27: xpb[14] = 1024'd104004128847087174803570074437805457451566631097602904982208999142409355282318266731891589443734549219212085307298285867372077674376017700000277315302574593974938717895040705314106195844789530496010626274178276834864220834740438567386361383108619373935862146341141186496173763051195518801656629128258112239190;
            5'd28: xpb[14] = 1024'd48120317178697009493169482518369080850473559929567312808745846671954159574810839357880317727185837485747312826200169986551494257466393750029284563083695744413344641913211626792806680524606784426343146917331764199017092308142985994010125826709605912212425235302534498796351129647126011008290468438707200533371;
            5'd29: xpb[14] = 1024'd116303201194431585581567818003747136994078915887267404763414549266475859204612550893884117225294800061725689752559547540309974681397990134613451935881147935785441240500953765609137404395941244077985865168872491409534324631766430193598868839993821899755808227678044869126635024316985136232042997575781883311883;
            5'd30: xpb[14] = 1024'd60419389526041420271167226084310760392985844719231812589951396796020663497105123519872845508746088328260917271461431659489391264488366184642459183662269086223847164519124687087837889075758498008318385812025978773687196105168977620222633283594808438032371316639438181426812390912915628438676836886230971606064;
            5'd31: xpb[14] = 1024'd4535577857651254960766634164874383791892773551196220416488244325565467789597696145861573792197376594796144790363315778668807847578742234671466431443390236662253088537295608566538373755575751938650906455179466137840067578571525046846397727195794976308934405600831493726989757508846120645310676196680059900245;
        endcase
    end

    always_comb begin
        case(flag[5][5:0])
            6'd0: xpb[15] = 1024'd0;
            6'd1: xpb[15] = 1024'd98392578778755286223981948527533436340098278317315998249644400992532031378354273295940222252482006740108835562090093383503176056175779476905396964628586734484020180847304482360249668409213708655801911157553716597360830376207933009700059655081620206559568650695229461043690090126316939443090947580190168581544;
            6'd2: xpb[15] = 1024'd72718461873385831049164969650252439935498129508896312371156946920087167419399407681865373290306339170774521716722693332427288271510338619255633804240842428034349687125037747382869097626910211590293624706720193348357299902194969246435140740480010963852317397976341864057273652178705245869063205333754742678757;
            6'd3: xpb[15] = 1024'd47044344968016375874347990772971443530897980700476626492669492847642303460444542067790524328130671601440207871355293281351400486844897761605870643853098121584679193402771012405488526844606714524785338255886670099353769428182005483170221825878401721145066145257454267070857214231093552295035463087319316775970;
            6'd4: xpb[15] = 1024'd21370228062646920699531011895690447126297831892056940614182038775197439501489676453715675365955004032105894025987893230275512702179456903956107483465353815135008699680504277428107956062303217459277051805053146850350238954169041719905302911276792478437814892538566670084440776283481858721007720840883890873183;
            6'd5: xpb[15] = 1024'd119762806841402206923512960423223883466396110209372938863826439767729470879843949749655897618437010772214729588077986613778688758355236380861504448093940549619028880527808759788357624471516926115078962962606863447711069330376974729605362566358412684997383543233796131128130866409798798164098668421074059454727;
            6'd6: xpb[15] = 1024'd94088689936032751748695981545942887061795961400953252985338985695284606920889084135581048656261343202880415742710586562702800973689795523211741287706196243169358386805542024810977053689213429049570676511773340198707538856364010966340443651756803442290132290514908534141714428462187104590070926174638633551940;
            6'd7: xpb[15] = 1024'd68414573030663296573879002668661890657195812592533567106851531622839742961934218521506199694085675633546101897343186511626913189024354665561978127318451936719687893083275289833596482906909931984062390060939816949704008382351047203075524737155194199582881037796020937155297990514575411016043183928203207649153;
            6'd8: xpb[15] = 1024'd42740456125293841399062023791380894252595663784113881228364077550394879002979352907431350731910008064211788051975786460551025404358913807912214966930707630270017399361008554856215912124606434918554103610106293700700477908338083439810605822553584956875629785077133340168881552566963717442015441681767781746366;
            6'd9: xpb[15] = 1024'd17066339219924386224245044914099897847995514975694195349876623477950015044024487293356501769734340494877474206608386409475137619693472950262451806542963323820346905638741819878835341342302937853045817159272770451696947434325119676545686907951975714168378532358245743182465114619352023867987699435332355843579;
            6'd10: xpb[15] = 1024'd115458917998679672448226993441633334188093793293010193599521024470482046422378760589296724022216347234986309768698479792978313675869252427167848771171550058304367086486046302239085009751516646508847728316826487049057777810533052686245746563033595920727947183053475204226155204745668963311078647015522524425123;
            6'd11: xpb[15] = 1024'd89784801093310217273410014564352337783493644484590507721033570398037182463423894975221875060040679665651995923331079741902425891203811569518085610783805751854696592763779567261704438969213149443339441865992963800054247336520088922980827648431986678020695930334587607239738766798057269737050904769087098522336;
            6'd12: xpb[15] = 1024'd64110684187940762098593035687071341378893495676170821842546116325592318504469029361147026097865012096317682077963679690826538106538370711868322450396061445405026099041512832284323868186909652377831155415159440551050716862507125159715908733830377435313444677615700010253322328850445576163023162522651672619549;
            6'd13: xpb[15] = 1024'd38436567282571306923776056809790344974293346867751135964058662253147454545514163747072177135689344526983368232596279639750650321872929854218559290008317138955355605319246097306943297404606155312322868964325917302047186388494161396450989819228768192606193424896812413266905890902833882588995420276216246716762;
            6'd14: xpb[15] = 1024'd12762450377201851748959077932509348569693198059331450085571208180702590586559298132997328173513676957649054387228879588674762537207488996568796129620572832505685111596979362329562726622302658246814582513492394053043655914481197633186070904627158949898942172177924816280489452955222189014967678029780820813975;
            6'd15: xpb[15] = 1024'd111155029155957137972941026460042784909791476376647448335215609173234621964913571428937550425995683697757889949318972972177938593383268473474193094249159566989705292444283844689812395031516366902616493671046110650404486290689130642886130559708779156458510822873154277324179543081539128458058625609970989395519;
            6'd16: xpb[15] = 1024'd85480912250587682798124047582761788505191327568227762456728155100789758005958705814862701463820016128423576103951572921102050808717827615824429933861415260540034798722017109712431824249212869837108207220212587401400955816676166879621211645107169913751259570154266680337763105133927434884030883363535563492732;
            6'd17: xpb[15] = 1024'd59806795345218227623307068705480792100591178759808076578240701028344894047003840200787852501644348559089262258584172870026163024052386758174666773473670954090364304999750374735051253466909372771599920769379064152397425342663203116356292730505560671044008317435379083351346667186315741310003141117100137589945;
            6'd18: xpb[15] = 1024'd34132678439848772448490089828199795695991029951388390699753246955900030088048974586713003539468680989754948413216772818950275239386945900524903613085926647640693811277483639757670682684605875706091634318545540903393894868650239353091373815903951428336757064716491486364930229238704047735975398870664711687158;
            6'd19: xpb[15] = 1024'd8458561534479317273673110950918799291390881142968704821265792883455166129094108972638154577293013420420634567849372767874387454721505042875140452698182341191023317555216904780290111902302378640583347867712017654390364394637275589826454901302342185629505811997603889378513791291092354161947656624229285784371;
            6'd20: xpb[15] = 1024'd106851140313234603497655059478452235631489159460284703070910193875987197507448382268578376829775020160529470129939466151377563510897284519780537417326769075675043498402521387140539780311516087296385259025265734251751194770845208599526514556383962392189074462692833350422203881417409293605038604204419454365915;
            6'd21: xpb[15] = 1024'd81177023407865148322838080601171239226889010651865017192422739803542333548493516654503527867599352591195156284572066100301675726231843662130774256939024769225373004680254652163159209529212590230876972574432211002747664296832244836261595641782353149481823209973945753435787443469797600031010861957984028463128;
            6'd22: xpb[15] = 1024'd55502906502495693148021101723890242822288861843445331313935285731097469589538651040428678905423685021860842439204666049225787941566402804481011096551280462775702510957987917185778638746909093165368686123598687753744133822819281072996676727180743906774571957255058156449371005522185906456983119711548602560341;
            6'd23: xpb[15] = 1024'd29828789597126237973204122846609246417688713035025645435447831658652605630583785426353829943248017452526528593837265998149900156900961946831247936163536156326032017235721182208398067964605596099860399672765164504740603348806317309731757812579134664067320704536170559462954567574574212882955377465113176657554;
            6'd24: xpb[15] = 1024'd4154672691756782798387143969328250013088564226605959556960377586207741671628919812278980981072349883192214748469865947074012372235521089181484775775791849876361523513454447231017497182302099034352113221931641255737072874793353546466838897977525421360069451817282962476538129626962519308927635218677750754767;
            6'd25: xpb[15] = 1024'd102547251470512069022369092496861686353186842543921957806604778578739773049983193108219203233554356623301050310559959330577188428411300566086881740404378584360381704360758929591267165591515807690154024379485357853097903251001286556166898553059145627919638102512512423520228219753279458752018582798867919336311;
            6'd26: xpb[15] = 1024'd76873134565142613847552113619580689948586693735502271928117324506294909091028327494144354271378689053966736465192559279501300643745859708437118580016634277910711210638492194613886594809212310624645737928651834604094372776988322792901979638457536385212386849793624826533811781805667765177990840552432493433524;
            6'd27: xpb[15] = 1024'd51199017659773158672735134742299693543986544927082586049629870433850045132073461880069505309203021484632422619825159228425412859080418850787355419628889971461040716916225459636506024026908813559137451477818311355090842302975359029637060723855927142505135597074737229547395343858056071603963098305997067530737;
            6'd28: xpb[15] = 1024'd25524900754403703497918155865018697139386396118662900171142416361405181173118596265994656347027353915298108774457759177349525074414977993137592259241145665011370223193958724659125453244605316493629165026984788106087311828962395266372141809254317899797884344355849632560978905910444378029935356059561641627950;
            6'd29: xpb[15] = 1024'd123917479533158989721900104392552133479484674435978898420786817353937212551472869561934878599509360655406944336547852560852701130590757470042989223869732399495390404041263207019375121653819025149431076184538504703448142205170328276072201464335938106357452995051079093604668996036761317473026303639751810209494;
            6'd30: xpb[15] = 1024'd98243362627789534547083125515271137074884525627559212542299363281492348592518003947860029637333693086072630491180452509776813345925316612393226063481988093045719910318996472041994550871515528083922789733704981454444611731157364512807282549734328863650201742332191496618252558089149623898998561393316384306707;
            6'd31: xpb[15] = 1024'd72569245722420079372266146637990140670284376819139526663811909209047484633563138333785180675158025516738316645813052458700925561259875754743462903094243786596049416596729737064613980089212031018414503282871458205441081257144400749542363635132719620942950489613303899631836120141537930324970819146880958403920;
            6'd32: xpb[15] = 1024'd46895128817050624197449167760709144265684228010719840785324455136602620674608272719710331712982357947404002800445652407625037776594434897093699742706499480146378922874463002087233409306908533952906216832037934956437550783131436986277444720531110378235699236894416302645419682193926236750943076900445532501133;
            6'd33: xpb[15] = 1024'd21221011911681169022632188883428147861084079202300154906837001064157756715653407105635482750806690378069688955078252356549149991928994039443936582318755173696708429152196267109852838524605036887397930381204411707434020309118473223012525805929501135528447984175528705659003244246314543176915334654010106598346;
            6'd34: xpb[15] = 1024'd119613590690436455246614137410961584201182357519616153156481402056689788094007680401575705003288697118178524517168345740052326048104773516349333546947341908180728609999500749470102506933818745543199841538758128304794850685326406232712585461011121342088016634870758166702693334372631482620006282234200275179890;
            6'd35: xpb[15] = 1024'd93939473785067000071797158533680587796582208711196467277993947984244924135052814787500856041113029548844210671800945688976438263439332658699570386559597601731058116277234014492721936151515248477691555087924605055791320211313442469447666546409512099380765382151870569716276896425019789045978539987764849277103;
            6'd36: xpb[15] = 1024'd68265356879697544896980179656399591391982059902776781399506493911800060176097949173426007078937361979509896826433545637900550478773891801049807226171853295281387622554967279515341365369211751412183268637091081806787789737300478706182747631807902856673514129432982972729860458477408095471950797741329423374316;
            6'd37: xpb[15] = 1024'd42591239974328089722163200779118594987381911094357095521019039839355196217143083559351158116761694410175582981066145586824662694108450943400044065784108988831717128832700544537960794586908254346674982186257558557784259263287514942917828717206293613966262876714095375743444020529796401897923055494893997471529;
            6'd38: xpb[15] = 1024'd16917123068958634547346221901837598582781762285937409642531585766910332258188217945276309154586026840841269135698745535748774909443010085750280905396364682382046635110433809560580223804604757281166695735424035308780728789274551179652909802604684371259011623995207778757027582582184708323895313248458571568742;
            6'd39: xpb[15] = 1024'd115309701847713920771328170429371034922880040603253407892175986759442363636542491241216531407068033580950104697788838919251950965618789562655677870024951416866066815957738291920829892213818465936968606892977751906141559165482484189352969457686304577818580274690437239800717672708501647766986260828648740150286;
            6'd40: xpb[15] = 1024'd89635584942344465596511191552090038518279891794833722013688532686997499677587625627141682444892366011615790852421438868176063180953348705005914709637207110416396322235471556943449321431514968871460320442144228657138028691469520426088050543084695335111329021971549642814301234760889954192958518582213314247499;
            6'd41: xpb[15] = 1024'd63961468036975010421694212674809042113679742986414036135201078614552635718632760013066833482716698442281477007054038817100175396287907847356151549249462803966725828513204821966068750649211471805952033991310705408134498217456556662823131628483086092404077769252662045827884796813278260618930776335777888344712;
            6'd42: xpb[15] = 1024'd38287351131605555246877233797528045709079594177994350256713624542107771759677894398991984520541030872947163161686638766024287611622466989706388388861718497517055334790938086988688179866907974740443747540477182159130967743443592899558212713881476849696826516533774448841468358865666567044903034089342462441925;
            6'd43: xpb[15] = 1024'd12613234226236100072060254920247049304479445369574664378226170469662907800723028784917135558365363303612849316319238714948399826957026132056625228473974191067384841068671352011307609084604477674935461089643658910127437269430629136293293799279867606989575263814886851855051920918054873470875291842907036539138;
            6'd44: xpb[15] = 1024'd111005813004991386296042203447780485644577723686890662627870571462194939179077302080857357810847370043721684878409332098451575883132805608962022193102560925551405021915975834371557277493818186330737372247197375507488267645638562145993353454361487813549143914510116312898742011044371812913966239423097205120682;
            6'd45: xpb[15] = 1024'd85331696099621931121225224570499489239977574878470976749383117389750075220122436466782508848671702474387371033041932047375688098467364751312259032714816619101734528193709099394176706711514689265229085796363852258484737171625598382728434539759878570841892661791228715912325573096760119339938497176661779217895;
            6'd46: xpb[15] = 1024'd59657579194252475946408245693218492835377426070051290870895663317305211261167570852707659886496034905053057187674531996299800313801923893662495872327072312652064034471442364416796135929211192199720799345530329009481206697612634619463515625158269328134641409072341118925909135149148425765910754930226353315108;
            6'd47: xpb[15] = 1024'd33983462288883020771591266815937496430777277261631604992408209244860347302212705238632810924320367335718743342307131945223912529136483036012732711939328006202393540749175629439415565146907695134212512894696805760477676223599670856198596710556660085427390156353453521939492697201536732191883012683790927412321;
            6'd48: xpb[15] = 1024'd8309345383513565596774287938656500026177128453211919113920755172415483343257839624557961962144699766384429496939731894148024744471042178362969551551583699752723047026908894462034994364604198068704226443863282511474145749586707092933677795955050842720138903634565924953076259253925038617855270437355501509534;
            6'd49: xpb[15] = 1024'd106701924162268851820756236466189936366275406770527917363565156164947514721612112920498184214626706506493265059029825277651200800646821655268366516180170434236743227874213376822284662773817906724506137601416999108834976125794640102633737451036671049279707554329795385996766349380241978060946218017545670091078;
            6'd50: xpb[15] = 1024'd81027807256899396645939257588908939961675257962108231485077702092502650762657247306423335252451038937158951213662425226575313015981380797618603355792426127787072734151946641844904091991514409658997851150583475859831445651781676339368818536435061806572456301610907789010349911432630284486918475771110244188291;
            6'd51: xpb[15] = 1024'd55353690351529941471122278711627943557075109153688545606590248020057786803702381692348486290275371367824637368295025175499425231315939939968840195404681821337402240429679906867523521209210912593489564699749952610827915177768712576103899621833452563865205048892020192023933473485018590912890733524674818285504;
            6'd52: xpb[15] = 1024'd29679573446160486296305299834346947152474960345268859728102793947612922844747516078273637328099703798490323522927625124423537446650499082319077035016937514887731746707413171890142950426907415527981278248916429361824384703755748812838980707231843321157953796173132595037517035537406897338862991278239392382717;
            6'd53: xpb[15] = 1024'd4005456540791031121488320957065950747874811536849173849615339875168058885792650464198788365924036229156009677560225073347649661985058224669313874629193208438061252985146436912762379644603918462472991798082906112820854229742785049574061792630234078450702543454244998051100597589795203764835249031803966479930;
            6'd54: xpb[15] = 1024'd102398035319546317345470269484599387087973089854165172099259740867700090264146923760139010618406042969264845239650318456850825718160837701574710839257779942922081433832450919273012048053817627118274902955636622710181684605950718059274121447711854285010271194149474459094790687716112143207926196611994135061474;
            6'd55: xpb[15] = 1024'd76723918414176862170653290607318390683372941045745486220772286795255226305192058146064161656230375399930531394282918405774937933495396843924947678870035636472410940110184184295631477271514130052766616504803099461178154131937754296009202533110245042303019941430586862108374249768500449633898454365558709158687;
            6'd56: xpb[15] = 1024'd51049801508807406995836311730037394278772792237325800342284832722810362346237192531989312694054707830596217548915518354699050148829955986275184518482291330022740446387917449318250906489210632987258330053969576212174623657924790532744283618508635799595768688711699265121957811820888756059870712119123283255900;
            6'd57: xpb[15] = 1024'd25375684603437951821019332852756397874172643428906114463797378650365498387282326917914463731879040261261903703548118303623162364164515128625421358094547023573069952665650714340870335706907135921750043603136052963171093183911826769479364703907026556888517435992811668135541373873277062485842969872687857353113;
            6'd58: xpb[15] = 1024'd123768263382193238045001281380289834214270921746222112713441779642897529765636600213854685984361047001370739265638211687126338420340294605530818322723133758057090133512955196701120004116120844577551954760689769560531923560119759779179424358988646763448086086688041129179231463999594001928933917452878025934657;
            6'd59: xpb[15] = 1024'd98094146476823782870184302503008837809670772937802426834954325570452665806681734599779837022185379432036425420270811636050450635674853747881055162335389451607419639790688461723739433333817347512043668309856246311528393086106796015914505444387037520740834833969153532192815026051982308354906175206442600031870;
            6'd60: xpb[15] = 1024'd72420029571454327695367323625727841405070624129382740956466871498007801847726868985704988060009711862702111574903411584974562851009412890231292001947645145157749146068421726746358862551513850446535381859022723062524862612093832252649586529785428278033583581250265935206398588104370614780878432960007174129083;
            6'd61: xpb[15] = 1024'd46745912666084872520550344748446845000470475320963055077979417425562937888772003371630139097834044293367797729536011533898675066343972032581528841559900838708078652346154991768978291769210353381027095408189199813521332138080868489384667615183819035326332328531378338219982150156758921206850690713571748226296;
            6'd62: xpb[15] = 1024'd21071795760715417345733365871165848595870326512543369199491963353118073929817137757555290135658376724033483884168611482822787281678531174931765681172156532258408158623888256791597720986906856315518808957355676564517801664067904726119748700582209792619081075812490741233565712209147227632822948467136322323509;
            6'd63: xpb[15] = 1024'd119464374539470703569715314398699284935968604829859367449136364345650105308171411053495512388140383464142319446258704866325963337854310651837162645800743266742428339471192739151847389396120564971320720114909393161878632040275837735819808355663829999178649726507720202277255802335464167075913896047326490905053;
        endcase
    end

    always_comb begin
        case(flag[5][11:6])
            6'd0: xpb[16] = 1024'd0;
            6'd1: xpb[16] = 1024'd93790257634101248394898335521418288531368456021439681570648910273205241349216545439420663425964715894808005600891304815250075553188869794187399485412998960292757845748926004174466818613817067905812433664075869912875101566262873972554889441062220756471398473788832605290839364387852473501886153800891065002266;
            6'd2: xpb[16] = 1024'd63513819584077755390997743638022144318038484917143679013165965481433587361123951968826255637271757480172861794325116195921087265536519253819638845809666879651825016928280791011303398036116930090314669719764499979385842282304851172144800312441212063675977044163548152551572200701776313986653617775156535520201;
            6'd3: xpb[16] = 1024'd33237381534054262387097151754626000104708513812847676455683020689661933373031358498231847848578799065537717987758927576592098977884168713451878206206334799010892188107635577848139977458416792274816905775453130045896582998346828371734711183820203370880555614538263699812305037015700154471421081749422006038136;
            6'd4: xpb[16] = 1024'd2960943484030769383196559871229855891378542708551673898200075897890279384938765027637440059885840650902574181192738957263110690231818173084117566603002718369959359286990364684976556880716654459319141831141760112407323714388805571324622055199194678085134184912979247073037873329623994956188545723687476556071;
            6'd5: xpb[16] = 1024'd96751201118132017778094895392648144422746998729991355468848986171095520734155310467058103485850556545710579782084043772513186243420687967271517052016001678662717205035916368859443375494533722365131575495217630025282425280651679543879511496261415434556532658701811852363877237717476468458074699524578541558337;
            6'd6: xpb[16] = 1024'd66474763068108524774194303509252000209417027625695352911366041379323866746062716996463695697157598131075435975517855153184197955768337426903756412412669598021784376215271155696279954916833584549633811550906260091793165996693656743469422367640406741761111229076527399624610074031400308942842163498844012076272;
            6'd7: xpb[16] = 1024'd36198325018085031770293711625855855996087056521399350353883096587552212757970123525869287908464639716440292168951666533855209668115986886535995772809337517380851547394625942533116534339133446734136047606594890158303906712735633943059333239019398048965689799451242946885342910345324149427609627473109482594207;
            6'd8: xpb[16] = 1024'd5921886968061538766393119742459711782757085417103347796400151795780558769877530055274880119771681301805148362385477914526221380463636346168235133206005436739918718573980729369953113761433308918638283662283520224814647428777611142649244110398389356170268369825958494146075746659247989912377091447374953112142;
            6'd9: xpb[16] = 1024'd99712144602162787161291455263878000314125541438543029367049062068985800119094075494695543545736397196613153963276782729776296933652506140355634618619004397032676564322906733544419932375250376824450717326359390137689748995040485115204133551460610112641666843614791099436915111047100463414263245248266018114408;
            6'd10: xpb[16] = 1024'd69435706552139294157390863380481856100795570334247026809566117277214146131001482024101135757043438781978010156710594110447308646000155599987873979015672316391743735502261520381256511797550239008952953382048020204200489711082462314794044422839601419846245413989506646697647947361024303899030709222531488632343;
            6'd11: xpb[16] = 1024'd39159268502115801153490271497085711887465599229951024252083172485442492142908888553506727968350480367342866350144405491118320358347805059620113339412340235750810906681616307218093091219850101193455189437736650270711230427124439514383955294218592727050823984364222193958380783674948144383798173196796959150278;
            6'd12: xpb[16] = 1024'd8882830452092308149589679613689567674135628125655021694600227693670838154816295082912320179657521952707722543578216871789332070695454519252352699809008155109878077860971094054929670642149963377957425493425280337221971143166416713973866165597584034255402554738937741219113619988871984868565637171062429668213;
            6'd13: xpb[16] = 1024'd102673088086193556544488015135107856205504084147094703265249137966876079504032840522332983605622237847515728144469521687039407623884324313439752185222007115402635923609897098229396489255967031283769859157501150250097072709429290686528755606659804790726801028527770346509952984376724458370451790971953494670479;
            6'd14: xpb[16] = 1024'd72396650036170063540587423251711711992174113042798700707766193175104425515940247051738575816929279432880584337903333067710419336231973773071991545618675034761703094789251885066233068678266893468272095213189780316607813425471267886118666478038796097931379598902485893770685820690648298855219254946218965188414;
            6'd15: xpb[16] = 1024'd42120211986146570536686831368315567778844141938502698150283248383332771527847653581144168028236321018245440531337144448381431048579623232704230906015342954120770265968606671903069648100566755652774331268878410383118554141513245085708577349417787405135958169277201441031418657004572139339986718920484435706349;
            6'd16: xpb[16] = 1024'd11843773936123077532786239484919423565514170834206695592800303591561117539755060110549760239543362603610296724770955829052442760927272692336470266412010873479837437147961458739906227522866617837276567324567040449629294857555222285298488220796778712340536739651916988292151493318495979824754182894749906224284;
            6'd17: xpb[16] = 1024'd105634031570224325927684575006337712096882626855646377163449213864766358888971605549970423665508078498418302325662260644302518314116142486523869751825009833772595282896887462914373046136683685743089000988642910362504396423818096257853377661858999468811935213440749593582990857706348453326640336695640971226550;
            6'd18: xpb[16] = 1024'd75357593520200832923783983122941567883552655751350374605966269072994704900879012079376015876815120083783158519096072024973530026463791946156109112221677753131662454076242249751209625558983547927591237044331540429015137139860073457443288533237990776016513783815465140843723694020272293811407800669906441744485;
            6'd19: xpb[16] = 1024'd45081155470177339919883391239545423670222684647054372048483324281223050912786418608781608088122161669148014712529883405644541738811441405788348472618345672490729625255597036588046204981283410112093473100020170495525877855902050657033199404616982083221092354190180688104456530334196134296175264644171912262420;
            6'd20: xpb[16] = 1024'd14804717420153846915982799356149279456892713542758369491000379489451396924693825138187200299429203254512870905963694786315553451159090865420587833015013591849796796434951823424882784403583272296595709155708800562036618571944027856623110275995973390425670924564896235365189366648119974780942728618437382780355;
            6'd21: xpb[16] = 1024'd108594975054255095310881134877567567988261169564198051061649289762656638273910370577607863725393919149320876506854999601565629004347960659607987318428012552142554642183877827599349603017400340202408142819784670474911720138206901829177999717058194146897069398353728840656028731035972448282828882419328447782621;
            6'd22: xpb[16] = 1024'd78318537004231602306980542994171423774931198459902048504166344970884984285817777107013455936700960734685732700288810982236640716695610119240226678824680471501621813363232614436186182439700202386910378875473300541422460854248879028767910588437185454101647968728444387916761567349896288767596346393593918300556;
            6'd23: xpb[16] = 1024'd48042098954208109303079951110775279561601227355606045946683400179113330297725183636419048148008002320050588893722622362907652429043259578872466039221348390860688984542587401273022761862000064571412614931161930607933201570290856228357821459816176761306226539103159935177494403663820129252363810367859388818491;
            6'd24: xpb[16] = 1024'd17765660904184616299179359227379135348271256251310043389200455387341676309632590165824640359315043905415445087156433743578664141390909038504705399618016310219756155721942188109859341284299926755914850986850560674443942286332833427947732331195168068510805109477875482438227239977743969737131274342124859336426;
            6'd25: xpb[16] = 1024'd111555918538285864694077694748797423879639712272749724959849365660546917658849135605245303785279759800223450688047738558828739694579778832692104885031015270512514001470868192284326159898116994661727284650926430587319043852595707400502621772257388824982203583266708087729066604365596443239017428143015924338692;
            6'd26: xpb[16] = 1024'd81279480488262371690177102865401279666309741168453722402366420868775263670756542134650895996586801385588306881481549939499751406927428292324344245427683189871581172650222979121162739320416856846229520706615060653829784568637684600092532643636380132186782153641423634989799440679520283723784892117281394856627;
            6'd27: xpb[16] = 1024'd51003042438238878686276510982005135452979770064157719844883476077003609682663948664056488207893842970953163074915361320170763119275077751956583605824351109230648343829577765957999318742716719030731756762303690720340525284679661799682443515015371439391360724016139182250532276993444124208552356091546865374562;
            6'd28: xpb[16] = 1024'd20726604388215385682375919098608991239649798959861717287400531285231955694571355193462080419200884556318019268349172700841774831622727211588822966221019028589715515008932552794835898165016581215233992817992320786851266000721638999272354386394362746595939294390854729511265113307367964693319820065812335892497;
            6'd29: xpb[16] = 1024'd114516862022316634077274254620027279771018254981301398858049441558437197043787900632882743845165600451126024869240477516091850384811597005776222451634017988882473360757858556969302716778833649121046426482068190699726367566984512971827243827456583503067337768179687334802104477695220438195205973866703400894763;
            6'd30: xpb[16] = 1024'd84240423972293141073373662736631135557688283877005396300566496766665543055695307162288336056472642036490881062674288896762862097159246465408461812030685908241540531937213343806139296201133511305548662537756820766237108283026490171417154698835574810271916338554402882062837314009144278679973437840968871412698;
            6'd31: xpb[16] = 1024'd53963985922269648069473070853234991344358312772709393743083551974893889067602713691693928267779683621855737256108100277433873809506895925040701172427353827600607703116568130642975875623433373490050898593445450832747848999068467371007065570214566117476494908929118429323570150323068119164740901815234341930633;
            6'd32: xpb[16] = 1024'd23687547872246155065572478969838847131028341668413391185600607183122235079510120221099520479086725207220593449541911658104885521854545384672940532824021746959674874295922917479812455045733235674553134649134080899258589715110444570596976441593557424681073479303833976584302986636991959649508365789499812448568;
            6'd33: xpb[16] = 1024'd117477805506347403460470814491257135662396797689853072756249517456327476428726665660520183905051441102028599050433216473354961075043415178860340018237020707252432720044848921654279273659550303580365568313209950812133691281373318543151865882655778181152471953092666581875142351024844433151394519590390877450834;
            6'd34: xpb[16] = 1024'd87201367456323910456570222607860991449066826585557070198766572664555822440634072189925776116358482687393455243867027854025972787391064638492579378633688626611499891224203708491115853081850165764867804368898580878644431997415295742741776754034769488357050523467382129135875187338768273636161983564656347968769;
            6'd35: xpb[16] = 1024'd56924929406300417452669630724464847235736855481261067641283627872784168452541478719331368327665524272758311437300839234696984499738714098124818739030356545970567062403558495327952432504150027949370040424587210945155172713457272942331687625413760795561629093842097676396608023652692114120929447538921818486704;
            6'd36: xpb[16] = 1024'd26648491356276924448769038841068703022406884376965065083800683081012514464448885248736960538972565858123167630734650615367996212086363557757058099427024465329634233582913282164789011926449890133872276480275841011665913429499250141921598496792752102766207664216813223657340859966615954605696911513187289004639;
            6'd37: xpb[16] = 1024'd120438748990378172843667374362486991553775340398404746654449593354217755813665430688157623964937281752931173231625955430618071765275233351944457584840023425622392079331839286339255830540266958039684710144351710924541014995762124114476487937854972859237606138005645828948180224354468428107583065314078354006905;
            6'd38: xpb[16] = 1024'd90162310940354679839766782479090847340445369294108744096966648562446101825572837217563216176244323338296029425059766811289083477622882811576696945236691344981459250511194073176092409962566820224186946200040340991051755711804101314066398809233964166442184708380361376208913060668392268592350529288343824524840;
            6'd39: xpb[16] = 1024'd59885872890331186835866190595694703127115398189812741539483703770674447837480243746968808387551364923660885618493578191960095189970532271208936305633359264340526421690548860012928989384866682408689182255728971057562496427846078513656309680612955473646763278755076923469645896982316109077117993262609295042775;
            6'd40: xpb[16] = 1024'd29609434840307693831965598712298558913785427085516738982000758978902793849387650276374400598858406509025741811927389572631106902318181730841175666030027183699593592869903646849765568807166544593191418311417601124073237143888055713246220551991946780851341849129792470730378733296239949561885457236874765560710;
            6'd41: xpb[16] = 1024'd123399692474408942226863934233716847445153883106956420552649669252108035198604195715795064024823122403833747412818694387881182455507051525028575151443026143992351438618829651024232387420983612499003851975493471036948338710150929685801109993054167537322740322918625076021218097684092423063771611037765830562976;
            6'd42: xpb[16] = 1024'd93123254424385449222963342350320703231823912002660417995166724460336381210511602245200656236130163989198603606252505768552194167854700984660814511839694063351418609798184437861068966843283474683506088031182101103459079426192906885391020864433158844527318893293340623281950933998016263548539075012031301080911;
            6'd43: xpb[16] = 1024'd62846816374361956219062750466924559018493940898364415437683779668564727222419008774606248447437205574563459799686317149223205880202350444293053872236361982710485780977539224697905546265583336868008324086870731169969820142234884084980931735812150151731897463668056170542683770311940104033306538986296771598846;
            6'd44: xpb[16] = 1024'd32570378324338463215162158583528414805163969794068412880200834876793073234326415304011840658744247159928315993120128529894217592549999903925293232633029902069552952156894011534742125687883199052510560142559361236480560858276861284570842607191141458936476034042771717803416606625863944518074002960562242116781;
            6'd45: xpb[16] = 1024'd2293940274314970211261566700132270591833998689772410322717890085021419246233821833417432870051288745293172186553939910565229304897649363557532593029697821428620123336248798371578705110183061237012796198247991302991301574318838484160753478570132766141054604417487265064149442939787785002841466934827712634716;
            6'd46: xpb[16] = 1024'd96084197908416218606159902221550559123202454711212091893366800358226660595450367272838096296016004640101177787445244725815304858086519157744932078442696781721377969085174802546045523724000129142825229862323861215866403140581712456715642919632353522612453078206319870354988807327640258504727620735718777636982;
            6'd47: xpb[16] = 1024'd65807759858392725602259310338154414909872483606916089335883855566455006607357773802243688507323046225466033980879056106486316570434168617377171438839364701080445140264529589382882103146299991327327465918012491282377143856623689656305553791011344829817031648581035417615721643641564098989495084709984248154917;
            6'd48: xpb[16] = 1024'd35531321808369232598358718454758270696542512502620086778400910774683352619265180331649280718630087810830890174312867487157328282781818077009410799236032620439512311443884376219718682568599853511829701973701121348887884572665666855895464662390336137021610218955750964876454479955487939474262548684249718672852;
            6'd49: xpb[16] = 1024'd5254883758345739594458126571362126483212541398324084220917965982911698631172586861054872929937129396195746367746678867828339995129467536641650159632700539798579482623239163056555261990899715696331938029389751415398625288707644055485375533769327444226188789330466512137187316269411779959030012658515189190787;
            6'd50: xpb[16] = 1024'd99045141392446987989356462092780415014580997419763765791566876256116939980389132300475536355901845291003751968637983683078415548318337330829049645045699500091337328372165167231022080604716783602144371693465621328273726854970518028040264974831548200697587263119299117428026680657264253460916166459406254193053;
            6'd51: xpb[16] = 1024'd68768703342423494985455870209384270801251026315467763234083931464345285992296538829881128567208886876368608162071795063749427260665986790461289005442367419450404499551519954067858660027016645786646607749154251394784467571012495227630175846210539507902165833494014664688759516971188093945683630433671724710988;
            6'd52: xpb[16] = 1024'd38492265292400001981555278325988126587921055211171760676600986672573632004203945359286720778515928461733464355505606444420438973013636250093528365839035338809471670730874740904695239449316507971148843804842881461295208287054472427220086717589530815106744403868730211949492353285111934430451094407937195228923;
            6'd53: xpb[16] = 1024'd8215827242376508977654686442591982374591084106875758119118041880801978016111351888692312989822970047098320548939417825091450685361285709725767726235703258168538841910229527741531818871616370155651079860531511527805949003096449626809997588968522122311322974243445759210225189599035774915218558382202665746858;
            6'd54: xpb[16] = 1024'd102006084876477757372553021964010270905959540128315439689766952154007219365327897328112976415787685941906326149830722640341526238550155503913167211648702218461296687659155531915998637485433438061463513524607381440681050569359323599364887030030742878782721448032278364501064553986888248417104712183093730749124;
            6'd55: xpb[16] = 1024'd71729646826454264368652430080614126692629569024019437132284007362235565377235303857518568627094727527271182343264534021012537950897804963545406572045370137820363858838510318752835216907733300245965749580296011507191791285401300798954797901409734185987300018406993911761797390300812088901872176157359201267059;
            6'd56: xpb[16] = 1024'd41453208776430771364751838197217982479299597919723434574801062570463911389142710386924160838401769112636038536698345401683549663245454423177645932442038057179431030017865105589671796330033162430467985635984641573702532001443277998544708772788725493191878588781709459022530226614735929386639640131624671784994;
            6'd57: xpb[16] = 1024'd11176770726407278360851246313821838265969626815427432017318117778692257401050116916329753049708810698000894730132156782354561375593103882809885292838705976538498201197219892426508375752333024614970221691673271640213272717485255198134619644167716800396457159156425006283263062928659769871407104105890142302929;
            6'd58: xpb[16] = 1024'd104967028360508526755749581835240126797338082836867113587967028051897498750266662355750416475673526592808900331023461597604636928781973676997284778251704936831256046946145896600975194366150092520782655355749141553088374283748129170689509085229937556867855632945257611574102427316512243373293257906781207305195;
            6'd59: xpb[16] = 1024'd74690590310485033751848989951843982584008111732571111030484083260125844762174068885156008686980568178173756524457272978275648641129623136629524138648372856190323218125500683437811773788449954705284891411437771619599114999790106370279419956608928864072434203319973158834835263630436083858060721881046677823130;
            6'd60: xpb[16] = 1024'd44414152260461540747948398068447838370678140628275108473001138468354190774081475414561600898287609763538612717891084358946660353477272596261763499045040775549390389304855470274648353210749816889787127467126401686109855715832083569869330827987920171277012773694688706095568099944359924342828185855312148341065;
            6'd61: xpb[16] = 1024'd14137714210438047744047806185051694157348169523979105915518193676582536785988881943967193109594651348903468911324895739617672065824922055894002859441708694908457560484210257111484932633049679074289363522815031752620596431874060769459241699366911478481591344069404253356300936258283764827595649829577618859000;
            6'd62: xpb[16] = 1024'd107927971844539296138946141706469982688716625545418787486167103949787778135205427383387856535559367243711474512216200554867747619013791850081402344854707655201215406233136261285951751246866746980101797186890901665495697998136934742014131140429132234952989817858236858647140300646136238329481803630468683861266;
            6'd63: xpb[16] = 1024'd77651533794515803135045549823073838475386654441122784928684159158016124147112833912793448746866408829076330705650011935538759331361441309713641705251375574560282577412491048122788330669166609164604033242579531732006438714178911941604042011808123542157568388232952405907873136960060078814249267604734154379201;
        endcase
    end

    always_comb begin
        case(flag[5][16:12])
            5'd0: xpb[17] = 1024'd0;
            5'd1: xpb[17] = 1024'd47375095744492310131144957939677694262056683336826782371201214366244470159020240442199040958173450414441186899083823316209771043709090769345881065648043493919349748591845834959624910091466471349106269298268161798517179430220889141193952883187114849362146958607667953168605973273983919299016731578999624897136;
            5'd2: xpb[17] = 1024'd94750191488984620262289915879355388524113366673653564742402428732488940318040480884398081916346900828882373798167646632419542087418181538691762131296086987838699497183691669919249820182932942698212538596536323597034358860441778282387905766374229698724293917215335906337211946547967838598033463157999249794272;
            5'd3: xpb[17] = 1024'd18058591549352188994635946414218650041471622884744662985471788033756515139751582416582051659862676933880411289793976514050249290286051973482483071927799440824358571205966287541244491082882208326008610286417245549187177440441770650616880079878115098819620972408886801475711391748023124879931504910373280207077;
            5'd4: xpb[17] = 1024'd65433687293844499125780904353896344303528306221571445356673002400000985298771822858781092618036127348321598188877799830260020333995142742828364137575842934743708319797812122500869401174348679675114879584685407347704356870662659791810832963065229948181767931016554754644317365022007044178948236489372905104213;
            5'd5: xpb[17] = 1024'd112808783038336809256925862293574038565584989558398227727874216766245455457792063300980133576209577762762785087961623146469791377704233512174245203223886428663058068389657957460494311265815151024221148882953569146221536300883548933004785846252344797543914889624222707812923338295990963477964968068372530001349;
            5'd6: xpb[17] = 1024'd36117183098704377989271892828437300082943245769489325970943576067513030279503164833164103319725353867760822579587953028100498580572103946964966143855598881648717142411932575082488982165764416652017220572834491098374354880883541301233760159756230197639241944817773602951422783496046249759863009820746560414154;
            5'd7: xpb[17] = 1024'd83492278843196688120416850768114994344999929106316108342144790433757500438523405275363144277898804282202009478671776344310269624281194716310847209503642375568066891003778410042113892257230888001123489871102652896891534311104430442427713042943345047001388903425441556120028756770030169058879741399746185311290;
            5'd8: xpb[17] = 1024'd6800678903564256852762881302978255862358185317407206585214149735025075260234506807547114021414580387200046970298106225940976827149065151101568150135354828553725965026053027664108563157180153628919561560983574849044352891104422810656687356447230447096715958618992451258528201970085455340777783152120215724095;
            5'd9: xpb[17] = 1024'd54175774648056566983907839242655950124414868654233988956415364101269545419254747249746154979588030801641233869381929542150747870858155920447449215783398322473075713617898862623733473248646624978025830859251736647561532321325311951850640239634345296458862917226660404427134175244069374639794514731119840621231;
            5'd10: xpb[17] = 1024'd101550870392548877115052797182333644386471551991060771327616578467514015578274987691945195937761481216082420768465752858360518914567246689793330281431441816392425462209744697583358383340113096327132100157519898446078711751546201093044593122821460145821009875834328357595740148518053293938811246310119465518367;
            5'd11: xpb[17] = 1024'd24859270452916445847398827717196905903829808202151869570685937768781590399986089224129165681277257321080458260092082739991226117435117124584051222063154269378084536232019315205353054240062361954928171847400820398231530331546193461273567436325345545916336931027879252734239593718108580220709288062493495931172;
            5'd12: xpb[17] = 1024'd72234366197408755978543785656874600165886491538978651941887152135026060559006329666328206639450707735521645159175906056200997161144207893929932287711197763297434284823865150164977964331528833304034441145668982196748709761767082602467520319512460395278483889635547205902845566992092499519726019641493120828308;
            5'd13: xpb[17] = 1024'd119609461941901066109688743596552294427943174875805434313088366501270530718026570108527247597624158149962832058259729372410768204853298663275813353359241257216784033415710985124602874422995304653140710443937143995265889191987971743661473202699575244640630848243215159071451540266076418818742751220492745725444;
            5'd14: xpb[17] = 1024'd42917862002268634842034774131415555945301431086896532556157725802538105539737671640711217341139934254960869549886059254041475407721169098066534293990953710202443107437985602746597545322944570280936782133818065947418707771987964111890447516203460644735957903436766054209950985466131705100640792972866776138249;
            5'd15: xpb[17] = 1024'd90292957746760944973179732071093250207358114423723314927358940168782575698757912082910258299313384669402056448969882570251246451430259867412415359638997204121792856029831437706222455414411041630043051432086227745935887202208853253084400399390575494098104862044434007378556958740115624399657524551866401035385;
            5'd16: xpb[17] = 1024'd13601357807128513705525762605956511724716370634814413170428299470050150520469013615094228042829160774400093940596212451881953654298130302203136300270709657107451930052106055328217126314360307257839123121967149698088705782208845621313374712894460894193431917237984902517056403940170910681555566304240431448190;
            5'd17: xpb[17] = 1024'd60976453551620823836670720545634205986773053971641195541629513836294620679489254057293269001002611188841280839680035768091724698007221071549017365918753151026801678643951890287842036405826778606945392420235311496605885212429734762507327596081575743555578875845652855685662377214154829980572297883240056345326;
            5'd18: xpb[17] = 1024'd108351549296113133967815678485311900248829737308467977912830728202539090838509494499492309959176061603282467738763859084301495741716311840894898431566796644946151427235797725247466946497293249956051661718503473295123064642650623903701280479268690592917725834453320808854268350488138749279589029462239681242462;
            5'd19: xpb[17] = 1024'd31659949356480702700161709020175161766187993519559076155900087503806665660220596031676279702691837708280505230390188965932202944584182275685619372198509097931810501258072342869461617397242515583847733408384395247275883222650616271930254792772575993013052889646871703992767795688194035561487071214613711655267;
            5'd20: xpb[17] = 1024'd79035045100973012831306666959852856028244676856385858527101301870051135819240836473875320660865288122721692129474012282141973988293273045031500437846552591851160249849918177829086527488708986932954002706652557045793062652871505413124207675959690842375199848254539657161373768962177954860503802793613336552403;
            5'd21: xpb[17] = 1024'd2343445161340581563652697494716117545602933067476956770170661171318710640951938006059290404381064227719729621100342163772681191161143479822221378478265044836819323872192795451081198388658252560750074396533478997945881232871497781353181989463576242470526903448090552299873214162233241142401844545987366965208;
            5'd22: xpb[17] = 1024'd49718540905832891694797655434393811807659616404303739141371875537563180799972178448258331362554514642160916520184165479982452234870234249168102444126308538756169072464038630410706108480124723909856343694801640796463060663092386922547134872650691091832673862055758505468479187436217160441418576124986991862344;
            5'd23: xpb[17] = 1024'd97093636650325201825942613374071506069716299741130521512573089903807650958992418890457372320727965056602103419267988796192223278579325018513983509774352032675518821055884465370331018571591195258962612993069802594980240093313276063741087755837805941194820820663426458637085160710201079740435307703986616759480;
            5'd24: xpb[17] = 1024'd20402036710692770558288643908934767587074555952221619755642449205075225780703520422641342064243741161600140910894318677822930481447195453304704450406064485661177895078159082992325689471540460886758684682950724547133058673313268431970062069341691341290147875856977353775584605910256366022333349456360647172285;
            5'd25: xpb[17] = 1024'd67777132455185080689433601848612461849131239289048402126843663571319695939723760864840383022417191576041327809978141994032701525156286222650585516054107979580527643670004917951950599563006932235864953981218886345650238103534157573164014952528806190652294834464645306944190579184240285321350081035360272069421;
            5'd26: xpb[17] = 1024'd115152228199677390820578559788290156111187922625875184498044877937564166098744001307039423980590641990482514709061965310242472568865376991996466581702151473499877392261850752911575509654473403584971223279487048144167417533755046714357967835715921040014441793072313260112796552458224204620366812614359896966557;
            5'd27: xpb[17] = 1024'd38460628260044959552924590323153417628546178836966282741114237238831740920455102839223393724106418095480552200688295191873179771733247426787187522333863926485536466284125370533570180554422669212767294969367970096320236113755039082586942149219806440109768848265864155251295997658279490902264854366733927379362;
            5'd28: xpb[17] = 1024'd85835724004537269684069548262831111890602862173793065112315451605076211079475343281422434682279868509921739099772118508082950815442338196133068587981907420404886214875971205493195090645889140561873564267636131894837415543975928223780895032406921289471915806873532108419901970932263410201281585945733552276498;
            5'd29: xpb[17] = 1024'd9144124064904838416415578797694373407961118384884163355384810906343785901186444813606404425795644614919776591398448389713658018310208630923789528613619873390545288898245823115189761545838406189669635957517053846990234123975920592009869345910806689567242862067083003558401416132318696483179627698107582689303;
            5'd30: xpb[17] = 1024'd56519219809397148547560536737372067670017801721710945726586025272588256060206685255805445383969095029360963490482271705923429062019299400269670594261663367309895037490091658074814671637304877538775905255785215645507413554196809733203822229097921538929389820674750956727007389406302615782196359277107207586439;
            5'd31: xpb[17] = 1024'd103894315553889458678705494677049761932074485058537728097787239638832726219226925698004486342142545443802150389566095022133200105728390169615551659909706861229244786081937493034439581728771348887882174554053377444024592984417698874397775112285036388291536779282418909895613362680286535081213090856106832483575;
        endcase
    end

    always_comb begin
        case(flag[6][5:0])
            6'd0: xpb[18] = 1024'd0;
            6'd1: xpb[18] = 1024'd13601357807128513705525762605956511724716370634814413170428299470050150520469013615094228042829160774400093940596212451881953654298130302203136300270709657107451930052106055328217126314360307257839123121967149698088705782208845621313374712894460894193431917237984902517056403940170910681555566304240431448190;
            6'd2: xpb[18] = 1024'd27202715614257027411051525211913023449432741269628826340856598940100301040938027230188456085658321548800187881192424903763907308596260604406272600541419314214903860104212110656434252628720614515678246243934299396177411564417691242626749425788921788386863834475969805034112807880341821363111132608480862896380;
            6'd3: xpb[18] = 1024'd40804073421385541116577287817869535174149111904443239511284898410150451561407040845282684128487482323200281821788637355645860962894390906609408900812128971322355790156318165984651378943080921773517369365901449094266117346626536863940124138683382682580295751713954707551169211820512732044666698912721294344570;
            6'd4: xpb[18] = 1024'd54405431228514054822103050423826046898865482539257652681713197880200602081876054460376912171316643097600375762384849807527814617192521208812545201082838628429807720208424221312868505257441229031356492487868598792354823128835382485253498851577843576773727668951939610068225615760683642726222265216961725792760;
            6'd5: xpb[18] = 1024'd68006789035642568527628813029782558623581853174072065852141497350250752602345068075471140214145803872000469702981062259409768271490651511015681501353548285537259650260530276641085631571801536289195615609835748490443528911044228106566873564472304470967159586189924512585282019700854553407777831521202157240950;
            6'd6: xpb[18] = 1024'd81608146842771082233154575635739070348298223808886479022569796820300903122814081690565368256974964646400563643577274711291721925788781813218817801624257942644711580312636331969302757886161843547034738731802898188532234693253073727880248277366765365160591503427909415102338423641025464089333397825442588689140;
            6'd7: xpb[18] = 1024'd95209504649899595938680338241695582073014594443700892192998096290351053643283095305659596299804125420800657584173487163173675580086912115421954101894967599752163510364742387297519884200522150804873861853770047886620940475461919349193622990261226259354023420665894317619394827581196374770888964129683020137330;
            6'd8: xpb[18] = 1024'd108810862457028109644206100847652093797730965078515305363426395760401204163752108920753824342633286195200751524769699615055629234385042417625090402165677256859615440416848442625737010514882458062712984975737197584709646257670764970506997703155687153547455337903879220136451231521367285452444530433923451585520;
            6'd9: xpb[18] = 1024'd122412220264156623349731863453608605522447335713329718533854695230451354684221122535848052385462446969600845465365912066937582888683172719828226702436386913967067370468954497953954136829242765320552108097704347282798352039879610591820372416050148047740887255141864122653507635461538196134000096738163883033710;
            6'd10: xpb[18] = 1024'd11946882387160395656458698654750684502465279222408447576151139635524609867380997240927209213633933434557789998504631084240472702140082687476202877690765530140828625951489335944541023952085866857081033611284257134522696971867559440168768559261379492667499268965731967140457511327780473798436973215778719997569;
            6'd11: xpb[18] = 1024'd25548240194288909361984461260707196227181649857222860746579439105574760387850010856021437256463094208957883939100843536122426356438212989679339177961475187248280556003595391272758150266446174114920156733251406832611402754076405061482143272155840386860931186203716869657513915267951384479992539520019151445759;
            6'd12: xpb[18] = 1024'd39149598001417423067510223866663707951898020492037273917007738575624910908319024471115665299292254983357977879697055988004380010736343291882475478232184844355732486055701446600975276580806481372759279855218556530700108536285250682795517985050301281054363103441701772174570319208122295161548105824259582893949;
            6'd13: xpb[18] = 1024'd52750955808545936773035986472620219676614391126851687087436038045675061428788038086209893342121415757758071820293268439886333665034473594085611778502894501463184416107807501929192402895166788630598402977185706228788814318494096304108892697944762175247795020679686674691626723148293205843103672128500014342139;
            6'd14: xpb[18] = 1024'd66352313615674450478561749078576731401330761761666100257864337515725211949257051701304121384950576532158165760889480891768287319332603896288748078773604158570636346159913557257409529209527095888437526099152855926877520100702941925422267410839223069441226937917671577208683127088464116524659238432740445790329;
            6'd15: xpb[18] = 1024'd79953671422802964184087511684533243126047132396480513428292636985775362469726065316398349427779737306558259701485693343650240973630734198491884379044313815678088276212019612585626655523887403146276649221120005624966225882911787546735642123733683963634658855155656479725739531028635027206214804736980877238519;
            6'd16: xpb[18] = 1024'd93555029229931477889613274290489754850763503031294926598720936455825512990195078931492577470608898080958353642081905795532194627928864500695020679315023472785540206264125667913843781838247710404115772343087155323054931665120633168049016836628144857828090772393641382242795934968805937887770371041221308686709;
            6'd17: xpb[18] = 1024'd107156387037059991595139036896446266575479873666109339769149235925875663510664092546586805513438058855358447582678118247414148282226994802898156979585733129892992136316231723242060908152608017661954895465054305021143637447329478789362391549522605752021522689631626284759852338908976848569325937345461740134899;
            6'd18: xpb[18] = 1024'd120757744844188505300664799502402778300196244300923752939577535395925814031133106161681033556267219629758541523274330699296101936525125105101293279856442787000444066368337778570278034466968324919794018587021454719232343229538324410675766262417066646214954606869611187276908742849147759250881503649702171583089;
            6'd19: xpb[18] = 1024'd10292406967192277607391634703544857280214187810002481981873979800999069214292980866760190384438706094715486056413049716598991749982035072749269455110821403174205321850872616560864921589811426456322944100601364570956688161526273259024162405628298091141566620693479031763858618715390036915318380127317008546948;
            6'd20: xpb[18] = 1024'd23893764774320791312917397309501369004930558444816895152302279271049219734761994481854418427267866869115579997009262168480945404280165374952405755381531060281657251902978671889082047904171733714162067222568514269045393943735118880337537118522758985334998537931463934280915022655560947596873946431557439995138;
            6'd21: xpb[18] = 1024'd37495122581449305018443159915457880729646929079631308322730578741099370255231008096948646470097027643515673937605474620362899058578295677155542055652240717389109181955084727217299174218532040972001190344535663967134099725943964501650911831417219879528430455169448836797971426595731858278429512735797871443328;
            6'd22: xpb[18] = 1024'd51096480388577818723968922521414392454363299714445721493158878211149520775700021712042874512926188417915767878201687072244852712876425979358678355922950374496561112007190782545516300532892348229840313466502813665222805508152810122964286544311680773721862372407433739315027830535902768959985079040038302891518;
            6'd23: xpb[18] = 1024'd64697838195706332429494685127370904179079670349260134663587177681199671296169035327137102555755349192315861818797899524126806367174556281561814656193660031604013042059296837873733426847252655487679436588469963363311511290361655744277661257206141667915294289645418641832084234476073679641540645344278734339708;
            6'd24: xpb[18] = 1024'd78299196002834846135020447733327415903796040984074547834015477151249821816638048942231330598584509966715955759394111976008760021472686583764950956464369688711464972111402893201950553161612962745518559710437113061400217072570501365591035970100602562108726206883403544349140638416244590323096211648519165787898;
            6'd25: xpb[18] = 1024'd91900553809963359840546210339283927628512411618888961004443776621299972337107062557325558641413670741116049699990324427890713675770816885968087256735079345818916902163508948530167679475973270003357682832404262759488922854779346986904410682995063456302158124121388446866197042356415501004651777952759597236088;
            6'd26: xpb[18] = 1024'd105501911617091873546071972945240439353228782253703374174872076091350122857576076172419786684242831515516143640586536879772667330068947188171223557005789002926368832215615003858384805790333577261196805954371412457577628636988192608217785395889524350495590041359373349383253446296586411686207344257000028684278;
            6'd27: xpb[18] = 1024'd119103269424220387251597735551196951077945152888517787345300375561400273378045089787514014727071992289916237581182749331654620984367077490374359857276498660033820762267721059186601932104693884519035929076338562155666334419197038229531160108783985244689021958597358251900309850236757322367762910561240460132468;
            6'd28: xpb[18] = 1024'd8637931547224159558324570752339030057963096397596516387596819966473528561204964492593171555243478754873182114321468348957510797823987458022336032530877276207582017750255897177188819227536986055564854589918472007390679351184987077879556251995216689615633972421226096387259726102999600032199787038855297096327;
            6'd29: xpb[18] = 1024'd22239289354352673263850333358295541782679467032410929558025119436523679081673978107687399598072639529273276054917680800839464452122117760225472332801586933315033947802361952505405945541897293313403977711885621705479385133393832699192930964889677583809065889659210998904316130043170510713755353343095728544517;
            6'd30: xpb[18] = 1024'd35840647161481186969376095964252053507395837667225342728453418906573829602142991722781627640901800303673369995513893252721418106420248062428608633072296590422485877854468007833623071856257600571243100833852771403568090915602678320506305677784138478002497806897195901421372533983341421395310919647336159992707;
            6'd31: xpb[18] = 1024'd49442004968609700674901858570208565232112208302039755898881718376623980122612005337875855683730961078073463936110105704603371760718378364631744933343006247529937807906574063161840198170617907829082223955819921101656796697811523941819680390678599372195929724135180803938428937923512332076866485951576591440897;
            6'd32: xpb[18] = 1024'd63043362775738214380427621176165076956828578936854169069310017846674130643081018952970083726560121852473557876706318156485325415016508666834881233613715904637389737958680118490057324484978215086921347077787070799745502480020369563133055103573060266389361641373165706455485341863683242758422052255817022889087;
            6'd33: xpb[18] = 1024'd76644720582866728085953383782121588681544949571668582239738317316724281163550032568064311769389282626873651817302530608367279069314638969038017533884425561744841668010786173818274450799338522344760470199754220497834208262229215184446429816467521160582793558611150608972541745803854153439977618560057454337277;
            6'd34: xpb[18] = 1024'd90246078389995241791479146388078100406261320206482995410166616786774431684019046183158539812218443401273745757898743060249232723612769271241153834155135218852293598062892229146491577113698829602599593321721370195922914044438060805759804529361982054776225475849135511489598149744025064121533184864297885785467;
            6'd35: xpb[18] = 1024'd103847436197123755497004908994034612130977690841297408580594916256824582204488059798252767855047604175673839698494955512131186377910899573444290134425844875959745528114998284474708703428059136860438716443688519894011619826646906427073179242256442948969657393087120414006654553684195974803088751168538317233657;
            6'd36: xpb[18] = 1024'd117448794004252269202530671599991123855694061476111821751023215726874732724957073413346995897876764950073933639091167964013140032209029875647426434696554533067197458167104339802925829742419444118277839565655669592100325608855752048386553955150903843163089310325105316523710957624366885484644317472778748681847;
            6'd37: xpb[18] = 1024'd6983456127256041509257506801133202835712004985190550793319660131947987908116948118426152726048251415030878172229886981316029845665939843295402609950933149240958713649639177793512716865262545654806765079235579443824670540843700896734950098362135288089701324148973161010660833490609163149081193950393585645706;
            6'd38: xpb[18] = 1024'd20584813934384555214783269407089714560428375620004963963747959601998138428585961733520380768877412189430972112826099433197983499964070145498538910221642806348410643701745233121729843179622852912645888201202729141913376323052546518048324811256596182283133241386958063527717237430780073830636760254634017093896;
            6'd39: xpb[18] = 1024'd34186171741513068920309032013046226285144746254819377134176259072048288949054975348614608811706572963831066053422311885079937154262200447701675210492352463455862573753851288449946969493983160170485011323169878840002082105261392139361699524151057076476565158624942966044773641370950984512192326558874448542086;
            6'd40: xpb[18] = 1024'd47787529548641582625834794619002738009861116889633790304604558542098439469523988963708836854535733738231159994018524336961890808560330749904811510763062120563314503805957343778164095808343467428324134445137028538090787887470237760675074237045517970669997075862927868561830045311121895193747892863114879990276;
            6'd41: xpb[18] = 1024'd61388887355770096331360557224959249734577487524448203475032858012148589989993002578803064897364894512631253934614736788843844462858461052107947811033771777670766433858063399106381222122703774686163257567104178236179493669679083381988448949939978864863428993100912771078886449251292805875303459167355311438466;
            6'd42: xpb[18] = 1024'd74990245162898610036886319830915761459293858159262616645461157482198740510462016193897292940194055287031347875210949240725798117156591354311084111304481434778218363910169454434598348437064081944002380689071327934268199451887929003301823662834439759056860910338897673595942853191463716556859025471595742886656;
            6'd43: xpb[18] = 1024'd88591602970027123742412082436872273184010228794077029815889456952248891030931029808991520983023216061431441815807161692607751771454721656514220411575191091885670293962275509762815474751424389201841503811038477632356905234096774624615198375728900653250292827576882576112999257131634627238414591775836174334846;
            6'd44: xpb[18] = 1024'd102192960777155637447937845042828784908726599428891442986317756422299041551400043424085749025852376835831535756403374144489705425752851958717356711845900748993122224014381565091032601065784696459680626933005627330445611016305620245928573088623361547443724744814867478630055661071805537919970158080076605783036;
            6'd45: xpb[18] = 1024'd115794318584284151153463607648785296633442970063705856156746055892349192071869057039179977068681537610231629696999586596371659080050982260920493012116610406100574154066487620419249727380145003717519750054972777028534316798514465867241947801517822441637156662052852381147112065011976448601525724384317037231226;
            6'd46: xpb[18] = 1024'd5328980707287923460190442849927375613460913572784585199042500297422447255028931744259133896853024075188574230138305613674548893507892228568469187370989022274335409549022458409836614502988105254048675568552686880258661730502414715590343944729053886563768675876720225634061940878218726265962600861931874195085;
            6'd47: xpb[18] = 1024'd18930338514416437165716205455883887338177284207598998369470799767472597775497945359353361939682184849588668170734518065556502547806022530771605487641698679381787339601128513738053740817348412511887798690519836578347367512711260336903718657623514780757200593114705128151118344818389636947518167166172305643275;
            6'd48: xpb[18] = 1024'd32531696321544950871241968061840399062893654842413411539899099237522748295966958974447589982511345623988762111330730517438456202104152832974741787912408336489239269653234569066270867131708719769726921812486986276436073294920105958217093370517975674950632510352690030668174748758560547629073733470412737091465;
            6'd49: xpb[18] = 1024'd46133054128673464576767730667796910787610025477227824710327398707572898816435972589541818025340506398388856051926942969320409856402283135177878088183117993596691199705340624394487993446069027027566044934454135974524779077128951579530468083412436569144064427590674933185231152698731458310629299774653168539655;
            6'd50: xpb[18] = 1024'd59734411935801978282293493273753422512326396112042237880755698177623049336904986204636046068169667172788949992523155421202363510700413437381014388453827650704143129757446679722705119760429334285405168056421285672613484859337797200843842796306897463337496344828659835702287556638902368992184866078893599987845;
            6'd51: xpb[18] = 1024'd73335769742930491987819255879709934237042766746856651051183997647673199857373999819730274110998827947189043933119367873084317164998543739584150688724537307811595059809552735050922246074789641543244291178388435370702190641546642822157217509201358357530928262066644738219343960579073279673740432383134031436035;
            6'd52: xpb[18] = 1024'd86937127550059005693345018485666445961759137381671064221612297117723350377843013434824502153827988721589137873715580324966270819296674041787286988995246964919046989861658790379139372389149948801083414300355585068790896423755488443470592222095819251724360179304629640736400364519244190355295998687374462884225;
            6'd53: xpb[18] = 1024'd100538485357187519398870781091622957686475508016485477392040596587773500898312027049918730196657149495989231814311792776848224473594804343990423289265956622026498919913764845707356498703510256058922537422322734766879602205964334064783966934990280145917792096542614543253456768459415101036851564991614894332415;
            6'd54: xpb[18] = 1024'd114139843164316033104396543697579469411191878651299890562468896057823651418781040665012958239486310270389325754908005228730178127892934646193559589536666279133950849965870901035573625017870563316761660544289884464968307988173179686097341647884741040111224013780599445770513172399586011718407131295855325780605;
            6'd55: xpb[18] = 1024'd3674505287319805411123378898721548391209822160378619604765340462896906601940915370092115067657796735346270288046724246033067941349844613841535764791044895307712105448405739026160512140713664853290586057869794316692652920161128534445737791095972485037836027604467290257463048265828289382844007773470162744464;
            6'd56: xpb[18] = 1024'd17275863094448319116649141504678060115926192795193032775193639932947057122409928985186343110486957509746364228642936697915021595647974916044672065061754552415164035500511794354377638455073972111129709179836944014781358702369974155759112503990433379231267944842452192774519452205999200064399574077710594192654;
            6'd57: xpb[18] = 1024'd30877220901576832822174904110634571840642563430007445945621939402997207642878942600280571153316118284146458169239149149796975249946105218247808365332464209522615965552617849682594764769434279368968832301804093712870064484578819777072487216884894273424699862080437095291575856146170110745955140381951025640844;
            6'd58: xpb[18] = 1024'd44478578708705346527700666716591083565358934064821859116050238873047358163347956215374799196145279058546552109835361601678928904244235520450944665603173866630067895604723905010811891083794586626807955423771243410958770266787665398385861929779355167618131779318421997808632260086341021427510706686191457089034;
            6'd59: xpb[18] = 1024'd58079936515833860233226429322547595290075304699636272286478538343097508683816969830469027238974439832946646050431574053560882558542365822654080965873883523737519825656829960339029017398154893884647078545738393109047476048996511019699236642673816061811563696556406900325688664026511932109066272990431888537224;
            6'd60: xpb[18] = 1024'd71681294322962373938752191928504107014791675334450685456906837813147659204285983445563255281803600607346739991027786505442836212840496124857217266144593180844971755708936015667246143712515201142486201667705542807136181831205356641012611355568276956004995613794391802842745067966682842790621839294672319985414;
            6'd61: xpb[18] = 1024'd85282652130090887644277954534460618739508045969265098627335137283197809724754997060657483324632761381746833931623998957324789867138626427060353566415302837952423685761042070995463270026875508400325324789672692505224887613414202262325986068462737850198427531032376705359801471906853753472177405598912751433604;
            6'd62: xpb[18] = 1024'd98884009937219401349803717140417130464224416604079511797763436753247960245224010675751711367461922156146927872220211409206743521436756729263489866686012495059875615813148126323680396341235815658164447911639842203313593395623047883639360781357198744391859448270361607876857875847024664153732971903153182881794;
            6'd63: xpb[18] = 1024'd112485367744347915055329479746373642188940787238893924968191736223298110765693024290845939410291082930547021812816423861088697175734887031466626166956722152167327545865254181651897522655596122916003571033606991901402299177831893504952735494251659638585291365508346510393914279787195574835288538207393614329984;
        endcase
    end

    always_comb begin
        case(flag[6][11:6])
            6'd0: xpb[19] = 1024'd0;
            6'd1: xpb[19] = 1024'd2020029867351687362056314947515721168958730747972654010488180628371365948852898995925096238462569395503966345955142878391586989191796999114602342211100768341088801347789019642484409778439224452532496547186901753126644109819842353301131637462891083511903379332214354880864155653437852499725414685008451293843;
            6'd2: xpb[19] = 1024'd4040059734703374724112629895031442337917461495945308020976361256742731897705797991850192476925138791007932691910285756783173978383593998229204684422201536682177602695578039284968819556878448905064993094373803506253288219639684706602263274925782167023806758664428709761728311306875704999450829370016902587686;
            6'd3: xpb[19] = 1024'd6060089602055062086168944842547163506876192243917962031464541885114097846558696987775288715387708186511899037865428635174760967575390997343807026633302305023266404043367058927453229335317673357597489641560705259379932329459527059903394912388673250535710137996643064642592466960313557499176244055025353881529;
            6'd4: xpb[19] = 1024'd8080119469406749448225259790062884675834922991890616041952722513485463795411595983700384953850277582015865383820571513566347956767187996458409368844403073364355205391156078569937639113756897810129986188747607012506576439279369413204526549851564334047613517328857419523456622613751409998901658740033805175372;
            6'd5: xpb[19] = 1024'd10100149336758436810281574737578605844793653739863270052440903141856829744264494979625481192312846977519831729775714391957934945958984995573011711055503841705444006738945098212422048892196122262662482735934508765633220549099211766505658187314455417559516896661071774404320778267189262498627073425042256469215;
            6'd6: xpb[19] = 1024'd12120179204110124172337889685094327013752384487835924062929083770228195693117393975550577430775416373023798075730857270349521935150781994687614053266604610046532808086734117854906458670635346715194979283121410518759864658919054119806789824777346501071420275993286129285184933920627114998352488110050707763058;
            6'd7: xpb[19] = 1024'd14140209071461811534394204632610048182711115235808578073417264398599561641970292971475673669237985768527764421686000148741108924342578993802216395477705378387621609434523137497390868449074571167727475830308312271886508768738896473107921462240237584583323655325500484166049089574064967498077902795059159056901;
            6'd8: xpb[19] = 1024'd16160238938813498896450519580125769351669845983781232083905445026970927590823191967400769907700555164031730767641143027132695913534375992916818737688806146728710410782312157139875278227513795620259972377495214025013152878558738826409053099703128668095227034657714839046913245227502819997803317480067610350744;
            6'd9: xpb[19] = 1024'd18180268806165186258506834527641490520628576731753886094393625655342293539676090963325866146163124559535697113596285905524282902726172992031421079899906915069799212130101176782359688005953020072792468924682115778139796988378581179710184737166019751607130413989929193927777400880940672497528732165076061644587;
            6'd10: xpb[19] = 1024'd20200298673516873620563149475157211689587307479726540104881806283713659488528989959250962384625693955039663459551428783915869891917969991146023422111007683410888013477890196424844097784392244525324965471869017531266441098198423533011316374628910835119033793322143548808641556534378524997254146850084512938430;
            6'd11: xpb[19] = 1024'd22220328540868560982619464422672932858546038227699194115369986912085025437381888955176058623088263350543629805506571662307456881109766990260625764322108451751976814825679216067328507562831468977857462019055919284393085208018265886312448012091801918630937172654357903689505712187816377496979561535092964232273;
            6'd12: xpb[19] = 1024'd24240358408220248344675779370188654027504768975671848125858167540456391386234787951101154861550832746047596151461714540699043870301563989375228106533209220093065616173468235709812917341270693430389958566242821037519729317838108239613579649554693002142840551986572258570369867841254229996704976220101415526116;
            6'd13: xpb[19] = 1024'd26260388275571935706732094317704375196463499723644502136346348168827757335087686947026251100013402141551562497416857419090630859493360988489830448744309988434154417521257255352297327119709917882922455113429722790646373427657950592914711287017584085654743931318786613451234023494692082496430390905109866819959;
            6'd14: xpb[19] = 1024'd28280418142923623068788409265220096365422230471617156146834528797199123283940585942951347338475971537055528843372000297482217848685157987604432790955410756775243218869046274994781736898149142335454951660616624543773017537477792946215842924480475169166647310651000968332098179148129934996155805590118318113802;
            6'd15: xpb[19] = 1024'd30300448010275310430844724212735817534380961219589810157322709425570489232793484938876443576938540932559495189327143175873804837876954986719035133166511525116332020216835294637266146676588366787987448207803526296899661647297635299516974561943366252678550689983215323212962334801567787495881220275126769407645;
            6'd16: xpb[19] = 1024'd32320477877626997792901039160251538703339691967562464167810890053941855181646383934801539815401110328063461535282286054265391827068751985833637475377612293457420821564624314279750556455027591240519944754990428050026305757117477652818106199406257336190454069315429678093826490455005639995606634960135220701488;
            6'd17: xpb[19] = 1024'd34340507744978685154957354107767259872298422715535118178299070682313221130499282930726636053863679723567427881237428932656978816260548984948239817588713061798509622912413333922234966233466815693052441302177329803152949866937320006119237836869148419702357448647644032974690646108443492495332049645143671995331;
            6'd18: xpb[19] = 1024'd36360537612330372517013669055282981041257153463507772188787251310684587079352181926651732292326249119071394227192571811048565805452345984062842159799813830139598424260202353564719376011906040145584937849364231556279593976757162359420369474332039503214260827979858387855554801761881344995057464330152123289174;
            6'd19: xpb[19] = 1024'd38380567479682059879069984002798702210215884211480426199275431939055953028205080922576828530788818514575360573147714689440152794644142983177444502010914598480687225607991373207203785790345264598117434396551133309406238086577004712721501111794930586726164207312072742736418957415319197494782879015160574583017;
            6'd20: xpb[19] = 1024'd40400597347033747241126298950314423379174614959453080209763612567427318977057979918501924769251387910079326919102857567831739783835939982292046844222015366821776026955780392849688195568784489050649930943738035062532882196396847066022632749257821670238067586644287097617283113068757049994508293700169025876860;
            6'd21: xpb[19] = 1024'd42420627214385434603182613897830144548133345707425734220251793195798684925910878914427021007713957305583293265058000446223326773027736981406649186433116135162864828303569412492172605347223713503182427490924936815659526306216689419323764386720712753749970965976501452498147268722194902494233708385177477170703;
            6'd22: xpb[19] = 1024'd44440657081737121965238928845345865717092076455398388230739973824170050874763777910352117246176526701087259611013143324614913762219533980521251528644216903503953629651358432134657015125662937955714924038111838568786170416036531772624896024183603837261874345308715807379011424375632754993959123070185928464546;
            6'd23: xpb[19] = 1024'd46460686949088809327295243792861586886050807203371042241228154452541416823616676906277213484639096096591225956968286203006500751411330979635853870855317671845042430999147451777141424904102162408247420585298740321912814525856374125926027661646494920773777724640930162259875580029070607493684537755194379758389;
            6'd24: xpb[19] = 1024'd48480716816440496689351558740377308055009537951343696251716335080912782772469575902202309723101665492095192302923429081398087740603127978750456213066418440186131232346936471419625834682541386860779917132485642075039458635676216479227159299109386004285681103973144517140739735682508459993409952440202831052232;
            6'd25: xpb[19] = 1024'd50500746683792184051407873687893029223968268699316350262204515709284148721322474898127405961564234887599158648878571959789674729794924977865058555277519208527220033694725491062110244460980611313312413679672543828166102745496058832528290936572277087797584483305358872021603891335946312493135367125211282346075;
            6'd26: xpb[19] = 1024'd52520776551143871413464188635408750392926999447289004272692696337655514670175373894052502200026804283103124994833714838181261718986721976979660897488619976868308835042514510704594654239419835765844910226859445581292746855315901185829422574035168171309487862637573226902468046989384164992860781810219733639918;
            6'd27: xpb[19] = 1024'd54540806418495558775520503582924471561885730195261658283180876966026880619028272889977598438489373678607091340788857716572848708178518976094263239699720745209397636390303530347079064017859060218377406774046347334419390965135743539130554211498059254821391241969787581783332202642822017492586196495228184933761;
            6'd28: xpb[19] = 1024'd56560836285847246137576818530440192730844460943234312293669057594398246567881171885902694676951943074111057686744000594964435697370315975208865581910821513550486437738092549989563473796298284670909903321233249087546035074955585892431685848960950338333294621302001936664196358296259869992311611180236636227604;
            6'd29: xpb[19] = 1024'd58580866153198933499633133477955913899803191691206966304157238222769612516734070881827790915414512469615024032699143473356022686562112974323467924121922281891575239085881569632047883574737509123442399868420150840672679184775428245732817486423841421845198000634216291545060513949697722492037025865245087521447;
            6'd30: xpb[19] = 1024'd60600896020550620861689448425471635068761922439179620314645418851140978465586969877752887153877081865118990378654286351747609675753909973438070266333023050232664040433670589274532293353176733575974896415607052593799323294595270599033949123886732505357101379966430646425924669603135574991762440550253538815290;
            6'd31: xpb[19] = 1024'd62620925887902308223745763372987356237720653187152274325133599479512344414439868873677983392339651260622956724609429230139196664945706972552672608544123818573752841781459608917016703131615958028507392962793954346925967404415112952335080761349623588869004759298645001306788825256573427491487855235261990109133;
            6'd32: xpb[19] = 1024'd64640955755253995585802078320503077406679383935124928335621780107883710363292767869603079630802220656126923070564572108530783654137503971667274950755224586914841643129248628559501112910055182481039889509980856100052611514234955305636212398812514672380908138630859356187652980910011279991213269920270441402976;
            6'd33: xpb[19] = 1024'd66660985622605682947858393268018798575638114683097582346109960736255076312145666865528175869264790051630889416519714986922370643329300970781877292966325355255930444477037648201985522688494406933572386057167757853179255624054797658937344036275405755892811517963073711068517136563449132490938684605278892696819;
            6'd34: xpb[19] = 1024'd68681015489957370309914708215534519744596845431070236356598141364626442260998565861453272107727359447134855762474857865313957632521097969896479635177426123597019245824826667844469932466933631386104882604354659606305899733874640012238475673738296839404714897295288065949381292216886984990664099290287343990662;
            6'd35: xpb[19] = 1024'd70701045357309057671971023163050240913555576179042890367086321992997808209851464857378368346189928842638822108430000743705544621712894969011081977388526891938108047172615687486954342245372855838637379151541561359432543843694482365539607311201187922916618276627502420830245447870324837490389513975295795284505;
            6'd36: xpb[19] = 1024'd72721075224660745034027338110565962082514306927015544377574502621369174158704363853303464584652498238142788454385143622097131610904691968125684319599627660279196848520404707129438752023812080291169875698728463112559187953514324718840738948664079006428521655959716775711109603523762689990114928660304246578348;
            6'd37: xpb[19] = 1024'd74741105092012432396083653058081683251473037674988198388062683249740540107557262849228560823115067633646754800340286500488718600096488967240286661810728428620285649868193726771923161802251304743702372245915364865685832063334167072141870586126970089940425035291931130591973759177200542489840343345312697872191;
            6'd38: xpb[19] = 1024'd76761134959364119758139968005597404420431768422960852398550863878111906056410161845153657061577637029150721146295429378880305589288285966354889004021829196961374451215982746414407571580690529196234868793102266618812476173154009425443002223589861173452328414624145485472837914830638394989565758030321149166034;
            6'd39: xpb[19] = 1024'd78781164826715807120196282953113125589390499170933506409039044506483272005263060841078753300040206424654687492250572257271892578480082965469491346232929965302463252563771766056891981359129753648767365340289168371939120282973851778744133861052752256964231793956359840353702070484076247489291172715329600459877;
            6'd40: xpb[19] = 1024'd80801194694067494482252597900628846758349229918906160419527225134854637954115959837003849538502775820158653838205715135663479567671879964584093688444030733643552053911560785699376391137568978101299861887476070125065764392793694132045265498515643340476135173288574195234566226137514099989016587400338051753720;
            6'd41: xpb[19] = 1024'd82821224561419181844308912848144567927307960666878814430015405763226003902968858832928945776965345215662620184160858014055066556863676963698696030655131501984640855259349805341860800916008202553832358434662971878192408502613536485346397135978534423988038552620788550115430381790951952488742002085346503047563;
            6'd42: xpb[19] = 1024'd84841254428770869206365227795660289096266691414851468440503586391597369851821757828854042015427914611166586530116000892446653546055473962813298372866232270325729656607138824984345210694447427006364854981849873631319052612433378838647528773441425507499941931953002904996294537444389804988467416770354954341406;
            6'd43: xpb[19] = 1024'd86861284296122556568421542743176010265225422162824122450991767019968735800674656824779138253890484006670552876071143770838240535247270961927900715077333038666818457954927844626829620472886651458897351529036775384445696722253221191948660410904316591011845311285217259877158693097827657488192831455363405635249;
            6'd44: xpb[19] = 1024'd88881314163474243930477857690691731434184152910796776461479947648340101749527555820704234492353053402174519222026286649229827524439067961042503057288433807007907259302716864269314030251325875911429848076223677137572340832073063545249792048367207674523748690617431614758022848751265509987918246140371856929092;
            6'd45: xpb[19] = 1024'd90901344030825931292534172638207452603142883658769430471968128276711467698380454816629330730815622797678485567981429527621414513630864960157105399499534575348996060650505883911798440029765100363962344623410578890698984941892905898550923685830098758035652069949645969638887004404703362487643660825380308222935;
            6'd46: xpb[19] = 1024'd92921373898177618654590487585723173772101614406742084482456308905082833647233353812554426969278192193182451913936572406013001502822661959271707741710635343690084861998294903554282849808204324816494841170597480643825629051712748251852055323292989841547555449281860324519751160058141214987369075510388759516778;
            6'd47: xpb[19] = 1024'd94941403765529306016646802533238894941060345154714738492944489533454199596086252808479523207740761588686418259891715284404588492014458958386310083921736112031173663346083923196767259586643549269027337717784382396952273161532590605153186960755880925059458828614074679400615315711579067487094490195397210810621;
            6'd48: xpb[19] = 1024'd96961433632880993378703117480754616110019075902687392503432670161825565544939151804404619446203330984190384605846858162796175481206255957500912426132836880372262464693872942839251669365082773721559834264971284150078917271352432958454318598218772008571362207946289034281479471365016919986819904880405662104464;
            6'd49: xpb[19] = 1024'd98981463500232680740759432428270337278977806650660046513920850790196931493792050800329715684665900379694350951802001041187762470398052956615514768343937648713351266041661962481736079143521998174092330812158185903205561381172275311755450235681663092083265587278503389162343627018454772486545319565414113398307;
            6'd50: xpb[19] = 1024'd101001493367584368102815747375786058447936537398632700524409031418568297442644949796254811923128469775198317297757143919579349459589849955730117110555038417054440067389450982124220488921961222626624827359345087656332205490992117665056581873144554175595168966610717744043207782671892624986270734250422564692150;
            6'd51: xpb[19] = 1024'd103021523234936055464872062323301779616895268146605354534897212046939663391497848792179908161591039170702283643712286797970936448781646954844719452766139185395528868737240001766704898700400447079157323906531989409458849600811960018357713510607445259107072345942932098924071938325330477485996148935431015985993;
            6'd52: xpb[19] = 1024'd105041553102287742826928377270817500785853998894578008545385392675311029340350747788105004400053608566206249989667429676362523437973443953959321794977239953736617670085029021409189308478839671531689820453718891162585493710631802371658845148070336342618975725275146453804936093978768329985721563620439467279836;
            6'd53: xpb[19] = 1024'd107061582969639430188984692218333221954812729642550662555873573303682395289203646784030100638516177961710216335622572554754110427165240953073924137188340722077706471432818041051673718257278895984222317000905792915712137820451644724959976785533227426130879104607360808685800249632206182485446978305447918573679;
            6'd54: xpb[19] = 1024'd109081612836991117551041007165848943123771460390523316566361753932053761238056545779955196876978747357214182681577715433145697416357037952188526479399441490418795272780607060694158128035718120436754813548092694668838781930271487078261108422996118509642782483939575163566664405285644034985172392990456369867522;
            6'd55: xpb[19] = 1024'd111101642704342804913097322113364664292730191138495970576849934560425127186909444775880293115441316752718149027532858311537284405548834951303128821610542258759884074128396080336642537814157344889287310095279596421965426040091329431562240060459009593154685863271789518447528560939081887484897807675464821161365;
            6'd56: xpb[19] = 1024'd113121672571694492275153637060880385461688921886468624587338115188796493135762343771805389353903886148222115373488001189928871394740631950417731163821643027100972875476185099979126947592596569341819806642466498175092070149911171784863371697921900676666589242604003873328392716592519739984623222360473272455208;
            6'd57: xpb[19] = 1024'd115141702439046179637209952008396106630647652634441278597826295817167859084615242767730485592366455543726081719443144068320458383932428949532333506032743795442061676823974119621611357371035793794352303189653399928218714259731014138164503335384791760178492621936218228209256872245957592484348637045481723749051;
            6'd58: xpb[19] = 1024'd117161732306397866999266266955911827799606383382413932608314476445539225033468141763655581830829024939230048065398286946712045373124225948646935848243844563783150478171763139264095767149475018246884799736840301681345358369550856491465634972847682843690396001268432583090121027899395444984074051730490175042894;
            6'd59: xpb[19] = 1024'd119181762173749554361322581903427548968565114130386586618802657073910590982321040759580678069291594334734014411353429825103632362316022947761538190454945332124239279519552158906580176927914242699417296284027203434472002479370698844766766610310573927202299380600646937970985183552833297483799466415498626336737;
            6'd60: xpb[19] = 1024'd121201792041101241723378896850943270137523844878359240629290837702281956931173939755505774307754163730237980757308572703495219351507819946876140532666046100465328080867341178549064586706353467151949792831214105187598646589190541198067898247773465010714202759932861292851849339206271149983524881100507077630580;
            6'd61: xpb[19] = 1024'd123221821908452929085435211798458991306482575626331894639779018330653322880026838751430870546216733125741947103263715581886806340699616945990742874877146868806416882215130198191548996484792691604482289378401006940725290699010383551369029885236356094226106139265075647732713494859709002483250295785515528924423;
            6'd62: xpb[19] = 1024'd1175156091679875048692599341160279730742879248568864522135343894047793491570598837340895570021628211802764041761365025699329489050193610550185092071916596213815008993348000496403167071714710335704588317200668847487573958609329131705182953016017728471189615183172944583471122439218221965857020643898385733935;
            6'd63: xpb[19] = 1024'd3195185959031562410748914288676000899701609996541518532623524522419159440423497833265991808484197607306730387716507904090916478241990609664787434283017364554903810341137020138887576850153934788237084864387570600614218068429171485006314590478908811983092994515387299464335278092656074465582435328906837027778;
        endcase
    end

    always_comb begin
        case(flag[6][16:12])
            5'd0: xpb[20] = 1024'd0;
            5'd1: xpb[20] = 1024'd5215215826383249772805229236191722068660340744514172543111705150790525389276396829191088046946767002810696733671650782482503467433787608779389776494118132895992611688926039781371986628593159240769581411574472353740862178249013838307446227941799895494996373847601654345199433746093926965307850013915288321621;
            5'd2: xpb[20] = 1024'd10430431652766499545610458472383444137320681489028345086223410301581050778552793658382176093893534005621393467343301564965006934867575217558779552988236265791985223377852079562743973257186318481539162823148944707481724356498027676614892455883599790989992747695203308690398867492187853930615700027830576643242;
            5'd3: xpb[20] = 1024'd15645647479149749318415687708575166205981022233542517629335115452371576167829190487573264140840301008432090201014952347447510402301362826338169329482354398687977835066778119344115959885779477722308744234723417061222586534747041514922338683825399686484989121542804963035598301238281780895923550041745864964863;
            5'd4: xpb[20] = 1024'd20860863305532999091220916944766888274641362978056690172446820603162101557105587316764352187787068011242786934686603129930013869735150435117559105976472531583970446755704159125487946514372636963078325646297889414963448712996055353229784911767199581979985495390406617380797734984375707861231400055661153286484;
            5'd5: xpb[20] = 1024'd26076079131916248864026146180958610343301703722570862715558525753952626946381984145955440234733835014053483668358253912412517337168938043896948882470590664479963058444630198906859933142965796203847907057872361768704310891245069191537231139708999477474981869238008271725997168730469634826539250069576441608105;
            5'd6: xpb[20] = 1024'd31291294958299498636831375417150332411962044467085035258670230904743152335658380975146528281680602016864180402029904694895020804602725652676338658964708797375955670133556238688231919771558955444617488469446834122445173069494083029844677367650799372969978243085609926071196602476563561791847100083491729929726;
            5'd7: xpb[20] = 1024'd36506510784682748409636604653342054480622385211599207801781936055533677724934777804337616328627369019674877135701555477377524272036513261455728435458826930271948281822482278469603906400152114685387069881021306476186035247743096868152123595592599268464974616933211580416396036222657488757154950097407018251347;
            5'd8: xpb[20] = 1024'd41721726611065998182441833889533776549282725956113380344893641206324203114211174633528704375574136022485573869373206259860027739470300870235118211952945063167940893511408318250975893028745273926156651292595778829926897425992110706459569823534399163959970990780813234761595469968751415722462800111322306572968;
            5'd9: xpb[20] = 1024'd46936942437449247955247063125725498617943066700627552888005346357114728503487571462719792422520903025296270603044857042342531206904088479014507988447063196063933505200334358032347879657338433166926232704170251183667759604241124544767016051476199059454967364628414889106794903714845342687770650125237594894589;
            5'd10: xpb[20] = 1024'd52152158263832497728052292361917220686603407445141725431117051507905253892763968291910880469467670028106967336716507824825034674337876087793897764941181328959926116889260397813719866285931592407695814115744723537408621782490138383074462279417998954949963738476016543451994337460939269653078500139152883216210;
            5'd11: xpb[20] = 1024'd57367374090215747500857521598108942755263748189655897974228756658695779282040365121101968516414437030917664070388158607307538141771663696573287541435299461855918728578186437595091852914524751648465395527319195891149483960739152221381908507359798850444960112323618197797193771207033196618386350153068171537831;
            5'd12: xpb[20] = 1024'd62582589916598997273662750834300664823924088934170070517340461809486304671316761950293056563361204033728360804059809389790041609205451305352677317929417594751911340267112477376463839543117910889234976938893668244890346138988166059689354735301598745939956486171219852142393204953127123583694200166983459859452;
            5'd13: xpb[20] = 1024'd67797805742982247046467980070492386892584429678684243060452166960276830060593158779484144610307971036539057537731460172272545076639238914132067094423535727647903951956038517157835826171711070130004558350468140598631208317237179897996800963243398641434952860018821506487592638699221050549002050180898748181073;
            5'd14: xpb[20] = 1024'd73013021569365496819273209306684108961244770423198415603563872111067355449869555608675232657254738039349754271403110954755048544073026522911456870917653860543896563644964556939207812800304229370774139762042612952372070495486193736304247191185198536929949233866423160832792072445314977514309900194814036502694;
            5'd15: xpb[20] = 1024'd78228237395748746592078438542875831029905111167712588146675577261857880839145952437866320704201505042160451005074761737237552011506814131690846647411771993439889175333890596720579799428897388611543721173617085306112932673735207574611693419126998432424945607714024815177991506191408904479617750208729324824315;
            5'd16: xpb[20] = 1024'd83443453222131996364883667779067553098565451912226760689787282412648406228422349267057408751148272044971147738746412519720055478940601740470236423905890126335881787022816636501951786057490547852313302585191557659853794851984221412919139647068798327919941981561626469523190939937502831444925600222644613145936;
            5'd17: xpb[20] = 1024'd88658669048515246137688897015259275167225792656740933232898987563438931617698746096248496798095039047781844472418063302202558946374389349249626200400008259231874398711742676283323772686083707093082883996766030013594657030233235251226585875010598223414938355409228123868390373683596758410233450236559901467557;
            5'd18: xpb[20] = 1024'd93873884874898495910494126251450997235886133401255105776010692714229457006975142925439584845041806050592541206089714084685062413808176958029015976894126392127867010400668716064695759314676866333852465408340502367335519208482249089534032102952398118909934729256829778213589807429690685375541300250475189789178;
            5'd19: xpb[20] = 1024'd99089100701281745683299355487642719304546474145769278319122397865019982396251539754630672891988573053403237939761364867167565881241964566808405753388244525023859622089594755846067745943270025574622046819914974721076381386731262927841478330894198014404931103104431432558789241175784612340849150264390478110799;
            5'd20: xpb[20] = 1024'd104304316527664995456104584723834441373206814890283450862234103015810507785527936583821760938935340056213934673433015649650069348675752175587795529882362657919852233778520795627439732571863184815391628231489447074817243564980276766148924558835997909899927476952033086903988674921878539306157000278305766432420;
            5'd21: xpb[20] = 1024'd109519532354048245228909813960026163441867155634797623405345808166601033174804333413012848985882107059024631407104666432132572816109539784367185306376480790815844845467446835408811719200456344056161209643063919428558105743229290604456370786777797805394923850799634741249188108667972466271464850292221054754041;
            5'd22: xpb[20] = 1024'd114734748180431495001715043196217885510527496379311795948457513317391558564080730242203937032828874061835328140776317214615076283543327393146575082870598923711837457156372875190183705829049503296930791054638391782298967921478304442763817014719597700889920224647236395594387542414066393236772700306136343075662;
            5'd23: xpb[20] = 1024'd119949964006814744774520272432409607579187837123825968491569218468182083953357127071395025079775641064646024874447967997097579750977115001925964859364717056607830068845298914971555692457642662537700372466212864136039830099727318281071263242661397596384916598494838049939586976160160320202080550320051631397283;
            5'd24: xpb[20] = 1024'd1098484149073253148526574263786896903149750742604456906549068553995714005324384990571041912064733758013572200662125345001019377569682276150194510842504148570132005964653737415297439894718616057159756269400096643416331427755435346413730900919968042613093068928322646254679881832325614150269710507341325234573;
            5'd25: xpb[20] = 1024'd6313699975456502921331803499978618971810091487118629449660773704786239394600781819762129959011500760824268934333776127483522845003469884929584287336622281466124617653579777196669426523311775297929337680974568997157193606004449184721177128861767938108089442775924300599879315578419541115577560521256613556194;
            5'd26: xpb[20] = 1024'd11528915801839752694137032736170341040470432231632801992772478855576764783877178648953218005958267763634965668005426909966026312437257493708974063830740414362117229342505816978041413151904934538698919092549041350898055784253463023028623356803567833603085816623525954945078749324513468080885410535171901877815;
            5'd27: xpb[20] = 1024'd16744131628223002466942261972362063109130772976146974535884184006367290173153575478144306052905034766445662401677077692448529779871045102488363840324858547258109841031431856759413399780498093779468500504123513704638917962502476861336069584745367729098082190471127609290278183070607395046193260549087190199436;
            5'd28: xpb[20] = 1024'd21959347454606252239747491208553785177791113720661147078995889157157815562429972307335394099851801769256359135348728474931033247304832711267753616818976680154102452720357896540785386409091253020238081915697986058379780140751490699643515812687167624593078564318729263635477616816701322011501110563002478521057;
            5'd29: xpb[20] = 1024'd27174563280989502012552720444745507246451454465175319622107594307948340951706369136526482146798568772067055869020379257413536714738620320047143393313094813050095064409283936322157373037684412261007663327272458412120642319000504537950962040628967520088074938166330917980677050562795248976808960576917766842678;
            5'd30: xpb[20] = 1024'd32389779107372751785357949680937229315111795209689492165219299458738866340982765965717570193745335774877752602692030039896040182172407928826533169807212945946087676098209976103529359666277571501777244738846930765861504497249518376258408268570767415583071312013932572325876484308889175942116810590833055164299;
            5'd31: xpb[20] = 1024'd37604994933756001558163178917128951383772135954203664708331004609529391730259162794908658240692102777688449336363680822378543649606195537605922946301331078842080287787136015884901346294870730742546826150421403119602366675498532214565854496512567311078067685861534226671075918054983102907424660604748343485920;
        endcase
    end

    always_comb begin
        case(flag[7][5:0])
            6'd0: xpb[21] = 1024'd0;
            6'd1: xpb[21] = 1024'd83443453222131996364883667779067553098565451912226760689787282412648406228422349267057408751148272044971147738746412519720055478940601740470236423905890126335881787022816636501951786057490547852313302585191557659853794851984221412919139647068798327919941981561626469523190939937502831444925600222644613145936;
            6'd2: xpb[21] = 1024'd42820210760139251330968408153320673452432476698717837251442709760319917119535559624099746287638869780499146070035331604861047117039983146385312722795449211738072899476062055666273332923463889983316407561995875473343228853747546052873300724454367206573064059709135881016275351801077029872732510618663631807541;
            6'd3: xpb[21] = 1024'd2196968298146506297053148527573793806299501485208913813098137107991428010648769981142083824129467516027144401324250690002038755139364552300389021685008297140264011929307474830594879789437232114319512538800193286832662855510870692827461801839936085226186137856645292509359763664651228300539421014682650469146;
            6'd4: xpb[21] = 1024'd85640421520278502661936816306641346904864953397435674502885419520639834239071119248199492575277739560998292140070663209722094234079966292770625445590898423476145798952124111332546665846927779966632815123991750946686457707495092105746601448908734413146128119418271762032550703602154059745465021237327263615082;
            6'd5: xpb[21] = 1024'd45017179058285757628021556680894467258731978183926751064540846868311345130184329605241830111768337296526290471359582294863085872179347698685701744480457508878336911405369530496868212712901122097635920100796068760175891709258416745700762526294303291799250197565781173525635115465728258173271931633346282276687;
            6'd6: xpb[21] = 1024'd4393936596293012594106297055147587612599002970417827626196274215982856021297539962284167648258935032054288802648501380004077510278729104600778043370016594280528023858614949661189759578874464228639025077600386573665325711021741385654923603679872170452372275713290585018719527329302456601078842029365300938292;
            6'd7: xpb[21] = 1024'd87837389818425008958989964834215140711164454882644588315983556628631262249719889229341576399407207077025436541394913899724132989219330845071014467275906720616409810881431586163141545636365012080952327662791944233519120563005962798574063250748670498372314257274917054541910467266805288046004442252009914084228;
            6'd8: xpb[21] = 1024'd47214147356432263925074705208468261065031479669135664877638983976302773140833099586383913935897804812553434872683832984865124627318712250986090766165465806018600923334677005327463092502338354211955432639596262047008554564769287438528224328134239377025436335422426466034994879130379486473811352648028932745833;
            6'd9: xpb[21] = 1024'd6590904894439518891159445582721381418898504455626741439294411323974284031946309943426251472388402548081433203972752070006116265418093656901167065055024891420792035787922424491784639368311696342958537616400579860497988566532612078482385405519808255678558413569935877528079290993953684901618263044047951407438;
            6'd10: xpb[21] = 1024'd90034358116571515256043113361788934517463956367853502129081693736622690260368659210483660223536674593052580942719164589726171744358695397371403488960915017756673822810739060993736425425802244195271840201592137520351783418516833491401525052588606583598500395131562347051270230931456516346543863266692564553374;
            6'd11: xpb[21] = 1024'd49411115654578770222127853736042054871330981154344578690737121084294201151481869567525997760027272328580579274008083674867163382458076803286479787850474103158864935263984480158057972291775586326274945178396455333841217420280158131355686129974175462251622473279071758544354642795030714774350773662711583214979;
            6'd12: xpb[21] = 1024'd8787873192586025188212594110295175225198005940835655252392548431965712042595079924568335296517870064108577605297002760008155020557458209201556086740033188561056047717229899322379519157748928457278050155200773147330651422043482771309847207359744340904744551426581170037439054658604913202157684058730601876584;
            6'd13: xpb[21] = 1024'd92231326414718021553096261889362728323763457853062415942179830844614118271017429191625744047666142109079725344043415279728210499498059949671792510645923314896937834740046535824331305215239476309591352740392330807184446274027704184228986854428542668824686532988207639560629994596107744647083284281375215022520;
            6'd14: xpb[21] = 1024'd51608083952725276519181002263615848677630482639553492503835258192285629162130639548668081584156739844607723675332334364869202137597441355586868809535482400299128947193291954988652852081212818440594457717196648620673880275791028824183147931814111547477808611135717051053714406459681943074890194677394233684125;
            6'd15: xpb[21] = 1024'd10984841490732531485265742637868969031497507426044569065490685539957140053243849905710419120647337580135722006621253450010193775696822761501945108425041485701320059646537374152974398947186160571597562694000966434163314277554353464137309009199680426130930689283226462546798818323256141502697105073413252345730;
            6'd16: xpb[21] = 1024'd94428294712864527850149410416936522130062959338271329755277967952605546281666199172767827871795609625106869745367665969730249254637424501972181532330931612037201846669354010654926185004676708423910865279192524094017109129538574877056448656268478754050872670844852932069989758260758972947622705296057865491666;
            6'd17: xpb[21] = 1024'd53805052250871782816234150791189642483929984124762406316933395300277057172779409529810165408286207360634868076656585054871240892736805907887257831220490697439392959122599429819247731870650050554913970255996841907506543131301899517010609733654047632703994748992362343563074170124333171375429615692076884153271;
            6'd18: xpb[21] = 1024'd13181809788879037782318891165442762837797008911253482878588822647948568063892619886852502944776805096162866407945504140012232530836187313802334130110049782841584071575844848983569278736623392685917075232801159720995977133065224156964770811039616511357116827139871755056158581987907369803236526088095902814876;
            6'd19: xpb[21] = 1024'd96625263011011034147202558944510315936362460823480243568376105060596974292314969153909911695925077141134014146691916659732288009776789054272570554015939909177465858598661485485521064794113940538230377817992717380849771985049445569883910458108414839277058808701498224579349521925410201248162126310740515960812;
            6'd20: xpb[21] = 1024'd56002020549018289113287299318763436290229485609971320130031532408268485183428179510952249232415674876662012477980835744873279647876170460187646852905498994579656971051906904649842611660087282669233482794797035194339205986812770209838071535493983717930180886849007636072433933788984399675969036706759534622417;
            6'd21: xpb[21] = 1024'd15378778087025544079372039693016556644096510396462396691686959755939996074541389867994586768906272612190010809269754830014271285975551866102723151795058079981848083505152323814164158526060624800236587771601353007828639988576094849792232612879552596583302964996517047565518345652558598103775947102778553284022;
            6'd22: xpb[21] = 1024'd98822231309157540444255707472084109742661962308689157381474242168588402302963739135051995520054544657161158548016167349734326764916153606572959575700948206317729870527968960316115944583551172652549890356792910667682434840560316262711372259948350924503244946558143517088709285590061429548701547325423166429958;
            6'd23: xpb[21] = 1024'd58198988847164795410340447846337230096528987095180233943129669516259913194076949492094333056545142392689156879305086434875318403015535012488035874590507291719920982981214379480437491449524514783552995333597228481171868842323640902665533337333919803156367024705652928581793697453635627976508457721442185091563;
            6'd24: xpb[21] = 1024'd17575746385172050376425188220590350450396011881671310504785096863931424085190159849136670593035740128217155210594005520016310041114916418403112173480066377122112095434459798644759038315497856914556100310401546294661302844086965542619694414719488681809489102853162340074878109317209826404315368117461203753168;
            6'd25: xpb[21] = 1024'd101019199607304046741308855999657903548961463793898071194572379276579830313612509116194079344184012173188302949340418039736365520055518158873348597385956503457993882457276435146710824372988404766869402895593103954515097696071186955538834061788287009729431084414788809598069049254712657849240968340105816899104;
            6'd26: xpb[21] = 1024'd60395957145311301707393596373911023902828488580389147756227806624251341204725719473236416880674609908716301280629337124877357158154899564788424896275515588860184994910521854311032371238961746897872507872397421768004531697834511595492995139173855888382553162562298221091153461118286856277047878736124835560709;
            6'd27: xpb[21] = 1024'd19772714683318556673478336748164144256695513366880224317883233971922852095838929830278754417165207644244299611918256210018348796254280970703501195165074674262376107363767273475353918104935089028875612849201739581493965699597836235447156216559424767035675240709807632584237872981861054704854789132143854222314;
            6'd28: xpb[21] = 1024'd103216167905450553038362004527231697355260965279106985007670516384571258324261279097336163168313479689215447350664668729738404275194882711173737619070964800598257894386583909977305704162425636881188915434393297241347760551582057648366295863628223094955617222271434102107428812919363886149780389354788467368250;
            6'd29: xpb[21] = 1024'd62592925443457808004446744901484817709127990065598061569325943732242769215374489454378500704804077424743445681953587814879395913294264117088813917960523886000449006839829329141627251028398979012192020411197615054837194553345382288320456941013791973608739300418943513600513224782938084577587299750807486029855;
            6'd30: xpb[21] = 1024'd21969682981465062970531485275737938062995014852089138130981371079914280106487699811420838241294675160271444013242506900020387551393645523003890216850082971402640119293074748305948797894372321143195125388001932868326628555108706928274618018399360852261861378566452925093597636646512283005394210146826504691460;
            6'd31: xpb[21] = 1024'd105413136203597059335415153054805491161560466764315898820768653492562686334910049078478246992442947205242591751988919419740443030334247263474126640755973097738521906315891384807900583951862868995508427973193490528180423407092928341193757665468159180181803360128079394616788576584015114450319810369471117837396;
            6'd32: xpb[21] = 1024'd64789893741604314301499893429058611515427491550806975382424080840234197226023259435520584528933544940770590083277838504881434668433628669389202939645532183140713018769136803972222130817836211126511532949997808341669857408856252981147918742853728058834925438275588806109872988447589312878126720765490136499001;
            6'd33: xpb[21] = 1024'd24166651279611569267584633803311731869294516337298051944079508187905708117136469792562922065424142676298588414566757590022426306533010075304279238535091268542904131222382223136543677683809553257514637926802126155159291410619577621102079820239296937488047516423098217602957400311163511305933631161509155160606;
            6'd34: xpb[21] = 1024'd107610104501743565632468301582379284967859968249524812633866790600554114345558819059620330816572414721269736153313170109742481785473611815774515662440981394878785918245198859638495463741300101109827940511993683815013086262603799034021219467308095265407989497984724687126148340248666342750859231384153768306542;
            6'd35: xpb[21] = 1024'd66986862039750820598553041956632405321726993036015889195522217948225625236672029416662668353063012456797734484602089194883473423572993221689591961330540480280977030698444278802817010607273443240831045488798001628502520264367123673975380544693664144061111576132234098619232752112240541178666141780172786968147;
            6'd36: xpb[21] = 1024'd26363619577758075564637782330885525675594017822506965757177645295897136127785239773705005889553610192325732815891008280024465061672374627604668260220099565683168143151689697967138557473246785371834150465602319441991954266130448313929541622079233022714233654279743510112317163975814739606473052176191805629752;
            6'd37: xpb[21] = 1024'd109807072799890071929521450109953078774159469734733726446964927708545542356207589040762414640701882237296880554637420799744520540612976368074904684125989692019049930174506334469090343530737333224147453050793877101845749118114669726848681269148031350634175635841369979635508103913317571051398652398836418775688;
            6'd38: xpb[21] = 1024'd69183830337897326895606190484206199128026494521224803008620355056217053247320799397804752177192479972824878885926339884885512178712357773989980983015548777421241042627751753633411890396710675355150558027598194915335183119877994366802842346533600229287297713988879391128592515776891769479205562794855437437293;
            6'd39: xpb[21] = 1024'd28560587875904581861690930858459319481893519307715879570275782403888564138434009754847089713683077708352877217215258970026503816811739179905057281905107862823432155080997172797733437262684017486153663004402512728824617121641319006757003423919169107940419792136388802621676927640465967907012473190874456098898;
            6'd40: xpb[21] = 1024'd112004041098036578226574598637526872580458971219942640260063064816536970366856359021904498464831349753324024955961671489746559295752340920375293705810997989159313942103813809299685223320174565338466965589594070388678411973625540419676143070987967435860361773698015272144867867577968799351938073413519069244834;
            6'd41: xpb[21] = 1024'd71380798636043833192659339011779992934325996006433716821718492164208481257969569378946836001321947488852023287250590574887550933851722326290370004700557074561505054557059228464006770186147907469470070566398388202167845975388865059630304148373536314513483851845524683637952279441542997779744983809538087906439;
            6'd42: xpb[21] = 1024'd30757556174051088158744079386033113288193020792924793383373919511879992149082779735989173537812545224380021618539509660028542571951103732205446303590116159963696167010304647628328317052121249600473175543202706015657279977152189699584465225759105193166605929993034095131036691305117196207551894205557106568044;
            6'd43: xpb[21] = 1024'd114201009396183084523627747165100666386758472705151554073161201924528398377505129003046582288960817269351169357285922179748598050891705472675682727496006286299577954033121284130280103109611797452786478128394263675511074829136411112503604872827903521086547911554660564654227631242620027652477494428201719713980;
            6'd44: xpb[21] = 1024'd73577766934190339489712487539353786740625497491642630634816629272199909268618339360088919825451415004879167688574841264889589688991086878590759026385565371701769066486366703294601649975585139583789583105198581489000508830899735752457765950213472399739669989702169976147312043106194226080284404824220738375585;
            6'd45: xpb[21] = 1024'd32954524472197594455797227913606907094492522278133707196472056619871420159731549717131257361942012740407166019863760350030581327090468284505835325275124457103960178939612122458923196841558481714792688082002899302489942832663060392411927027599041278392792067849679387640396454969768424508091315220239757037190;
            6'd46: xpb[21] = 1024'd116397977694329590820680895692674460193057974190360467886259339032519826388153898984188666113090284785378313758610172869750636806031070024976071749181014583439841965962428758960874982899049029567105990667194456962343737684647281805331066674667839606312734049411305857163587394907271255953016915442884370183126;
            6'd47: xpb[21] = 1024'd75774735232336845786765636066927580546924998976851544447914766380191337279267109341231003649580882520906312089899091954891628444130451430891148048070573668842033078415674178125196529765022371698109095643998774775833171686410606445285227752053408484965856127558815268656671806770845454380823825838903388844731;
            6'd48: xpb[21] = 1024'd35151492770344100752850376441180700900792023763342621009570193727862848170380319698273341186071480256434310421188011040032620082229832836806224346960132754244224190868919597289518076630995713829112200620803092589322605688173931085239388829438977363618978205706324680149756218634419652808630736234922407506336;
            6'd49: xpb[21] = 1024'd118594945992476097117734044220248253999357475675569381699357476140511254398802668965330749937219752301405458159934423559752675561170434577276460770866022880580105977891736233791469862688486261681425503205994650249176400540158152498158528476507775691538920187267951149672947158571922484253556336457567020652272;
            6'd50: xpb[21] = 1024'd77971703530483352083818784594501374353224500462060458261012903488182765289915879322373087473710350036933456491223342644893667199269815983191537069755581965982297090344981652955791409554459603812428608182798968062665834541921477138112689553893344570192042265415460561166031570435496682681363246853586039313877;
            6'd51: xpb[21] = 1024'd37348461068490607049903524968754494707091525248551534822668330835854276181029089679415425010200947772461454822512261730034658837369197389106613368645141051384488202798227072120112956420432945943431713159603285876155268543684801778066850631278913448845164343562969972659115982299070881109170157249605057975482;
            6'd52: xpb[21] = 1024'd120791914290622603414787192747822047805656977160778295512455613248502682409451438946472833761349219817432602561258674249754714316309799129576849792551031177720369989821043708622064742477923493795745015744794843536009063395669023190985990278347711776765106325124596442182306922236573712554095757472249671121418;
            6'd53: xpb[21] = 1024'd80168671828629858380871933122075168159524001947269372074111040596174193300564649303515171297839817552960600892547593334895705954409180535491926091440590263122561102274289127786386289343896835926748120721599161349498497397432347830940151355733280655418228403272105853675391334100147910981902667868268689783023;
            6'd54: xpb[21] = 1024'd39545429366637113346956673496328288513391026733760448635766467943845704191677859660557508834330415288488599223836512420036697592508561941407002390330149348524752214727534546950707836209870178057751225698403479162987931399195672470894312433118849534071350481419615265168475745963722109409709578264287708444628;
            6'd55: xpb[21] = 1024'd122988882588769109711840341275395841611956478645987209325553750356494110420100208927614917585478687333459746962582924939756753071449163681877238814236039474860634001750351183452659622267360725910064528283595036822841726251179893883813452080187647861991292462981241734691666685901224940854635178486932321590564;
            6'd56: xpb[21] = 1024'd82365640126776364677925081649648961965823503432478285887209177704165621311213419284657255121969285068987745293871844024897744709548545087792315113125598560262825114203596602616981169133334068041067633260399354636331160252943218523767613157573216740644414541128751146184751097764799139282442088882951340252169;
            6'd57: xpb[21] = 1024'd41742397664783619644009822023902082319690528218969362448864605051837132202326629641699592658459882804515743625160763110038736347647926493707391412015157645665016226656842021781302715999307410172070738237203672449820594254706543163721774234958785619297536619276260557677835509628373337710248999278970358913774;
            6'd58: xpb[21] = 1024'd1119155202790874610094562398155202673557553005460439010520032399508643093439839998741930194950480540043741956449682195179727985747307899622467710904716731067207339110087440945624262865280752303073843214007990263310028256469867803675935312344354497950658697423769969170919921491947536138055909674989377575379;
            6'd59: xpb[21] = 1024'd84562608424922870974978230177222755772123004917687199700307314812157049321862189265799338946098752585014889695196094714899783464687909640092704134810606857403089126132904077447576048922771300155387145799199547923163823108454089216595074959413152825870600678985396438694110861429450367582981509897633990721315;
            6'd60: xpb[21] = 1024'd43939365962930125941062970551475876125990029704178276261962742159828560212975399622841676482589350320542888026485013800040775102787291046007780433700165942805280238586149496611897595788744642286390250776003865736653257110217413856549236036798721704523722757132905850187195273293024566010788420293653009382920;
            6'd61: xpb[21] = 1024'd3316123500937380907147710925728996479857054490669352823618169507500071104088609979884014019079948056070886357773932885181766740886672451922856732589725028207471351039394915776219142654717984417393355752808183550142691111980738496503397114184290583176844835280415261680279685156598764438595330689672028044525;
            6'd62: xpb[21] = 1024'd86759576723069377272031378704796549578422506402896113513405451920148477332510959246941422770228220101042034096520345404901822219827274192393093156495615154543353138062211552278170928712208532269706658337999741209996485963964959909422536761253088911096786816842041731203470625094101595883520930912316641190461;
            6'd63: xpb[21] = 1024'd46136334261076632238116119079049669932289531189387190075060879267819988223624169603983760306718817836570032427809264490042813857926655598308169455385174239945544250515456971442492475578181874400709763314804059023485919965728284549376697838638657789749908894989551142696555036957675794311327841308335659852066;
        endcase
    end

    always_comb begin
        case(flag[7][11:6])
            6'd0: xpb[22] = 1024'd0;
            6'd1: xpb[22] = 1024'd5513091799083887204200859453302790286156555975878266636716306615491499114737379961026097843209415572098030759098183575183805496026037004223245754274733325347735362968702390606814022444155216531712868291608376836975353967491609189330858916024226668403030973137060554189639448821249992739134751704354678513671;
            6'd2: xpb[22] = 1024'd11026183598167774408401718906605580572313111951756533273432613230982998229474759922052195686418831144196061518196367150367610992052074008446491508549466650695470725937404781213628044888310433063425736583216753673950707934983218378661717832048453336806061946274121108379278897642499985478269503408709357027342;
            6'd3: xpb[22] = 1024'd16539275397251661612602578359908370858469667927634799910148919846474497344212139883078293529628246716294092277294550725551416488078111012669737262824199976043206088906107171820442067332465649595138604874825130510926061902474827567992576748072680005209092919411181662568918346463749978217404255113064035541013;
            6'd4: xpb[22] = 1024'd22052367196335548816803437813211161144626223903513066546865226461965996458949519844104391372837662288392123036392734300735221984104148016892983017098933301390941451874809562427256089776620866126851473166433507347901415869966436757323435664096906673612123892548242216758557795284999970956539006817418714054684;
            6'd5: xpb[22] = 1024'd27565458995419436021004297266513951430782779879391333183581533077457495573686899805130489216047077860490153795490917875919027480130185021116228771373666626738676814843511953034070112220776082658564341458041884184876769837458045946654294580121133342015154865685302770948197244106249963695673758521773392568355;
            6'd6: xpb[22] = 1024'd33078550794503323225205156719816741716939335855269599820297839692948994688424279766156587059256493432588184554589101451102832976156222025339474525648399952086412177812214343640884134664931299190277209749650261021852123804949655135985153496145360010418185838822363325137836692927499956434808510226128071082026;
            6'd7: xpb[22] = 1024'd38591642593587210429406016173119532003095891831147866457014146308440493803161659727182684902465909004686215313687285026286638472182259029562720279923133277434147540780916734247698157109086515721990078041258637858827477772441264325316012412169586678821216811959423879327476141748749949173943261930482749595697;
            6'd8: xpb[22] = 1024'd44104734392671097633606875626422322289252447807026133093730452923931992917899039688208782745675324576784246072785468601470443968208296033785966034197866602781882903749619124854512179553241732253702946332867014695802831739932873514646871328193813347224247785096484433517115590569999941913078013634837428109368;
            6'd9: xpb[22] = 1024'd49617826191754984837807735079725112575409003782904399730446759539423492032636419649234880588884740148882276831883652176654249464234333038009211788472599928129618266718321515461326201997396948785415814624475391532778185707424482703977730244218040015627278758233544987706755039391249934652212765339192106623039;
            6'd10: xpb[22] = 1024'd55130917990838872042008594533027902861565559758782666367163066154914991147373799610260978432094155720980307590981835751838054960260370042232457542747333253477353629687023906068140224441552165317128682916083768369753539674916091893308589160242266684030309731370605541896394488212499927391347517043546785136710;
            6'd11: xpb[22] = 1024'd60644009789922759246209453986330693147722115734660933003879372770406490262111179571287076275303571293078338350080019327021860456286407046455703297022066578825088992655726296674954246885707381848841551207692145206728893642407701082639448076266493352433340704507666096086033937033749920130482268747901463650381;
            6'd12: xpb[22] = 1024'd66157101589006646450410313439633483433878671710539199640595679385897989376848559532313174118512986865176369109178202902205665952312444050678949051296799904172824355624428687281768269329862598380554419499300522043704247609899310271970306992290720020836371677644726650275673385854999912869617020452256142164052;
            6'd13: xpb[22] = 1024'd71670193388090533654611172892936273720035227686417466277311986001389488491585939493339271961722402437274399868276386477389471448338481054902194805571533229520559718593131077888582291774017814912267287790908898880679601577390919461301165908314946689239402650781787204465312834676249905608751772156610820677723;
            6'd14: xpb[22] = 1024'd77183285187174420858812032346239064006191783662295732914028292616880987606323319454365369804931818009372430627374570052573276944364518059125440559846266554868295081561833468495396314218173031443980156082517275717654955544882528650632024824339173357642433623918847758654952283497499898347886523860965499191394;
            6'd15: xpb[22] = 1024'd82696376986258308063012891799541854292348339638173999550744599232372486721060699415391467648141233581470461386472753627757082440390555063348686314120999880216030444530535859102210336662328247975693024374125652554630309512374137839962883740363400026045464597055908312844591732318749891087021275565320177705065;
            6'd16: xpb[22] = 1024'd88209468785342195267213751252844644578504895614052266187460905847863985835798079376417565491350649153568492145570937202940887936416592067571932068395733205563765807499238249709024359106483464507405892665734029391605663479865747029293742656387626694448495570192968867034231181139999883826156027269674856218736;
            6'd17: xpb[22] = 1024'd93722560584426082471414610706147434864661451589930532824177212463355484950535459337443663334560064725666522904669120778124693432442629071795177822670466530911501170467940640315838381550638681039118760957342406228581017447357356218624601572411853362851526543330029421223870629961249876565290778974029534732407;
            6'd18: xpb[22] = 1024'd99235652383509969675615470159450225150818007565808799460893519078846984065272839298469761177769480297764553663767304353308498928468666076018423576945199856259236533436643030922652403994793897570831629248950783065556371414848965407955460488436080031254557516467089975413510078782499869304425530678384213246078;
            6'd19: xpb[22] = 1024'd104748744182593856879816329612753015436974563541687066097609825694338483180010219259495859020978895869862584422865487928492304424494703080241669331219933181606971896405345421529466426438949114102544497540559159902531725382340574597286319404460306699657588489604150529603149527603749862043560282382738891759749;
            6'd20: xpb[22] = 1024'd110261835981677744084017189066055805723131119517565332734326132309829982294747599220521956864188311441960615181963671503676109920520740084464915085494666506954707259374047812136280448883104330634257365832167536739507079349832183786617178320484533368060619462741211083792788976424999854782695034087093570273420;
            6'd21: xpb[22] = 1024'd115774927780761631288218048519358596009287675493443599371042438925321481409484979181548054707397727014058645941061855078859915416546777088688160839769399832302442622342750202743094471327259547165970234123775913576482433317323792975948037236508760036463650435878271637982428425246249847521829785791448248787091;
            6'd22: xpb[22] = 1024'd121288019579845518492418907972661386295444231469321866007758745540812980524222359142574152550607142586156676700160038654043720912572814092911406594044133157650177985311452593349908493771414763697683102415384290413457787284815402165278896152532986704866681409015332192172067874067499840260964537495802927300762;
            6'd23: xpb[22] = 1024'd2734415694804664297820840021149743836902360319464448516343197091327584301650600193585179179158883848811558051800728794648462567757630762579492223302535442064222673710583766619092277024052774508085773098605427404068780402086114581644776498873983924002892478738275688331600794814821199982980599373532011330102;
            6'd24: xpb[22] = 1024'd8247507493888551502021699474452534123058916295342715153059503706819083416387980154611277022368299420909588810898912369832268063783667766802737977577268767411958036679286157225906299468207991039798641390213804241044134369577723770975635414898210592405923451875336242521240243636071192722115351077886689843773;
            6'd25: xpb[22] = 1024'd13760599292972438706222558927755324409215472271220981789775810322310582531125360115637374865577714993007619569997095945016073559809704771025983731852002092759693399647988547832720321912363207571511509681822181078019488337069332960306494330922437260808954425012396796710879692457321185461250102782241368357444;
            6'd26: xpb[22] = 1024'd19273691092056325910423418381058114695372028247099248426492116937802081645862740076663472708787130565105650329095279520199879055835741775249229486126735418107428762616690938439534344356518424103224377973430557914994842304560942149637353246946663929211985398149457350900519141278571178200384854486596046871115;
            6'd27: xpb[22] = 1024'd24786782891140213114624277834360904981528584222977515063208423553293580760600120037689570551996546137203681088193463095383684551861778779472475240401468743455164125585393329046348366800673640634937246265038934751970196272052551338968212162970890597615016371286517905090158590099821170939519606190950725384786;
            6'd28: xpb[22] = 1024'd30299874690224100318825137287663695267685140198855781699924730168785079875337499998715668395205961709301711847291646670567490047887815783695720994676202068802899488554095719653162389244828857166650114556647311588945550239544160528299071078995117266018047344423578459279798038921071163678654357895305403898457;
            6'd29: xpb[22] = 1024'd35812966489307987523025996740966485553841696174734048336641036784276578990074879959741766238415377281399742606389830245751295543913852787918966748950935394150634851522798110259976411688984073698362982848255688425920904207035769717629929995019343934421078317560639013469437487742321156417789109599660082412128;
            6'd30: xpb[22] = 1024'd41326058288391874727226856194269275839998252150612314973357343399768078104812259920767864081624792853497773365488013820935101039939889792142212503225668719498370214491500500866790434133139290230075851139864065262896258174527378906960788911043570602824109290697699567659076936563571149156923861304014760925799;
            6'd31: xpb[22] = 1024'd46839150087475761931427715647572066126154808126490581610073650015259577219549639881793961924834208425595804124586197396118906535965926796365458257500402044846105577460202891473604456577294506761788719431472442099871612142018988096291647827067797271227140263834760121848716385384821141896058613008369439439470;
            6'd32: xpb[22] = 1024'd52352241886559649135628575100874856412311364102368848246789956630751076334287019842820059768043623997693834883684380971302712031991963800588704011775135370193840940428905282080418479021449723293501587723080818936846966109510597285622506743092023939630171236971820676038355834206071134635193364712724117953141;
            6'd33: xpb[22] = 1024'd57865333685643536339829434554177646698467920078247114883506263246242575449024399803846157611253039569791865642782564546486517528018000804811949766049868695541576303397607672687232501465604939825214456014689195773822320077002206474953365659116250608033202210108881230227995283027321127374328116417078796466812;
            6'd34: xpb[22] = 1024'd63378425484727423544030294007480436984624476054125381520222569861734074563761779764872255454462455141889896401880748121670323024044037809035195520324602020889311666366310063294046523909760156356927324306297572610797674044493815664284224575140477276436233183245941784417634731848571120113462868121433474980483;
            6'd35: xpb[22] = 1024'd68891517283811310748231153460783227270781032030003648156938876477225573678499159725898353297671870713987927160978931696854128520070074813258441274599335346237047029335012453900860546353915372888640192597905949447773028011985424853615083491164703944839264156383002338607274180669821112852597619825788153494154;
            6'd36: xpb[22] = 1024'd74404609082895197952432012914086017556937588005881914793655183092717072793236539686924451140881286286085957920077115272037934016096111817481687028874068671584782392303714844507674568798070589420353060889514326284748381979477034042945942407188930613242295129520062892796913629491071105591732371530142832007825;
            6'd37: xpb[22] = 1024'd79917700881979085156632872367388807843094143981760181430371489708208571907973919647950548984090701858183988679175298847221739512122148821704932783148801996932517755272417235114488591242225805952065929181122703121723735946968643232276801323213157281645326102657123446986553078312321098330867123234497510521496;
            6'd38: xpb[22] = 1024'd85430792681062972360833731820691598129250699957638448067087796323700071022711299608976646827300117430282019438273482422405545008148185825928178537423535322280253118241119625721302613686381022483778797472731079958699089914460252421607660239237383950048357075794184001176192527133571091070001874938852189035167;
            6'd39: xpb[22] = 1024'd90943884480146859565034591273994388415407255933516714703804102939191570137448679570002744670509533002380050197371665997589350504174222830151424291698268647627988481209822016328116636130536239015491665764339456795674443881951861610938519155261610618451388048931244555365831975954821083809136626643206867548838;
            6'd40: xpb[22] = 1024'd96456976279230746769235450727297178701563811909394981340520409554683069252186059531028842513718948574478080956469849572773156000200259834374670045973001972975723844178524406934930658574691455547204534055947833632649797849443470800269378071285837286854419022068305109555471424776071076548271378347561546062509;
            6'd41: xpb[22] = 1024'd101970068078314633973436310180599968987720367885273247977236716170174568366923439492054940356928364146576111715568033147956961496226296838597915800247735298323459207147226797541744681018846672078917402347556210469625151816935079989600236987310063955257449995205365663745110873597321069287406130051916224576180;
            6'd42: xpb[22] = 1024'd107483159877398521177637169633902759273876923861151514613953022785666067481660819453081038200137779718674142474666216723140766992252333842821161554522468623671194570115929188148558703463001888610630270639164587306600505784426689178931095903334290623660480968342426217934750322418571062026540881756270903089851;
            6'd43: xpb[22] = 1024'd112996251676482408381838029087205549560033479837029781250669329401157566596398199414107136043347195290772173233764400298324572488278370847044407308797201949018929933084631578755372725907157105142343138930772964143575859751918298368261954819358517292063511941479486772124389771239821054765675633460625581603522;
            6'd44: xpb[22] = 1024'd118509343475566295586038888540508339846190035812908047887385636016649065711135579375133233886556610862870203992862583873508377984304407851267653063071935274366665296053333969362186748351312321674056007222381340980551213719409907557592813735382743960466542914616547326314029220061071047504810385164980260117193;
            6'd45: xpb[22] = 1024'd124022435274650182790239747993811130132346591788786314524101942632140564825872959336159331729766026434968234751960767448692183480330444855490898817346668599714400659022036359969000770795467538205768875513989717817526567686901516746923672651406970628869573887753607880503668668882321040243945136869334938630864;
            6'd46: xpb[22] = 1024'd5468831389609328595641680042299487673804720638928897032686394182655168603301200387170358358317767697623116103601457589296925135515261525158984446605070884128445347421167533238184554048105549016171546197210854808137560804172229163289552997747967848005784957476551376663201589629642399965961198747064022660204;
            6'd47: xpb[22] = 1024'd10981923188693215799842539495602277959961276614807163669402700798146667718038580348196456201527183269721146862699641164480730631541298529382230200879804209476180710389869923844998576492260765547884414488819231645112914771663838352620411913772194516408815930613611930852841038450892392705095950451418701173875;
            6'd48: xpb[22] = 1024'd16495014987777103004043398948905068246117832590685430306119007413638166832775960309222554044736598841819177621797824739664536127567335533605475955154537534823916073358572314451812598936415982079597282780427608482088268739155447541951270829796421184811846903750672485042480487272142385444230702155773379687546;
            6'd49: xpb[22] = 1024'd22008106786860990208244258402207858532274388566563696942835314029129665947513340270248651887946014413917208380896008314848341623593372537828721709429270860171651436327274705058626621380571198611310151072035985319063622706647056731282129745820647853214877876887733039232119936093392378183365453860128058201217;
            6'd50: xpb[22] = 1024'd27521198585944877412445117855510648818430944542441963579551620644621165062250720231274749731155429986015239139994191890032147119619409542051967463704004185519386799295977095665440643824726415143023019363644362156038976674138665920612988661844874521617908850024793593421759384914642370922500205564482736714888;
            6'd51: xpb[22] = 1024'd33034290385028764616645977308813439104587500518320230216267927260112664176988100192300847574364845558113269899092375465215952615645446546275213217978737510867122162264679486272254666268881631674735887655252738993014330641630275109943847577869101190020939823161854147611398833735892363661634957268837415228559;
            6'd52: xpb[22] = 1024'd38547382184112651820846836762116229390744056494198496852984233875604163291725480153326945417574261130211300658190559040399758111671483550498458972253470836214857525233381876879068688713036848206448755946861115829989684609121884299274706493893327858423970796298914701801038282557142356400769708973192093742230;
            6'd53: xpb[22] = 1024'd44060473983196539025047696215419019676900612470076763489700540491095662406462860114353043260783676702309331417288742615583563607697520554721704726528204161562592888202084267485882711157192064738161624238469492666965038576613493488605565409917554526827001769435975255990677731378392349139904460677546772255901;
            6'd54: xpb[22] = 1024'd49573565782280426229248555668721809963057168445955030126416847106587161521200240075379141103993092274407362176386926190767369103723557558944950480802937486910328251170786658092696733601347281269874492530077869503940392544105102677936424325941781195230032742573035810180317180199642341879039212381901450769572;
            6'd55: xpb[22] = 1024'd55086657581364313433449415122024600249213724421833296763133153722078660635937620036405238947202507846505392935485109765951174599749594563168196235077670812258063614139489048699510756045502497801587360821686246340915746511596711867267283241966007863633063715710096364369956629020892334618173964086256129283243;
            6'd56: xpb[22] = 1024'd60599749380448200637650274575327390535370280397711563399849460337570159750674999997431336790411923418603423694583293341134980095775631567391441989352404137605798977108191439306324778489657714333300229113294623177891100479088321056598142157990234532036094688847156918559596077842142327357308715790610807796914;
            6'd57: xpb[22] = 1024'd66112841179532087841851134028630180821526836373589830036565766953061658865412379958457434633621338990701454453681476916318785591801668571614687743627137462953534340076893829913138800933812930865013097404903000014866454446579930245929001074014461200439125661984217472749235526663392320096443467494965486310585;
            6'd58: xpb[22] = 1024'd71625932978615975046051993481932971107683392349468096673282073568553157980149759919483532476830754562799485212779660491502591087827705575837933497901870788301269703045596220519952823377968147396725965696511376851841808414071539435259859990038687868842156635121278026938874975484642312835578219199320164824256;
            6'd59: xpb[22] = 1024'd77139024777699862250252852935235761393839948325346363309998380184044657094887139880509630320040170134897515971877844066686396583853742580061179252176604113649005066014298611126766845822123363928438833988119753688817162381563148624590718906062914537245187608258338581128514424305892305574712970903674843337927;
            6'd60: xpb[22] = 1024'd82652116576783749454453712388538551679996504301224629946714686799536156209624519841535728163249585706995546730976027641870202079879779584284425006451337438996740428983001001733580868266278580460151702279728130525792516349054757813921577822087141205648218581395399135318153873127142298313847722608029521851598;
            6'd61: xpb[22] = 1024'd88165208375867636658654571841841341966153060277102896583430993415027655324361899802561826006459001279093577490074211217054007575905816588507670760726070764344475791951703392340394890710433796991864570571336507362767870316546367003252436738111367874051249554532459689507793321948392291052982474312384200365269;
            6'd62: xpb[22] = 1024'd93678300174951523862855431295144132252309616252981163220147300030519154439099279763587923849668416851191608249172394792237813071931853592730916515000804089692211154920405782947208913154589013523577438862944884199743224284037976192583295654135594542454280527669520243697432770769642283792117226016738878878940;
            6'd63: xpb[22] = 1024'd99191391974035411067056290748446922538466172228859429856863606646010653553836659724614021692877832423289639008270578367421618567957890596954162269275537415039946517889108173554022935598744230055290307154553261036718578251529585381914154570159821210857311500806580797887072219590892276531251977721093557392611;
        endcase
    end

    always_comb begin
        case(flag[7][16:12])
            5'd0: xpb[23] = 1024'd0;
            5'd1: xpb[23] = 1024'd104704483773119298271257150201749712824622728204737696493579913261502152668574039685640119536087247995387669767368761942605424063983927601177408023550270740387681880857810564160836958042899446587003175446161637873693932219021194571245013486184047879260342473943641352076711668412142269270386729425448235906282;
            5'd2: xpb[23] = 1024'd85342271862113855143715372998684992904547029283739708859027971458027409999838940461265167857516821681332190127280030450631784287126634867799655922084210439841673087146049910984043676894281687452696153283936035901023503587821492369525048402684866309253865044473165646123316808750355905523654769024270877328233;
            5'd3: xpb[23] = 1024'd65980059951108412016173595795620272984471330362741721224476029654552667331103841236890216178946395367276710487191298958658144510269342134421903820618150139295664293434289257807250395745663928318389131121710433928353074956621790167805083319185684739247387615002689940169921949088569541776922808623093518750184;
            5'd4: xpb[23] = 1024'd46617848040102968888631818592555553064395631441743733589924087851077924662368742012515264500375969053221230847102567466684504733412049401044151719152089838749655499722528604630457114597046169184082108959484831955682646325422087966085118235686503169240910185532214234216527089426783178030190848221916160172135;
            5'd5: xpb[23] = 1024'd27255636129097525761090041389490833144319932520745745955372146047603181993633642788140312821805542739165751207013835974710864956554756667666399617686029538203646706010767951453663833448428410049775086797259229983012217694222385764365153152187321599234432756061738528263132229764996814283458887820738801594086;
            5'd6: xpb[23] = 1024'd7893424218092082633548264186426113224244233599747758320820204244128439324898543563765361143235116425110271566925104482737225179697463934288647516219969237657637912299007298276870552299810650915468064635033628010341789063022683562645188068688140029227955326591262822309737370103210450536726927419561443016037;
            5'd7: xpb[23] = 1024'd112597907991211380904805414388175826048866961804485454814400117505630591993472583249405480679322364420497941334293866425342649243681391535466055539770239978045319793156817862437707510342710097502471240081195265884035721282043878133890201554872187908488297800534904174386449038515352719807113656845009678922319;
            5'd8: xpb[23] = 1024'd93235696080205937777263637185111106128791262883487467179848175702155849324737484025030529000751938106442461694205134933369009466824098802088303438304179677499310999445057209260914229194092338368164217918969663911365292650844175932170236471373006338481820371064428468433054178853566356060381696443832320344270;
            5'd9: xpb[23] = 1024'd73873484169200494649721859982046386208715563962489479545296233898681106656002384800655577322181511792386982054116403441395369689966806068710551336838119376953302205733296556084120948045474579233857195756744061938694864019644473730450271387873824768475342941593952762479659319191779992313649736042654961766221;
            5'd10: xpb[23] = 1024'd54511272258195051522180082778981666288639865041491491910744292095206363987267285576280625643611085478331502414027671949421729913109513335332799235372059076407293412021535902907327666896856820099550173594518459966024435388444771528730306304374643198468865512123477056526264459529993628566917775641477603188172;
            5'd11: xpb[23] = 1024'd35149060347189608394638305575916946368564166120493504276192350291731621318532186351905673965040659164276022773938940457448090136252220601955047133905998775861284618309775249730534385748239060965243151432292857993354006757245069327010341220875461628462388082653001350572869599868207264820185815240300244610123;
            5'd12: xpb[23] = 1024'd15786848436184165267096528372852226448488467199495516641640408488256878649797087127530722286470232850220543133850208965474450359394927868577295032439938475315275824598014596553741104599621301830936129270067256020683578126045367125290376137376280058455910653182525644619474740206420901073453854839122886032074;
            5'd13: xpb[23] = 1024'd120491332209303463538353678574601939273111195404233213135220321749759031318371126813170841822557480845608212901218970908079874423378855469754703055990209215702957705455825160714578062642520748417939304716228893894377510345066561696535389623560327937716253127126166996696186408618563170343840584264571121938356;
            5'd14: xpb[23] = 1024'd101129120298298020410811901371537219353035496483235225500668379946284288649636027588795890143987054531552733261130239416106234646521562736376950954524148915156948911744064507537784781493902989283632282554003291921707081713866859494815424540061146367709775697655691290742791548956776806597108623863393763360307;
            5'd15: xpb[23] = 1024'd81766908387292577283270124168472499432959797562237237866116438142809545980900928364420938465416628217497253621041507924132594869664270002999198853058088614610940118032303854360991500345285230149325260391777689949036653082667157293095459456561964797703298268185215584789396689294990442850376663462216404782258;
            5'd16: xpb[23] = 1024'd62404696476287134155728346965407779512884098641239250231564496339334803312165829140045986786846201903441773980952776432158955092806977269621446751592028314064931324320543201184198219196667471015018238229552087976366224451467455091375494373062783227696820838714739878836001829633204079103644703061039046204209;
            5'd17: xpb[23] = 1024'd43042484565281691028186569762343059592808399720241262597012554535860060643430729915671035108275775589386294340864044940185315315949684536243694650125968013518922530608782548007404938048049711880711216067326486003695795820267752889655529289563601657690343409244264172882606969971417715356912742659861687626160;
            5'd18: xpb[23] = 1024'd23680272654276247900644792559278339672732700799243274962460612732385317974695630691296083429705349275330814700775313448211675539092391802865942548659907712972913736897021894830611656899431952746404193905100884031025367189068050687935564206064420087683865979773788466929212110309631351610180782258684329048111;
            5'd19: xpb[23] = 1024'd4318060743270804773103015356213619752657001878245287327908670928910575305960531466921131751134922961275335060686581956238035762235099069488190447193847412426904943185261241653818375750814193612097171742875282058354938557868348486215599122565238517677388550303312760975817250647844987863448821857506970470062;
            5'd20: xpb[23] = 1024'd109022544516390103044360165557963332577279730082982983821488584190412727974534571152561251287222170956663004828055343898843459826219026670665598470744118152814586824043071805814655333793713640199100347189036919932048870776889543057460612608749286396937731024246954113052528919059987257133835551282955206376344;
            5'd21: xpb[23] = 1024'd89660332605384659916818388354898612657204031161984996186936642386937985305799471928186299608651744642607525187966612406869820049361733937287846369278057852268578030331311152637862052645095881064793325026811317959378442145689840855740647525250104826931253594776478407099134059398200893387103590881777847798295;
            5'd22: xpb[23] = 1024'd70298120694379216789276611151833892737128332240987008552384700583463242637064372703811347930081318328552045547877880914896180272504441203910094267811997551722569236619550499461068771496478121930486302864585715986708013514490138654020682441750923256924776165306002701145739199736414529640371630480600489220246;
            5'd23: xpb[23] = 1024'd50935908783373773661734833948769172817052633319989020917832758779988499968329273479436396251510892014496565907789149422922540495647148470532342166345937251176560442907789846284275490347860362796179280702360114014037584883290436452300717358251741686918298735835526995192344340074628165893639670079423130642197;
            5'd24: xpb[23] = 1024'd31573696872368330534193056745704452896976934398991033283280816976513757299594174255061444572940465700441086267700417930948900718789855737154590064879876950630551649196029193107482209199242603661872258540134512041367156252090734250580752274752560116911821306365051289238949480412841802146907709678245772064148;
            5'd25: xpb[23] = 1024'd12211484961362887406651279542639732976901235477993045648728875173039014630859075030686492894370039386385606627611686438975260941932563003776837963413816650084542855484268539930688928050624844527565236377908910068696727620891032048860787191253378546905343876894575583285554620751055438400175749277068413486099;
            5'd26: xpb[23] = 1024'd116915968734482185677908429744389445801523963682730742142308788434541167299433114716326612430457287381773276394980448381580685005916490604954245986964087390472224736342079104091525886093524291114568411824070547942390659839912226620105800677437426426165686350838216935362266289163197707670562478702516649392381;
            5'd27: xpb[23] = 1024'd97553756823476742550366652541324725881448264761732754507756846631066424630698015491951660751886861067717796754891716889607045229059197871576493885498027089926215942630318450914732604944906531980261389661844945969720231208712524418385835593938244856159208921367741229408871429501411343923830518301339290814332;
            5'd28: xpb[23] = 1024'd78191544912471299422824875338260005961372565840734766873204904827591681961962916267576709073316434753662317114802985397633405452201905138198741784031966789380207148918557797737939323796288772845954367499619343997049802577512822216665870510439063286152731491897265523455476569839624980177098557900161932236283;
            5'd29: xpb[23] = 1024'd58829333001465856295283098135195286041296866919736779238652963024116939293227817043201757394746008439606837474714253905659765675344612404820989682565906488834198355206797144561146042647671013711647345337393742024379373946313120014945905426939881716146254062426789817502081710177838616430366597498984573658234;
            5'd30: xpb[23] = 1024'd39467121090460413167741320932130566121221167998738791604101021220642196624492717818826805716175582125551357834625522413686125898487319671443237581099846188288189561495036491384352761499053254577340323175168140051708945315113417813225940343440700146139776632956314111548686850516052252683634637097807215080185;
            5'd31: xpb[23] = 1024'd20104909179454970040199543729065846201145469077740803969549079417167453955757618594451854037605155811495878194536790921712486121630026938065485479633785887742180767783275838207559480350435495443033301012942538079038516683913715611505975259941518576133299203485838405595291990854265888936902676696629856502136;
        endcase
    end

    always_comb begin
        case(flag[8][5:0])
            6'd0: xpb[24] = 1024'd0;
            6'd1: xpb[24] = 1024'd62404696476287134155728346965407779512884098641239250231564496339334803312165829140045986786846201903441773980952776432158955092806977269621446751592028314064931324320543201184198219196667471015018238229552087976366224451467455091375494373062783227696820838714739878836001829633204079103644703061039046204209;
            6'd2: xpb[24] = 1024'd742697268449526912657766526001126281069770156742816334997137613692711287022519370076902359034729497440398554448059429738846344772734204687733378167725587196171974071515185030766199201817736308726278850716936106368088052714013409786010176442337006126821774015362699641897131192479525190170716295452497924087;
            6'd3: xpb[24] = 1024'd63147393744736661068386113491408905793953868797982066566561633953027514599188348510122889145880931400882172535400835861897801437579711474309180129759753901261103298392058386214964418398485207323744517080269024082734312504181468501161504549505120233823642612730102578477898960825683604293815419356491544128296;
            6'd4: xpb[24] = 1024'd1485394536899053825315533052002252562139540313485632669994275227385422574045038740153804718069458994880797108896118859477692689545468409375466756335451174392343948143030370061532398403635472617452557701433872212736176105428026819572020352884674012253643548030725399283794262384959050380341432590904995848174;
            6'd5: xpb[24] = 1024'd63890091013186187981043880017410032075023638954724882901558771566720225886210867880199791504915660898322571089848895291636647782352445678996913507927479488457275272463573571245730617600302943632470795930985960189102400556895481910947514725947457239950464386745465278119796092018163129483986135651944042052383;
            6'd6: xpb[24] = 1024'd2228091805348580737973299578003378843209310470228449004991412841078133861067558110230707077104188492321195663344178289216539034318202614063200134503176761588515922214545555092298597605453208926178836552150808319104264158142040229358030529327011018380465322046088098925691393577438575570512148886357493772261;
            6'd7: xpb[24] = 1024'd64632788281635714893701646543411158356093409111467699236555909180412937173233387250276693863950390395762969644296954721375494127125179883684646886095205075653447246535088756276496816802120679941197074781702896295470488609609495320733524902389794246077286160760827977761693223210642654674156851947396539976470;
            6'd8: xpb[24] = 1024'd2970789073798107650631066104004505124279080626971265339988550454770845148090077480307609436138917989761594217792237718955385379090936818750933512670902348784687896286060740123064796807270945234905115402867744425472352210856053639144040705769348024507287096061450798567588524769918100760682865181809991696348;
            6'd9: xpb[24] = 1024'd65375485550085241806359413069412284637163179268210515571553046794105648460255906620353596222985119893203368198745014151114340471897914088372380264262930662849619220606603941307263016003938416249923353632419832401838576662323508730519535078832131252204107934776190677403590354403122179864327568242849037900557;
            6'd10: xpb[24] = 1024'd3713486342247634563288832630005631405348850783714081674985688068463556435112596850384511795173647487201992772240297148694231723863671023438666890838627935980859870357575925153830996009088681543631394253584680531840440263570067048930050882211685030634108870076813498209485655962397625950853581477262489620435;
            6'd11: xpb[24] = 1024'd66118182818534768719017179595413410918232949424953331906550184407798359747278425990430498582019849390643766753193073580853186816670648293060113642430656250045791194678119126338029215205756152558649632483136768508206664715037522140305545255274468258330929708791553377045487485595601705054498284538301535824644;
            6'd12: xpb[24] = 1024'd4456183610697161475946599156006757686418620940456898009982825682156267722135116220461414154208376984642391326688356578433078068636405228126400269006353523177031844429091110184597195210906417852357673104301616638208528316284080458716061058654022036760930644092176197851382787154877151141024297772714987544522;
            6'd13: xpb[24] = 1024'd66860880086984295631674946121414537199302719581696148241547322021491071034300945360507400941054578888084165307641133010592033161443382497747847020598381837241963168749634311368795414407573888867375911333853704614574752767751535550091555431716805264457751482806916076687384616788081230244669000833754033748731;
            6'd14: xpb[24] = 1024'd5198880879146688388604365682007883967488391097199714344979963295848979009157635590538316513243106482082789881136416008171924413409139432814133647174079110373203818500606295215363394412724154161083951955018552744576616368998093868502071235096359042887752418107538897493279918347356676331195014068167485468609;
            6'd15: xpb[24] = 1024'd67603577355433822544332712647415663480372489738438964576544459635183782321323464730584303300089308385524563862089192440330879506216116702435580398766107424438135142821149496399561613609391625176102190184570640720942840820465548959877565608159142270584573256822278776329281747980560755434839717129206531672818;
            6'd16: xpb[24] = 1024'd5941578147596215301262132208009010248558161253942530679977100909541690296180154960615218872277835979523188435584475437910770758181873637501867025341804697569375792572121480246129593614541890469810230805735488850944704421712107278288081411538696049014574192122901597135177049539836201521365730363619983392696;
            6'd17: xpb[24] = 1024'd68346274623883349456990479173416789761442259895181780911541597248876493608345984100661205659124037882964962416537251870069725850988850907123313776933833011634307116892664681430327812811209361484828469035287576827310928873179562369663575784601479276711395030837641475971178879173040280625010433424659029596905;
            6'd18: xpb[24] = 1024'd6684275416045742213919898734010136529627931410685347014974238523234401583202674330692121231312565476963586990032534867649617102954607842189600403509530284765547766643636665276895792816359626778536509656452424957312792474426120688074091587981033055141395966138264296777074180732315726711536446659072481316783;
            6'd19: xpb[24] = 1024'd69088971892332876369648245699417916042512030051924597246538734862569204895368503470738108018158767380405360970985311299808572195761585111811047155101558598830479090964179866461094012013027097793554747886004512933679016925893575779449585961043816282838216804853004175613076010365519805815181149720111527520992;
            6'd20: xpb[24] = 1024'd7426972684495269126577665260011262810697701567428163349971376136927112870225193700769023590347294974403985544480594297388463447727342046877333781677255871961719740715151850307661992018177363087262788507169361063680880527140134097860101764423370061268217740153626996418971311924795251901707162954524979240870;
            6'd21: xpb[24] = 1024'd69831669160782403282306012225419042323581800208667413581535872476261916182391022840815010377193496877845759525433370729547418540534319316498780533269284186026651065035695051491860211214844834102281026736721449040047104978607589189235596137486153288965038578868366875254973141557999331005351866015564025445079;
            6'd22: xpb[24] = 1024'd8169669952944796039235431786012389091767471724170979684968513750619824157247713070845925949382024471844384098928653727127309792500076251565067159844981459157891714786667035338428191219995099395989067357886297170048968579854147507646111940865707067395039514168989696060868443117274777091877879249977477164957;
            6'd23: xpb[24] = 1024'd70574366429231930194963778751420168604651570365410229916533010089954627469413542210891912736228226375286158079881430159286264885307053521186513911437009773222823039107210236522626410416662570411007305587438385146415193031321602599021606313928490295091860352883729574896870272750478856195522582311016523369166;
            6'd24: xpb[24] = 1024'd8912367221394322951893198312013515372837241880913796019965651364312535444270232440922828308416753969284782653376713156866156137272810456252800538012707046354063688858182220369194390421812835704715346208603233276417056632568160917432122117308044073521861288184352395702765574309754302282048595545429975089044;
            6'd25: xpb[24] = 1024'd71317063697681457107621545277421294885721340522153046251530147703647338756436061580968815095262955872726556634329489589025111230079787725874247289604735360418995013178725421553392609618480306719733584438155321252783281084035616008807616490370827301218682126899092274538767403942958381385693298606469021293253;
            6'd26: xpb[24] = 1024'd9655064489843849864550964838014641653907012037656612354962788978005246731292751810999730667451483466725181207824772586605002482045544660940533916180432633550235662929697405399960589623630572013441625059320169382785144685282174327218132293750381079648683062199715095344662705502233827472219311840882473013131;
            6'd27: xpb[24] = 1024'd72059760966130984020279311803422421166791110678895862586527285317340050043458580951045717454297685370166955188777549018763957574852521930561980667772460947615166987250240606584158808820298043028459863288872257359151369136749629418593626666813164307345503900914454974180664535135437906575864014901921519217340;
            6'd28: xpb[24] = 1024'd10397761758293376777208731364015767934976782194399428689959926591697958018315271181076633026486212964165579762272832016343848826818278865628267294348158220746407637001212590430726788825448308322167903910037105489153232737996187737004142470192718085775504836215077794986559836694713352662390028136334970937218;
            6'd29: xpb[24] = 1024'd72802458234580510932937078329423547447860880835638678921524422931032761330481100321122619813332414867607353743225608448502803919625256135249714045940186534811338961321755791614925008022115779337186142139589193465519457189463642828379636843255501313472325674929817673822561666327917431766034731197374017141427;
            6'd30: xpb[24] = 1024'd11140459026742903689866497890016894216046552351142245024957064205390669305337790551153535385520942461605978316720891446082695171591013070316000672515883807942579611072727775461492988027266044630894182760754041595521320790710201146790152646635055091902326610230440494628456967887192877852560744431787468861305;
            6'd31: xpb[24] = 1024'd73545155503030037845594844855424673728930650992381495256521560544725472617503619691199522172367144365047752297673667878241650264397990339937447424107912122007510935393270976645691207223933515645912420990306129571887545242177656238165647019697838319599147448945180373464458797520396956956205447492826515065514;
            6'd32: xpb[24] = 1024'd11883156295192430602524264416018020497116322507885061359954201819083380592360309921230437744555671959046376871168950875821541516363747275003734050683609395138751585144242960492259187229083780939620461611470977701889408843424214556576162823077392098029148384245803194270354099079672403042731460727239966785392;
            6'd33: xpb[24] = 1024'd74287852771479564758252611381425800010000421149124311591518698158418183904526139061276424531401873862488150852121727307980496609170724544625180802275637709203682909464786161676457406425751251954638699841023065678255633294891669647951657196140175325725969222960543073106355928712876482146376163788279012989601;
            6'd34: xpb[24] = 1024'd12625853563641957515182030942019146778186092664627877694951339432776091879382829291307340103590401456486775425617010305560387861136481479691467428851334982334923559215758145523025386430901517248346740462187913808257496896138227966362172999519729104155970158261165893912251230272151928232902177022692464709479;
            6'd35: xpb[24] = 1024'd75030550039929091670910377907426926291070191305867127926515835772110895191548658431353326890436603359928549406569786737719342953943458749312914180443363296399854883536301346707223605627568988263364978691740001784623721347605683057737667372582512331852790996975905772748253059905356007336546880083731510913688;
            6'd36: xpb[24] = 1024'd13368550832091484427839797468020273059255862821370694029948477046468803166405348661384242462625130953927173980065069735299234205909215684379200807019060569531095533287273330553791585632719253557073019312904849914625584948852241376148183175962066110282791932276528593554148361464631453423072893318144962633566;
            6'd37: xpb[24] = 1024'd75773247308378618583568144433428052572139961462609944261512973385803606478571177801430229249471332857368947961017846167458189298716192954000647558611088883596026857607816531737989804829386724572091257542456937890991809400319696467523677549024849337979612770991268472390150191097835532526717596379184008837775;
            6'd38: xpb[24] = 1024'd14111248100541011340497563994021399340325632978113510364945614660161514453427868031461144821659860451367572534513129165038080550681949889066934185186786156727267507358788515584557784834536989865799298163621786020993673001566254785934193352404403116409613706291891293196045492657110978613243609613597460557653;
            6'd39: xpb[24] = 1024'd76515944576828145496225910959429178853209731619352760596510110999496317765593697171507131608506062354809346515465905597197035643488927158688380936778814470792198831679331716768756004031204460880817536393173873997359897453033709877309687725467186344106434545006631172032047322290315057716888312674636506761862;
            6'd40: xpb[24] = 1024'd14853945368990538253155330520022525621395403134856326699942752273854225740450387401538047180694589948807971088961188594776926895454684093754667563354511743923439481430303700615323984036354726174525577014338722127361761054280268195720203528846740122536435480307253992837942623849590503803414325909049958481740;
            6'd41: xpb[24] = 1024'd77258641845277672408883677485430305134279501776095576931507248613189029052616216541584033967540791852249745069913965026935881988261661363376114314946540057988370805750846901799522203233022197189543815243890810103727985505747723287095697901909523350233256319021993871673944453482794582907059028970089004685949;
            6'd42: xpb[24] = 1024'd15596642637440065165813097046023651902465173291599143034939889887546937027472906771614949539729319446248369643409248024515773240227418298442400941522237331119611455501818885646090183238172462483251855865055658233729849106994281605506213705289077128663257254322616692479839755042070028993585042204502456405827;
            6'd43: xpb[24] = 1024'd78001339113727199321541444011431431415349271932838393266504386226881740339638735911660936326575521349690143624362024456674728333034395568063847693114265645184542779822362086830288402434839933498270094094607746210096073558461736696881708078351860356360078093037356571315841584675274108097229745265541502610036;
            6'd44: xpb[24] = 1024'd16339339905889592078470863572024778183534943448341959369937027501239648314495426141691851898764048943688768197857307454254619585000152503130134319689962918315783429573334070676856382439990198791978134715772594340097937159708295015292223881731414134790079028337979392121736886234549554183755758499954954329914;
            6'd45: xpb[24] = 1024'd78744036382176726234199210537432557696419042089581209601501523840574451626661255281737838685610250847130542178810083886413574677807129772751581071281991232380714753893877271861054601636657669806996372945324682316464161611175750106667718254794197362486899867052719270957738715867753633287400461560994000534123;
            6'd46: xpb[24] = 1024'd17082037174339118991128630098025904464604713605084775704934165114932359601517945511768754257798778441129166752305366883993465929772886707817867697857688505511955403644849255707622581641807935100704413566489530446466025212422308425078234058173751140916900802353342091763634017427029079373926474795407452254001;
            6'd47: xpb[24] = 1024'd79486733650626253146856977063433683977488812246324025936498661454267162913683774651814741044644980344570940733258143316152421022579863977439314449449716819576886727965392456891820800838475406115722651796041618422832249663889763516453728431236534368613721641068081970599635847060233158477571177856446498458210;
            6'd48: xpb[24] = 1024'd17824734442788645903786396624027030745674483761827592039931302728625070888540464881845656616833507938569565306753426313732312274545620912505601076025414092708127377716364440738388780843625671409430692417206466552834113265136321834864244234616088147043722576368704791405531148619508604564097191090859950178088;
            6'd49: xpb[24] = 1024'd80229430919075780059514743589434810258558582403066842271495799067959874200706294021891643403679709842011339287706202745891267367352598182127047827617442406773058702036907641922587000040293142424448930646758554529200337716603776926239738607678871374740543415083444670241532978252712683667741894151898996382297;
            6'd50: xpb[24] = 1024'd18567431711238172816444163150028157026744253918570408374928440342317782175562984251922558975868237436009963861201485743471158619318355117193334454193139679904299351787879625769154980045443407718156971267923402659202201317850335244650254411058425153170544350384067491047428279811988129754267907386312448102175;
            6'd51: xpb[24] = 1024'd80972128187525306972172510115435936539628352559809658606492936681652585487728813391968545762714439339451737842154262175630113712125332386814781205785167993969230676108422826953353199242110878733175209497475490635568425769317790336025748784121208380867365189098807369883430109445192208857912610447351494306384;
            6'd52: xpb[24] = 1024'd19310128979687699729101929676029283307814024075313224709925577956010493462585503621999461334902966933450362415649545173210004964091089321881067832360865267100471325859394810799921179247261144026883250118640338765570289370564348654436264587500762159297366124399430190689325411004467654944438623681764946026262;
            6'd53: xpb[24] = 1024'd81714825455974833884830276641437062820698122716552474941490074295345296774751332762045448121749168836892136396602321605368960056898066591502514583952893581165402650179938011984119398443928615041901488348192426741936513822031803745811758960563545386994186963114170069525327240637671734048083326742803992230471;
            6'd54: xpb[24] = 1024'd20052826248137226641759696202030409588883794232056041044922715569703204749608022992076363693937696430890760970097604602948851308863823526568801210528590854296643299930909995830687378449078880335609528969357274871938377423278362064222274763943099165424187898414792890331222542196947180134609339977217443950349;
            6'd55: xpb[24] = 1024'd82457522724424360797488043167438189101767892873295291276487211909038008061773852132122350480783898334332534951050381035107806401670800796190247962120619168361574624251453197014885597645746351350627767198909362848304601874745817155597769137005882393121008737129532769167224371830151259238254043038256490154558;
            6'd56: xpb[24] = 1024'd20795523516586753554417462728031535869953564388798857379919853183395916036630542362153266052972425928331159524545664032687697653636557731256534588696316441492815274002425180861453577650896616644335807820074210978306465475992375474008284940385436171551009672430155589973119673389426705324780056272669941874436;
            6'd57: xpb[24] = 1024'd83200219992873887710145809693439315382837663030038107611484349522730719348796371502199252839818627831772933505498440464846652746443535000877981340288344755557746598322968382045651796847564087659354046049626298954672689927459830565383779313448219399247830511144895468809121503022630784428424759333708988078645;
            6'd58: xpb[24] = 1024'd21538220785036280467075229254032662151023334545541673714916990797088627323653061732230168412007155425771558078993723462426543998409291935944267966864042028688987248073940365892219776852714352953062086670791147084674553528706388883794295116827773177677831446445518289615016804581906230514950772568122439798523;
            6'd59: xpb[24] = 1024'd83942917261323414622803576219440441663907433186780923946481487136423430635818890872276155198853357329213332059946499894585499091216269205565714718456070342753918572394483567076417996049381823968080324900343235061040777980173843975169789489890556405374652285160258168451018634215110309618595475629161486002732;
            6'd60: xpb[24] = 1024'd22280918053485807379732995780033788432093104702284490049914128410781338610675581102307070771041884923211956633441782892165390343182026140632001345031767615885159222145455550922985976054532089261788365521508083191042641581420402293580305293270110183804653220460880989256913935774385755705121488863574937722610;
            6'd61: xpb[24] = 1024'd84685614529772941535461342745441567944977203343523740281478624750116141922841410242353057557888086826653730614394559324324345435989003410253448096623795929950090546465998752107184195251199560276806603751060171167408866032887857384955799666332893411501474059175620868092915765407589834808766191924613983926819;
            6'd62: xpb[24] = 1024'd23023615321935334292390762306034914713162874859027306384911266024474049897698100472383973130076614420652355187889842321904236687954760345319734723199493203081331196216970735953752175256349825570514644372225019297410729634134415703366315469712447189931474994476243688898811066966865280895292205159027435646697;
            6'd63: xpb[24] = 1024'd85428311798222468448119109271442694226046973500266556616475762363808853209863929612429959916922816324094129168842618754063191780761737614941181474791521517146262520537513937137950394453017296585532882601777107273776954085601870794741809842775230417628295833190983567734812896600069359998936908220066481850906;
        endcase
    end

    always_comb begin
        case(flag[8][11:6])
            6'd0: xpb[25] = 1024'd0;
            6'd1: xpb[25] = 1024'd23766312590384861205048528832036040994232645015770122719908403638166761184720619842460875489111343918092753742337901751643083032727494550007468101367218790277503170288485920984518374458167561879240923222941955403778817686848429113152325646154784196058296768491606388540708198159344806085462921454479933570784;
            6'd2: xpb[25] = 1024'd47532625180769722410097057664072081988465290031540245439816807276333522369441239684921750978222687836185507484675803503286166065454989100014936202734437580555006340576971841969036748916335123758481846445883910807557635373696858226304651292309568392116593536983212777081416396318689612170925842908959867141568;
            6'd3: xpb[25] = 1024'd71298937771154583615145586496108122982697935047310368159725210914500283554161859527382626467334031754278261227013705254929249098182483650022404304101656370832509510865457762953555123374502685637722769668825866211336453060545287339456976938464352588174890305474819165622124594478034418256388764363439800712352;
            6'd4: xpb[25] = 1024'd95065250361539444820194115328144163976930580063080490879633614552667044738882479369843501956445375672371014969351607006572332130909978200029872405468875161110012681153943683938073497832670247516963692891767821615115270747393716452609302584619136784233187073966425554162832792637379224341851685817919734283136;
            6'd5: xpb[25] = 1024'd118831562951924306025242644160180204971163225078850613599542018190833805923603099212304377445556719590463768711689508758215415163637472750037340506836093951387515851442429604922591872290837809396204616114709777018894088434242145565761628230773920980291483842458031942703540990796724030427314607272399667853920;
            6'd6: xpb[25] = 1024'd18531179858184425831492245587401813220697442968885052191318566764023671771014580144750181720010389199113373046569917075279434355523746965489648483186981700731328347161344308569480007557488165554135341729264492576308545270869677905948975307245475727082960707535521273214142660882140203495658838900254006940373;
            6'd7: xpb[25] = 1024'd42297492448569287036540774419437854214930087984655174911226970402190432955735199987211057209121733117206126788907818826922517388251241515497116584554200491008831517449830229553998382015655727433376264952206447980087362957718107019101300953400259923141257476027127661754850859041485009581121760354733940511157;
            6'd8: xpb[25] = 1024'd66063805038954148241589303251473895209162733000425297631135374040357194140455819829671932698233077035298880531245720578565600420978736065504584685921419281286334687738316150538516756473823289312617188175148403383866180644566536132253626599555044119199554244518734050295559057200829815666584681809213874081941;
            6'd9: xpb[25] = 1024'd89830117629339009446637832083509936203395378016195420351043777678523955325176439672132808187344420953391634273583622330208683453706230615512052787288638071563837858026802071523035130931990851191858111398090358787644998331414965245405952245709828315257851013010340438836267255360174621752047603263693807652725;
            6'd10: xpb[25] = 1024'd113596430219723870651686360915545977197628023031965543070952181316690716509897059514593683676455764871484388015921524081851766486433725165519520888655856861841341028315287992507553505390158413071099034621032314191423816018263394358558277891864612511316147781501946827376975453519519427837510524718173741223509;
            6'd11: xpb[25] = 1024'd13296047125983990457935962342767585447162240921999981662728729889880582357308540447039487950909434480133992350801932398915785678319999380971828865006744611185153524034202696154441640656808769229029760235587029748838272854890926698745624968336167258107624646579436157887577123604935600905854756346028080309962;
            6'd12: xpb[25] = 1024'd37062359716368851662984491174803626441394885937770104382637133528047343542029160289500363440020778398226746093139834150558868711047493930979296966373963401462656694322688617138960015114976331108270683458528985152617090541739355811897950614490951454165921415071042546428285321764280406991317677800508013880746;
            6'd13: xpb[25] = 1024'd60828672306753712868033020006839667435627530953540227102545537166214104726749780131961238929132122316319499835477735902201951743774988480986765067741182191740159864611174538123478389573143892987511606681470940556395908228587784925050276260645735650224218183562648934968993519923625213076780599254987947451530;
            6'd14: xpb[25] = 1024'd84594984897138574073081548838875708429860175969310349822453940804380865911470399974422114418243466234412253577815637653845034776502483030994233169108400982017663034899660459107996764031311454866752529904412895960174725915436214038202601906800519846282514952054255323509701718082970019162243520709467881022314;
            6'd15: xpb[25] = 1024'd108361297487523435278130077670911749424092820985080472542362344442547627096191019816882989907354810152505007320153539405488117809229977581001701270475619772295166205188146380092515138489479016745993453127354851363953543602284643151354927552955304042340811720545861712050409916242314825247706442163947814593098;
            6'd16: xpb[25] = 1024'd8060914393783555084379679098133357673627038875114911134138893015737492943602500749328794181808479761154611655033947722552137001116251796454009246826507521638978700907061083739403273756129372903924178741909566921368000438912175491542274629426858789132288585623351042561011586327730998316050673791802153679551;
            6'd17: xpb[25] = 1024'd31827226984168416289428207930169398667859683890885033854047296653904254128323120591789669670919823679247365397371849474195220033843746346461477348193726311916481871195547004723921648214296934783165101964851522325146818125760604604694600275581642985190585354114957431101719784487075804401513595246282087250335;
            6'd18: xpb[25] = 1024'd55593539574553277494476736762205439662092328906655156573955700292071015313043740434250545160031167597340119139709751225838303066571240896468945449560945102193985041484032925708440022672464496662406025187793477728925635812609033717846925921736427181248882122606563819642427982646420610486976516700762020821119;
            6'd19: xpb[25] = 1024'd79359852164938138699525265594241480656324973922425279293864103930237776497764360276711420649142511515432872882047652977481386099298735446476413550928163892471488211772518846692958397130632058541646948410735433132704453499457462830999251567891211377307178891098170208183136180805765416572439438155241954391903;
            6'd20: xpb[25] = 1024'd103126164755322999904573794426277521650557618938195402013772507568404537682484980119172296138253855433525626624385554729124469132026229996483881652295382682748991382061004767677476771588799620420887871633677388536483271186305891944151577214045995573365475659589776596723844378965110222657902359609721887962687;
            6'd21: xpb[25] = 1024'd2825781661583119710823395853499129900091836828229840605549056141594403529896461051618100412707525042175230959265963046188488323912504211936189628646270432092803877779919471324364906855449976578818597248232104093897728022933424284338924290517550320156952524667265927234446049050526395726246591237576227049140;
            6'd22: xpb[25] = 1024'd26592094251967980915871924685535170894324481843999963325457459779761164714617080894078975901818868960267984701603864797831571356639998761943657730013489222370307048068405392308883281313617538458059520471174059497676545709781853397491249936672334516215249293158872315775154247209871201811709512692056160619924;
            6'd23: xpb[25] = 1024'd50358406842352842120920453517571211888557126859770086045365863417927925899337700736539851390930212878360738443941766549474654389367493311951125831380708012647810218356891313293401655771785100337300443694116014901455363396630282510643575582827118712273546061650478704315862445369216007897172434146536094190708;
            6'd24: xpb[25] = 1024'd74124719432737703325968982349607252882789771875540208765274267056094687084058320579000726880041556796453492186279668301117737422094987861958593932747926802925313388645377234277920030229952662216541366917057970305234181083478711623795901228981902908331842830142085092856570643528560813982635355601016027761492;
            6'd25: xpb[25] = 1024'd97891032023122564531017511181643293877022416891310331485182670694261448268778940421461602369152900714546245928617570052760820454822482411966062034115145593202816558933863155262438404688120224095782290139999925709012998770327140736948226875136687104390139598633691481397278841687905620068098277055495961332276;
            6'd26: xpb[25] = 1024'd121657344613507425736066040013679334871255061907080454205091074332428209453499560263922477858264244632638999670955471804403903487549976961973530135482364383480319729222349076246956779146287785975023213362941881112791816457175569850100552521291471300448436367125297869937987039847250426153561198509975894903060;
            6'd27: xpb[25] = 1024'd21356961519767545542315641440900943120789279797114892796867622905618075300911041196368282132717914241288604005835880121467922679436251177425838111833252132824132224941263779893844914412938142132953938977496596670206273293803102190287899597763026047239913232202787200448588709932666599221905430137830233989513;
            6'd28: xpb[25] = 1024'd45123274110152406747364170272936984115021924812885015516776026543784836485631661038829157621829258159381357748173781873111005712163745727433306213200470923101635395229749700878363288871105704012194862200438552073985090980651531303440225243917810243298210000694393588989296908092011405307368351592310167560297;
            6'd29: xpb[25] = 1024'd68889586700537267952412699104973025109254569828655138236684430181951597670352280881290033110940602077474111490511683624754088744891240277440774314567689713379138565518235621862881663329273265891435785423380507477763908667499960416592550890072594439356506769185999977530005106251356211392831273046790101131081;
            6'd30: xpb[25] = 1024'd92655899290922129157461227937009066103487214844425260956592833820118358855072900723750908600051945995566865232849585376397171777618734827448242415934908503656641735806721542847400037787440827770676708646322462881542726354348389529744876536227378635414803537677606366070713304410701017478294194501270034701865;
            6'd31: xpb[25] = 1024'd116422211881306990362509756769045107097719859860195383676501237458285120039793520566211784089163289913659618975187487128040254810346229377455710517302127293934144906095207463831918412245608389649917631869264418285321544041196818642897202182382162831473100306169212754611421502570045823563757115955749968272649;
            6'd32: xpb[25] = 1024'd16121828787567110168759358196266715347254077750229822268277786031474985887205001498657588363616959522309223310067895445104274002232503592908018493653015043277957401814122167478806547512258745807848357483819133842736000877824350983084549258853717578264577171246702085122023172655461996632101347583604307359102;
            6'd33: xpb[25] = 1024'd39888141377951971373807887028302756341486722765999944988186189669641747071925621341118463852728303440401977052405797196747357034959998142915486595020233833555460572102608088463324921970426307687089280706761089246514818564672780096236874905008501774322873939738308473662731370814806802717564269038084240929886;
            6'd34: xpb[25] = 1024'd63654453968336832578856415860338797335719367781770067708094593307808508256646241183579339341839647358494730794743698948390440067687492692922954696387452623832963742391094009447843296428593869566330203929703044650293636251521209209389200551163285970381170708229914862203439568974151608803027190492564174500670;
            6'd35: xpb[25] = 1024'd87420766558721693783904944692374838329952012797540190428002996945975269441366861026040214830950991276587484537081600700033523100414987242930422797754671414110466912679579930432361670886761431445571127152645000054072453938369638322541526197318070166439467476721521250744147767133496414888490111947044108071454;
            6'd36: xpb[25] = 1024'd111187079149106554988953473524410879324184657813310313147911400584142030626087480868501090320062335194680238279419502451676606133142481792937890899121890204387970082968065851416880045344928993324812050375586955457851271625218067435693851843472854362497764245213127639284855965292841220973953033401524041642238;
            6'd37: xpb[25] = 1024'd10886696055366674795203074951632487573718875703344751739687949157331896473498961800946894594516004803329842614299910768740625325028756008390198875472777953731782578686980555063768180611579349482742775990141671015265728461845599775881198919944409109289241110290616969795457635378257394042297265029378380728691;
            6'd38: xpb[25] = 1024'd34653008645751536000251603783668528567951520719114874459596352795498657658219581643407770083627348721422596356637812520383708357756250558397666976839996744009285748975466476048286555069746911361983699213083626419044546148694028889033524566099193305347537878782223358336165833537602200127760186483858314299475;
            6'd39: xpb[25] = 1024'd58419321236136397205300132615704569562184165734884997179504756433665418842940201485868645572738692639515350098975714272026791390483745108405135078207215534286788919263952397032804929527914473241224622436025581822823363835542458002185850212253977501405834647273829746876874031696947006213223107938338247870259;
            6'd40: xpb[25] = 1024'd82185633826521258410348661447740610556416810750655119899413160071832180027660821328329521061850036557608103841313616023669874423211239658412603179574434324564292089552438318017323303986082035120465545658967537226602181522390887115338175858408761697464131415765436135417582229856291812298686029392818181441043;
            6'd41: xpb[25] = 1024'd105951946416906119615397190279776651550649455766425242619321563709998941212381441170790396550961380475700857583651517775312957455938734208420071280941653114841795259840924239001841678444249596999706468881909492630380999209239316228490501504563545893522428184257042523958290428015636618384148950847298115011827;
            6'd42: xpb[25] = 1024'd5651563323166239421646791706998259800183673656459681211098112283188807059792922103236200825415050084350461918531926092376976647825008423872379257292540864185607755559838942648729813710899953157637194496464208187795456045866848568677848581035100640313905049334531854468892098101052791452493182475152454098280;
            6'd43: xpb[25] = 1024'd29417875913551100626695320539034300794416318672229803931006515921355568244513541945697076314526394002443215660869827844020059680552502973879847358659759654463110925848324863633248188169067515036878117719406163591574273732715277681830174227189884836372201817826138243009600296260397597537956103929632387669064;
            6'd44: xpb[25] = 1024'd53184188503935961831743849371070341788648963687999926650914919559522329429234161788157951803637737920535969403207729595663142713279997523887315460026978444740614096136810784617766562627235076916119040942348118995353091419563706794982499873344669032430498586317744631550308494419742403623419025384112321239848;
            6'd45: xpb[25] = 1024'd76950501094320823036792378203106382782881608703770049370823323197689090613954781630618827292749081838628723145545631347306225746007492073894783561394197235018117266425296705602284937085402638795359964165290074399131909106412135908134825519499453228488795354809351020091016692579087209708881946838592254810632;
            6'd46: xpb[25] = 1024'd100716813684705684241840907035142423777114253719540172090731726835855851798675401473079702781860425756721476887883533098949308778734986623902251662761416025295620436713782626586803311543570200674600887388232029802910726793260565021287151165654237424547092123300957408631724890738432015794344868293072188381416;
            6'd47: xpb[25] = 1024'd416430590965804048090508462364032026648471609574610682508275409045717646086882405525507056314095365371081222763941416013327970621260839354559639112303774639432932432697330233691446810220556832531613002786745360325183629888097361474498242125792171338568988378446739142326560823848188862689099920926527467869;
            6'd48: xpb[25] = 1024'd24182743181350665253139037294400073020881116625344733402416679047212478830807502247986382545425439283463834965101843167656411003348755389362027740479522564916936102721183251218209821268388118711772536225728700764104001316736526474626823888280576367396865756870053127683034758983192994948152021375406461038653;
            6'd49: xpb[25] = 1024'd47949055771735526458187566126436114015113761641114856122325082685379240015528122090447258034536783201556588707439744919299494036076249939369495841846741355194439273009669172202728195726555680591013459448670656167882819003584955587779149534435360563455162525361659516223742957142537801033614942829886394609437;
            6'd50: xpb[25] = 1024'd71715368362120387663236094958472155009346406656884978842233486323546001200248741932908133523648127119649342449777646670942577068803744489376963943213960145471942443298155093187246570184723242470254382671612611571661636690433384700931475180590144759513459293853265904764451155301882607119077864284366328180221;
            6'd51: xpb[25] = 1024'd95481680952505248868284623790508196003579051672655101562141889961712762384969361775369009012759471037742096192115548422585660101531239039384432044581178935749445613586641014171764944642890804349495305894554566975440454377281813814083800826744928955571756062344872293305159353461227413204540785738846261751005;
            6'd52: xpb[25] = 1024'd119247993542890110073333152622544236997811696688425224282050293599879523569689981617829884501870814955834849934453450174228743134258733589391900145948397726026948783875126935156283319101058366228736229117496522379219272064130242927236126472899713151630052830836478681845867551620572219290003707193326195321789;
            6'd53: xpb[25] = 1024'd18947610449150229879582754049765845247345914578459662873826842173069389417101462550275688776324484564484454269333858491292762326145007804844208122299285475370761279594041638803171454367708722386666954732051237936633728900757775267423473549371267898421529695913968012356469221705988392358347938821180534408242;
            6'd54: xpb[25] = 1024'd42713923039535091084631282881801886241578559594229785593735245811236150601822082392736564265435828482577208011671760242935845358872502354851676223666504265648264449882527559787689828825876284265907877954993193340412546587606204380575799195526052094479826464405574400897177419865333198443810860275660467979026;
            6'd55: xpb[25] = 1024'd66480235629919952289679811713837927235811204609999908313643649449402911786542702235197439754547172400669961754009661994578928391599996904859144325033723055925767620171013480772208203284043846145148801177935148744191364274454633493728124841680836290538123232897180789437885618024678004529273781730140401549810;
            6'd56: xpb[25] = 1024'd90246548220304813494728340545873968230043849625770031033552053087569672971263322077658315243658516318762715496347563746222011424327491454866612426400941846203270790459499401756726577742211408024389724400877104147970181961303062606880450487835620486596420001388787177978593816184022810614736703184620335120594;
            6'd57: xpb[25] = 1024'd114012860810689674699776869377910009224276494641540153753460456725736434155983941920119190732769860236855469238685465497865094457054986004874080527768160636480773960747985322741244952200378969903630647623819059551748999648151491720032776133990404682654716769880393566519302014343367616700199624639100268691378;
            6'd58: xpb[25] = 1024'd13712477716949794506026470805131617473810712531574592345237005298926300003395422852564995007223529845505073573565873814929113648941260220326388504119048385824586456466900026388133087467029326061561373238373775109163456484779024060220123210461959429446193634957882897029903684428783789768543856266954607777831;
            6'd59: xpb[25] = 1024'd37478790307334655711074999637167658468043357547344715065145408937093061188116042695025870496334873763597827315903775566572196681668754770333856605486267176102089626755385947372651461925196887940802296461315730512942274171627453173372448856616743625504490403449489285570611882588128595854006777721434541348615;
            6'd60: xpb[25] = 1024'd61245102897719516916123528469203699462276002563114837785053812575259822372836662537486745985446217681690581058241677318215279714396249320341324706853485966379592797043871868357169836383364449820043219684257685916721091858475882286524774502771527821562787171941095674111320080747473401939469699175914474919399;
            6'd61: xpb[25] = 1024'd85011415488104378121172057301239740456508647578884960504962216213426583557557282379947621474557561599783334800579579069858362747123743870348792808220704756657095967332357789341688210841532011699284142907199641320499909545324311399677100148926312017621083940432702062652028278906818208024932620630394408490183;
            6'd62: xpb[25] = 1024'd108777728078489239326220586133275781450741292594655083224870619851593344742277902222408496963668905517876088542917480821501445779851238420356260909587923546934599137620843710326206585299699573578525066130141596724278727232172740512829425795081096213679380708924308451192736477066163014110395542084874342060967;
            6'd63: xpb[25] = 1024'd8477344984749359132470187560497389700275510484689521816647168424783210589689383154854301238122575126525692877797889138565464971737512635808568885938811296278411633339758413973094720566349929736455791744696312281693184068800272853016772871552650960470857574001797781703338147151579187178739773712728681147420;
        endcase
    end

    always_comb begin
        case(flag[8][16:12])
            5'd0: xpb[26] = 1024'd0;
            5'd1: xpb[26] = 1024'd32243657575134220337518716392533430694508155500459644536555572062949971774410002997315176727233919044618446620135790890208548004465007185816036987306030086555914803628244334957613095024517491615696714967638267685472001755648701966169098517707435156529154342493404170244046345310923993264202695167208614718204;
            5'd2: xpb[26] = 1024'd64487315150268440675037432785066861389016311000919289073111144125899943548820005994630353454467838089236893240271581780417096008930014371632073974612060173111829607256488669915226190049034983231393429935276535370944003511297403932338197035414870313058308684986808340488092690621847986528405390334417229436408;
            5'd3: xpb[26] = 1024'd96730972725402661012556149177600292083524466501378933609666716188849915323230008991945530181701757133855339860407372670625644013395021557448110961918090259667744410884733004872839285073552474847090144902914803056416005266946105898507295553122305469587463027480212510732139035932771979792608085501625844154612;
            5'd4: xpb[26] = 1024'd4907934616412139951275938165319290033334194876102894018090433186822991760330873079245635694278001869030637073085670126255128177018808408708987824207789305289968539943406122492822140906552760741476662262165830895523646172373911091711415501146511176849797466559499622946078853169767340039692090842208864388485;
            5'd5: xpb[26] = 1024'd37151592191546360288794654557852720727842350376562538554646005249772963534740876076560812421511920913649083693221461016463676181483815594525024811513819391845883343571650457450435235931070252357173377229804098580995647928022613057880514018853946333378951809052903793190125198480691333303894786009417479106689;
            5'd6: xpb[26] = 1024'd69395249766680580626313370950386151422350505877022183091201577312722935309150879073875989148745839958267530313357251906672224185948822780341061798819849478401798147199894792408048330955587743972870092197442366266467649683671315024049612536561381489908106151546307963434171543791615326568097481176626093824893;
            5'd7: xpb[26] = 1024'd101638907341814800963832087342919582116858661377481827627757149375672907083560882071191165875979759002885976933493042796880772190413829966157098786125879564957712950828139127365661425980105235588566807165080633951939651439320016990218711054268816646437260494039712133678217889102539319832300176343834708543097;
            5'd8: xpb[26] = 1024'd9815869232824279902551876330638580066668389752205788036180866373645983520661746158491271388556003738061274146171340252510256354037616817417975648415578610579937079886812244985644281813105521482953324524331661791047292344747822183422831002293022353699594933118999245892157706339534680079384181684417728776970;
            5'd9: xpb[26] = 1024'd42059526807958500240070592723172010761176545252665432572736438436595955295071749155806448115789922782679720766307131142718804358502624003234012635721608697135851883515056579943257376837623013098650039491969929476519294100396524149591929520000457510228749275612403416136204051650458673343586876851626343495174;
            5'd10: xpb[26] = 1024'd74303184383092720577589309115705441455684700753125077109292010499545927069481752153121624843023841827298167386442922032927352362967631189050049623027638783691766687143300914900870471862140504714346754459608197161991295856045226115761028037707892666757903618105807586380250396961382666607789572018834958213378;
            5'd11: xpb[26] = 1024'd106546841958226940915108025508238872150192856253584721645847582562495898843891755150436801570257760871916614006578712923135900367432638374866086610333668870247681490771545249858483566886657996330043469427246464847463297611693928081930126555415327823287057960599211756624296742272306659871992267186043572931582;
            5'd12: xpb[26] = 1024'd14723803849236419853827814495957870100002584628308682054271299560468975280992619237736907082834005607091911219257010378765384531056425226126963472623367915869905619830218367478466422719658282224429986786497492686570938517121733275134246503439533530549392399678498868838236559509302020119076272526626593165455;
            5'd13: xpb[26] = 1024'd46967461424370640191346530888491300794510740128768326590826871623418947055402622235052083810067924651710357839392801268973932535521432411943000459929398002425820423458462702436079517744175773840126701754135760372042940272770435241303345021146968687078546742171903039082282904820226013383278967693835207883659;
            5'd14: xpb[26] = 1024'd79211118999504860528865247281024731489018895629227971127382443686368918829812625232367260537301843696328804459528592159182480539986439597759037447235428088981735227086707037393692612768693265455823416721774028057514942028419137207472443538854403843607701084665307209326329250131150006647481662861043822601863;
            5'd15: xpb[26] = 1024'd111454776574639080866383963673558162183527051129687615663938015749318890604222628229682437264535762740947251079664383049391028544451446783575074434541458175537650030714951372351305707793210757071520131689412295742986943784067839173641542056561839000136855427158711379570375595442073999911684358028252437320067;
            5'd16: xpb[26] = 1024'd19631738465648559805103752661277160133336779504411576072361732747291967041323492316982542777112007476122548292342680505020512708075233634835951296831157221159874159773624489971288563626211042965906649048663323582094584689495644366845662004586044707399189866237998491784315412679069360158768363368835457553940;
            5'd17: xpb[26] = 1024'd51875396040782780142622469053810590827844935004871220608917304810241938815733495314297719504345926520740994912478471395229060712540240820651988284137187307715788963401868824928901658650728534581603364016301591267566586445144346333014760522293479863928344208731402662028361757989993353422971058536044072272144;
            5'd18: xpb[26] = 1024'd84119053615917000480141185446344021522353090505330865145472876873191910590143498311612896231579845565359441532614262285437608717005248006468025271443217394271703767030113159886514753675246026197300078983939858953038588200793048299183859040000915020457498551224806832272408103300917346687173753703252686990348;
            5'd19: xpb[26] = 1024'd116362711191051220817659901838877452216861246005790509682028448936141882364553501308928072958813764609977888152750053175646156721470255192284062258749247480827618570658357494844127848699763517812996793951578126638510589956441750265352957557708350176986652893718211002516454448611841339951376448870461301708552;
            5'd20: xpb[26] = 1024'd24539673082060699756379690826596450166670974380514470090452165934114958801654365396228178471390009345153185365428350631275640885094042043544939121038946526449842699717030612464110704532763803707383311310829154477618230861869555458557077505732555884248987332797498114730394265848836700198460454211044321942425;
            5'd21: xpb[26] = 1024'd56783330657194920093898407219129880861179129880974114627007737997064930576064368393543355198623928389771631985564141521484188889559049229360976108344976613005757503345274947421723799557281295323080026278467422163090232617518257424726176023439991040778141675290902284974440611159760693462663149378252936660629;
            5'd22: xpb[26] = 1024'd89026988232329140431417123611663311555687285381433759163563310060014902350474371390858531925857847434390078605699932411692736894024056415177013095651006699561672306973519282379336894581798786938776741246105689848562234373166959390895274541147426197307296017784306455218486956470684686726865844545461551378833;
            5'd23: xpb[26] = 1024'd121270645807463360768935840004196742250195440881893403700118882122964874124884374388173708653091766479008525225835723301901284898489063600993050082957036786117587110601763617336949989606316278554473456213743957534034236128815661357064373058854861353836450360277710625462533301781608679991068539712670166097037;
            5'd24: xpb[26] = 1024'd29447607698472839707655628991915740200005169256617364108542599120937950561985238475473814165668011214183822438514020757530769062112850452253926945246735831739811239660436734956932845439316564448859973572994985373141877034243466550268493006879067061098784799356997737676473119018604040238152545053253186330910;
            5'd25: xpb[26] = 1024'd61691265273607060045174345384449170894513324757077008645098171183887922336395241472788990892901930258802269058649811647739317066577857638069963932552765918295726043288681069914545940463834056064556688540633253058613878789892168516437591524586502217627939141850401907920519464329528033502355240220461801049114;
            5'd26: xpb[26] = 1024'd93934922848741280382693061776982601589021480257536653181653743246837894110805244470104167620135849303420715678785602537947865071042864823886000919858796004851640846916925404872159035488351547680253403508271520744085880545540870482606690042293937374157093484343806078164565809640452026766557935387670415767318;
            5'd27: xpb[26] = 1024'd2111884739750759321412850764701599538831208632260613590077460244810970547906108557404273132712094038596012891463899993577349234666651675146877782148495050473864975975598522492141891321351833574639920867522548583193521450968675675810809990318143081419427923423093190378505626877447387013641940728253436001191;
            5'd28: xpb[26] = 1024'd34355542314884979658931567157235030233339364132720258126633032307760942322316111554719449859946013083214459511599690883785897239131658860962914769454525137029779779603842857449754986345869325190336635835160816268665523206617377641979908508025578237948582265916497360622551972188371380277844635895462050719395;
            5'd29: xpb[26] = 1024'd66599199890019199996450283549768460927847519633179902663188604370710914096726114552034626587179932127832906131735481773994445243596666046778951756760555223585694583232087192407368081370386816806033350802799083954137524962266079608149007025733013394477736608409901530866598317499295373542047331062670665437599;
            5'd30: xpb[26] = 1024'd98842857465153420333968999942301891622355675133639547199744176433660885871136117549349803314413851172451352751871272664202993248061673232594988744066585310141609386860331527364981176394904308421730065770437351639609526717914781574318105543440448551006890950903305701110644662810219366806250026229879280155803;
            5'd31: xpb[26] = 1024'd7019819356162899272688788930020889572165403508363507608167893431633962308236981636649908826990095907626649964549570119832477411685460083855865606356284355763833515919004644984964032227904594316116583129688379478717167623342586767522225491464654258269225389982592813324584480047214727053334031570462300389676;
        endcase
    end

    always_comb begin
        case(flag[9][5:0])
            6'd0: xpb[27] = 1024'd0;
            6'd1: xpb[27] = 1024'd19631738465648559805103752661277160133336779504411576072361732747291967041323492316982542777112007476122548292342680505020512708075233634835951296831157221159874159773624489971288563626211042965906649048663323582094584689495644366845662004586044707399189866237998491784315412679069360158768363368835457553940;
            6'd2: xpb[27] = 1024'd39263476931297119610207505322554320266673559008823152144723465494583934082646984633965085554224014952245096584685361010041025416150467269671902593662314442319748319547248979942577127252422085931813298097326647164189169378991288733691324009172089414798379732475996983568630825358138720317536726737670915107880;
            6'd3: xpb[27] = 1024'd58895215396945679415311257983831480400010338513234728217085198241875901123970476950947628331336022428367644877028041515061538124225700904507853890493471663479622479320873469913865690878633128897719947145989970746283754068486933100536986013758134122197569598713995475352946238037208080476305090106506372661820;
            6'd4: xpb[27] = 1024'd78526953862594239220415010645108640533347118017646304289446930989167868165293969267930171108448029904490193169370722020082050832300934539343805187324628884639496639094497959885154254504844171863626596194653294328378338757982577467382648018344178829596759464951993967137261650716277440635073453475341830215760;
            6'd5: xpb[27] = 1024'd98158692328242799025518763306385800666683897522057880361808663736459835206617461584912713885560037380612741461713402525102563540376168174179756484155786105799370798868122449856442818131055214829533245243316617910472923447478221834228310022930223536995949331189992458921577063395346800793841816844177287769700;
            6'd6: xpb[27] = 1024'd117790430793891358830622515967662960800020677026469456434170396483751802247940953901895256662672044856735289754056083030123076248451401809015707780986943326959244958641746939827731381757266257795439894291979941492567508136973866201073972027516268244395139197427990950705892476074416160952610180213012745323640;
            6'd7: xpb[27] = 1024'd13355473575415177236927341224125688188659029405145348378400274166066873951955307308862728225126378023414688638941270100564525115685415109296498952801769507185428443845800212461389706191960095040036345732256025228297731976248613794954655462419083502527509160251872384460101360679556888094259853755222608393249;
            6'd8: xpb[27] = 1024'd32987212041063737042031093885402848321995808909556924450762006913358840993278799625845271002238385499537236931283950605585037823760648744132450249632926728345302603619424702432678269818171138005942994780919348810392316665744258161800317467005128209926699026489870876244416773358626248253028217124058065947189;
            6'd9: xpb[27] = 1024'd52618950506712296847134846546680008455332588413968500523123739660650808034602291942827813779350392975659785223626631110605550531835882378968401546464083949505176763393049192403966833444382180971849643829582672392486901355239902528645979471591172917325888892727869368028732186037695608411796580492893523501129;
            6'd10: xpb[27] = 1024'd72250688972360856652238599207957168588669367918380076595485472407942775075925784259810356556462400451782333515969311615626063239911116013804352843295241170665050923166673682375255397070593223937756292878245995974581486044735546895491641476177217624725078758965867859813047598716764968570564943861728981055069;
            6'd11: xpb[27] = 1024'd91882427438009416457342351869234328722006147422791652667847205155234742117249276576792899333574407927904881808311992120646575947986349648640304140126398391824925082940298172346543960696804266903662941926909319556676070734231191262337303480763262332124268625203866351597363011395834328729333307230564438609009;
            6'd12: xpb[27] = 1024'd111514165903657976262446104530511488855342926927203228740208937902526709158572768893775442110686415404027430100654672625667088656061583283476255436957555612984799242713922662317832524323015309869569590975572643138770655423726835629182965485349307039523458491441864843381678424074903688888101670599399896162949;
            6'd13: xpb[27] = 1024'd7079208685181794668750929786974216243981279305879120684438815584841780862587122300742913673140748570706828985539859696108537523295596583757046608772381793210982727917975934951490848757709147114166042415848726874500879263001583223063648920252122297655828454265746277135887308680044416029751344141609759232558;
            6'd14: xpb[27] = 1024'd26710947150830354473854682448251376377318058810290696756800548332133747903910614617725456450252756046829377277882540201129050231370830218592997905603539014370856887691600424922779412383920190080072691464512050456595463952497227589909310924838167005055018320503744768920202721359113776188519707510445216786498;
            6'd15: xpb[27] = 1024'd46342685616478914278958435109528536510654838314702272829162281079425714945234106934707999227364763522951925570225220706149562939446063853428949202434696235530731047465224914894067976010131233045979340513175374038690048641992871956754972929424211712454208186741743260704518134038183136347288070879280674340438;
            6'd16: xpb[27] = 1024'd65974424082127474084062187770805696643991617819113848901524013826717681986557599251690542004476770999074473862567901211170075647521297488264900499265853456690605207238849404865356539636342276011885989561838697620784633331488516323600634934010256419853398052979741752488833546717252496506056434248116131894378;
            6'd17: xpb[27] = 1024'd85606162547776033889165940432082856777328397323525424973885746574009649027881091568673084781588778475197022154910581716190588355596531123100851796097010677850479367012473894836645103262553318977792638610502021202879218020984160690446296938596301127252587919217740244273148959396321856664824797616951589448318;
            6'd18: xpb[27] = 1024'd105237901013424593694269693093360016910665176827937001046247479321301616069204583885655627558700785951319570447253262221211101063671764757936803092928167899010353526786098384807933666888764361943699287659165344784973802710479805057291958943182345834651777785455738736057464372075391216823593160985787047002258;
            6'd19: xpb[27] = 1024'd802943794948412100574518349822744299303529206612892990477357003616687773218937292623099121155119117998969332138449291652549930905778058217594264742994079236537011990151657441591991323458199188295739099441428520704026549754552651172642378085161092784147748279620169811673256680531943965242834527996910071867;
            6'd20: xpb[27] = 1024'd20434682260596971905678271011099904432640308711024469062839089750908654814542429609605641898267126594121517624481129796673062638981011693053545561574151300396411171763776147412880554949669242154202388148104752102798611239250197018018304382671205800183337614517618661595988669359601304124011197896832367625807;
            6'd21: xpb[27] = 1024'd40066420726245531710782023672377064565977088215436045135200822498200621855865921926588184675379134070244065916823810301693575347056245327889496858405308521556285331537400637384169118575880285120109037196768075684893195928745841384863966387257250507582527480755617153380304082038670664282779561265667825179747;
            6'd22: xpb[27] = 1024'd59698159191894091515885776333654224699313867719847621207562555245492588897189414243570727452491141546366614209166490806714088055131478962725448155236465742716159491311025127355457682202091328086015686245431399266987780618241485751709628391843295214981717346993615645164619494717740024441547924634503282733687;
            6'd23: xpb[27] = 1024'd79329897657542651320989528994931384832650647224259197279924287992784555938512906560553270229603149022489162501509171311734600763206712597561399452067622963876033651084649617326746245828302371051922335294094722849082365307737130118555290396429339922380907213231614136948934907396809384600316288003338740287627;
            6'd24: xpb[27] = 1024'd98961636123191211126093281656208544965987426728670773352286020740076522979836398877535813006715156498611710793851851816755113471281946232397350748898780185035907810858274107298034809454513414017828984342758046431176949997232774485400952401015384629780097079469612628733250320075878744759084651372174197841567;
            6'd25: xpb[27] = 1024'd118593374588839770931197034317485705099324206233082349424647753487368490021159891194518355783827163974734259086194532321775626179357179867233302045729937406195781970631898597269323373080724456983735633391421370013271534686728418852246614405601429337179286945707611120517565732754948104917853014741009655395507;
            6'd26: xpb[27] = 1024'd14158417370363589337501859573948432487962558611758241368877631169683561725174244601485827346281497141413657971079719392217075046591193167514093217544763586421965455835951869902981697515418294228332084831697453749001758526003166446127297840504244595311656908531492554271774617360088832059502688283219518465116;
            6'd27: xpb[27] = 1024'd33790155836012149142605612235225592621299338116169817441239363916975528766497736918468370123393504617536206263422399897237587754666426802350044514375920807581839615609576359874270261141629337194238733880360777331096343215498810812972959845090289302710846774769491046056090030039158192218271051652054976019056;
            6'd28: xpb[27] = 1024'd53421894301660708947709364896502752754636117620581393513601096664267495807821229235450912900505512093658754555765080402258100462741660437185995811207078028741713775383200849845558824767840380160145382929024100913190927904994455179818621849676334010110036641007489537840405442718227552377039415020890433572996;
            6'd29: xpb[27] = 1024'd73053632767309268752813117557779912887972897124992969585962829411559462849144721552433455677617519569781302848107760907278613170816894072021947108038235249901587935156825339816847388394051423126052031977687424495285512594490099546664283854262378717509226507245488029624720855397296912535807778389725891126936;
            6'd30: xpb[27] = 1024'd92685371232957828557916870219057073021309676629404545658324562158851429890468213869415998454729527045903851140450441412299125878892127706857898404869392471061462094930449829788135952020262466091958681026350748077380097283985743913509945858848423424908416373483486521409036268076366272694576141758561348680876;
            6'd31: xpb[27] = 1024'd112317109698606388363020622880334233154646456133816121730686294906143396931791706186398541231841534522026399432793121917319638586967361341693849701700549692221336254704074319759424515646473509057865330075014071659474681973481388280355607863434468132307606239721485013193351680755435632853344505127396806234816;
            6'd32: xpb[27] = 1024'd7882152480130206769325448136796960543284808512492013674916172588458468635806059593366012794295867688705798317678308987761087454201374641974640873515375872447519739908127592393082840081167346302461781515290155395204905812756135874236291298337283390439976202545366446947560565360576359994994178669606669304425;
            6'd33: xpb[27] = 1024'd27513890945778766574429200798074120676621588016903589747277905335750435677129551910348555571407875164828346610020989492781600162276608276810592170346533093607393899681752082364371403707378389268368430563953478977299490502251780241081953302923328097839166068783364938731875978039645720153762542038442126858365;
            6'd34: xpb[27] = 1024'd47145629411427326379532953459351280809958367521315165819639638083042402718453044227331098348519882640950894902363669997802112870351841911646543467177690314767268059455376572335659967333589432234275079612616802559394075191747424607927615307509372805238355935021363430516191390718715080312530905407277584412305;
            6'd35: xpb[27] = 1024'd66777367877075886184636706120628440943295147025726741892001370830334369759776536544313641125631890117073443194706350502822625578427075546482494764008847535927142219229001062306948530959800475200181728661280126141488659881243068974773277312095417512637545801259361922300506803397784440471299268776113041966245;
            6'd36: xpb[27] = 1024'd86409106342724445989740458781905601076631926530138317964363103577626336801100028861296183902743897593195991487049031007843138286502309181318446060840004757087016379002625552278237094586011518166088377709943449723583244570738713341618939316681462220036735667497360414084822216076853800630067632144948499520185;
            6'd37: xpb[27] = 1024'd106040844808373005794844211443182761209968706034549894036724836324918303842423521178278726679855905069318539779391711512863650994577542816154397357671161978246890538776250042249525658212222561131995026758606773305677829260234357708464601321267506927435925533735358905869137628755923160788835995513783957074125;
            6'd38: xpb[27] = 1024'd1605887589896824201149036699645488598607058413225785980954714007233375546437874585246198242310238235997938664276898583305099861811556116435188529485988158473074023980303314883183982646916398376591478198882857041408053099509105302345284756170322185568295496559240339623346513361063887930485669055993820143734;
            6'd39: xpb[27] = 1024'd21237626055545384006252789360922648731943837917637362053316446754525342587761366902228741019422245712120486956619579088325612569886789751271139826317145379632948183753927804854472546273127441342498127247546180623502637789004749669190946760756366892967485362797238831407661926040133248089254032424829277697674;
            6'd40: xpb[27] = 1024'd40869364521193943811356542022199808865280617422048938125678179501817309629084859219211283796534253188243035248962259593346125277962023386107091123148302600792822343527552294825761109899338484308404776296209504205597222478500394036036608765342411600366675229035237323191977338719202608248022395793664735251614;
            6'd41: xpb[27] = 1024'd60501102986842503616460294683476968998617396926460514198039912249109276670408351536193826573646260664365583541304940098366637986037257020943042419979459821952696503301176784797049673525549527274311425344872827787691807167996038402882270769928456307765865095273235814976292751398271968406790759162500192805554;
            6'd42: xpb[27] = 1024'd80132841452491063421564047344754129131954176430872090270401644996401243711731843853176369350758268140488131833647620603387150694112490655778993716810617043112570663074801274768338237151760570240218074393536151369786391857491682769727932774514501015165054961511234306760608164077341328565559122531335650359494;
            6'd43: xpb[27] = 1024'd99764579918139623226667800006031289265290955935283666342763377743693210753055336170158912127870275616610680125990301108407663402187724290614945013641774264272444822848425764739626800777971613206124723442199474951880976546987327136573594779100545722564244827749232798544923576756410688724327485900171107913434;
            6'd44: xpb[27] = 1024'd119396318383788183031771552667308449398627735439695242415125110490985177794378828487141454904982283092733228418332981613428176110262957925450896310472931485432318982622050254710915364404182656172031372490862798533975561236482971503419256783686590429963434693987231290329238989435480048883095849269006565467374;
            6'd45: xpb[27] = 1024'd14961361165312001438076377923771176787266087818371134359354988173300249498393181894108926467436616259412627303218168683869624977496971225731687482287757665658502467826103527344573688838876493416627823931138882269705785075757719097299940218589405688095804656811112724083447874040620776024745522811216428536983;
            6'd46: xpb[27] = 1024'd34593099630960561243180130585048336920602867322782710431716720920592216539716674211091469244548623735535175595560849188890137685572204860567638779118914886818376627599728017315862252465087536382534472979802205851800369765253363464145602223175450395494994523049111215867763286719690136183513886180051886090923;
            6'd47: xpb[27] = 1024'd54224838096609121048283883246325497053939646827194286504078453667884183581040166528074012021660631211657723887903529693910650393647438495403590075950072107978250787373352507287150816091298579348441122028465529433894954454749007830991264227761495102894184389287109707652078699398759496342282249548887343644863;
            6'd48: xpb[27] = 1024'd73856576562257680853387635907602657187276426331605862576440186415176150622363658845056554798772638687780272180246210198931163101722672130239541372781229329138124947146976997258439379717509622314347771077128853015989539144244652197836926232347539810293374255525108199436394112077828856501050612917722801198803;
            6'd49: xpb[27] = 1024'd93488315027906240658491388568879817320613205836017438648801919162468117663687151162039097575884646163902820472588890703951675809797905765075492669612386550297999106920601487229727943343720665280254420125792176598084123833740296564682588236933584517692564121763106691220709524756898216659818976286558258752743;
            6'd50: xpb[27] = 1024'd113120053493554800463595141230156977453949985340429014721163651909760084705010643479021640352996653640025368764931571208972188517873139399911443966443543771457873266694225977201016506969931708246161069174455500180178708523235940931528250241519629225091753988001105183005024937435967576818587339655393716306683;
            6'd51: xpb[27] = 1024'd8685096275078618869899966486619704842588337719104906665393529592075156409024996885989111915450986806704767649816758279413637385107152700192235138258369951684056751898279249834674831404625545490757520614731583915908932362510688525408933676422444483224123950824986616759233822041108303960237013197603579376292;
            6'd52: xpb[27] = 1024'd28316834740727178675003719147896864975925117223516482737755262339367123450348489202971654692562994282827315942159438784434150093182386335028186435089527172843930911671903739805963395030836588456664169663394907498003517052006332892254595681008489190623313817062985108543549234720177664119005376566439036930232;
            6'd53: xpb[27] = 1024'd47948573206375738480107471809174025109261896727928058810116995086659090491671981519954197469675001758949864234502119289454662801257619969864137731920684394003805071445528229777251958657047631422570818712058231080098101741501977259100257685594533898022503683300983600327864647399247024277773739935274494484172;
            6'd54: xpb[27] = 1024'd67580311672024298285211224470451185242598676232339634882478727833951057532995473836936740246787009235072412526844799794475175509332853604700089028751841615163679231219152719748540522283258674388477467760721554662192686430997621625945919690180578605421693549538982092112180060078316384436542103304109952038112;
            6'd55: xpb[27] = 1024'd87212050137672858090314977131728345375935455736751210954840460581243024574318966153919283023899016711194960819187480299495688217408087239536040325582998836323553390992777209719829085909469717354384116809384878244287271120493265992791581694766623312820883415776980583896495472757385744595310466672945409592052;
            6'd56: xpb[27] = 1024'd106843788603321417895418729793005505509272235241162787027202193328534991615642458470901825801011024187317509111530160804516200925483320874371991622414156057483427550766401699691117649535680760320290765858048201826381855809988910359637243699352668020220073282014979075680810885436455104754078830041780867145992;
            6'd57: xpb[27] = 1024'd2408831384845236301723555049468232897910587619838678971432071010850063319656811877869297363465357353996907996415347874957649792717334174652782794228982237709611035970454972324775973970374597564887217298324285562112079649263657953517927134255483278352443244838860509435019770041595831895728503583990730215601;
            6'd58: xpb[27] = 1024'd22040569850493796106827307710745393031247367124250255043793803758142030360980304194851840140577364830119456288758028379978162500792567809488734091060139458869485195744079462296064537596585640530793866346987609144206664338759302320363589138841527985751633111076859001219335182720665192054496866952826187769541;
            6'd59: xpb[27] = 1024'd41672308316142355911931060372022553164584146628661831116155536505433997402303796511834382917689372306242004581100708884998675208867801444324685387891296680029359355517703952267353101222796683496700515395650932726301249028254946687209251143427572693150822977314857493003650595399734552213265230321661645323481;
            6'd60: xpb[27] = 1024'd61304046781790915717034813033299713297920926133073407188517269252725964443627288828816925694801379782364552873443389390019187916943035079160636684722453901189233515291328442238641664849007726462607164444314256308395833717750591054054913148013617400550012843552855984787966008078803912372033593690497102877421;
            6'd61: xpb[27] = 1024'd80935785247439475522138565694576873431257705637484983260879002000017931484950781145799468471913387258487101165786069895039700625018268713996587981553611122349107675064952932209930228475218769428513813492977579890490418407246235420900575152599662107949202709790854476572281420757873272530801957059332560431361;
            6'd62: xpb[27] = 1024'd100567523713088035327242318355854033564594485141896559333240734747309898526274273462782011249025394734609649458128750400060213333093502348832539278384768343508981834838577422181218792101429812394420462541640903472585003096741879787746237157185706815348392576028852968356596833436942632689570320428168017985301;
            6'd63: xpb[27] = 1024'd120199262178736595132346071017131193697931264646308135405602467494601865567597765779764554026137402210732197750471430905080726041168735983668490575215925564668855994612201912152507355727640855360327111590304227054679587786237524154591899161771751522747582442266851460140912246116011992848338683797003475539241;
        endcase
    end

    always_comb begin
        case(flag[9][11:6])
            6'd0: xpb[28] = 1024'd0;
            6'd1: xpb[28] = 1024'd15764304960260413538650896273593921086569617024984027349832345176916937271612119186732025588591735377411596635356617975522174908402749283949281747030751744895039479816255184786165680162334692604923563030580310790409811625512271748472582596674566780879952405090732893895121130721152719989988357339213338608850;
            6'd2: xpb[28] = 1024'd31528609920520827077301792547187842173139234049968054699664690353833874543224238373464051177183470754823193270713235951044349816805498567898563494061503489790078959632510369572331360324669385209847126061160621580819623251024543496945165193349133561759904810181465787790242261442305439979976714678426677217700;
            6'd3: xpb[28] = 1024'd47292914880781240615952688820781763259708851074952082049497035530750811814836357560196076765775206132234789906069853926566524725208247851847845241092255234685118439448765554358497040487004077814770689091740932371229434876536815245417747790023700342639857215272198681685363392163458159969965072017640015826550;
            6'd4: xpb[28] = 1024'd63057219841041654154603585094375684346278468099936109399329380707667749086448476746928102354366941509646386541426471902088699633610997135797126988123006979580157919265020739144662720649338770419694252122321243161639246502049086993890330386698267123519809620362931575580484522884610879959953429356853354435400;
            6'd5: xpb[28] = 1024'd78821524801302067693254481367969605432848085124920136749161725884584686358060595933660127942958676887057983176783089877610874542013746419746408735153758724475197399081275923930828400811673463024617815152901553952049058127561358742362912983372833904399762025453664469475605653605763599949941786696066693044250;
            6'd6: xpb[28] = 1024'd94585829761562481231905377641563526519417702149904164098994071061501623629672715120392153531550412264469579812139707853133049450416495703695690482184510469370236878897531108716994080974008155629541378183481864742458869753073630490835495580047400685279714430544397363370726784326916319939930144035280031653100;
            6'd7: xpb[28] = 1024'd110350134721822894770556273915157447605987319174888191448826416238418560901284834307124179120142147641881176447496325828655224358819244987644972229215262214265276358713786293503159761136342848234464941214062175532868681378585902239308078176721967466159666835635130257265847915048069039929918501374493370261950;
            6'd8: xpb[28] = 1024'd2047743997958566910408242783936935947858509074136534670526906350358602835587814583841133494076208709849623675395450369598335426380773937039093851229682918226625163960470260951695202107160335118078306636255246476914132153877277214815682203713304797772799337311746093130862517695293126902788168887081114386469;
            6'd9: xpb[28] = 1024'd17812048958218980449059139057530857034428126099120562020359251527275540107199933770573159082667944087261220310752068345120510334783523220988375598260434663121664643776725445737860882269495027723001869666835557267323943779389548963288264800387871578652751742402478987025983648416445846892776526226294452995319;
            6'd10: xpb[28] = 1024'd33576353918479393987710035331124778120997743124104589370191596704192477378812052957305184671259679464672816946108686320642685243186272504937657345291186408016704123592980630524026562431829720327925432697415868057733755404901820711760847397062438359532704147493211880921104779137598566882764883565507791604169;
            6'd11: xpb[28] = 1024'd49340658878739807526360931604718699207567360149088616720023941881109414650424172144037210259851414842084413581465304296164860151589021788886939092321938152911743603409235815310192242594164412932848995727996178848143567030414092460233429993737005140412656552583944774816225909858751286872753240904721130213019;
            6'd12: xpb[28] = 1024'd65104963839000221065011827878312620294136977174072644069856287058026351922036291330769235848443150219496010216821922271687035059991771072836220839352689897806783083225491000096357922756499105537772558758576489638553378655926364208706012590411571921292608957674677668711347040579904006862741598243934468821869;
            6'd13: xpb[28] = 1024'd80869268799260634603662724151906541380706594199056671419688632234943289193648410517501261437034885596907606852178540247209209968394520356785502586383441642701822563041746184882523602918833798142696121789156800428963190281438635957178595187086138702172561362765410562606468171301056726852729955583147807430719;
            6'd14: xpb[28] = 1024'd96633573759521048142313620425500462467276211224040698769520977411860226465260529704233287025626620974319203487535158222731384876797269640734784333414193387596862042858001369668689283081168490747619684819737111219373001906950907705651177783760705483052513767856143456501589302022209446842718312922361146039569;
            6'd15: xpb[28] = 1024'd112397878719781461680964516699094383553845828249024726119353322588777163736872648890965312614218356351730800122891776198253559785200018924684066080444945132491901522674256554454854963243503183352543247850317422009782813532463179454123760380435272263932466172946876350396710432743362166832706670261574484648419;
            6'd16: xpb[28] = 1024'd4095487995917133820816485567873871895717018148273069341053812700717205671175629167682266988152417419699247350790900739196670852761547874078187702459365836453250327920940521903390404214320670236156613272510492953828264307754554429631364407426609595545598674623492186261725035390586253805576337774162228772938;
            6'd17: xpb[28] = 1024'd19859792956177547359467381841467792982286635173257096690886157877634142942787748354414292576744152797110843986147518714718845761164297158027469449490117581348289807737195706689556084376655362841080176303090803744238075933266826178103947004101176376425551079714225080156846166111738973795564695113375567381788;
            6'd18: xpb[28] = 1024'd35624097916437960898118278115061714068856252198241124040718503054551080214399867541146318165335888174522440621504136690241020669567046441976751196520869326243329287553450891475721764538990055446003739333671114534647887558779097926576529600775743157305503484804957974051967296832891693785553052452588905990638;
            6'd19: xpb[28] = 1024'd51388402876698374436769174388655635155425869223225151390550848231468017486011986727878343753927623551934037256860754665763195577969795725926032943551621071138368767369706076261887444701324748050927302364251425325057699184291369675049112197450309938185455889895690867947088427554044413775541409791802244599488;
            6'd20: xpb[28] = 1024'd67152707836958787975420070662249556241995486248209178740383193408384954757624105914610369342519358929345633892217372641285370486372545009875314690582372816033408247185961261048053124863659440655850865394831736115467510809803641423521694794124876719065408294986423761842209558275197133765529767131015583208338;
            6'd21: xpb[28] = 1024'd82917012797219201514070966935843477328565103273193206090215538585301892029236225101342394931111094306757230527573990616807545394775294293824596437613124560928447727002216445834218805025994133260774428425412046905877322435315913171994277390799443499945360700077156655737330688996349853755518124470228921817188;
            6'd22: xpb[28] = 1024'd98681317757479615052721863209437398415134720298177233440047883762218829300848344288074420519702829684168827162930608592329720303178043577773878184643876305823487206818471630620384485188328825865697991455992357696287134060828184920466859987474010280825313105167889549632451819717502573745506481809442260426038;
            6'd23: xpb[28] = 1024'd114445622717740028591372759483031319501704337323161260789880228939135766572460463474806446108294565061580423798287226567851895211580792861723159931674628050718526686634726815406550165350663518470621554486572668486696945686340456668939442584148577061705265510258622443527572950438655293735494839148655599034888;
            6'd24: xpb[28] = 1024'd6143231993875700731224728351810807843575527222409604011580719051075808506763443751523400482228626129548871026186351108795006279142321811117281553689048754679875491881410782855085606321481005354234919908765739430742396461631831644447046611139914393318398011935238279392587553085879380708364506661243343159407;
            6'd25: xpb[28] = 1024'd21907536954136114269875624625404728930145144247393631361413064227992745778375562938255426070820361506960467661542969084317181187545071095066563300719800499574914971697665967641251286483815697959158482939346050221152208087144103392919629207814481174198350417025971173287708683807032100698352864000456681768257;
            6'd26: xpb[28] = 1024'd37671841914396527808526520898998650016714761272377658711245409404909683049987682124987451659412096884372064296899587059839356095947820379015845047750552244469954451513921152427416966646150390564082045969926361011562019712656375141392211804489047955078302822116704067182829814528184820688341221339670020377107;
            6'd27: xpb[28] = 1024'd53436146874656941347177417172592571103284378297361686061077754581826620321599801311719477248003832261783660932256205035361531004350569662965126794781303989364993931330176337213582646808485083169005609000506671801971831338168646889864794401163614735958255227207436961077950945249337540678329578678883358985957;
            6'd28: xpb[28] = 1024'd69200451834917354885828313446186492189853995322345713410910099758743557593211920498451502836595567639195257567612823010883705912753318946914408541812055734260033411146431521999748326970819775773929172031086982592381642963680918638337376997838181516838207632298169854973072075970490260668317936018096697594807;
            6'd29: xpb[28] = 1024'd84964756795177768424479209719780413276423612347329740760742444935660494864824039685183528425187303016606854202969440986405880821156068230863690288842807479155072890962686706785914007133154468378852735061667293382791454589193190386809959594512748297718160037388902748868193206691642980658306293357310036203657;
            6'd30: xpb[28] = 1024'd100729061755438181963130105993374334362993229372313768110574790112577432136436158871915554013779038394018450838326058961928055729558817514812972035873559224050112370778941891572079687295489160983776298092247604173201266214705462135282542191187315078598112442479635642763314337412795700648294650696523374812507;
            6'd31: xpb[28] = 1024'd116493366715698595501781002266968255449562846397297795460407135289494369408048278058647579602370773771430047473682676937450230637961566798762253782904310968945151850595197076358245367457823853588699861122827914963611077840217733883755124787861881859478064847570368536658435468133948420638283008035736713421357;
            6'd32: xpb[28] = 1024'd8190975991834267641632971135747743791434036296546138682107625401434411342351258335364533976304834839398494701581801478393341705523095748156375404918731672906500655841881043806780808428641340472313226545020985907656528615509108859262728814853219191091197349246984372523450070781172507611152675548324457545876;
            6'd33: xpb[28] = 1024'd23955280952094681180283867409341664878003653321530166031939970578351348613963377522096559564896570216810091336938419453915516613925845032105657151949483417801540135658136228592946488590976033077236789575601296698066340241021380607735311411527785971971149754337717266418571201502325227601141032887537796154726;
            6'd34: xpb[28] = 1024'd39719585912355094718934763682935585964573270346514193381772315755268285885575496708828585153488305594221687972295037429437691522328594316054938898980235162696579615474391413379112168753310725682160352606181607488476151866533652356207894008202352752851102159428450160313692332223477947591129390226751134763576;
            6'd35: xpb[28] = 1024'd55483890872615508257585659956529507051142887371498220731604660932185223157187615895560610742080040971633284607651655404959866430731343600004220646010986907591619095290646598165277848915645418287083915636761918278885963492045924104680476604876919533731054564519183054208813462944630667581117747565964473372426;
            6'd36: xpb[28] = 1024'd71248195832875921796236556230123428137712504396482248081437006109102160428799735082292636330671776349044881243008273380482041339134092883953502393041738652486658575106901782951443529077980110892007478667342229069295775117558195853153059201551486314611006969609915948103934593665783387571106104905177811981276;
            6'd37: xpb[28] = 1024'd87012500793136335334887452503717349224282121421466275431269351286019097700411854269024661919263511726456477878364891356004216247536842167902784140072490397381698054923156967737609209240314803496931041697922539859705586743070467601625641798226053095490959374700648841999055724386936107561094462244391150590126;
            6'd38: xpb[28] = 1024'd102776805753396748873538348777311270310851738446450302781101696462936034972023973455756687507855247103868074513721509331526391155939591451852065887103242142276737534739412152523774889402649496101854604728502850650115398368582739350098224394900619876370911779791381735894176855108088827551082819583604489198976;
            6'd39: xpb[28] = 1024'd118541110713657162412189245050905191397421355471434330130934041639852972243636092642488713096446982481279671149078127307048566064342340735801347634133993887171777014555667337309940569564984188706778167759083161440525209994095011098570806991575186657250864184882114629789297985829241547541071176922817827807826;
            6'd40: xpb[28] = 1024'd10238719989792834552041213919684679739292545370682673352634531751793014177939072919205667470381043549248118376977251847991677131903869685195469256148414591133125819802351304758476010535801675590391533181276232384570660769386386074078411018566523988863996686558730465654312588476465634513940844435405571932345;
            6'd41: xpb[28] = 1024'd26003024950053248090692110193278600825862162395666700702466876928709951449551192105937693058972778926659715012333869823513852040306618969144751003179166336028165299618606489544641690698136368195315096211856543174980472394898657822550993615241090769743949091649463359549433719197618354503929201774618910541195;
            6'd42: xpb[28] = 1024'd41767329910313661629343006466872521912431779420650728052299222105626888721163311292669718647564514304071311647690487799036026948709368253094032750209918080923204779434861674330807370860471060800238659242436853965390284020410929571023576211915657550623901496740196253444554849918771074493917559113832249150045;
            6'd43: xpb[28] = 1024'd57531634870574075167993902740466442999001396445634755402131567282543825992775430479401744236156249681482908283047105774558201857112117537043314497240669825818244259251116859116973051022805753405162222273017164755800095645923201319496158808590224331503853901830929147339675980639923794483905916453045587758895;
            6'd44: xpb[28] = 1024'd73295939830834488706644799014060364085571013470618782751963912459460763264387549666133769824747985058894504918403723750080376765514866820992596244271421570713283739067372043903138731185140446010085785303597475546209907271435473067968741405264791112383806306921662041234797111361076514473894273792258926367745;
            6'd45: xpb[28] = 1024'd89060244791094902245295695287654285172140630495602810101796257636377700535999668852865795413339720436306101553760341725602551673917616104941877991302173315608323218883627228689304411347475138615009348334177786336619718896947744816441324001939357893263758712012394935129918242082229234463882631131472264976595;
            6'd46: xpb[28] = 1024'd104824549751355315783946591561248206258710247520586837451628602813294637807611788039597821001931455813717698189116959701124726582320365388891159738332925060503362698699882413475470091509809831219932911364758097127029530522460016564913906598613924674143711117103127829025039372803381954453870988470685603585445;
            6'd47: xpb[28] = 1024'd120588854711615729322597487834842127345279864545570864801460947990211575079223907226329846590523191191129294824473577676646901490723114672840441485363676805398402178516137598261635771672144523824856474395338407917439342147972288313386489195288491455023663522193860722920160503524534674443859345809898942194295;
            6'd48: xpb[28] = 1024'd12286463987751401462449456703621615687151054444819208023161438102151617013526887503046800964457252259097742052372702217590012558284643622234563107378097509359750983762821565710171212642962010708469839817531478861484792923263663288894093222279828786636796023870476558785175106171758761416729013322486686318814;
            6'd49: xpb[28] = 1024'd28050768948011815001100352977215536773720671469803235372993783279068554285139006689778826553048987636509338687729320193112187466687392906183844854408849254254790463579076750496336892805296703313393402848111789651894604548775935037366675818954395567516748428961209452680296236892911481406717370661700024927664;
            6'd50: xpb[28] = 1024'd43815073908272228539751249250809457860290288494787262722826128455985491556751125876510852141640723013920935323085938168634362375090142190133126601439600999149829943395331935282502572967631395918316965878692100442304416174288206785839258415628962348396700834051942346575417367614064201396705728000913363536514;
            6'd51: xpb[28] = 1024'd59579378868532642078402145524403378946859905519771290072658473632902428828363245063242877730232458391332531958442556144156537283492891474082408348470352744044869423211587120068668253129966088523240528909272411232714227799800478534311841012303529129276653239142675240470538498335216921386694085340126702145364;
            6'd52: xpb[28] = 1024'd75343683828793055617053041797997300033429522544755317422490818809819366099975364249974903318824193768744128593799174119678712191895640758031690095501104488939908903027842304854833933292300781128164091939852722023124039425312750282784423608978095910156605644233408134365659629056369641376682442679340040754214;
            6'd53: xpb[28] = 1024'd91107988789053469155703938071591221119999139569739344772323163986736303371587483436706928907415929146155725229155792095200887100298390041980971842531856233834948382844097489640999613454635473733087654970433032813533851050825022031257006205652662691036558049324141028260780759777522361366670800018553379363064;
            6'd54: xpb[28] = 1024'd106872293749313882694354834345185142206568756594723372122155509163653240643199602623438954496007664523567321864512410070723062008701139325930253589562607978729987862660352674427165293616970166338011218001013343603943662676337293779729588802327229471916510454414873922155901890498675081356659157357766717971914;
            6'd55: xpb[28] = 1024'd122636598709574296233005730618779063293138373619707399471987854340570177914811721810170980084599399900978918499869028046245236917103888609879535336593359723625027342476607859213330973779304858942934781031593654394353474301849565528202171399001796252796462859505606816051023021219827801346647514696980056580764;
            6'd56: xpb[28] = 1024'd14334207985709968372857699487558551635009563518955742693688344452510219849114702086887934458533460968947365727768152587188347984665417559273656958607780427586376147723291826661866414750122345826548146453786725338398925077140940503709775425993133584409595361182222651916037623867051888319517182209567800705283;
            6'd57: xpb[28] = 1024'd30098512945970381911508595761152472721579180543939770043520689629427157120726821273619960047125196346358962363124770562710522893068166843222938705638532172481415627539547011448032094912457038431471709484367036128808736702653212252182358022667700365289547766272955545811158754588204608309505539548781139314133;
            6'd58: xpb[28] = 1024'd45862817906230795450159492034746393808148797568923797393353034806344094392338940460351985635716931723770558998481388538232697801470916127172220452669283917376455107355802196234197775074791731036395272514947346919218548328165484000654940619342267146169500171363688439706279885309357328299493896887994477922983;
            6'd59: xpb[28] = 1024'd61627122866491208988810388308340314894718414593907824743185379983261031663951059647084011224308667101182155633838006513754872709873665411121502199700035662271494587172057381020363455237126423641318835545527657709628359953677755749127523216016833927049452576454421333601401016030510048289482254227207816531833;
            6'd60: xpb[28] = 1024'd77391427826751622527461284581934235981288031618891852093017725160177968935563178833816036812900402478593752269194624489277047618276414695070783946730787407166534066988312565806529135399461116246242398576107968500038171579190027497600105812691400707929404981545154227496522146751662768279470611566421155140683;
            6'd61: xpb[28] = 1024'd93155732787012036066112180855528157067857648643875879442850070337094906207175298020548062401492137856005348904551242464799222526679163979020065693761539152061573546804567750592694815561795808851165961606688279290447983204702299246072688409365967488809357386635887121391643277472815488269458968905634493749533;
            6'd62: xpb[28] = 1024'd108920037747272449604763077129122078154427265668859906792682415514011843478787417207280087990083873233416945539907860440321397435081913262969347440792290896956613026620822935378860495724130501456089524637268590080857794830214570994545271006040534269689309791726620015286764408193968208259447326244847832358383;
            6'd63: xpb[28] = 1024'd617647023408121744615045997901566496298455568108250014382905625951885413090397483997042364017934301385392767806984981264508502643442212363469062806711600917961831867506902827395936694947988339702890059461661024903245605505945970052875033031871601302442293403235851151779010841192295232316993757435576482902;
        endcase
    end

    always_comb begin
        case(flag[9][16:12])
            5'd0: xpb[29] = 1024'd0;
            5'd1: xpb[29] = 1024'd16381951983668535283265942271495487582868072593092277364215250802868822684702516670729067952609669678796989403163602956786683411046191496312750809837463345813001311683762087613561616857282680944626453090041971815313057231018217718525457629706438382182394698493968745046900141562345015222305351096648915091752;
            5'd2: xpb[29] = 1024'd32763903967337070566531884542990975165736145186184554728430501605737645369405033341458135905219339357593978806327205913573366822092382992625501619674926691626002623367524175227123233714565361889252906180083943630626114462036435437050915259412876764364789396987937490093800283124690030444610702193297830183504;
            5'd3: xpb[29] = 1024'd49145855951005605849797826814486462748604217779276832092645752408606468054107550012187203857829009036390968209490808870360050233138574488938252429512390037439003935051286262840684850571848042833879359270125915445939171693054653155576372889119315146547184095481906235140700424687035045666916053289946745275256;
            5'd4: xpb[29] = 1024'd65527807934674141133063769085981950331472290372369109456861003211475290738810066682916271810438678715187957612654411827146733644184765985251003239349853383252005246735048350454246467429130723778505812360167887261252228924072870874101830518825753528729578793975874980187600566249380060889221404386595660367008;
            5'd5: xpb[29] = 1024'd81909759918342676416329711357477437914340362965461386821076254014344113423512583353645339763048348393984947015818014783933417055230957481563754049187316729065006558418810438067808084286413404723132265450209859076565286155091088592627288148532191910911973492469843725234500707811725076111526755483244575458760;
            5'd6: xpb[29] = 1024'd98291711902011211699595653628972925497208435558553664185291504817212936108215100024374407715658018072781936418981617740720100466277148977876504859024780074878007870102572525681369701143696085667758718540251830891878343386109306311152745778238630293094368190963812470281400849374070091333832106579893490550512;
            5'd7: xpb[29] = 1024'd114673663885679746982861595900468413080076508151645941549506755620081758792917616695103475668267687751578925822145220697506783877323340474189255668862243420691009181786334613294931318000978766612385171630293802707191400617127524029678203407945068675276762889457781215328300990936415106556137457676542405642264;
            5'd8: xpb[29] = 1024'd6988920185223540867328610767149467918246153619002534785590151357973686140310994455817472406219683120932765817851330219714403447528311635946846353683375725570319818900525483570862695666744241835701427111948534676140096997924844975238682467968277608192337684537632902345094604424831488761324118946565726249685;
            5'd9: xpb[29] = 1024'd23370872168892076150594553038644955501114226212094812149805402160842508825013511126546540358829352799729755221014933176501086858574503132259597163520839071383321130584287571184424312524026922780327880201990506491453154228943062693764140097674715990374732383031601647391994745987176503983629470043214641341437;
            5'd10: xpb[29] = 1024'd39752824152560611433860495310140443083982298805187089514020652963711331509716027797275608311439022478526744624178536133287770269620694628572347973358302417196322442268049658797985929381309603724954333292032478306766211459961280412289597727381154372557127081525570392438894887549521519205934821139863556433189;
            5'd11: xpb[29] = 1024'd56134776136229146717126437581635930666850371398279366878235903766580154194418544468004676264048692157323734027342139090074453680666886124885098783195765763009323753951811746411547546238592284669580786382074450122079268690979498130815055357087592754739521780019539137485795029111866534428240172236512471524941;
            5'd12: xpb[29] = 1024'd72516728119897682000392379853131418249718443991371644242451154569448976879121061138733744216658361836120723430505742046861137091713077621197849593033229108822325065635573834025109163095874965614207239472116421937392325921997715849340512986794031136921916478513507882532695170674211549650545523333161386616693;
            5'd13: xpb[29] = 1024'd88898680103566217283658322124626905832586516584463921606666405372317799563823577809462812169268031514917712833669345003647820502759269117510600402870692454635326377319335921638670779953157646558833692562158393752705383153015933567865970616500469519104311177007476627579595312236556564872850874429810301708445;
            5'd14: xpb[29] = 1024'd105280632087234752566924264396122393415454589177556198970881656175186622248526094480191880121877701193714702236832947960434503913805460613823351212708155800448327689003098009252232396810440327503460145652200365568018440384034151286391428246206907901286705875501445372626495453798901580095156225526459216800197;
            5'd15: xpb[29] = 1024'd121662584070903287850190206667617880998322661770648476335096906978055444933228611150920948074487370872511691639996550917221187324851652110136102022545619146261329000686860096865794013667723008448086598742242337383331497615052369004916885875913346283469100573995414117673395595361246595317461576623108131891949;
            5'd16: xpb[29] = 1024'd13977840370447081734657221534298935836492307238005069571180302715947372280621988911634944812439366241865531635702660439428806895056623271893692707366751451140639637801050967141725391333488483671402854223897069352280193995849689950477364935936555216384675369075265804690189208849662977522648237893131452499370;
            5'd17: xpb[29] = 1024'd30359792354115617017923163805794423419360379831097346935395553518816194965324505582364012765049035920662521038866263396215490306102814768206443517204214796953640949484813054755287008190771164616029307313939041167593251226867907669002822565642993598567070067569234549737089350412007992744953588989780367591122;
            5'd18: xpb[29] = 1024'd46741744337784152301189106077289911002228452424189624299610804321685017650027022253093080717658705599459510442029866353002173717149006264519194327041678142766642261168575142368848625048053845560655760403981012982906308457886125387528280195349431980749464766063203294783989491974353007967258940086429282682874;
            5'd19: xpb[29] = 1024'd63123696321452687584455048348785398585096525017281901663826055124553840334729538923822148670268375278256499845193469309788857128195197760831945136879141488579643572852337229982410241905336526505282213494022984798219365688904343106053737825055870362931859464557172039830889633536698023189564291183078197774626;
            5'd20: xpb[29] = 1024'd79505648305121222867720990620280886167964597610374179028041305927422663019432055594551216622878044957053489248357072266575540539241389257144695946716604834392644884536099317595971858762619207449908666584064956613532422919922560824579195454762308745114254163051140784877789775099043038411869642279727112866378;
            5'd21: xpb[29] = 1024'd95887600288789758150986932891776373750832670203466456392256556730291485704134572265280284575487714635850478651520675223362223950287580753457446756554068180205646196219861405209533475619901888394535119674106928428845480150940778543104653084468747127296648861545109529924689916661388053634174993376376027958130;
            5'd22: xpb[29] = 1024'd112269552272458293434252875163271861333700742796558733756471807533160308388837088936009352528097384314647468054684278180148907361333772249770197566391531526018647507903623492823095092477184569339161572764148900244158537381958996261630110714175185509479043560039078274971590058223733068856480344473024943049882;
            5'd23: xpb[29] = 1024'd4584808572002087318719890029952916171870388263915326992555203271052235736230466696723349266049379684001308050390387702356526931538743411527788251212663830897958145017814363099026470142950044562477828245803632213107233762756317207190589774198394442394618355118929961988383671712149451061667005743048263657303;
            5'd24: xpb[29] = 1024'd20966760555670622601985832301448403754738460857007604356770454073921058420932983367452417218659049362798297453553990659143210342584934907840539061050127176710959456701576450712588087000232725507104281335845604028420290993774534925716047403904832824577013053612898707035283813274494466283972356839697178749055;
            5'd25: xpb[29] = 1024'd37348712539339157885251774572943891337606533450099881720985704876789881105635500038181485171268719041595286856717593615929893753631126404153289870887590522523960768385338538326149703857515406451730734425887575843733348224792752644241505033611271206759407752106867452082183954836839481506277707936346093840807;
            5'd26: xpb[29] = 1024'd53730664523007693168517716844439378920474606043192159085200955679658703790338016708910553123878388720392276259881196572716577164677317900466040680725053868336962080069100625939711320714798087396357187515929547659046405455810970362766962663317709588941802450600836197129084096399184496728583059032995008932559;
            5'd27: xpb[29] = 1024'd70112616506676228451783659115934866503342678636284436449416206482527526475040533379639621076488058399189265663044799529503260575723509396778791490562517214149963391752862713553272937572080768340983640605971519474359462686829188081292420293024147971124197149094804942175984237961529511950888410129643924024311;
            5'd28: xpb[29] = 1024'd86494568490344763735049601387430354086210751229376713813631457285396349159743050050368689029097728077986255066208402486289943986769700893091542300399980559962964703436624801166834554429363449285610093696013491289672519917847405799817877922730586353306591847588773687222884379523874527173193761226292839116063;
            5'd29: xpb[29] = 1024'd102876520474013299018315543658925841669078823822468991177846708088265171844445566721097756981707397756783244469372005443076627397815892389404293110237443905775966015120386888780396171286646130230236546786055463104985577148865623518343335552437024735488986546082742432269784521086219542395499112322941754207815;
            5'd30: xpb[29] = 1024'd119258472457681834301581485930421329251946896415561268542061958891133994529148083391826824934317067435580233872535608399863310808862083885717043920074907251588967326804148976393957788143928811174862999876097434920298634379883841236868793182143463117671381244576711177316684662648564557617804463419590669299567;
            5'd31: xpb[29] = 1024'd11573728757225628186048500797102384090116541882917861778145354629025921876541461152540821672269062804934073868241717922070930379067055047474634604896039556468277963918339846669889165809694286398179255357752166889247330760681162182429272242166672050586956039656562864333478276136980939822991124689613989906988;
        endcase
    end

    always_comb begin
        case(flag[10][5:0])
            6'd0: xpb[30] = 1024'd0;
            6'd1: xpb[30] = 1024'd13977840370447081734657221534298935836492307238005069571180302715947372280621988911634944812439366241865531635702660439428806895056623271893692707366751451140639637801050967141725391333488483671402854223897069352280193995849689950477364935936555216384675369075265804690189208849662977522648237893131452499370;
            6'd2: xpb[30] = 1024'd27955680740894163469314443068597871672984614476010139142360605431894744561243977823269889624878732483731063271405320878857613790113246543787385414733502902281279275602101934283450782666976967342805708447794138704560387991699379900954729871873110432769350738150531609380378417699325955045296475786262904998740;
            6'd3: xpb[30] = 1024'd41933521111341245203971664602896807509476921714015208713540908147842116841865966734904834437318098725596594907107981318286420685169869815681078122100254353421918913403152901425176174000465451014208562671691208056840581987549069851432094807809665649154026107225797414070567626548988932567944713679394357498110;
            6'd4: xpb[30] = 1024'd55911361481788326938628886137195743345969228952020278284721210863789489122487955646539779249757464967462126542810641757715227580226493087574770829467005804562558551204203868566901565333953934685611416895588277409120775983398759801909459743746220865538701476301063218760756835398651910090592951572525809997480;
            6'd5: xpb[30] = 1024'd69889201852235408673286107671494679182461536190025347855901513579736861403109944558174724062196831209327658178513302197144034475283116359468463536833757255703198189005254835708626956667442418357014271119485346761400969979248449752386824679682776081923376845376329023450946044248314887613241189465657262496850;
            6'd6: xpb[30] = 1024'd83867042222682490407943329205793615018953843428030417427081816295684233683731933469809668874636197451193189814215962636572841370339739631362156244200508706843837826806305802850352348000930902028417125343382416113681163975098139702864189615619331298308052214451594828141135253097977865135889427358788714996220;
            6'd7: xpb[30] = 1024'd97844882593129572142600550740092550855446150666035486998262119011631605964353922381444613687075563693058721449918623076001648265396362903255848951567260157984477464607356769992077739334419385699819979567279485465961357970947829653341554551555886514692727583526860632831324461947640842658537665251920167495590;
            6'd8: xpb[30] = 1024'd111822722963576653877257772274391486691938457904040556569442421727578978244975911293079558499514929934924253085621283515430455160452986175149541658934011609125117102408407737133803130667907869371222833791176554818241551966797519603818919487492441731077402952602126437521513670797303820181185903145051619994960;
            6'd9: xpb[30] = 1024'd1733867649898994213116066403875989783732338016309942012490869378549455188288761294699432097296621867346635313866450520280198214668389112488074241284432019332066065639887486937898282809879147321315490406686384324157385112426312781331305853745767498195258418263275184181596351573038164686715451211557478009999;
            6'd10: xpb[30] = 1024'd15711708020346075947773287938174925620224645254315011583671172094496827468910750206334376909735988109212166949569110959709005109725012384381766948651183470472705703440938454079623674143367630992718344630583453676437579108276002731808670789682322714579933787338540988871785560422701142209363689104688930509369;
            6'd11: xpb[30] = 1024'd29689548390793157682430509472473861456716952492320081154851474810444199749532739117969321722175354351077698585271771399137812004781635656275459656017934921613345341241989421221349065476856114664121198854480523028717773104125692682286035725618877930964609156413806793561974769272364119732011926997820383008739;
            6'd12: xpb[30] = 1024'd43667388761240239417087731006772797293209259730325150726031777526391572030154728029604266534614720592943230220974431838566618899838258928169152363384686372753984979043040388363074456810344598335524053078377592380997967099975382632763400661555433147349284525489072598252163978122027097254660164890951835508109;
            6'd13: xpb[30] = 1024'd57645229131687321151744952541071733129701566968330220297212080242338944310776716941239211347054086834808761856677092277995425794894882200062845070751437823894624616844091355504799848143833082006926907302274661733278161095825072583240765597491988363733959894564338402942353186971690074777308402784083288007479;
            6'd14: xpb[30] = 1024'd71623069502134402886402174075370668966193874206335289868392382958286316591398705852874156159493453076674293492379752717424232689951505471956537778118189275035264254645142322646525239477321565678329761526171731085558355091674762533718130533428543580118635263639604207632542395821353052299956640677214740506849;
            6'd15: xpb[30] = 1024'd85600909872581484621059395609669604802686181444340359439572685674233688872020694764509100971932819318539825128082413156853039585008128743850230485484940726175903892446193289788250630810810049349732615750068800437838549087524452484195495469365098796503310632714870012322731604671016029822604878570346193006219;
            6'd16: xpb[30] = 1024'd99578750243028566355716617143968540639178488682345429010752988390181061152642683676144045784372185560405356763785073596281846480064752015743923192851692177316543530247244256929976022144298533021135469973965869790118743083374142434672860405301654012887986001790135817012920813520679007345253116463477645505589;
            6'd17: xpb[30] = 1024'd113556590613475648090373838678267476475670795920350498581933291106128433433264672587778990596811551802270888399487734035710653375121375287637615900218443628457183168048295224071701413477787016692538324197862939142398937079223832385150225341238209229272661370865401621703110022370341984867901354356609098004959;
            6'd18: xpb[30] = 1024'd3467735299797988426232132807751979567464676032619884024981738757098910376577522589398864194593243734693270627732901040560396429336778224976148482568864038664132131279774973875796565619758294642630980813372768648314770224852625562662611707491534996390516836526550368363192703146076329373430902423114956019998;
            6'd19: xpb[30] = 1024'd17445575670245070160889354342050915403956983270624953596162041473046282657199511501033809007032609976558802263435561479989203324393401496869841189935615489804771769080825941017521956953246778314033835037269838000594964220702315513139976643428090212775192205601816173053381911995739306896079140316246408519368;
            6'd20: xpb[30] = 1024'd31423416040692151895546575876349851240449290508630023167342344188993654937821500412668753819471976218424333899138221919418010219450024768763533897302366940945411406881876908159247348286735261985436689261166907352875158216552005463617341579364645429159867574677081977743571120845402284418727378209377861018738;
            6'd21: xpb[30] = 1024'd45401256411139233630203797410648787076941597746635092738522646904941027218443489324303698631911342460289865534840882358846817114506648040657226604669118392086051044682927875300972739620223745656839543485063976705155352212401695414094706515301200645544542943752347782433760329695065261941375616102509313518108;
            6'd22: xpb[30] = 1024'd59379096781586315364861018944947722913433904984640162309702949620888399499065478235938643444350708702155397170543542798275624009563271312550919312035869843226690682483978842442698130953712229328242397708961046057435546208251385364572071451237755861929218312827613587123949538544728239464023853995640766017478;
            6'd23: xpb[30] = 1024'd73356937152033397099518240479246658749926212222645231880883252336835771779687467147573588256790074944020928806246203237704430904619894584444612019402621294367330320285029809584423522287200712999645251932858115409715740204101075315049436387174311078313893681902879391814138747394391216986672091888772218516848;
            6'd24: xpb[30] = 1024'd87334777522480478834175462013545594586418519460650301452063555052783144060309456059208533069229441185886460441948863677133237799676517856338304726769372745507969958086080776726148913620689196671048106156755184761995934199950765265526801323110866294698569050978145196504327956244054194509320329781903671016218;
            6'd25: xpb[30] = 1024'd101312617892927560568832683547844530422910826698655371023243857768730516340931444970843477881668807427751992077651524116562044694733141128231997434136124196648609595887131743867874304954177680342450960380652254114276128195800455216004166259047421511083244420053411001194517165093717172031968567675035123515588;
            6'd26: xpb[30] = 1024'd115290458263374642303489905082143466259403133936660440594424160484677888621553433882478422694108173669617523713354184555990851589789764400125690141502875647789249233688182711009599696287666164013853814604549323466556322191650145166481531194983976727467919789128676805884706373943380149554616805568166576014958;
            6'd27: xpb[30] = 1024'd5201602949696982639348199211627969351197014048929826037472608135648365564866283884098296291889865602039905941599351560840594644005167337464222723853296057996198196919662460813694848429637441963946471220059152972472155337278938343993917561237302494585775254789825552544789054719114494060146353634672434029997;
            6'd28: xpb[30] = 1024'd19179443320144064374005420745926905187689321286934895608652910851595737845488272795733241104329231843905437577302012000269401539061790609357915431220047509136837834720713427955420239763125925635349325443956222324752349333128628294471282497173857710970450623865091357234978263568777471582794591527803886529367;
            6'd29: xpb[30] = 1024'd33157283690591146108662642280225841024181628524939965179833213567543110126110261707368185916768598085770969213004672439698208434118413881251608138586798960277477472521764395097145631096614409306752179667853291677032543328978318244948647433110412927355125992940357161925167472418440449105442829420935339028737;
            6'd30: xpb[30] = 1024'd47135124061038227843319863814524776860673935762945034751013516283490482406732250619003130729207964327636500848707332879127015329175037153145300845953550411418117110322815362238871022430102892978155033891750361029312737324828008195426012369046968143739801362015622966615356681268103426628091067314066791528107;
            6'd31: xpb[30] = 1024'd61112964431485309577977085348823712697166243000950104322193818999437854687354239530638075541647330569502032484409993318555822224231660425038993553320301862558756748123866329380596413763591376649557888115647430381592931320677698145903377304983523360124476731090888771305545890117766404150739305207198244027477;
            6'd32: xpb[30] = 1024'd75090804801932391312634306883122648533658550238955173893374121715385226967976228442273020354086696811367564120112653757984629119288283696932686260687053313699396385924917296522321805097079860320960742339544499733873125316527388096380742240920078576509152100166154575995735098967429381673387543100329696526847;
            6'd33: xpb[30] = 1024'd89068645172379473047291528417421584370150857476960243464554424431332599248598217353907965166526063053233095755815314197413436014344906968826378968053804764840036023725968263664047196430568343992363596563441569086153319312377078046858107176856633792893827469241420380685924307817092359196035780993461149026217;
            6'd34: xpb[30] = 1024'd103046485542826554781948749951720520206643164714965313035734727147279971529220206265542909978965429295098627391517974636842242909401530240720071675420556215980675661527019230805772587764056827663766450787338638438433513308226767997335472112793189009278502838316686185376113516666755336718684018886592601525587;
            6'd35: xpb[30] = 1024'd117024325913273636516605971486019456043135471952970382606915029863227343809842195177177854791404795536964159027220635076271049804458153512613764382787307667121315299328070197947497979097545311335169305011235707790713707304076457947812837048729744225663178207391951990066302725516418314241332256779724054024957;
            6'd36: xpb[30] = 1024'd6935470599595976852464265615503959134929352065239768049963477514197820753155045178797728389186487469386541255465802081120792858673556449952296965137728077328264262559549947751593131239516589285261961626745537296629540449705251125325223414983069992781033673053100736726385406292152658746861804846229912039996;
            6'd37: xpb[30] = 1024'd20913310970043058587121487149802894971421659303244837621143780230145193033777034090432673201625853711252072891168462520549599753730179721845989672504479528468903900360600914893318522573005072956664815850642606648909734445554941075802588350919625209165709042128366541416574615141815636269510042739361364539366;
            6'd38: xpb[30] = 1024'd34891151340490140321778708684101830807913966541249907192324082946092565314399023002067618014065219953117604526871122959978406648786802993739682379871230979609543538161651882035043913906493556628067670074539676001189928441404631026279953286856180425550384411203632346106763823991478613792158280632492817038736;
            6'd39: xpb[30] = 1024'd48868991710937222056435930218400766644406273779254976763504385662039937595021011913702562826504586194983136162573783399407213543843426265633375087237982430750183175962702849176769305239982040299470524298436745353470122437254320976757318222792735641935059780278898150796953032841141591314806518525624269538106;
            6'd40: xpb[30] = 1024'd62846832081384303791093151752699702480898581017260046334684688377987309875643000825337507638943952436848667798276443838836020438900049537527067794604733881890822813763753816318494696573470523970873378522333814705750316433104010927234683158729290858319735149354163955487142241690804568837454756418755722037476;
            6'd41: xpb[30] = 1024'd76824672451831385525750373286998638317390888255265115905864991093934682156264989736972452451383318678714199433979104278264827333956672809420760501971485333031462451564804783460220087906959007642276232746230884058030510428953700877712048094665846074704410518429429760177331450540467546360102994311887174536846;
            6'd42: xpb[30] = 1024'd90802512822278467260407594821297574153883195493270185477045293809882054436886978648607397263822684920579731069681764717693634229013296081314453209338236784172102089365855750601945479240447491313679086970127953410310704424803390828189413030602401291089085887504695564867520659390130523882751232205018627036216;
            6'd43: xpb[30] = 1024'd104780353192725548995064816355596509990375502731275255048225596525829426717508967560242342076262051162445262705384425157122441124069919353208145916704988235312741727166906717743670870573935974985081941194025022762590898420653080778666777966538956507473761256579961369557709868239793501405399470098150079535586;
            6'd44: xpb[30] = 1024'd118758193563172630729722037889895445826867809969280324619405899241776798998130956471877286888701417404310794341087085596551248019126542625101838624071739686453381364967957684885396261907424458656484795417922092114871092416502770729144142902475511723858436625655227174247899077089456478928047707991281532034956;
            6'd45: xpb[30] = 1024'd8669338249494971065580332019379948918661690081549710062454346892747275941443806473497160486483109336733176569332252601400991073341945562440371206422160096660330328199437434689491414049395736606577452033431921620786925562131563906656529268728837490976292091316375920907981757865190823433577256057787390049995;
            6'd46: xpb[30] = 1024'd22647178619942052800237553553678884755153997319554779633634649608694648222065795385132105298922475578598708205034913040829797968398568834334063913788911547800969966000488401831216805382884220277980306257328990973067119557981253857133894204665392707360967460391641725598170966714853800956225493950918842549365;
            6'd47: xpb[30] = 1024'd36625018990389134534894775087977820591646304557559849204814952324642020502687784296767050111361841820464239840737573480258604863455192106227756621155662998941609603801539368972942196716372703949383160481226060325347313553830943807611259140601947923745642829466907530288360175564516778478873731844050295048735;
            6'd48: xpb[30] = 1024'd50602859360836216269551996622276756428138611795564918775995255040589392783309773208401994923801208062329771476440233919687411758511815378121449328522414450082249241602590336114667588049861187620786014705123129677627507549680633758088624076538503140130318198542173334978549384414179756001521969737181747548105;
            6'd49: xpb[30] = 1024'd64580699731283298004209218156575692264630919033569988347175557756536765063931762120036939736240574304195303112142894359116218653568438650015142035889165901222888879403641303256392979383349671292188868929020199029907701545530323708565989012475058356514993567617439139668738593263842733524170207630313200047475;
            6'd50: xpb[30] = 1024'd78558540101730379738866439690874628101123226271575057918355860472484137344553751031671884548679940546060834747845554798545025548625061921908834743255917352363528517204692270398118370716838154963591723152917268382187895541380013659043353948411613572899668936692704944358927802113505711046818445523444652546845;
            6'd51: xpb[30] = 1024'd92536380472177461473523661225173563937615533509580127489536163188431509625175739943306829361119306787926366383548215237973832443681685193802527450622668803504168155005743237539843762050326638634994577376814337734468089537229703609520718884348168789284344305767970749049117010963168688569466683416576105046215;
            6'd52: xpb[30] = 1024'd106514220842624543208180882759472499774107840747585197060716465904378881905797728854941774173558673029791898019250875677402639338738308465696220157989420254644807792806794204681569153383815122306397431600711407086748283533079393559998083820284724005669019674843236553739306219812831666092114921309707557545585;
            6'd53: xpb[30] = 1024'd120492061213071624942838104293771435610600147985590266631896768620326254186419717766576718985998039271657429654953536116831446233794931737589912865356171705785447430607845171823294544717303605977800285824608476439028477528929083510475448756221279222053695043918502358429495428662494643614763159202839010044955;
            6'd54: xpb[30] = 1024'd10403205899393965278696398423255938702394028097859652074945216271296731129732567768196592583779731204079811883198703121681189288010334674928445447706592115992396393839324921627389696859274883927892942440118305944944310674557876687987835122474604989171550509579651105089578109438228988120292707269344868059994;
            6'd55: xpb[30] = 1024'd24381046269841047013353619957554874538886335335864721646125518987244103410354556679831537396219097445945343518901363561109996183066957946822138155073343567133036031640375888769115088192763367599295796664015375297224504670407566638465200058411160205556225878654916909779767318287891965642940945162476320559364;
            6'd56: xpb[30] = 1024'd38358886640288128748010841491853810375378642573869791217305821703191475690976545591466482208658463687810875154604024000538803078123581218715830862440095018273675669441426855910840479526251851270698650887912444649504698666257256588942564994347715421940901247730182714469956527137554943165589183055607773058734;
            6'd57: xpb[30] = 1024'd52336727010735210482668063026152746211870949811874860788486124419138847971598534503101427021097829929676406790306684439967609973180204490609523569806846469414315307242477823052565870859740334942101505111809514001784892662106946539419929930284270638325576616805448519160145735987217920688237420948739225558104;
            6'd58: xpb[30] = 1024'd66314567381182292217325284560451682048363257049879930359666427135086220252220523414736371833537196171541938426009344879396416868236827762503216277173597920554954945043528790194291262193228818613504359335706583354065086657956636489897294866220825854710251985880714323850334944836880898210885658841870678057474;
            6'd59: xpb[30] = 1024'd80292407751629373951982506094750617884855564287884999930846729851033592532842512326371316645976562413407470061712005318825223763293451034396908984540349371695594582844579757336016653526717302284907213559603652706345280653806326440374659802157381071094927354955980128540524153686543875733533896735002130556844;
            6'd60: xpb[30] = 1024'd94270248122076455686639727629049553721347871525890069502027032566980964813464501238006261458415928655273001697414665758254030658350074306290601691907100822836234220645630724477742044860205785956310067783500722058625474649656016390852024738093936287479602724031245933230713362536206853256182134628133583056214;
            6'd61: xpb[30] = 1024'd108248088492523537421296949163348489557840178763895139073207335282928337094086490149641206270855294897138533333117326197682837553406697578184294399273852273976873858446681691619467436193694269627712922007397791410905668645505706341329389674030491503864278093106511737920902571385869830778830372521265035555584;
            6'd62: xpb[30] = 1024'd122225928862970619155954170697647425394332486001900208644387637998875709374708479061276151083294661139004064968819986637111644448463320850077987106640603725117513496247732658761192827527182753299115776231294860763185862641355396291806754609967046720248953462181777542611091780235532808301478610414396488054954;
            6'd63: xpb[30] = 1024'd12137073549292959491812464827131928486126366114169594087436085649846186318021329062896024681076353071426447197065153641961387502678723787416519688991024135324462459479212408565287979669154031249208432846804690269101695786984189469319140976220372487366808927842926289271174461011267152807008158480902346069993;
        endcase
    end

    always_comb begin
        case(flag[10][11:6])
            6'd0: xpb[31] = 1024'd0;
            6'd1: xpb[31] = 1024'd26114913919740041226469686361430864322618673352174663658616388365793558598643317974530969493515719313291978832767814081390194397735347059310212396357775586465102097280263375707013371002642514920611287070701759621381889782833879419796505912156927703751484296918192093961363669860930130329656396374033798569363;
            6'd2: xpb[31] = 1024'd52229827839480082452939372722861728645237346704349327317232776731587117197286635949061938987031438626583957665535628162780388795470694118620424792715551172930204194560526751414026742005285029841222574141403519242763779565667758839593011824313855407502968593836384187922727339721860260659312792748067597138726;
            6'd3: xpb[31] = 1024'd78344741759220123679409059084292592967856020056523990975849165097380675795929953923592908480547157939875936498303442244170583193206041177930637189073326759395306291840790127121040113007927544761833861212105278864145669348501638259389517736470783111254452890754576281884091009582790390988969189122101395708089;
            6'd4: xpb[31] = 1024'd104459655678960164905878745445723457290474693408698654634465553463174234394573271898123877974062877253167915331071256325560777590941388237240849585431102345860408389121053502828053484010570059682445148282807038485527559131335517679186023648627710815005937187672768375845454679443720521318625585496135194277452;
            6'd5: xpb[31] = 1024'd6507873914575464733549504402339888868394939635137634164950086763990897655907450962639776252920922257016744756381576972371908147835514961995901856772546891391819811831745661197436615821695368881746237745121558260545088063948500326017550991101409069490601581176843411776711821230722018631163292043543398362484;
            6'd6: xpb[31] = 1024'd32622787834315505960019190763770753191013612987312297823566475129784456254550768937170745746436641570308723589149391053762102545570862021306114253130322477856921909112009036904449986824337883802357524815823317881926977846782379745814056903258336773242085878095035505738075491091652148960819688417577196931847;
            6'd7: xpb[31] = 1024'd58737701754055547186488877125201617513632286339486961482182863495578014853194086911701715239952360883600702421917205135152296943306209080616326649488098064322024006392272412611463357826980398722968811886525077503308867629616259165610562815415264476993570175013227599699439160952582279290476084791610995501210;
            6'd8: xpb[31] = 1024'd84852615673795588412958563486632481836250959691661625140799251861371573451837404886232684733468080196892681254685019216542491341041556139926539045845873650787126103672535788318476728829622913643580098957226837124690757412450138585407068727572192180745054471931419693660802830813512409620132481165644794070573;
            6'd9: xpb[31] = 1024'd110967529593535629639428249848063346158869633043836288799415640227165132050480722860763654226983799510184660087452833297932685738776903199236751442203649237252228200952799164025490099832265428564191386027928596746072647195284018005203574639729119884496538768849611787622166500674442539949788877539678592639936;
            6'd10: xpb[31] = 1024'd13015747829150929467099008804679777736789879270275268329900173527981795311814901925279552505841844514033489512763153944743816295671029923991803713545093782783639623663491322394873231643390737763492475490243116521090176127897000652035101982202818138981203162353686823553423642461444037262326584087086796724968;
            6'd11: xpb[31] = 1024'd39130661748890970693568695166110642059408552622449931988516561893775353910458219899810521999357563827325468345530968026134010693406376983302016109902869369248741720943754698101886602646033252684103762560944876142472065910730880071831607894359745842732687459271878917514787312322374167591982980461120595294331;
            6'd12: xpb[31] = 1024'd65245575668631011920038381527541506382027225974624595647132950259568912509101537874341491492873283140617447178298782107524205091141724042612228506260644955713843818224018073808899973648675767604715049631646635763853955693564759491628113806516673546484171756190071011476150982183304297921639376835154393863694;
            6'd13: xpb[31] = 1024'd91360489588371053146508067888972370704645899326799259305749338625362471107744855848872460986389002453909426011066596188914399488877071101922440902618420542178945915504281449515913344651318282525326336702348395385235845476398638911424619718673601250235656053108263105437514652044234428251295773209188192433057;
            6'd14: xpb[31] = 1024'd117475403508111094372977754250403235027264572678973922964365726991156029706388173823403430479904721767201404843834410270304593886612418161232653298976196128644048012784544825222926715653960797445937623773050155006617735259232518331221125630830528953987140350026455199398878321905164558580952169583221991002420;
            6'd15: xpb[31] = 1024'd19523621743726394200648513207019666605184818905412902494850260291972692967722352887919328758762766771050234269144730917115724443506544885987705570317640674175459435495236983592309847465086106645238713235364674781635264191845500978052652973304227208471804743530530235330135463692166055893489876130630195087452;
            6'd16: xpb[31] = 1024'd45638535663466435427118199568450530927803492257587566153466648657766251566365670862450298252278486084342213101912544998505918841241891945297917966675416260640561532775500359299323218467728621565850000306066434403017153974679380397849158885461154912223289040448722329291499133553096186223146272504663993656815;
            6'd17: xpb[31] = 1024'd71753449583206476653587885929881395250422165609762229812083037023559810165008988836981267745794205397634191934680359079896113238977239004608130363033191847105663630055763735006336589470371136486461287376768194024399043757513259817645664797618082615974773337366914423252862803414026316552802668878697792226178;
            6'd18: xpb[31] = 1024'd97868363502946517880057572291312259573040838961936893470699425389353368763652306811512237239309924710926170767448173161286307636712586063918342759390967433570765727336027110713349960473013651407072574447469953645780933540347139237442170709775010319726257634285106517214226473274956446882459065252731590795541;
            6'd19: xpb[31] = 1024'd123983277422686559106527258652743123895659512314111557129315813755146927362295624786043206732825644024218149600215987242676502034447933123228555155748743020035867824616290486420363331475656166327683861518171713267162823323181018657238676621931938023477741931203298611175590143135886577212115461626765389364904;
            6'd20: xpb[31] = 1024'd26031495658301858934198017609359555473579758540550536659800347055963590623629803850559105011683689028066979025526307889487632591342059847983607427090187565567279247326982644789746463286781475526984950980486233042180352255794001304070203964405636277962406324707373647106847284922888074524653168174173593449936;
            6'd21: xpb[31] = 1024'd52146409578041900160667703970790419796198431892725200318416735421757149222273121825090074505199408341358957858294121970877826989077406907293819823447963152032381344607246020496759834289423990447596238051187992663562242038627880723866709876562563981713890621625565741068210954783818204854309564548207392019299;
            6'd22: xpb[31] = 1024'd78261323497781941387137390332221284118817105244899863977033123787550707820916439799621043998715127654650936691061936052268021386812753966604032219805738738497483441887509396203773205292066505368207525121889752284944131821461760143663215788719491685465374918543757835029574624644748335183965960922241190588662;
            6'd23: xpb[31] = 1024'd104376237417521982613607076693652148441435778597074527635649512153344266419559757774152013492230846967942915523829750133658215784548101025914244616163514324962585539167772771910786576294709020288818812192591511906326021604295639563459721700876419389216859215461949928990938294505678465513622357296274989158025;
            6'd24: xpb[31] = 1024'd6424455653137282441277835650268580019356024823513507166134045454160929680893936838667911771088891971791744949140070780469346341442227750669296887504958870493996961878464930280169708105834329488119901654906031681343550536908622210291249043350117643701523608966024964922195436292679962826160063843683193243057;
            6'd25: xpb[31] = 1024'd32539369572877323667747522011699444341974698175688170824750433819954488279537254813198881264604611285083723781907884861859540739177574809979509283862734456959099059158728305987183079108476844408731188725607791302725440319742501630087754955507045347453007905884217058883559106153610093155816460217716991812420;
            6'd26: xpb[31] = 1024'd58654283492617364894217208373130308664593371527862834483366822185748046878180572787729850758120330598375702614675698943249735136912921869289721680220510043424201156438991681694196450111119359329342475796309550924107330102576381049884260867663973051204492202802409152844922776014540223485472856591750790381783;
            6'd27: xpb[31] = 1024'd84769197412357406120686894734561172987212044880037498141983210551541605476823890762260820251636049911667681447443513024639929534648268928599934076578285629889303253719255057401209821113761874249953762867011310545489219885410260469680766779820900754955976499720601246806286445875470353815129252965784588951146;
            6'd28: xpb[31] = 1024'd110884111332097447347156581095992037309830718232212161800599598917335164075467208736791789745151769224959660280211327106030123932383615987910146472936061216354405350999518433108223192116404389170565049937713070166871109668244139889477272691977828458707460796638793340767650115736400484144785649339818387520509;
            6'd29: xpb[31] = 1024'd12932329567712747174827340052608468887750964458651141331084132218151827336801387801307688024009814228808489705521647752841254489277742712665198744277505761885816773710210591477606323927529698369866139400027589941888638600857122536308800034451526713192125190142868376698907257523401981457323355887226591605541;
            6'd30: xpb[31] = 1024'd39047243487452788401297026414039333210369637810825804989700520583945385935444705775838657517525533542100468538289461834231448887013089771975411140635281348350918870990473967184619694930172213290477426470729349563270528383691001956105305946608454416943609487061060470660270927384332111786979752261260390174904;
            6'd31: xpb[31] = 1024'd65162157407192829627766712775470197532988311163000468648316908949738944534088023750369627011041252855392447371057275915621643284748436831285623536993056934816020968270737342891633065932814728211088713541431109184652418166524881375901811858765382120695093783979252564621634597245262242116636148635294188744267;
            6'd32: xpb[31] = 1024'd91277071326932870854236399136901061855606984515175132306933297315532503132731341724900596504556972168684426203825089997011837682483783890595835933350832521281123065551000718598646436935457243131700000612132868806034307949358760795698317770922309824446578080897444658582998267106192372446292545009327987313630;
            6'd33: xpb[31] = 1024'd117391985246672912080706085498331926178225657867349795965549685681326061731374659699431565998072691481976405036592904078402032080219130949906048329708608107746225162831264094305659807938099758052311287682834628427416197732192640215494823683079237528198062377815636752544361936967122502775948941383361785882993;
            6'd34: xpb[31] = 1024'd19440203482288211908376844454948357756145904093788775496034218982142724992708838763947464276930736485825234461903224725213162637113257674661100601050052653277636585541956252675042939749225067251612377145149148202433726664805622862326351025552935782682726771319711788475619078754124000088486647930769989968025;
            6'd35: xpb[31] = 1024'd45555117402028253134846530816379222078764577445963439154650607347936283591352156738478433770446455799117213294671038806603357034848604733971312997407828239742738682822219628382056310751867582172223664215850907823815616447639502282122856937709863486434211068237903882436982748615054130418143044304803788537388;
            6'd36: xpb[31] = 1024'd71670031321768294361316217177810086401383250798138102813266995713729842189995474713009403263962175112409192127438852887993551432583951793281525393765603826207840780102483004089069681754510097092834951286552667445197506230473381701919362849866791190185695365156095976398346418475984260747799440678837587106751;
            6'd37: xpb[31] = 1024'd97784945241508335587785903539240950724001924150312766471883384079523400788638792687540372757477894425701170960206666969383745830319298852591737790123379412672942877382746379796083052757152612013446238357254427066579396013307261121715868762023718893937179662074288070359710088336914391077455837052871385676114;
            6'd38: xpb[31] = 1024'd123899859161248376814255589900671815046620597502487430130499772445316959387282110662071342250993613738993149792974481050773940228054645911901950186481154999138044974663009755503096423759795126934057525427956186687961285796141140541512374674180646597688663958992480164321073758197844521407112233426905184245477;
            6'd39: xpb[31] = 1024'd25948077396863676641926348857288246624540843728926409660984305746133622648616289726587240529851658742841979218284801697585070784948772636657002457822599544669456397373701913872479555570920436133358614890270706462978814728754123188343902016654344852173328352496555200252330899984846018719649939974313388330509;
            6'd40: xpb[31] = 1024'd52062991316603717868396035218719110947159517081101073319600694111927181247259607701118210023367378056133958051052615778975265182684119695967214854180375131134558494653965289579492926573562951053969901960972466084360704511588002608140407928811272555924812649414747294213694569845776149049306336348347186899872;
            6'd41: xpb[31] = 1024'd78177905236343759094865721580149975269778190433275736978217082477720739845902925675649179516883097369425936883820429860365459580419466755277427250538150717599660591934228665286506297576205465974581189031674225705742594294421882027936913840968200259676296946332939388175058239706706279378962732722380985469235;
            6'd42: xpb[31] = 1024'd104292819156083800321335407941580839592396863785450400636833470843514298444546243650180149010398816682717915716588243941755653978154813814587639646895926304064762689214492040993519668578847980895192476102375985327124484077255761447733419753125127963427781243251131482136421909567636409708619129096414784038598;
            6'd43: xpb[31] = 1024'd6341037391699100149006166898197271170317110011889380167318004144330961705880422714696047289256861686566745141898564588566784535048940539342691918237370849596174111925184199362902800389973290094493565564690505102142013009868744094564947095598826217912445636755206518067679051354637907021156835643822988123630;
            6'd44: xpb[31] = 1024'd32455951311439141375475853259628135492935783364064043825934392510124520304523740689227016782772580999858723974666378669956978932784287598652904314595146436061276209205447575069916171392615805015104852635392264723523902792702623514361453007755753921663929933673398612029042721215568037350813232017856786692993;
            6'd45: xpb[31] = 1024'd58570865231179182601945539621058999815554456716238707484550780875918078903167058663757986276288300313150702807434192751347173330519634657963116710952922022526378306485710950776929542395258319935716139706094024344905792575536502934157958919912681625415414230591590705990406391076498167680469628391890585262356;
            6'd46: xpb[31] = 1024'd84685779150919223828415225982489864138173130068413371143167169241711637501810376638288955769804019626442681640202006832737367728254981717273329107310697608991480403765974326483942913397900834856327426776795783966287682358370382353954464832069609329166898527509782799951770060937428298010126024765924383831719;
            6'd47: xpb[31] = 1024'd110800693070659265054884912343920728460791803420588034801783557607505196100453694612819925263319738939734660472969820914127562125990328776583541503668473195456582501046237702190956284400543349776938713847497543587669572141204261773750970744226537032918382824427974893913133730798358428339782421139958182401082;
            6'd48: xpb[31] = 1024'd12848911306274564882555671300537160038712049647027014332268090908321859361787873677335823542177783943583489898280141560938692682884455501338593775009917740987993923756929860560339416211668658976239803309812063362687101073817244420582498086700235287403047217932049929844390872585359925652320127687366386486114;
            6'd49: xpb[31] = 1024'd38963825226014606109025357661968024361330722999201677990884479274115417960431191651866793035693503256875468731047955642328887080619802560648806171367693327453096021037193236267352787214311173896851090380513822984068990856651123840379003998857162991154531514850242023805754542446290055981976524061400185055477;
            6'd50: xpb[31] = 1024'd65078739145754647335495044023398888683949396351376341649500867639908976559074509626397762529209222570167447563815769723719081478355149619959018567725468913918198118317456611974366158216953688817462377451215582605450880639485003260175509911014090694906015811768434117767118212307220186311632920435433983624840;
            6'd51: xpb[31] = 1024'd91193653065494688561964730384829753006568069703551005308117256005702535157717827600928732022724941883459426396583583805109275876090496679269230964083244500383300215597719987681379529219596203738073664521917342226832770422318882679972015823171018398657500108686626211728481882168150316641289316809467782194203;
            6'd52: xpb[31] = 1024'd117308566985234729788434416746260617329186743055725668966733644371496093756361145575459701516240661196751405229351397886499470273825843738579443360441020086848402312877983363388392900222238718658684951592619101848214660205152762099768521735327946102408984405604818305689845552029080446970945713183501580763566;
            6'd53: xpb[31] = 1024'd19356785220850029616105175702877048907106989282164648497218177672312757017695324639975599795098706200600234654661718533310600830719970463334495631782464632379813735588675521757776032033364027857986041054933621623232189137765744746600049077801644356893648799108893341621102693816081944283483419730909784848598;
            6'd54: xpb[31] = 1024'd45471699140590070842574862064307913229725662634339312155834566038106315616338642614506569288614425513892213487429532614700795228455317522644708028140240218844915832868938897464789403036006542778597328125635381244614078920599624166396554989958572060645133096027085435582466363677012074613139816104943583417961;
            6'd55: xpb[31] = 1024'd71586613060330112069044548425738777552344335986513975814450954403899874214981960589037538782130144827184192320197346696090989626190664581954920424498015805310017930149202273171802774038649057699208615196337140865995968703433503586193060902115499764396617392945277529543830033537942204942796212478977381987324;
            6'd56: xpb[31] = 1024'd97701526980070153295514234787169641874963009338688639473067342769693432813625278563568508275645864140476171152965160777481184023926011641265132820855791391775120027429465648878816145041291572619819902267038900487377858486267383005989566814272427468148101689863469623505193703398872335272452608853011180556687;
            6'd57: xpb[31] = 1024'd123816440899810194521983921148600506197581682690863303131683731135486991412268596538099477769161583453768149985732974858871378421661358700575345217213566978240222124709729024585829516043934087540431189337740660108759748269101262425786072726429355171899585986781661717466557373259802465602109005227044979126050;
            6'd58: xpb[31] = 1024'd25864659135425494349654680105216937775501928917302282662168264436303654673602775602615376048019628457616979411043295505682508978555485425330397488555011523771633547420421182955212647855059396739732278800055179883777277201714245072617600068903053426384250380285736753397814515046803962914646711774453183211082;
            6'd59: xpb[31] = 1024'd51979573055165535576124366466647802098120602269476946320784652802097213272246093577146345541535347770908958243811109587072703376290832484640609884912787110236735644700684558662226018857701911660343565870756939505159166984548124492414105981059981130135734677203928847359178184907734093244303108148486981780445;
            6'd60: xpb[31] = 1024'd78094486974905576802594052828078666420739275621651609979401041167890771870889411551677315035051067084200937076578923668462897774026179543950822281270562696701837741980947934369239389860344426580954852941458699126541056767382003912210611893216908833887218974122120941320541854768664223573959504522520780349808;
            6'd61: xpb[31] = 1024'd104209400894645618029063739189509530743357948973826273638017429533684330469532729526208284528566786397492915909346737749853092171761526603261034677628338283166939839261211310076252760862986941501566140012160458747922946550215883332007117805373836537638703271040313035281905524629594353903615900896554578919171;
            6'd62: xpb[31] = 1024'd6257619130260917856734498146125962321278195200265253168501962834500993730866908590724182807424831401341745334657058396664222728655653328016086948969782828698351261971903468445635892674112250700867229474474978522940475482828865978838645147847534792123367664544388071213162666416595851216153607443962783004203;
            6'd63: xpb[31] = 1024'd32372533050000959083204184507556826643896868552439916827118351200294552329510226565255152300940550714633724167424872478054417126391000387326299345327558415163453359252166844152649263676754765621478516545176738144322365265662745398635151060004462495874851961462580165174526336277525981545810003817996581573566;
        endcase
    end

    always_comb begin
        case(flag[10][16:12])
            5'd0: xpb[32] = 1024'd0;
            5'd1: xpb[32] = 1024'd58487446969741000309673870868987690966515541904614580485734739566088110928153544539786121794456270027925703000192686559444611524126347446636511741685334001628555456532430219859662634679397280542089803615878497765704255048496624818431656972161390199626336258380772259135890006138456111875466400192030380142929;
            5'd2: xpb[32] = 1024'd116974893939482000619347741737975381933031083809229160971469479132176221856307089079572243588912540055851406000385373118889223048252694893273023483370668003257110913064860439719325269358794561084179607231756995531408510096993249636863313944322780399252672516761544518271780012276912223750932800384060760285858;
            5'd3: xpb[32] = 1024'd51395645225098259530222685202148640154848198588108057329072363633287437447151494709343294168711135774333959593120566243754770731537822005354375100039670963951975695027719442241357664846674635904959213239248253450748404295268977682329992346800941149612188871728199719377563490341439702609280510749465545944456;
            5'd4: xpb[32] = 1024'd109883092194839259839896556071136331121363740492722637814807103199375548375305039249129415963167405802259662593313252803199382255664169451990886841725004965580531151560149662101020299526071916447049016855126751216452659343765602500761649318962331349238525130108971978513453496479895814484746910941495926087385;
            5'd5: xpb[32] = 1024'd44303843480455518750771499535309589343180855271601534172409987700486763966149444878900466542966001520742216186048445928064929938949296564072238458394007926275395933523008664623052695013951991267828622862618009135792553542041330546228327721440492099598041485075627179619236974544423293343094621306900711745983;
            5'd6: xpb[32] = 1024'd102791290450196519060445370404297280309696397176216114658144727266574874894302989418686588337422271548667919186241132487509541463075644010708750200079341927903951390055438884482715329693349271809918426478496506901496808590537955364659984693601882299224377743456399438755126980682879405218561021498931091888912;
            5'd7: xpb[32] = 1024'd37212041735812777971320313868470538531513511955095011015747611767686090485147395048457638917220867267150472778976325612375089146360771122790101816748344888598816172018297887004747725181229346630698032485987764820836702788813683410126663096080043049583894098423054639860910458747406884076908731864335877547510;
            5'd8: xpb[32] = 1024'd95699488705553778280994184737458229498029053859709591501482351333774201413300939588243760711677137295076175779169012171819700670487118569426613558433678890227371628550728106864410359860626627172787836101866262586540957837310308228558320068241433249210230356803826898996800464885862995952375132056366257690439;
            5'd9: xpb[32] = 1024'd30120239991170037191869128201631487719846168638588487859085235834885417004145345218014811291475733013558729371904205296685248353772245681507965175102681850922236410513587109386442755348506701993567442109357520505880852035586036274024998470719593999569746711770482100102583942950390474810722842421771043349037;
            5'd10: xpb[32] = 1024'd88607686960911037501542999070619178686361710543203068344819975400973527932298889757800933085932003041484432372096891856129859877898593128144476916788015852550791867046017329246105390027903982535657245725236018271585107084082661092456655442880984199196082970151254359238473949088846586686189242613801423491966;
            5'd11: xpb[32] = 1024'd23028438246527296412417942534792436908178825322081964702422859902084743523143295387571983665730598759966985964832084980995407561183720240225828533457018813245656649008876331768137785515784057356436851732727276190925001282358389137923333845359144949555599325117909560344257427153374065544536952979206209150564;
            5'd12: xpb[32] = 1024'd81515885216268296722091813403780127874694367226696545188157599468172854451296839927358105460186868787892688965024771540440019085310067686862340275142352814874212105541306551627800420195181337898526655348605773956629256330855013956354990817520535149181935583498681819480147433291830177420003353171236589293493;
            5'd13: xpb[32] = 1024'd15936636501884555632966756867953386096511482005575441545760483969284070042141245557129156039985464506375242557759964665305566768595194798943691891811355775569076887504165554149832815683061412719306261356097031875969150529130742001821669219998695899541451938465337020585930911356357656278351063536641374952091;
            5'd14: xpb[32] = 1024'd74424083471625555942640627736941077063027023910190022031495223535372180970294790096915277834441734534300945557952651224750178292721542245580203633496689777197632344036595774009495450362458693261396064971975529641673405577627366820253326192160086099167788196846109279721820917494813768153817463728671755095020;
            5'd15: xpb[32] = 1024'd8844834757241814853515571201114335284844138689068918389098108036483396561139195726686328414240330252783499150687844349615725976006669357661555250165692737892497125999454776531527845850338768082175670979466787561013299775903094865720004594638246849527304551812764480827604395559341247012165174094076540753618;
            5'd16: xpb[32] = 1024'd67332281726982815163189442070102026251359680593683498874832847602571507489292740266472450208696600280709202150880530909060337500133016804298066991851026739521052582531884996391190480529736048624265474595345285326717554824399719684151661566799637049153640810193536739963494401697797358887631574286106920896547;
            5'd17: xpb[32] = 1024'd1753033012599074074064385534275284473176795372562395232435732103682723080137145896243500788495195999191755743615724033925885183418143916379418608520029700215917364494743998913222876017616123445045080602836543246057449022675447729618339969277797799513157165160191941069277879762324837745979284651511706555145;
            5'd18: xpb[32] = 1024'd60240479982340074383738256403262975439692337277176975718170471669770834008290690436029622582951466027117458743808410593370496707544491363015930350205363701844472821027174218772885510697013403987134884218715041011761704071172072548049996941439187999139493423540964200205167885900780949621445684843542086698074;
            5'd19: xpb[32] = 1024'd118727926952081074693412127272250666406207879181791556203905211235858944936444234975815744377407736055043161744001097152815108231670838809652442091890697703473028277559604438632548145376410684529224687834593538777465959119668697366481653913600578198765829681921736459341057892039237061496912085035572466841003;
            5'd20: xpb[32] = 1024'd53148678237697333604287070736423924628024993960670452561508095736970160527288640605586794957206331773525715336736290277680655914955965921733793708559700664167893059522463441154580540864290759350004293842084796696805853317944425411948332316078738949125346036888391660446841370103764540355259795400977252499601;
            5'd21: xpb[32] = 1024'd111636125207438333913960941605411615594540535865285033047242835303058271455442185145372916751662601801451418336928976837125267439082313368370305450245034665796448516054893661014243175543688039892094097457963294462510108366441050230379989288240129148751682295269163919582731376242220652230726195593007632642530;
            5'd22: xpb[32] = 1024'd46056876493054592824835885069584873816357650644163929404845719804169487046286590775143967331461197519933971929664169961990815122367440480451657066914037626491313298017752663536275571031568114712873703465454552381850002564716778275846667690718289899111198650235819120688514854306748131089073905958412418301128;
            5'd23: xpb[32] = 1024'd104544323462795593134509755938572564782873192548778509890580459370257597974440135314930089125917467547859674929856856521435426646493787927088168808599371628119868754550182883395938205710965395254963507081333050147554257613213403094278324662879680098737534908616591379824404860445204242964540306150442798444057;
            5'd24: xpb[32] = 1024'd38965074748411852045384699402745823004690307327657406248183343871368813565284540944701139705716063266342228522592049646300974329778915039169520425268374588814733536513041885917970601198845470075743113088824308066894151811489131139745003065357840849097051263583246580930188338509731721822888016515847584102655;
            5'd25: xpb[32] = 1024'd97452521718152852355058570271733513971205849232271986733918083437456924493438085484487261500172333294267931522784736205745585853905262485806032166953708590443288993045472105777633235878242750617832916704702805832598406859985755958176660037519231048723387521964018840066078344648187833698354416707877964245584;
            5'd26: xpb[32] = 1024'd31873273003769111265933513735906772193022964011150883091520967938568140084282491114258312079970929012750485115519929330611133537190389597887383783622711551138153775008331108299665631366122825438612522712194063751938301058261484003643338439997391799082903876930674041171861822712715312556702127073282749904182;
            5'd27: xpb[32] = 1024'd90360719973510111575607384604894463159538505915765463577255707504656251012436035654044433874427199040676188115712615890055745061316737044523895525308045552766709231540761328159328266045520105980702326328072561517642556106758108822074995412158781998709240135311446300307751828851171424432168527265313130047111;
            5'd28: xpb[32] = 1024'd24781471259126370486482328069067721381355620694644359934858592005767466603280441283815484454225794759158741708447809014921292744601864156605247141977048513461574013503620330681360661533400180801481932335563819436982450305033836867541673814636942749068756490278101501413535306915698903290516237630717915705709;
            5'd29: xpb[32] = 1024'd83268918228867370796156198938055412347871162599258940420593331571855577531433985823601606248682064787084444708640495574365904268728211603241758883662382515090129470036050550541023296212797461343571735951442317202686705353530461685973330786798332948695092748658873760549425313054155015165982637822748295848638;
            5'd30: xpb[32] = 1024'd17689669514483629707031142402228670569688277378137836778196216072966793122278391453372656828480660505566998301375688699231451952013338715323110500331385475784994251998909553063055691700677536164351341958933575122026599551806189731440009189276493699054609103625528961655208791118682494024330348188153081507236;
            5'd31: xpb[32] = 1024'd76177116484224630016705013271216361536203819282752417263930955639054904050431935993158778622936930533492701301568375258676063476139686161959622242016719477413549708531339772922718326380074816706441145574812072887730854600302814549871666161437883898680945362006301220791098797257138605899796748380183461650165;
        endcase
    end

    always_comb begin
        case(flag[11][5:0])
            6'd0: xpb[33] = 1024'd0;
            6'd1: xpb[33] = 1024'd67332281726982815163189442070102026251359680593683498874832847602571507489292740266472450208696600280709202150880530909060337500133016804298066991851026739521052582531884996391190480529736048624265474595345285326717554824399719684151661566799637049153640810193536739963494401697797358887631574286106920896547;
            6'd2: xpb[33] = 1024'd10597867769840888927579956735389619758020934061631313621533840140166119641276341622929829202735526251975254894303568383541611159424813274040973858685722438108414490494198775444750721867954891527220751582303330807070748798578542595338344563916044649040461716972956421896882275321666084758144458745588247308763;
            6'd3: xpb[33] = 1024'd77930149496823704090769398805491646009380614655314812496366687742737627130569081889402279411432126532684457045184099292601948659557830078339040850536749177629467073026083771835941202397690940151486226177648616133788303622978262279490006130715681698194102527166493161860376677019463443645776033031695168205310;
            6'd4: xpb[33] = 1024'd21195735539681777855159913470779239516041868123262627243067680280332239282552683245859658405471052503950509788607136767083222318849626548081947717371444876216828980988397550889501443735909783054441503164606661614141497597157085190676689127832089298080923433945912843793764550643332169516288917491176494617526;
            6'd5: xpb[33] = 1024'd88528017266664593018349355540881265767401548716946126117900527882903746771845423512332108614167652784659711939487667676143559818982643352380014709222471615737881563520282547280691924265645831678706977759951946940859052421556804874828350694631726347234564244139449583757258952341129528403920491777283415514073;
            6'd6: xpb[33] = 1024'd31793603309522666782739870206168859274062802184893940864601520420498358923829024868789487608206578755925764682910705150624833478274439822122921576057167314325243471482596326334252165603864674581662254746909992421212246395735627786015033691748133947121385150918869265690646825964998254274433376236764741926289;
            6'd7: xpb[33] = 1024'd99125885036505481945929312276270885525422482778577439739434368023069866413121765135261937816903179036634966833791236059685170978407456626420988567908194053846296054014481322725442646133600723205927729342255277747929801220135347470166695258547770996275025961112406005654141227662795613162064950522871662822836;
            6'd8: xpb[33] = 1024'd42391471079363555710319826941558479032083736246525254486135360560664478565105366491719316810942105007901019577214273534166444637699253096163895434742889752433657961976795101779002887471819566108883006329213323228282995194314170381353378255664178596161846867891825687587529101286664339032577834982352989235052;
            6'd9: xpb[33] = 1024'd109723752806346370873509269011660505283443416840208753360968208163235986054398106758191767019638705288610221728094804443226782137832269900461962426593916491954710544508680098170193368001555614733148480924558608555000550018713890065505039822463815645315487678085362427551023502984461697920209409268459910131599;
            6'd10: xpb[33] = 1024'd52989338849204444637899783676948098790104670308156568107669200700830598206381708114649146013677631259876274471517841917708055797124066370204869293428612190542072452470993877223753609339774457636103757911516654035353743992892712976691722819580223245202308584864782109484411376608330423790722293727941236543815;
            6'd11: xpb[33] = 1024'd120321620576187259801089225747050125041464350901840066982502048303402105695674448381121596222374231540585476622398372826768393297257083174502936285279638930063125035002878873614944089869510506260369232506861939362071298817292432660843384386379860294355949395058318849447905778306127782678353868014048157440362;
            6'd12: xpb[33] = 1024'd63587206619045333565479740412337718548125604369787881729203040840996717847658049737578975216413157511851529365821410301249666956548879644245843152114334628650486942965192652668504331207729349163324509493819984842424492791471255572030067383496267894242770301837738531381293651929996508548866752473529483852578;
            6'd13: xpb[33] = 1024'd6852792661903407329870255077625312054786857837735696475904033378591329999641651094036354210452083483117582109244447775730940615840676113988750018949030327237848850927506431722064572545948192066279786480778030322777686765650078483216750380612675494129591208617158213314681525553865234419379636933010810264794;
            6'd14: xpb[33] = 1024'd74185074388886222493059697147727338306146538431419195350736880981162837488934391360508804419148683763826784260124978684791278115973692918286817010800057066758901433459391428113255053075684240690545261076123315649495241590049798167368411947412312543283232018810694953278175927251662593307011211219117731161341;
            6'd15: xpb[33] = 1024'd17450660431744296257450211813014931812807791899367010097437873518757449640917992716966183413187609735092837003548016159272551775265489388029723877634752765346263341421705207166815294413903083593500538063081361129848435564228621078555094944528720143170052925590114635211563800875531319177524095678599057573557;
            6'd16: xpb[33] = 1024'd84782942158727111420639653883116958064167472493050508972270721121328957130210732983438633621884210015802039154428547068332889275398506192327790869485779504867315923953590203558005774943639132217766012658426646456565990388628340762706756511328357192323693735783651375175058202573328678065155669964705978470104;
            6'd17: xpb[33] = 1024'd28048528201585185185030168548404551570828725960998323718971713658923569282194334339896012615923135987068091897851584542814162934690302662070697736320475203454677831915903982611566016281857975120721289645384691936919184362807163673893439508444764792210514642563071057108446076197197403935668554424187304882320;
            6'd18: xpb[33] = 1024'd95380809928568000348219610618506577822188406554681822593804561261495076771487074606368462824619736267777294048732115451874500434823319466368764728171501942975730414447788979002756496811594023744986764240729977263636739187206883358045101075244401841364155452756607797071940477894994762823300128710294225778867;
            6'd19: xpb[33] = 1024'd38646395971426074112610125283794171328849660022629637340505553799089688923470675962825841818658662239043346792155152926355774094115115936111671595006197641563092322410102758056316738149812866647942041227688022743989933161385706269231784072360809441250976359536027479005328351518863488693813013169775552191083;
            6'd20: xpb[33] = 1024'd105978677698408889275799567353896197580209340616313136215338401401661196412763416229298292027355262519752548943035683835416111594248132740409738586857224381084144904941987754447507218679548915272207515823033308070707487985785425953383445639160446490404617169729564218968822753216660847581444587455882473087630;
            6'd21: xpb[33] = 1024'd49244263741266963040190082019183791086870594084260950962039393939255808564747017585755671021394188491018601686458721309897385253539929210152645453691920079671506812904301533501067460017767758175162792809991353551060681959964248864570128636276854090291438076508983900902210626840529573451957471915363799499846;
            6'd22: xpb[33] = 1024'd116576545468249778203379524089285817338230274677944449836872241541827316054039757852228121230090788771727803837339252218957722753672946014450712445542946819192559395436186529892257940547503806799428267405336638877778236784363968548721790203076491139445078886702520640865705028538326932339589046201470720396393;
            6'd23: xpb[33] = 1024'd59842131511107851967770038754573410844891528145892264583573234079421928206023359208685500224129714742993856580762289693438996412964742484193619312377642517779921303398500308945818181885722649702383544392294684358131430758542791459908473200192898739331899793481940322799092902162195658210101930660952046808609;
            6'd24: xpb[33] = 1024'd3107717553965925732160553419861004351552781613840079330274226617016540358006960565142879218168640714259909324185327167920270072256538953936526179212338216367283211360814087999378423223941492605338821379252729838484624732721614371095156197309306339218720700261360004732480775786064384080614815120433373220825;
            6'd25: xpb[33] = 1024'd70439999280948740895349995489963030602912462207523578205107074219588047847299700831615329426865240994969111475065858076980607572389555758234593171063364955888335793892699084390568903753677541229604295974598015165202179557121334055246817764108943388372361510454896744695975177483861742968246389406540294117372;
            6'd26: xpb[33] = 1024'd13705585323806814659740510155250624109573715675471392951808066757182659999283302188072708420904166966235164218488895551461881231681352227977500037898060654475697701855012863444129145091896384132559572961556060645555373531300156966433500761225350988259182417234316426629363051107730468838759273866021620529588;
            6'd27: xpb[33] = 1024'd81037867050789629822929952225352650360933396269154891826640914359754167488576042454545158629600767246944366369369426460522218731814369032275567029749087393996750284386897859835319625621632432756825047556901345972272928355699876650585162328024988037412823227427853166592857452805527827726390848152128541426135;
            6'd28: xpb[33] = 1024'd24303453093647703587320466890640243867594649737102706573341906897348779640559643811002537623639693218210419112792463935003492391106165502018473896583783092584112192349211638888879866959851275659780324543859391452626122329878699561771845325141395637299644134207272848526245326429396553596903732611609867838351;
            6'd29: xpb[33] = 1024'd91635734820630518750509908960742270118954330330786205448174754499920287129852384077474987832336293498919621263672994844063829891239182306316540888434809832105164774881096635280070347489587324284045799139204676779343677154278419245923506891941032686453284944400809588489739728127193912484535306897716788734898;
            6'd30: xpb[33] = 1024'd34901320863488592514900423626029863625615583798734020194875747037514899281835985433932366826375219470185674007096032318545103550530978776059447755269505530692526682843410414333630588827806167187001076126162722259696871128457242157110189889057440286340105851180229270423127601751062638355048191357198115147114;
            6'd31: xpb[33] = 1024'd102233602590471407678089865696131889876975264392417519069708594640086406771128725700404817035071819750894876157976563227605441050663995580357514747120532270213579265375295410724821069357542215811266550721508007586414425952856961841261851455857077335493746661373766010386622003448859997242679765643305036043661;
            6'd32: xpb[33] = 1024'd45499188633329481442480380361419483383636517860365333816409587177681018923112327056862196029110745722160928901399600702086714709955792050100421613955227968800941173337609189778381310695761058714221827708466053066767619927035784752448534452973484935380567568153185692320009877072728723113192650102786362455877;
            6'd33: xpb[33] = 1024'd112831470360312296605669822431521509634996198454048832691242434780252526412405067323334646237807346002870131052280131611147052210088808854398488605806254708321993755869494186169571791225497107338487302303811338393485174751435504436600196019773121984534208378346722432283504278770526082000824224388893283352424;
            6'd34: xpb[33] = 1024'd56097056403170370370060337096809103141657451921996647437943427317847138564388668679792025231846271974136183795703169085628325869380605324141395472640950406909355663831807965223132032563715950241442579290769383873838368725614327347786879016889529584421029285126142114216892152394394807871337108848374609764640;
            6'd35: xpb[33] = 1024'd123429338130153185533249779166911129393017132515680146312776274920418646053681408946264475440542872254845385946583699994688663369513622128439462464491977146430408246363692961614322513093451998865708053886114669200555923550014047031938540583689166633574670095319678854180386554092192166758968683134481530661187;
            6'd36: xpb[33] = 1024'd66694924173011259297640293832198722899678385983627961059477267458013258205665010302721854434581798226111438690006737469169937028805418598182369331326672845017770154326006740667882754431670841768663330873072714680909117524192869943125223580805574233461491002099098536113774427716060892629481567593962857073403;
            6'd37: xpb[33] = 1024'd9960510215869333062030808497486316406339639451575775806178259995607870357648611659179233428620724197377491433429774943651210688097215067925276198161368543605132062288320519721442995769889684671618607860030760161262311498371692854311906577921981833348311908878518218047162301339929618499994452053444183485619;
            6'd38: xpb[33] = 1024'd77292791942852148225220250567588342657699320045259274681011107598179377846941351925651683637317324478086693584310305852711548188230231872223343190012395283126184644820205516112633476299625733295884082455376045487979866322771412538463568144721618882501952719072054958010656703037726977387626026339551104382166;
            6'd39: xpb[33] = 1024'd20558377985710221989610765232875936164360573513207089427712100135773989998924953282109062631356250449352746327733343327192821847522028341966250056847090981713546552782519295166193717637844576198839359442334090968333060296950235449650251141838026482388773625851474639944044576661595703258138910799032430794382;
            6'd40: xpb[33] = 1024'd87890659712693037152800207302977962415720254106890588302544947738345497488217693548581512840052850730061948478613874236253159347655045146264317048698117721234599135314404291557384198167580624823104834037679376295050615121349955133801912708637663531542414436045011379907538978359393062145770485085139351690929;
            6'd41: xpb[33] = 1024'd31156245755551110917190721968265555922381507574838403049245940275940109640201294905038891834091776701328001222036911710734433006946841616007223915532813419821961043276718070610944439505799467726060111024637421775403809095528778044988595705754071131429235342824431061840926851983261788016283369544620678103145;
            6'd42: xpb[33] = 1024'd98488527482533926080380164038367582173741188168521901924078787878511617129494035171511342042788376982037203372917442619794770507079858420305290907383840159343013625808603067002134920035535516350325585619982707102121363919928497729140257272553708180582876153017967801804421253681059146903914943830727598999692;
            6'd43: xpb[33] = 1024'd41754113525391999844770678703655175680402441636469716670779780416106229281477636527968721036827302953303256116340480094276044166371654890048197774218535857930375533770916846055695161373754359253280862606940752582474557894107320640326940269670115780469697059797387483737809127304927872774427828290208925411908;
            6'd44: xpb[33] = 1024'd109086395252374815007960120773757201931762122230153215545612628018677736770770376794441171245523903234012458267221011003336381666504671694346264766069562597451428116302801842446885641903490407877546337202286037909192112718507040324478601836469752829623337869990924223701303529002725231662059402576315846308455;
            6'd45: xpb[33] = 1024'd52351981295232888772350635439044795438423375698101030292313620556272348922753978150898550239562829205278511010644048477817655325796468164089171632904258296038790024265115621500445883241709250780501614189244083389545306692685863235665284833586160429510158776770343905634691402626593957532572287035797172720671;
            6'd46: xpb[33] = 1024'd119684263022215703935540077509146821689783056291784529167146468158843856412046718417371000448259429485987713161524579386877992825929484968387238624755285035559842606797000617891636363771445299404767088784589368716262861517085582919816946400385797478663799586963880645598185804324391316420203861321904093617218;
            6'd47: xpb[33] = 1024'd62949849065073777699930592174434415196444309759732343913847460696438468564030319773828379442298355457253765904947616861359266485221281438130145491589980734147204514759314396945196605109664142307722365771547414196616055491264405831003629397502205078550620493743300327531573677948260042290716745781385420029434;
            6'd48: xpb[33] = 1024'd6215435107931851464321106839722008703105563227680158660548453234033080716013921130285758436337281428519818648370654335840540144513077907873052358424676432734566422721628175998756846447882985210677642758505459676969249465443228742190312394618612678437441400522720009464961551572128768161229630240866746441650;
            6'd49: xpb[33] = 1024'd73547716834914666627510548909824034954465243821363657535381300836604588205306661396758208645033881709229020799251185244900877644646094712171119350275703172255619005253513172389947326977619033834943117353850745003686804289842948426341973961418249727591082210716256749428455953269926127048861204526973667338197;
            6'd50: xpb[33] = 1024'd16813302877772740391901063575111628461126497289311472282082293374199200357290262753215587639072807680495073542674222719382151303937891181914026217110398870842980913215826951443507568315837876737898394340808790484039998264021771337528656958534657327477903117495676431361843826893794852919374088986454993750413;
            6'd51: xpb[33] = 1024'd84145584604755555555090505645213654712486177882994971156915140976770707846583003019688037847769407961204275693554753628442488804070907986212093208961425610364033495747711947834698048845573925362163868936154075810757553088421491021680318525334294376631543927689213171325338228591592211807005663272561914646960;
            6'd52: xpb[33] = 1024'd27411170647613629319481020310501248219147431350942785903616133514365319998566604376145416841808333932470328436977791102923762463362704455955000075796121308951395403710025726888258290183792768265119145923112121291110747062600313932867001522450701976518364834468632853258726102215460937677518547732043241059176;
            6'd53: xpb[33] = 1024'd94743452374596444482670462380603274470507111944626284778448981116936827487859344642617867050504934213179530587858322011984099963495721260253067067647148048472447986241910723279448770713528816889384620518457406617828301887000033617018663089250339025672005644662169593222220503913258296565150122018150161955723;
            6'd54: xpb[33] = 1024'd38009038417454518247060977045890867977168365412574099525149973654531439639842945999075246044543860184445583331281359486465373622787517729995973934481843747059809894204224502333009012051747659792339897505415452098181495861178856528205346086366746625558826551441589275155608377537127022435663006477631488367939;
            6'd55: xpb[33] = 1024'd105341320144437333410250419115992894228528046006257598399982821257102947129135686265547696253240460465154785482161890395525711122920534534294040926332870486580862476736109498724199492581483708416605372100760737424899050685578576212357007653166383674712467361635126015119102779234924381323294580763738409264486;
            6'd56: xpb[33] = 1024'd48606906187295407174640933781280487735189299474205413146683813794697559281119287622005075247279386436420838225584927870006984782212331004036947793167566185168224384698423277777759733919702551319560649087718782905252244659757399123543690650282791274599288268414545697052490652858793107193807465223219735676702;
            6'd57: xpb[33] = 1024'd115939187914278222337830375851382513986548980067888912021516661397269066770412027888477525455975986717130040376465458779067322282345347808335014785018592924689276967230308274168950214449438599943826123683064068231969799484157118807695352217082428323752929078608082437015985054556590466081439039509326656573249;
            6'd58: xpb[33] = 1024'd59204773957136296102220890516670107493210233535836726768217653934863678922395629244934904450014912688396093119888496253548595941637144278077921651853288623276638875192622053222510455787657442846781400670022113712322993458335941718882035214198835923639749985387502118949372928180459191951951923968807982985465;
            6'd59: xpb[33] = 1024'd2470359999994369866611405181957700999871487003784541514918646472458291074379230601392283444053838659662145863311533728029869600928940747820828518687984321864000783154935832276070697125876285749736677656980159192676187432514764630068718211315243523526570892166921800882760801804327917822464808428289309397681;
            6'd60: xpb[33] = 1024'd69802641726977185029800847252059727251231167597468040389751494075029798563671970867864733652750438940371348014192064637090207101061957552118895510539011061385053365686820828667261177655612334374002152252325444519393742256914484314220379778114880572680211702360458540846255203502125276710096382714396230294228;
            6'd61: xpb[33] = 1024'd13068227769835258794191361917347320757892421065415855136452486612624410715655572224322112646789364911637400757615102111571480760353754021861802377373706759972415273649134607720821418993831177276957429239283489999746936231093307225407062775231288172567032609139878222779643077125994002580609267173877556706444;
            6'd62: xpb[33] = 1024'd80400509496818073957380803987449347009252101659099354011285334215195918204948312490794562855485965192346602908495633020631818260486770826159869369224733499493467856181019604112011899523567225901222903834628775326464491055493026909558724342030925221720673419333414962743137478823791361468240841459984477602991;
            6'd63: xpb[33] = 1024'd23666095539676147721771318652736940515913355127047168757986326752790530356931913847251941849524891163612655651918670495113091919778567295902776236059429198080829764143333383165572140861786068804178180821586820806817685029671849820745407339147332821607494326112834644676525352447660087338753725919465804015207;
        endcase
    end

    always_comb begin
        case(flag[11][11:6])
            6'd0: xpb[34] = 1024'd0;
            6'd1: xpb[34] = 1024'd90998377266658962884960760722838966767273035720730667632819174355362037846224654113724392058221491444321857802799201404173429419911584100200843227910455937601882346675218379556762621391522117428443655416932106133535239854071569504897068905946969870761135136306371384640019754145457446226385300205572724911754;
            6'd2: xpb[34] = 1024'd57930058849193184371122594040863500789847644315725651137506493645747180355140169317433712901785308579200566198140909373767794998981947865846526330804580834270074018780865541775895003591527029135577113225476972420706118857922242236829159242210710292255450369198625711249932980216986259435651910584519855339177;
            6'd3: xpb[34] = 1024'd24861740431727405857284427358888034812422252910720634642193812936132322864055684521143033745349125714079274593482617343362160578052311631492209433698705730938265690886512703995027385791531940842710571034021838707876997861772914968761249578474450713749765602090880037859846206288515072644918520963466985766600;
            6'd4: xpb[34] = 1024'd115860117698386368742245188081727001579695288631451302275012987291494360710280338634867425803570617158401132396281818747535589997963895731693052661609161668540148037561731083551790007183054058271154226450953944841412237715844484473658318484421420584510900738397251422499865960433972518871303821169039710678354;
            6'd5: xpb[34] = 1024'd82791799280920590228407021399751535602269897226446285779700306581879503219195853838576746647134434293279840791623526717129955577034259497338735764503286565208339709667378245770922389383058969978287684259498811128583116719695157205590408820685161006005215971289505749109779186505501332080570431547986841105777;
            6'd6: xpb[34] = 1024'd49723480863454811714568854717776069624844505821441269284387625872264645728111369042286067490698251428158549186965234686724321156104623262984418867397411461876531381773025407990054771583063881685421142068043677415753995723545829937522499156948901427499531204181760075719692412577030145289837041926933971533200;
            6'd7: xpb[34] = 1024'd16655162445989033200730688035800603647419114416436252789074945162649788237026884245995388334262068563037257582306942656318686735174987028630101970291536358544723053878672570209187153783068793392554599876588543702924874727396502669454589493212641848993846437074014402329605638648558958499103652305881101960623;
            6'd8: xpb[34] = 1024'd107653539712647996085691448758639570414692150137166920421894119518011826083251538359719780392483560007359115385106144060492116155086571128830945198201992296146605400553890949765949775174590910820998255293520649836460114581468072174351658399159611719754981573380385786969625392794016404725488952511453826872377;
            6'd9: xpb[34] = 1024'd74585221295182217571853282076664104437266758732161903926581438808396968592167053563429101236047377142237823780447852030086481734156934894476628301096117192814797072659538111985082157374595822528131713102065516123630993585318744906283748735423352141249296806272640113579538618865545217934755562890400957299800;
            6'd10: xpb[34] = 1024'd41516902877716439058015115394688638459841367327156887431268758098782111101082568767138422079611194277116532175789559999680847313227298660122311403990242089482988744765185274204214539574600734235265170910610382410801872589169417638215839071687092562743612039164894440189451844937074031144022173269348087727223;
            6'd11: xpb[34] = 1024'd8448584460250660544176948712713172482415975922151870935956077389167253609998083970847742923175011411995240571131267969275212892297662425767994506884366986151180416870832436423346921774605645942398628719155248697972751593020090370147929407950832984237927272057148766799365071008602844353288783648295218154646;
            6'd12: xpb[34] = 1024'd99446961726909623429137709435552139249689011642882538568775251744529291456222738084572134981396502856317098373930469373448642312209246525968837734794822923753062763546050815980109543166127763370842284136087354831507991447091659875044998313897802854999062408363520151439384825154060290579674083853867943066400;
            6'd13: xpb[34] = 1024'd66378643309443844915299542753576673272263620237877522073462571034914433965138253288281455824960319991195806769272177343043007891279610291614520837688947820421254435651697978199241925366132675077975741944632221118678870450942332606977088650161543276493377641255774478049298051225589103788940694232815073493823;
            6'd14: xpb[34] = 1024'd33310324891978066401461376071601207294838228832872505578149890325299576474053768491990776668524137126074515164613885312637373470349974057260203940583072717089446107757345140418374307566137586785109199753177087405849749454793005338909178986425283697987692874148028804659211277297117916998207304611762203921246;
            6'd15: xpb[34] = 1024'd242006474512287887623209389625741317412837427867489082837209615684718982969283695700097512087954260953223559955593282231739049420337822905887043477197613757637779862992302637506689766142498492242657561721953693020628458643678070841269322689024119482008107040283131269124503368646730207473914990709334348669;
            6'd16: xpb[34] = 1024'd91240383741171250772583970112464708084685873148598156715656383971046756829193937809424489570309445705275081362754794686405168469331921923106730271387653551359520126538210682194269311157664615920686312978654059826555868312715247575738338228635993990243143243346654515909144257514104176433859215196282059260423;
            6'd17: xpb[34] = 1024'd58172065323705472258745803430489242107260481743593140220343703261431899338109453013133810413873262840153789758096502655999534048402285688752413374281778448027711798643857844413401693357669527627819770787198926113726747316565920307670428564899734411737458476238908842519057483585632989643125825575229189687846;
            6'd18: xpb[34] = 1024'd25103746906239693744907636748513776129835090338588123725031022551817041847024968216843131257437079975032498153438210625593899627472649454398096477175903344695903470749505006632534075557674439334953228595743792400897626320416593039602518901163474833231773709131163169128970709657161802852392435954176320115269;
            6'd19: xpb[34] = 1024'd116102124172898656629868397471352742897108126059318791357850196907179079693249622330567523315658571419354355956237412029767329047384233554598939705086359282297785817424723386189296696949196556763396884012675898534432866174488162544499587807110444703992908845437534553768990463802619249078777736159749045027023;
            6'd20: xpb[34] = 1024'd83033805755432878116030230789377276919682734654313774862537516197564222202165137534276844159222388554233064351579119999361694626454597320244622807980484178965977489530370548408429079149201468470530341821220764821603745178338835276431678143374185125487224078329788880378903689874148062288044346538696175454446;
            6'd21: xpb[34] = 1024'd49965487337967099602192064107401810942257343249308758367224835487949364711080652737986165002786205689111772746920827968956060205524961085890305910874609075634169161636017710627561461349206380177663799629765631108774624182189508008363768479637925546981539311222043206988816915945676875497310956917643305881869;
            6'd22: xpb[34] = 1024'd16897168920501321088353897425426344964831951844303741871912154778334507219996167941695485846350022823990481142262535938550425784595324851535989013768733972302360833741664872846693843549211291884797257438310497395945503186040180740295858815901665968475854544114297533598730142017205688706577567296590436309292;
            6'd23: xpb[34] = 1024'd107895546187160283973314658148265311732104987565034409504731329133696545066220822055419877904571514268312338945061737342723855204506908951736832241679189909904243180416883252403456464940733409313240912855242603529480743040111750245192927721848635839236989680420668918238749896162663134932962867502163161221046;
            6'd24: xpb[34] = 1024'd74827227769694505459476491466289845754679596160029393009418648424081687575136337259129198748135331403191047340403445312318220783577272717382515344573314806572434852522530414622588847140738321020374370663787469816651622043962422977125018058112376260731304913312923244848663122234191948142229477881110291648469;
            6'd25: xpb[34] = 1024'd41758909352228726945638324784314379777254204755024376514105967714466830084051852462838519591699148538069755735745153281912586362647636483028198447467439703240626524628177576841721229340743232727507828472332336103822501047813095709057108394376116682225620146205177571458576348305720761351496088260057422075892;
            6'd26: xpb[34] = 1024'd8690590934762948431800158102338913799828813350019360018793287004851972592967367666547840435262965672948464131086861251506951941718000248673881550361564599908818196733824739060853611540748144434641286280877202390993380051663768440989198730639857103719935379097431898068489574377249574560762698639004552503315;
            6'd27: xpb[34] = 1024'd99688968201421911316760918825177880567101849070750027651612461360214010439192021780272232493484457117270321933886062655680381361629584348874724778272020537510700543409043118617616232932270261863084941697809308524528619905735337945886267636586826974481070515403803282708509328522707020787147998844577277415069;
            6'd28: xpb[34] = 1024'd66620649783956132802922752143202414589676457665745011156299780650599152948107536983981553337048274252149030329227770625274746940699948114520407881166145434178892215514690280836748615132275173570218399506354174811699498909586010677818357972850567395975385748296057609318422554594235833996414609223524407842492;
            6'd29: xpb[34] = 1024'd33552331366490354289084585461226948612251066260739994660987099940984295457023052187690874180612091387027738724569478594869112519770311880166090984060270330847083887620337443055880997332280085277351857314899041098870377913436683409750448309114307817469700981188311935928335780665764647205681219602471538269915;
            6'd30: xpb[34] = 1024'd484012949024575775246418779251482634825674855734978165674419231369437965938567391400195024175908521906447119911186564463478098840675645811774086954395227515275559725984605275013379532284996984485315123443907386041256917287356141682538645378048238964016214080566262538249006737293460414947829981418668697338;
            6'd31: xpb[34] = 1024'd91482390215683538660207179502090449402098710576465645798493593586731475812163221505124587082397399966228304922710387968636907518752259746012617314864851165117157906401202984831776000923807114412928970540376013519576496771358925646579607551325018109725151350386937647178268760882750906641333130186991393609092;
            6'd32: xpb[34] = 1024'd58414071798217760146369012820114983424673319171460629303180912877116618321078736708833907925961217101107013318052095938231273097822623511658300417758976061785349578506850147050908383123812026120062428348920879806747375775209598378511697887588758531219466583279191973788181986954279719850599740565938524036515;
            6'd33: xpb[34] = 1024'd25345753380751981632530846138139517447247927766455612807868232167501760829994251912543228769525034235985721713393803907825638676892987277303983520653100958453541250612497309270040765323816937827195886157465746093918254779060271110443788223852498952713781816171446300398095213025808533059866350944885654463938;
            6'd34: xpb[34] = 1024'd116344130647410944517491606860978484214520963487186280440687406522863798676218906026267620827746525680307579516193005311999068096804571377504826748563556896055423597287715688826803386715339055255639541574397852227453494633131840615340857129799468823474916952477817685038114967171265979286251651150458379375692;
            6'd35: xpb[34] = 1024'd83275812229945166003653440179003018237095572082181263945374725813248941185134421229976941671310342815186287911534713281593433675874935143150509851457681792723615269393362851045935768915343966962772999382942718514624373636982513347272947466063209244969232185370072011648028193242794792495518261529405509803115;
            6'd36: xpb[34] = 1024'd50207493812479387489815273497027552259670180677176247450062045103634083694049936433686262514874159950064996306876421251187799254945298908796192954351806689391806941499010013265068151115348878669906457191487584801795252640833186079205037802326949666463547418262326338257941419314323605704784871908352640230538;
            6'd37: xpb[34] = 1024'd17139175395013608975977106815052086282244789272171230954749364394019226202965451637395583358437977084943704702218129220782164834015662674441876057245931586059998613604657175484200533315353790377039915000032451088966131644683858811137128138590690087957862651154580664867854645385852418914051482287299770657961;
            6'd38: xpb[34] = 1024'd108137552661672571860937867537891053049517824992901898587568538749381264049190105751119975416659468529265562505017330624955594253927246774642719285156387523661880960279875555040963154706875907805483570416964557222501371498755428316034197044537659958718997787460952049507874399531309865140436782492872495569715;
            6'd39: xpb[34] = 1024'd75069234244206793347099700855915587072092433587896882092255858039766406558105620954829296260223285664144270900359038594549959832997610540288402388050512420330072632385522717260095536906880819512617028225509423509672250502606101047966287380801400380213313020353206376117787625602838678349703392871819625997138;
            6'd40: xpb[34] = 1024'd42000915826741014833261534173940121094667042182891865596943177330151549067021136158538617103787102799022979295700746564144325412067974305934085490944637316998264304491169879479227919106885731219750486034054289796843129506456773779898377717065140801707628253245460702727700851674367491558970003250766756424561;
            6'd41: xpb[34] = 1024'd8932597409275236319423367491964655117241650777886849101630496620536691575936651362247937947350919933901687691042454533738690991138338071579768593838762213666455976596817041698360301306890642926883943842599156084014008510307446511830468053328881223201943486137715029337614077745896304768236613629713886851984;
            6'd42: xpb[34] = 1024'd99930974675934199204384128214803621884514686498617516734449670975898729422161305475972330005572411378223545493841655937912120411049922171780611821749218151268338323272035421255122922698412760355327599259531262217549248364379016016727536959275851093963078622444086413977633831891353750994621913835286611763738;
            6'd43: xpb[34] = 1024'd66862656258468420690545961532828155907089295093612500239136990266283871931076820679681650849136228513102253889183363907506485990120285937426294924643343047936529995377682583474255304898417672062461057068076128504720127368229688748659627295539591515457393855336340740587547057962882564203888524214233742191161;
            6'd44: xpb[34] = 1024'd33794337841002642176707794850852689929663903688607483743824309556669014439992335883390971692700045647980962284525071877100851569190649703071978027537467944604721667483329745693387687098422583769594514876620994791891006372080361480591717631803331936951709088228595067197460284034411377413155134593180872618584;
            6'd45: xpb[34] = 1024'd726019423536863662869628168877223952238512283602467248511628847054156948907851087100292536263862782859670679866779846695217148261013468717661130431592841272913339588976907912520069298427495476727972685165861079061885375931034212523807968067072358446024321120849393807373510105940190622421744972128003046007;
            6'd46: xpb[34] = 1024'd91724396690195826547830388891716190719511548004333134881330803202416194795132505200824684594485354227181528482665981250868646568172597568918504358342048778874795686264195287469282690689949612905171628102097967212597125230002603717420876874014042229207159457427220778447393264251397636848807045177700727957761;
            6'd47: xpb[34] = 1024'd58656078272730048033992222209740724742086156599328118386018122492801337304048020404534005438049171362060236878007689220463012147242961334564187461236173675542987358369842449688415072889954524612305085910642833499768004233853276449352967210277782650701474690319475105057306490322926450058073655556647858385184;
            6'd48: xpb[34] = 1024'd25587759855264269520154055527765258764660765194323101890705441783186479812963535608243326281612988496938945273349397190057377726313325100209870564130298572211179030475489611907547455089959436319438543719187699786938883237703949181285057546541523072195789923211729431667219716394455263267340265935594988812607;
            6'd49: xpb[34] = 1024'd116586137121923232405114816250604225531933800915053769523524616138548517659188189721967718339834479941260803076148598594230807146224909200410713792040754509813061377150707991464310076481481553747882199136119805920474123091775518686182126452488492942956925059518100816307239470539912709493725566141167713724361;
            6'd50: xpb[34] = 1024'd83517818704457453891276649568628759554508409510048753028211935428933660168103704925677039183398297076139511471490306563825172725295272966056396894934879406481253049256355153683442458681486465455015656944664672207645002095626191418114216788752233364451240292410355142917152696611441522702992176520114844151784;
            6'd51: xpb[34] = 1024'd50449500286991675377438482886653293577083018105043736532899254719318802677019220129386360026962114211018219866832014533419538304365636731702079997829004303149444721362002315902574840881491377162149114753209538494815881099476864150046307125015973785945555525302609469527065922682970335912258786899061974579207;
            6'd52: xpb[34] = 1024'd17381181869525896863600316204677827599657626700038720037586574009703945185934735333095680870525931345896928262173722503013903883436000497347763100723129199817636393467649478121707223081496288869282572561754404781986760103327536881978397461279714207439870758194863796136979148754499149121525397278009105006630;
            6'd53: xpb[34] = 1024'd108379559136184859748561076927516794366930662420769387670405748365065983032159389446820072928747422790218786064972923907187333303347584597548606328633585137419518740142867857678469844473018406297726227978686510915521999957399106386875466367226684078201005894501235180776998902899956595347910697483581829918384;
            6'd54: xpb[34] = 1024'd75311240718719081234722910245541328389505271015764371175093067655451125541074904650529393772311239925097494460314631876781698882417948363194289431527710034087710412248515019897602226673023318004859685787231377202692878961249779118807556703490424499695321127393489507386912128971485408557177307862528960345807;
            6'd55: xpb[34] = 1024'd42242922301253302720884743563565862412079879610759354679780386945836268049990419854238714615875057059976202855656339846376064461488312128839972534421834930755902084354162182116734608873028229711993143595776243489863757965100451850739647039754164921189636360285743833996825355043014221766443918241476090773230;
            6'd56: xpb[34] = 1024'd9174603883787524207046576881590396434654488205754338184467706236221410558905935057948035459438874194854911250998047815970430040558675894485655637315959827424093756459809344335866991073033141419126601404321109777034636968951124582671737376017905342683951593177998160606738581114543034975710528620423221200653;
            6'd57: xpb[34] = 1024'd100172981150446487092007337604429363201927523926485005817286880591583448405130589171672427517660365639176769053797249220143859460470259994686498865226415765025976103135027723892629612464555258847570256821253215910569876823022694087568806281964875213445086729484369545246758335260000481202095828825995946112407;
            6'd58: xpb[34] = 1024'd67104662732980708578169170922453897224502132521479989321974199881968590914046104375381748361224182774055477449138957189738225039540623760332181968120540661694167775240674886111761994664560170554703714629798082197740755826873366819500896618228615634939401962376623871856671561331529294411362439204943076539830;
            6'd59: xpb[34] = 1024'd34036344315514930064331004240478431247076741116474972826661519172353733422961619579091069204787999908934185844480665159332590618610987525977865071014665558362359447346322048330894376864565082261837172438342948484911634830724039551432986954492356056433717195268878198466584787403058107620629049583890206967253;
            6'd60: xpb[34] = 1024'd968025898049151550492837558502965269651349711469956331348838462738875931877134782800390048351817043812894239822373128926956197681351291623548173908790455030551119451969210550026759064569993968970630246887814772082513834574712283365077290756096477928032428161132525076498013474586920829895659962837337394676;
            6'd61: xpb[34] = 1024'd91966403164708114435453598281341932036924385432200623964168012818100913778101788896524782106573308488134752042621574533100385617592935391824391401819246392632433466127187590106789380456092111397414285663819920905617753688646281788262146196703066348689167564467503909716517767620044367056280960168410062306430;
            6'd62: xpb[34] = 1024'd58898084747242335921615431599366466059498994027195607468855332108486056287017304100234102950137125623013460437963282502694751196663299157470074504713371289300625138232834752325921762656097023104547743472364787192788632692496954520194236532966806770183482797359758236326430993691573180265547570547357192733853;
            6'd63: xpb[34] = 1024'd25829766329776557407777264917391000082073602622190590973542651398871198795932819303943423793700942757892168833304990472289116775733662923115757607607496185968816810338481914545054144856101934811681201280909653479959511696347627252126326869230547191677798030252012562936344219763101993474814180926304323161276;
        endcase
    end

    always_comb begin
        case(flag[11][16:12])
            5'd0: xpb[35] = 1024'd0;
            5'd1: xpb[35] = 1024'd116828143596435520292738025640229966849346638342921258606361825754233236642157473417667815851922434202214026636104191876462546195645247023316600835517952123570699157013700294101816766247624052240124856697841759613494751550419196757023395775177517062438933166558383947576363973908559439701199481131877048073030;
            5'd2: xpb[35] = 1024'd109589591508746299186677123875645500953994849560106833084591796443489577947005807925320560489187194094984903864750890318346028550449273712078041546019573206207707639457829370866003293303730898758939515787296279380625142250617496741081812980671804675611046429702650837122621419743190246385280272437128501661729;
            5'd3: xpb[35] = 1024'd102351039421057078080616222111061035058643060777292407562821767132745919251854142432973305126451953987755781093397588760229510905253300400839482256521194288844716121901958447630189820359837745277754174876750799147755532950815796725140230186166092288783159692846917726668878865577821053069361063742379955250428;
            5'd4: xpb[35] = 1024'd95112487333367856974555320346476569163291271994477982041051737822002260556702476940626049763716713880526658322044287202112993260057327089600922967022815371481724604346087524394376347415944591796568833966205318914885923651014096709198647391660379901955272955991184616215136311412451859753441855047631408839127;
            5'd5: xpb[35] = 1024'd87873935245678635868494418581892103267939483211663556519281708511258601861550811448278794400981473773297535550690985643996475614861353778362363677524436454118733086790216601158562874472051438315383493055659838682016314351212396693257064597154667515127386219135451505761393757247082666437522646352882862427826;
            5'd6: xpb[35] = 1024'd80635383157989414762433516817307637372587694428849130997511679200514943166399145955931539038246233666068412779337684085879957969665380467123804388026057536755741569234345677922749401528158284834198152145114358449146705051410696677315481802648955128299499482279718395307651203081713473121603437658134316016525;
            5'd7: xpb[35] = 1024'd73396831070300193656372615052723171477235905646034705475741649889771284471247480463584283675510993558839290007984382527763440324469407155885245098527678619392750051678474754686935928584265131353012811234568878216277095751608996661373899008143242741471612745423985284853908648916344279805684228963385769605224;
            5'd8: xpb[35] = 1024'd66158278982610972550311713288138705581884116863220279953971620579027625776095814971237028312775753451610167236631080969646922679273433844646685809029299702029758534122603831451122455640371977871827470324023397983407486451807296645432316213637530354643726008568252174400166094750975086489765020268637223193923;
            5'd9: xpb[35] = 1024'd58919726894921751444250811523554239686532328080405854432201591268283967080944149478889772950040513344381044465277779411530405034077460533408126519530920784666767016566732908215308982696478824390642129413477917750537877152005596629490733419131817967815839271712519063946423540585605893173845811573888676782622;
            5'd10: xpb[35] = 1024'd51681174807232530338189909758969773791180539297591428910431561957540308385792483986542517587305273237151921693924477853413887388881487222169567230032541867303775499010861984979495509752585670909456788502932437517668267852203896613549150624626105580987952534856785953492680986420236699857926602879140130371321;
            5'd11: xpb[35] = 1024'd44442622719543309232129007994385307895828750514777003388661532646796649690640818494195262224570033129922798922571176295297369743685513910931007940534162949940783981454991061743682036808692517428271447592386957284798658552402196597607567830120393194160065798001052843038938432254867506542007394184391583960020;
            5'd12: xpb[35] = 1024'd37204070631854088126068106229800842000476961731962577866891503336052990995489153001848006861834793022693676151217874737180852098489540599692448651035784032577792463899120138507868563864799363947086106681841477051929049252600496581665985035614680807332179061145319732585195878089498313226088185489643037548719;
            5'd13: xpb[35] = 1024'd29965518544164867020007204465216376105125172949148152345121474025309332300337487509500751499099552915464553379864573179064334453293567288453889361537405115214800946343249215272055090920906210465900765771295996819059439952798796565724402241108968420504292324289586622131453323924129119910168976794894491137418;
            5'd14: xpb[35] = 1024'd22726966456475645913946302700631910209773384166333726823351444714565673605185822017153496136364312808235430608511271620947816808097593977215330072039026197851809428787378292036241617977013056984715424860750516586189830652997096549782819446603256033676405587433853511677710769758759926594249768100145944726117;
            5'd15: xpb[35] = 1024'd15488414368786424807885400936047444314421595383519301301581415403822014910034156524806240773629072701006307837157970062831299162901620665976770782540647280488817911231507368800428145033119903503530083950205036353320221353195396533841236652097543646848518850578120401223968215593390733278330559405397398314816;
            5'd16: xpb[35] = 1024'd8249862281097203701824499171462978419069806600704875779811386093078356214882491032458985410893832593777185065804668504714781517705647354738211493042268363125826393675636445564614672089226750022344743039659556120450612053393696517899653857591831260020632113722387290770225661428021539962411350710648851903515;
            5'd17: xpb[35] = 1024'd1011310193407982595763597406878512523718017817890450258041356782334697519730825540111730048158592486548062294451366946598263872509674043499652203543889445762834876119765522328801199145333596541159402129114075887581002753591996501958071063086118873192745376866654180316483107262652346646492142015900305492214;
            5'd18: xpb[35] = 1024'd117839453789843502888501623047108479373064656160811708864403182536567934161888298957779545900081026688762088930555558823060810068154921066816253039061841569333534033133465816430617965392957648781284258826955835501075754304011193258981466838263635935631678543425038127892847081171211786347691623147777353565244;
            5'd19: xpb[35] = 1024'd110600901702154281782440721282524013477712867377997283342633153225824275466736633465432290537345786581532966159202257264944292422958947755577693749563462651970542515577594893194804492449064495300098917916410355268206145004209493243039884043757923548803791806569305017439104527005842593031772414453028807153943;
            5'd20: xpb[35] = 1024'd103362349614465060676379819517939547582361078595182857820863123915080616771584967973085035174610546474303843387848955706827774777762974444339134460065083734607550998021723969958991019505171341818913577005864875035336535704407793227098301249252211161975905069713571906985361972840473399715853205758280260742642;
            5'd21: xpb[35] = 1024'd96123797526775839570318917753355081687009289812368432299093094604336958076433302480737779811875306367074720616495654148711257132567001133100575170566704817244559480465853046723177546561278188337728236095319394802466926404606093211156718454746498775148018332857838796531619418675104206399933997063531714331341;
            5'd22: xpb[35] = 1024'd88885245439086618464258015988770615791657501029554006777323065293593299381281636988390524449140066259845597845142352590594739487371027821862015881068325899881567962909982123487364073617385034856542895184773914569597317104804393195215135660240786388320131596002105686077876864509735013084014788368783167920040;
            5'd23: xpb[35] = 1024'd81646693351397397358197114224186149896305712246739581255553035982849640686129971496043269086404826152616475073789051032478221842175054510623456591569946982518576445354111200251550600673491881375357554274228434336727707805002693179273552865735074001492244859146372575624134310344365819768095579674034621508739;
            5'd24: xpb[35] = 1024'd74408141263708176252136212459601684000953923463925155733783006672105981990978306003696013723669586045387352302435749474361704196979081199384897302071568065155584927798240277015737127729598727894172213363682954103858098505200993163331970071229361614664358122290639465170391756178996626452176370979286075097438;
            5'd25: xpb[35] = 1024'd67169589176018955146075310695017218105602134681110730212012977361362323295826640511348758360934345938158229531082447916245186551783107888146338012573189147792593410242369353779923654785705574412986872453137473870988489205399293147390387276723649227836471385434906354716649202013627433136257162284537528686137;
            5'd26: xpb[35] = 1024'd59931037088329734040014408930432752210250345898296304690242948050618664600674975019001502998199105830929106759729146358128668906587134576907778723074810230429601892686498430544110181841812420931801531542591993638118879905597593131448804482217936841008584648579173244262906647848258239820337953589788982274836;
            5'd27: xpb[35] = 1024'd52692485000640512933953507165848286314898557115481879168472918739875005905523309526654247635463865723699983988375844800012151261391161265669219433576431313066610375130627507308296708897919267450616190632046513405249270605795893115507221687712224454180697911723440133809164093682889046504418744895040435863535;
            5'd28: xpb[35] = 1024'd45453932912951291827892605401263820419546768332667453646702889429131347210371644034306992272728625616470861217022543241895633616195187954430660144078052395703618857574756584072483235954026113969430849721501033172379661305994193099565638893206512067352811174867707023355421539517519853188499536200291889452234;
            5'd29: xpb[35] = 1024'd38215380825262070721831703636679354524194979549853028124932860118387688515219978541959736909993385509241738445669241683779115970999214643192100854579673478340627340018885660836669763010132960488245508810955552939510052006192493083624056098700799680524924438011973912901678985352150659872580327505543343040933;
            5'd30: xpb[35] = 1024'd30976828737572849615770801872094888628843190767038602603162830807644029820068313049612481547258145402012615674315940125662598325803241331953541565081294560977635822463014737600856290066239807007060167900410072706640442706390793067682473304195087293697037701156240802447936431186781466556661118810794796629632;
            5'd31: xpb[35] = 1024'd23738276649883628509709900107510422733491401984224177081392801496900371124916647557265226184522905294783492902962638567546080680607268020714982275582915643614644304907143814365042817122346653525874826989864592473770833406589093051740890509689374906869150964300507691994193877021412273240741910116046250218331;
        endcase
    end

    always_comb begin
        case(flag[12][5:0])
            6'd0: xpb[36] = 1024'd0;
            6'd1: xpb[36] = 1024'd8249862281097203701824499171462978419069806600704875779811386093078356214882491032458985410893832593777185065804668504714781517705647354738211493042268363125826393675636445564614672089226750022344743039659556120450612053393696517899653857591831260020632113722387290770225661428021539962411350710648851903515;
            6'd2: xpb[36] = 1024'd16499724562194407403648998342925956838139613201409751559622772186156712429764982064917970821787665187554370131609337009429563035411294709476422986084536726251652787351272891129229344178453500044689486079319112240901224106787393035799307715183662520041264227444774581540451322856043079924822701421297703807030;
            6'd3: xpb[36] = 1024'd24749586843291611105473497514388935257209419802114627339434158279235068644647473097376956232681497781331555197414005514144344553116942064214634479126805089377479181026909336693844016267680250067034229118978668361351836160181089553698961572775493780061896341167161872310676984284064619887234052131946555710545;
            6'd4: xpb[36] = 1024'd32999449124388814807297996685851913676279226402819503119245544372313424859529964129835941643575330375108740263218674018859126070822589418952845972169073452503305574702545782258458688356907000089378972158638224481802448213574786071598615430367325040082528454889549163080902645712086159849645402842595407614060;
            6'd5: xpb[36] = 1024'd41249311405486018509122495857314892095349033003524378899056930465391781074412455162294927054469162968885925329023342523573907588528236773691057465211341815629131968378182227823073360446133750111723715198297780602253060266968482589498269287959156300103160568611936453851128307140107699812056753553244259517575;
            6'd6: xpb[36] = 1024'd49499173686583222210946995028777870514418839604229254678868316558470137289294946194753912465362995562663110394828011028288689106233884128429268958253610178754958362053818673387688032535360500134068458237957336722703672320362179107397923145550987560123792682334323744621353968568129239774468104263893111421090;
            6'd7: xpb[36] = 1024'd57749035967680425912771494200240848933488646204934130458679702651548493504177437227212897876256828156440295460632679533003470623939531483167480451295878541880784755729455118952302704624587250156413201277616892843154284373755875625297577003142818820144424796056711035391579629996150779736879454974541963324605;
            6'd8: xpb[36] = 1024'd65998898248777629614595993371703827352558452805639006238491088744626849719059928259671883287150660750217480526437348037718252141645178837905691944338146905006611149405091564516917376713814000178757944317276448963604896427149572143197230860734650080165056909779098326161805291424172319699290805685190815228120;
            6'd9: xpb[36] = 1024'd74248760529874833316420492543166805771628259406343882018302474837705205933942419292130868698044493343994665592242016542433033659350826192643903437380415268132437543080728010081532048803040750201102687356936005084055508480543268661096884718326481340185689023501485616932030952852193859661702156395839667131635;
            6'd10: xpb[36] = 1024'd82498622810972037018244991714629784190698066007048757798113860930783562148824910324589854108938325937771850658046685047147815177056473547382114930422683631258263936756364455646146720892267500223447430396595561204506120533936965178996538575918312600206321137223872907702256614280215399624113507106488519035150;
            6'd11: xpb[36] = 1024'd90748485092069240720069490886092762609767872607753633577925247023861918363707401357048839519832158531549035723851353551862596694762120902120326423464951994384090330432000901210761392981494250245792173436255117324956732587330661696896192433510143860226953250946260198472482275708236939586524857817137370938665;
            6'd12: xpb[36] = 1024'd98998347373166444421893990057555741028837679208458509357736633116940274578589892389507824930725991125326220789656022056577378212467768256858537916507220357509916724107637346775376065070721000268136916475914673445407344640724358214795846291101975120247585364668647489242707937136258479548936208527786222842180;
            6'd13: xpb[36] = 1024'd107248209654263648123718489229018719447907485809163385137548019210018630793472383421966810341619823719103405855460690561292159730173415611596749409549488720635743117783273792339990737159947750290481659515574229565857956694118054732695500148693806380268217478391034780012933598564280019511347559238435074745695;
            6'd14: xpb[36] = 1024'd115498071935360851825542988400481697866977292409868260917359405303096987008354874454425795752513656312880590921265359066006941247879062966334960902591757083761569511458910237904605409249174500312826402555233785686308568747511751250595154006285637640288849592113422070783159259992301559473758909949083926649210;
            6'd15: xpb[36] = 1024'd123747934216458055527367487571944676286047099010573136697170791396175343223237365486884781163407488906657775987070027570721722765584710321073172395634025446887395905134546683469220081338401250335171145594893341806759180800905447768494807863877468900309481705835809361553384921420323099436170260659732778552725;
            6'd16: xpb[36] = 1024'd7931100813430517830393059338593221960418478485542328348850322424276804100810717609328695359643647190991811645417202640857440442449137341256223763659962769079531624240611911696204514236110794636205691026165658080845432004078247513429483151786070711063293916144079594293504054774416006381462921543756035971909;
            6'd17: xpb[36] = 1024'd16180963094527721532217558510056200379488285086247204128661708517355160315693208641787680770537479784768996711221871145572221960154784695994435256702231132205358017916248357260819186325337544658550434065825214201296044057471944031329137009377901971083926029866466885063729716202437546343874272254404887875424;
            6'd18: xpb[36] = 1024'd24430825375624925234042057681519178798558091686952079908473094610433516530575699674246666181431312378546181777026539650287003477860432050732646749744499495331184411591884802825433858414564294680895177105484770321746656110865640549228790866969733231104558143588854175833955377630459086306285622965053739778939;
            6'd19: xpb[36] = 1024'd32680687656722128935866556852982157217627898287656955688284480703511872745458190706705651592325144972323366842831208155001784995566079405470858242786767858457010805267521248390048530503791044703239920145144326442197268164259337067128444724561564491125190257311241466604181039058480626268696973675702591682454;
            6'd20: xpb[36] = 1024'd40930549937819332637691056024445135636697704888361831468095866796590228960340681739164637003218977566100551908635876659716566513271726760209069735829036221582837198943157693954663202593017794725584663184803882562647880217653033585028098582153395751145822371033628757374406700486502166231108324386351443585969;
            6'd21: xpb[36] = 1024'd49180412218916536339515555195908114055767511489066707247907252889668585175223172771623622414112810159877736974440545164431348030977374114947281228871304584708663592618794139519277874682244544747929406224463438683098492271046730102927752439745227011166454484756016048144632361914523706193519675097000295489484;
            6'd22: xpb[36] = 1024'd57430274500013740041340054367371092474837318089771583027718638982746941390105663804082607825006642753654922040245213669146129548683021469685492721913572947834489986294430585083892546771471294770274149264122994803549104324440426620827406297337058271187086598478403338914858023342545246155931025807649147392999;
            6'd23: xpb[36] = 1024'd65680136781110943743164553538834070893907124690476458807530025075825297604988154836541593235900475347432107106049882173860911066388668824423704214955841310960316379970067030648507218860698044792618892303782550923999716377834123138727060154928889531207718712200790629685083684770566786118342376518297999296514;
            6'd24: xpb[36] = 1024'd73929999062208147444989052710297049312976931291181334587341411168903653819870645869000578646794307941209292171854550678575692584094316179161915707998109674086142773645703476213121890949924794814963635343442107044450328431227819656626714012520720791228350825923177920455309346198588326080753727228946851200029;
            6'd25: xpb[36] = 1024'd82179861343305351146813551881760027732046737891886210367152797261982010034753136901459564057688140534986477237659219183290474101799963533900127201040378037211969167321339921777736563039151544837308378383101663164900940484621516174526367870112552051248982939645565211225535007626609866043165077939595703103544;
            6'd26: xpb[36] = 1024'd90429723624402554848638051053223006151116544492591086146964183355060366249635627933918549468581973128763662303463887688005255619505610888638338694082646400337795560996976367342351235128378294859653121422761219285351552538015212692426021727704383311269615053367952501995760669054631406005576428650244555007059;
            6'd27: xpb[36] = 1024'd98679585905499758550462550224685984570186351093295961926775569448138722464518118966377534879475805722540847369268556192720037137211258243376550187124914763463621954672612812906965907217605044881997864462420775405802164591408909210325675585296214571290247167090339792765986330482652945967987779360893406910574;
            6'd28: xpb[36] = 1024'd106929448186596962252287049396148962989256157694000837706586955541217078679400609998836520290369638316318032435073224697434818654916905598114761680167183126589448348348249258471580579306831794904342607502080331526252776644802605728225329442888045831310879280812727083536211991910674485930399130071542258814089;
            6'd29: xpb[36] = 1024'd115179310467694165954111548567611941408325964294705713486398341634295434894283101031295505701263470910095217500877893202149600172622552952852973173209451489715274742023885704036195251396058544926687350541739887646703388698196302246124983300479877091331511394535114374306437653338696025892810480782191110717604;
            6'd30: xpb[36] = 1024'd123429172748791369655936047739074919827395770895410589266209727727373791109165592063754491112157303503872402566682561706864381690328200307591184666251719852841101135699522149600809923485285294949032093581399443767154000751589998764024637158071708351352143508257501665076663314766717565855221831492839962621119;
            6'd31: xpb[36] = 1024'd7612339345763831958961619505723465501767150370379780917889258755475251986738944186198405308393461788206438225029736777000099367192627327774236034277657175033236854805587377827794356382994839250066639012671760041240251954762798508959312445980310162105955718565771897816782448120810472800514492376863220040303;
            6'd32: xpb[36] = 1024'd15862201626861035660786118677186443920836956971084656697700644848553608201621435218657390719287294381983623290834405281714880884898274682512447527319925538159063248481223823392409028472221589272411382052331316161690864008156495026858966303572141422126587832288159188587008109548832012762925843087512071943818;
            6'd33: xpb[36] = 1024'd24112063907958239362610617848649422339906763571789532477512030941631964416503926251116376130181126975760808356639073786429662402603922037250659020362193901284889642156860268957023700561448339294756125091990872282141476061550191544758620161163972682147219946010546479357233770976853552725337193798160923847333;
            6'd34: xpb[36] = 1024'd32361926189055443064435117020112400758976570172494408257323417034710320631386417283575361541074959569537993422443742291144443920309569391988870513404462264410716035832496714521638372650675089317100868131650428402592088114943888062658274018755803942167852059732933770127459432404875092687748544508809775750848;
            6'd35: xpb[36] = 1024'd40611788470152646766259616191575379178046376773199284037134803127788676846268908316034346951968792163315178488248410795859225438015216746727082006446730627536542429508133160086253044739901839339445611171309984523042700168337584580557927876347635202188484173455321060897685093832896632650159895219458627654363;
            6'd36: xpb[36] = 1024'd48861650751249850468084115363038357597116183373904159816946189220867033061151399348493332362862624757092363554053079300574006955720864101465293499488998990662368823183769605650867716829128589361790354210969540643493312221731281098457581733939466462209116287177708351667910755260918172612571245930107479557878;
            6'd37: xpb[36] = 1024'd57111513032347054169908614534501336016185989974609035596757575313945389276033890380952317773756457350869548619857747805288788473426511456203504992531267353788195216859406051215482388918355339384135097250629096763943924275124977616357235591531297722229748400900095642438136416688939712574982596640756331461393;
            6'd38: xpb[36] = 1024'd65361375313444257871733113705964314435255796575313911376568961407023745490916381413411303184650289944646733685662416310003569991132158810941716485573535716914021610535042496780097061007582089406479840290288652884394536328518674134256889449123128982250380514622482933208362078116961252537393947351405183364908;
            6'd39: xpb[36] = 1024'd73611237594541461573557612877427292854325603176018787156380347500102101705798872445870288595544122538423918751467084814718351508837806165679927978615804080039848004210678942344711733096808839428824583329948209004845148381912370652156543306714960242271012628344870223978587739544982792499805298062054035268423;
            6'd40: xpb[36] = 1024'd81861099875638665275382112048890271273395409776723662936191733593180457920681363478329274006437955132201103817271753319433133026543453520418139471658072443165674397886315387909326405186035589451169326369607765125295760435306067170056197164306791502291644742067257514748813400973004332462216648772702887171938;
            6'd41: xpb[36] = 1024'd90110962156735868977206611220353249692465216377428538716003119686258814135563854510788259417331787725978288883076421824147914544249100875156350964700340806291500791561951833473941077275262339473514069409267321245746372488699763687955851021898622762312276855789644805519039062401025872424627999483351739075453;
            6'd42: xpb[36] = 1024'd98360824437833072679031110391816228111535022978133414495814505779337170350446345543247244828225620319755473948881090328862696061954748229894562457742609169417327185237588279038555749364489089495858812448926877366196984542093460205855504879490454022332908969512032096289264723829047412387039350194000590978968;
            6'd43: xpb[36] = 1024'd106610686718930276380855609563279206530604829578838290275625891872415526565328836575706230239119452913532659014685758833577477579660395584632773950784877532543153578913224724603170421453715839518203555488586433486647596595487156723755158737082285282353541083234419387059490385257068952349450700904649442882483;
            6'd44: xpb[36] = 1024'd114860549000027480082680108734742184949674636179543166055437277965493882780211327608165215650013285507309844080490427338292259097366042939370985443827145895668979972588861170167785093542942589540548298528245989607098208648880853241654812594674116542374173196956806677829716046685090492311862051615298294785998;
            6'd45: xpb[36] = 1024'd123110411281124683784504607906205163368744442780248041835248664058572238995093818640624201060907118101087029146295095843007040615071690294109196936869414258794806366264497615732399765632169339562893041567905545727548820702274549759554466452265947802394805310679193968599941708113112032274273402325947146689513;
            6'd46: xpb[36] = 1024'd7293577878097146087530179672853709043115822255217233486928195086673699872667170763068115257143276385421064804642270913142758291936117314292248304895351580986942085370562843959384198529878883863927586999177862001635071905447349504489141740174549613148617520987464201340060841467204939219566063209970404108697;
            6'd47: xpb[36] = 1024'd15543440159194349789354678844316687462185628855922109266739581179752056087549661795527100668037108979198249870446939417857539809641764669030459797937619944112768479046199289523998870619105633886272330038837418122085683958841046022388795597766380873169249634709851492110286502895226479181977413920619256012212;
            6'd48: xpb[36] = 1024'd23793302440291553491179178015779665881255435456626985046550967272830412302432152827986086078930941572975434936251607922572321327347412023768671290979888307238594872721835735088613542708332383908617073078496974242536296012234742540288449455358212133189881748432238782880512164323248019144388764631268107915727;
            6'd49: xpb[36] = 1024'd32043164721388757193003677187242644300325242057331860826362353365908768517314643860445071489824774166752620002056276427287102845053059378506882784022156670364421266397472180653228214797559133930961816118156530362986908065628439058188103312950043393210513862154626073650737825751269559106800115341916959819242;
            6'd50: xpb[36] = 1024'd40293027002485960894828176358705622719395048658036736606173739458987124732197134892904056900718606760529805067860944932001884362758706733245094277064425033490247660073108626217842886886785883953306559157816086483437520119022135576087757170541874653231145975877013364420963487179291099069211466052565811722757;
            6'd51: xpb[36] = 1024'd48542889283583164596652675530168601138464855258741612385985125552065480947079625925363042311612439354306990133665613436716665880464354087983305770106693396616074053748745071782457558976012633975651302197475642603888132172415832093987411028133705913251778089599400655191189148607312639031622816763214663626272;
            6'd52: xpb[36] = 1024'd56792751564680368298477174701631579557534661859446488165796511645143837161962116957822027722506271948084175199470281941431447398170001442721517263148961759741900447424381517347072231065239383997996045237135198724338744225809528611887064885725537173272410203321787945961414810035334178994034167473863515529787;
            6'd53: xpb[36] = 1024'd65042613845777572000301673873094557976604468460151363945607897738222193376844607990281013133400104541861360265274950446146228915875648797459728756191230122867726841100017962911686903154466134020340788276794754844789356279203225129786718743317368433293042317044175236731640471463355718956445518184512367433302;
            6'd54: xpb[36] = 1024'd73292476126874775702126173044557536395674275060856239725419283831300549591727099022739998544293937135638545331079618950861010433581296152197940249233498485993553234775654408476301575243692884042685531316454310965239968332596921647686372600909199693313674430766562527501866132891377258918856868895161219336817;
            6'd55: xpb[36] = 1024'd81542338407971979403950672216020514814744081661561115505230669924378905806609590055198983955187769729415730396884287455575791951286943506936151742275766849119379628451290854040916247332919634065030274356113867085690580385990618165586026458501030953334306544488949818272091794319398798881268219605810071240332;
            6'd56: xpb[36] = 1024'd89792200689069183105775171387483493233813888262265991285042056017457262021492081087657969366081602323192915462688955960290573468992590861674363235318035212245206022126927299605530919422146384087375017395773423206141192439384314683485680316092862213354938658211337109042317455747420338843679570316458923143847;
            6'd57: xpb[36] = 1024'd98042062970166386807599670558946471652883694862970867064853442110535618236374572120116954776975434916970100528493624465005354986698238216412574728360303575371032415802563745170145591511373134109719760435432979326591804492778011201385334173684693473375570771933724399812543117175441878806090921027107775047362;
            6'd58: xpb[36] = 1024'd106291925251263590509424169730409450071953501463675742844664828203613974451257063152575940187869267510747285594298292969720136504403885571150786221402571938496858809478200190734760263600599884132064503475092535447042416546171707719284988031276524733396202885656111690582768778603463418768502271737756626950877;
            6'd59: xpb[36] = 1024'd114541787532360794211248668901872428491023308064380618624476214296692330666139554185034925598763100104524470660102961474434918022109532925888997714444840301622685203153836636299374935689826634154409246514752091567493028599565404237184641888868355993416834999378498981352994440031484958730913622448405478854392;
            6'd60: xpb[36] = 1024'd122791649813457997913073168073335406910093114665085494404287600389770686881022045217493911009656932698301655725907629979149699539815180280627209207487108664748511596829473081863989607779053384176753989554411647687943640652959100755084295746460187253437467113100886272123220101459506498693324973159054330757907;
            6'd61: xpb[36] = 1024'd6974816410430460216098739839983952584464494140054686055967131417872147758595397339937825205893090982635691384254805049285417216679607300810260575513045986940647315935538310090974040676762928477788534985683963962029891856131900500018971034368789064191279323409156504863339234813599405638617634043077588177091;
            6'd62: xpb[36] = 1024'd15224678691527663917923239011446931003534300740759561835778517510950503973477888372396810616786923576412876450059473554000198734385254655548472068555314350066473709611174755655588712765989678500133278025343520082480503909525597017918624891960620324211911437131543795633564896241620945601028984753726440080606;
            6'd63: xpb[36] = 1024'd23474540972624867619747738182909909422604107341464437615589903604028860188360379404855796027680756170190061515864142058714980252090902010286683561597582713192300103286811201220203384855216428522478021065003076202931115962919293535818278749552451584232543550853931086403790557669642485563440335464375291984121;
        endcase
    end

    always_comb begin
        case(flag[12][11:6])
            6'd0: xpb[37] = 1024'd0;
            6'd1: xpb[37] = 1024'd31724403253722071321572237354372887841673913942169313395401289697107216403242870437314781438574588763967246581668810563429761769796549365024895054639851076318126496962447646784818056944443178544822764104662632323381728016312990053717932607144282844253175664576318377174016219097664025525851686175024143887636;
            6'd2: xpb[37] = 1024'd63448806507444142643144474708745775683347827884338626790802579394214432806485740874629562877149177527934493163337621126859523539593098730049790109279702152636252993924895293569636113888886357089645528209325264646763456032625980107435865214288565688506351329152636754348032438195328051051703372350048287775272;
            6'd3: xpb[37] = 1024'd95173209761166213964716712063118663525021741826507940186203869091321649209728611311944344315723766291901739745006431690289285309389648095074685163919553228954379490887342940354454170833329535634468292313987896970145184048938970161153797821432848532759526993728955131522048657292992076577555058525072431662908;
            6'd4: xpb[37] = 1024'd2830917330763543887490022012677118621997228642941569453473303723451970275662342839244054539640680746425836919217748819139983238344977125544420093543073264338815313280219369801641988586255508457980858810263289447162551215031063441906751858893901927745882754891156450665958348316727469086288054873470981066213;
            6'd5: xpb[37] = 1024'd34555320584485615209062259367050006463671142585110882848874593420559186678905213276558835978215269510393083500886559382569745008141526490569315148182924340656941810242667016586460045530698687002803622914925921770544279231344053495624684466038184771999058419467474827839974567414391494612139741048495124953849;
            6'd6: xpb[37] = 1024'd66279723838207686530634496721422894305345056527280196244275883117666403082148083713873617416789858274360330082555369945999506777938075855594210202822775416975068307205114663371278102475141865547626387019588554093926007247657043549342617073182467616252234084043793205013990786512055520137991427223519268841485;
            6'd7: xpb[37] = 1024'd98004127091929757852206734075795782147018970469449509639677172814773619485390954151188398855364447038327576664224180509429268547734625220619105257462626493293194804167562310156096159419585044092449151124251186417307735263970033603060549680326750460505409748620111582188007005609719545663843113398543412729121;
            6'd8: xpb[37] = 1024'd5661834661527087774980044025354237243994457285883138906946607446903940551324685678488109079281361492851673838435497638279966476689954251088840187086146528677630626560438739603283977172511016915961717620526578894325102430062126883813503717787803855491765509782312901331916696633454938172576109746941962132426;
            6'd9: xpb[37] = 1024'd37386237915249159096552281379727125085668371228052452302347897144011156954567556115802890517855950256818920420104308201709728246486503616113735241725997604995757123522886386388102034116954195460784481725189211217706830446375116937531436324932086699744941174358631278505932915731118963698427795921966106020062;
            6'd10: xpb[37] = 1024'd69110641168971230418124518734100012927342285170221765697749186841118373357810426553117671956430539020786167001773118765139490016283052981138630296365848681313883620485334033172920091061397374005607245829851843541088558462688106991249368932076369543998116838934949655679949134828782989224279482096990249907698;
            6'd11: xpb[37] = 1024'd100835044422693301739696756088472900769016199112391079093150476538225589761053296990432453395005127784753413583441929328569251786079602346163525351005699757632010117447781679957738148005840552550430009934514475864470286479001097044967301539220652388251292503511268032853965353926447014750131168272014393795334;
            6'd12: xpb[37] = 1024'd8492751992290631662470066038031355865991685928824708360419911170355910826987028517732163618922042239277510757653246457419949715034931376633260280629219793016445939840658109404925965758766525373942576430789868341487653645093190325720255576681705783237648264673469351997875044950182407258864164620412943198639;
            6'd13: xpb[37] = 1024'd40217155246012702984042303392404243707665599870994021755821200867463127230229898955046945057496631003244757339322057020849711484831480741658155335269070869334572436803105756189744022703209703918765340535452500664869381661406180379438188183825988627490823929249787729171891264047846432784715850795437087086275;
            6'd14: xpb[37] = 1024'd71941558499734774305614540746777131549339513813163335151222490564570343633472769392361726496071219767212003920990867584279473254628030106683050389908921945652698933765553402974562079647652882463588104640115132988251109677719170433156120790970271471743999593826106106345907483145510458310567536970461230973911;
            6'd15: xpb[37] = 1024'd103665961753456845627186778101150019391013427755332648546623780261677560036715639829676507934645808531179250502659678147709235024424579471707945444548773021970825430728001049759380136592096061008410868744777765311632837694032160486874053398114554315997175258402424483519923702243174483836419223145485374861547;
            6'd16: xpb[37] = 1024'd11323669323054175549960088050708474487988914571766277813893214893807881102649371356976218158562722985703347676870995276559932953379908502177680374172293057355261253120877479206567954345022033831923435241053157788650204860124253767627007435575607710983531019564625802663833393266909876345152219493883924264852;
            6'd17: xpb[37] = 1024'd43048072576776246871532325405081362329662828513935591209294504590915097505892241794290999597137311749670594258539805839989694723176457867202575428812144133673387750083325125991386011289465212376746199345715790112031932876437243821344940042719890555236706684140944179837849612364573901871003905668908068152488;
            6'd18: xpb[37] = 1024'd74772475830498318193104562759454250171336742456104904604695794288022313909135112231605781035711900513637840840208616403419456492973007232227470483451995209991514247045772772776204068233908390921568963450378422435413660892750233875062872649864173399489882348717262557011865831462237927396855591843932212040124;
            6'd19: xpb[37] = 1024'd106496879084220389514676800113827138013010656398274218000097083985129530312377982668920562474286489277605087421877426966849218262769556597252365538091846286309640744008220419561022125178351569466391727555041054758795388909063223928780805257008456243743058013293580934185882050559901952922707278018956355927760;
            6'd20: xpb[37] = 1024'd14154586653817719437450110063385593109986143214707847267366518617259851378311714196220272698203403732129184596088744095699916191724885627722100467715366321694076566401096849008209942931277542289904294051316447235812756075155317209533759294469509638729413774455782253329791741583637345431440274367354905331065;
            6'd21: xpb[37] = 1024'd45878989907539790759022347417758480951660057156877160662767808314367067781554584633535054136777992496096431177757554659129677961521434992746995522355217398012203063363544495793027999875720720834727058155979079559194484091468307263251691901613792482982589439032100630503807960681301370957291960542379049218701;
            6'd22: xpb[37] = 1024'd77603393161261862080594584772131368793333971099046474058169098011474284184797455070849835575352581260063677759426365222559439731317984357771890576995068474330329560325992142577846056820163899379549822260641711882576212107781297316969624508758075327235765103608419007677824179778965396483143646717403193106337;
            6'd23: xpb[37] = 1024'd109327796414983933402166822126504256635007885041215787453570387708581500588040325508164617013927170024030924341095175785989201501114533722796785631634919550648456057288439789362664113764607077924372586365304344205957940124094287370687557115902358171488940768184737384851840398876629422008995332892427336993973;
            6'd24: xpb[37] = 1024'd16985503984581263324940132076062711731983371857649416720839822340711821653974057035464327237844084478555021515306492914839899430069862753266520561258439586032891879681316218809851931517533050747885152861579736682975307290186380651440511153363411566475296529346938703995750089900364814517728329240825886397278;
            6'd25: xpb[37] = 1024'd48709907238303334646512369430435599573657285799818730116241112037819038057216927472779108676418673242522268096975303478269661199866412118291415615898290662351018376643763865594669988461976229292707916966242369006357035306499370705158443760507694410728472193923257081169766308998028840043580015415850030284914;
            6'd26: xpb[37] = 1024'd80434310492025405968084606784808487415331199741988043511642401734926254460459797910093890114993262006489514678644114041699422969662961483316310670538141738669144873606211512379488045406419407837530681070905001329738763322812360758876376367651977254981647858499575458343782528095692865569431701590874174172550;
            6'd27: xpb[37] = 1024'd112158713745747477289656844139181375257005113684157356907043691432033470863702668347408671553567850770456761260312924605129184739459510848341205725177992814987271370568659159164306102350862586382353445175567633653120491339125350812594308974796260099234823523075893835517798747193356891095283387765898318060186;
            6'd28: xpb[37] = 1024'd19816421315344807212430154088739830353980600500590986174313126064163791929636399874708381777484765224980858434524241733979882668414839878810940654801512850371707192961535588611493920103788559205866011671843026130137858505217444093347263012257313494221179284238095154661708438217092283604016384114296867463491;
            6'd29: xpb[37] = 1024'd51540824569066878534002391443112718195654514442760299569714415761271008332879270312023163216059353988948105016193052297409644438211389243835835709441363926689833689923983235396311977048231737750688775776505658453519586521530434147065195619401596338474354948814413531835724657314756309129868070289321011351127;
            6'd30: xpb[37] = 1024'd83265227822788949855574628797485606037328428384929612965115705458378224736122140749337944654633942752915351597861862860839406208007938608860730764081215003007960186886430882181130033992674916295511539881168290776901314537843424200783128226545879182727530613390731909009740876412420334655719756464345155238763;
            6'd31: xpb[37] = 1024'd114989631076511021177146866151858493879002342327098926360516995155485441139365011186652726093208531516882598179530673424269167977804487973885625818721066079326086683848878528965948090937118094840334303985830923100283042554156414254501060833690162026980706277967050286183757095510084360181571442639369299126399;
            6'd32: xpb[37] = 1024'd22647338646108351099920176101416948975977829143532555627786429787615762205298742713952436317125445971406695353741990553119865906759817004355360748344586114710522506241754958413135908690044067663846870482106315577300409720248507535254014871151215421967062039129251605327666786533819752690304438987767848529704;
            6'd33: xpb[37] = 1024'd54371741899830422421492413455789836817651743085701869023187719484722978608541613151267217755700034735373941935410801116549627676556366369380255802984437191028649003204202605197953965634487246208669634586768947900682137736561497588971947478295498266220237703705569982501683005631483778216156125162791992417340;
            6'd34: xpb[37] = 1024'd86096145153552493743064650810162724659325657027871182418589009181830195011784483588581999194274623499341188517079611679979389446352915734405150857624288267346775500166650251982772022578930424753492398691431580224063865752874487642689880085439781110473413368281888359675699224729147803742007811337816136304976;
            6'd35: xpb[37] = 1024'd117820548407274565064636888164535612500999570970040495813990298878937411415027354025896780632849212263308435098748422243409151216149465099430045912264139343664901997129097898767590079523373603298315162796094212547445593769187477696407812692584063954726589032858206736849715443826811829267859497512840280192612;
            6'd36: xpb[37] = 1024'd25478255976871894987410198114094067597975057786474125081259733511067732480961085553196490856766126717832532272959739372259849145104794129899780841887659379049337819521974328214777897276299576121827729292369605024462960935279570977160766730045117349712944794020408055993625134850547221776592493861238829595917;
            6'd37: xpb[37] = 1024'd57202659230593966308982435468466955439648971728643438476661023208174948884203955990511272295340715481799778854628549935689610914901343494924675896527510455367464316484421974999595954220742754666650493397032237347844688951592561030878699337189400193966120458596726433167641353948211247302444180036262973483553;
            6'd38: xpb[37] = 1024'd88927062484316037630554672822839843281322885670812751872062312905282165287446826427826053733915304245767025436297360499119372684697892859949570951167361531685590813446869621784414011165185933211473257501694869671226416967905551084596631944333683038219296123173044810341657573045875272828295866211287117371189;
            6'd39: xpb[37] = 1024'd120651465738038108952126910177212731122996799612982065267463602602389381690689696865140835172489893009734272017966171062549134454494442224974466005807212608003717310409317268569232068109629111756296021606357501994608144984218541138314564551477965882472471787749363187515673792143539298354147552386311261258825;
            6'd40: xpb[37] = 1024'd28309173307635438874900220126771186219972286429415694534733037234519702756623428392440545396406807464258369192177488191399832383449771255444200935430732643388153132802193698016419885862555084579808588102632894471625512150310634419067518588939019277458827548911564506659583483167274690862880548734709810662130;
            6'd41: xpb[37] = 1024'd60033576561357510196472457481144074061646200371585007930134326931626919159866298829755326834981396228225615773846298754829594153246320620469095990070583719706279629764641344801237942806998263124631352207295526795007240166623624472785451196083302121712003213487882883833599702264938716388732234909733954549766;
            6'd42: xpb[37] = 1024'd91757979815079581518044694835516961903320114313754321325535616628734135563109169267070108273555984992192862355515109318259355923042869985493991044710434796024406126727088991586055999751441441669454116311958159118388968182936614526503383803227584965965178878064201261007615921362602741914583921084758098437402;
            6'd43: xpb[37] = 1024'd123482383068801652839616932189889849744994028255923634720936906325841351966352039704384889712130573756160108937183919881689117692839419350518886099350285872342532623689536638370874056695884620214276880416620791441770696199249604580221316410371867810218354542640519638181632140460266767440435607259782242325038;
            6'd44: xpb[37] = 1024'd31140090638398982762390242139448304841969515072357263988206340957971673032285771231684599936047488210684206111395237010539815621794748380988621028973805907726968446082413067818061874448810593037789446912896183918788063365341697860974270447832921205204710303802720957325541831484002159949168603608180791728343;
            6'd45: xpb[37] = 1024'd62864493892121054083962479493821192683643429014526577383607630655078889435528641668999381374622076974651452693064047573969577391591297746013516083613656984045094943044860714602879931393253771582612211017558816242169791381654687914692203054977204049457885968379039334499558050581666185475020289783204935615979;
            6'd46: xpb[37] = 1024'd94588897145843125405534716848194080525317342956695890779008920352186105838771512106314162813196665738618699274732858137399339161387847111038411138253508060363221440007308361387697988337696950127434975122221448565551519397967677968410135662121486893711061632955357711673574269679330211000871975958229079503615;
            6'd47: xpb[37] = 1024'd2246604715440455328308026797752535622292829773129520046278354984316426904705243633613873037113580193142796448944175266250037090343176141508146067877028095747657262400184790834885806090622922950947541618496841042568886564059771249163089699582540288697417394117559030817483960703065603509604972306627628906920;
            6'd48: xpb[37] = 1024'd33971007969162526649880264152125423463966743715298833441679644681423643307948114070928654475688168957110043030612985829679798860139725506533041122516879172065783759362632437619703863035066101495770305723159473365950614580372761302881022306726823132950593058693877407991500179800729629035456658481651772794556;
            6'd49: xpb[37] = 1024'd65695411222884597971452501506498311305640657657468146837080934378530859711190984508243435914262757721077289612281796393109560629936274871557936177156730248383910256325080084404521919979509280040593069827822105689332342596685751356598954913871105977203768723270195785165516398898393654561308344656675916682192;
            6'd50: xpb[37] = 1024'd97419814476606669293024738860871199147314571599637460232482224075638076114433854945558217352837346485044536193950606956539322399732824236582831231796581324702036753287527731189339976923952458585415833932484738012714070612998741410316887521015388821456944387846514162339532617996057680087160030831700060569828;
            6'd51: xpb[37] = 1024'd5077522046203999215798048810429654244290058416071089499751658707768397180367586472857927576754260939568633368161924085390020328688153267052566161420101360086472575680404160636527794676878431408928400428760130489731437779090834691069841558476442216443300149008715481483442309019793072595893027180098609973133;
            6'd52: xpb[37] = 1024'd36801925299926070537370286164802542085963972358240402895152948404875613583610456910172709015328849703535879949830734648819782098484702632077461216059952436404599072642851807421345851621321609953751164533422762813113165795403824744787774165620725060696475813585033858657458528117457098121744713355122753860769;
            6'd53: xpb[37] = 1024'd68526328553648141858942523519175429927637886300409716290554238101982829986853327347487490453903438467503126531499545212249543868281251997102356270699803512722725569605299454206163908565764788498573928638085395136494893811716814798505706772765007904949651478161352235831474747215121123647596399530146897748405;
            6'd54: xpb[37] = 1024'd100250731807370213180514760873548317769311800242579029685955527799090046390096197784802271892478027231470373113168355775679305638077801362127251325339654589040852066567747100990981965510207967043396692742748027459876621828029804852223639379909290749202827142737670613005490966312785149173448085705171041636041;
            6'd55: xpb[37] = 1024'd7908439376967543103288070823106772866287287059012658953224962431220367456029929312101982116394941685994470287379672904530003567033130392596986254963174624425287888960623530438169783263133939866909259239023419936893988994121898132976593417370344144189182903899871932149400657336520541682181082053569591039346;
            6'd56: xpb[37] = 1024'd39632842630689614424860308177479660707961201001181972348626252128327583859272799749416763554969530449961716869048483467959765336829679757621881309603025700743414385923071177222987840207577118411732023343686052260275717010434888186694526024514626988442358568476190309323416876434184567208032768228593734926982;
            6'd57: xpb[37] = 1024'd71357245884411685746432545531852548549635114943351285744027541825434800262515670186731544993544119213928963450717294031389527106626229122646776364242876777061540882885518824007805897152020296956554787448348684583657445026747878240412458631658909832695534233052508686497433095531848592733884454403617878814618;
            6'd58: xpb[37] = 1024'd103081649138133757068004782886225436391309028885520599139428831522542016665758540624046326432118707977896210032386104594819288876422778487671671418882727853379667379847966470792623954096463475501377551553011316907039173043060868294130391238803192676948709897628827063671449314629512618259736140578642022702254;
            6'd59: xpb[37] = 1024'd10739356707731086990778092835783891488284515701954228406698266154672337731692272151346036656035622432420307206597421723669986805378107518141406348506247888764103202240842900239811771849389448324890118049286709384056540209152961574883345276264246071935065658791028382815359005653248010768469136927040572105559;
            6'd60: xpb[37] = 1024'd42463759961453158312350330190156779329958429644123541802099555851779554134935142588660818094610211196387553788266232287099748575174656883166301403146098965082229699203290547024629828793832626869712882153949341707438268225465951628601277883408528916188241323367346759989375224750912036294320823102064715993195;
            6'd61: xpb[37] = 1024'd74188163215175229633922567544529667171632343586292855197500845548886770538178013025975599533184799960354800369935042850529510344971206248191196457785950041400356196165738193809447885738275805414535646258611974030819996241778941682319210490552811760441416987943665137163391443848576061820172509277088859880831;
            6'd62: xpb[37] = 1024'd105912566468897300955494804898902555013306257528462168592902135245993986941420883463290380971759388724322046951603853413959272114767755613216091512425801117718482693128185840594265942682718983959358410363274606354201724258091931736037143097697094604694592652519983514337407662946240087346024195452113003768467;
            6'd63: xpb[37] = 1024'd13570274038494630878268114848461010110281744344895797860171569878124308007354614990590091195676303178846144125815170542809970043723084643685826442049321153102918515521062270041453760435644956782870976859549998831219091424184025016790097135158147999680948413682184833481317353969975479854757191800511553171772;
        endcase
    end

    always_comb begin
        case(flag[12][16:12])
            5'd0: xpb[38] = 1024'd0;
            5'd1: xpb[38] = 1024'd45294677292216702199840352202833897951955658287065111255572859575231524410597485427904872634250891942813390707483981106239731813519634008710721496689172229421045012483509916826271817380088135327693740964212631154600819440497015070508029742302430843934124078258503210655333573067639505380608877975535697059408;
            5'd2: xpb[38] = 1024'd90589354584433404399680704405667795903911316574130222511145719150463048821194970855809745268501783885626781414967962212479463627039268017421442993378344458842090024967019833652543634760176270655387481928425262309201638880994030141016059484604861687868248156517006421310667146135279010761217755951071394118816;
            5'd3: xpb[38] = 1024'd11817336192525365200722129203687261111168547735459649638586723660717677894483317373699546688095001518997022714994449884140131599717681691577004365051185647329444362880958533141185212948747200261771025284250653617438097471270148438559110657224063082535552331361392573935894191128989883124707944099981496693893;
            5'd4: xpb[38] = 1024'd57112013484742067400562481406521159063124206022524760894159583235949202305080802801604419322345893461810413422478430990379863413237315700287725861740357876750489375364468449967457030328835335589464766248463284772038916911767163509067140399526493926469676409619895784591227764196629388505316822075517193753301;
            5'd5: xpb[38] = 1024'd102406690776958769600402833609355057015079864309589872149732442811180726715678288229509291956596785404623804129962412096619595226756949708998447358429530106171534387847978366793728847708923470917158507212675915926639736352264178579575170141828924770403800487878398995246561337264268893885925700051052890812709;
            5'd6: xpb[38] = 1024'd23634672385050730401444258407374522222337095470919299277173447321435355788966634747399093376190003037994045429988899768280263199435363383154008730102371294658888725761917066282370425897494400523542050568501307234876194942540296877118221314448126165071104662722785147871788382257979766249415888199962993387786;
            5'd7: xpb[38] = 1024'd68929349677267432601284610610208420174292753757984410532746306896666880199564120175303966010440894980807436137472880874519995012954997391864730226791543524079933738245426983108642243277582535851235791532713938389477014383037311947626251056750557009005228740981288358527121955325619271630024766175498690447194;
            5'd8: xpb[38] = 1024'd114224026969484134801124962813042318126248412045049521788319166471898404610161605603208838644691786923620826844956861980759726826474631400575451723480715753500978750728936899934914060657670671178929532496926569544077833823534327018134280799052987852939352819239791569182455528393258777010633644151034387506602;
            5'd9: xpb[38] = 1024'd35452008577576095602166387611061783333505643206378948915760170982153033683449952121098640064285004556991068144983349652420394799153045074731013095153556941988333088642875599423555638846241600785313075852751960852314292413810445315677331971672189247606656994084177721807682573386969649374123832299944490081679;
            5'd10: xpb[38] = 1024'd80746685869792797802006739813895681285461301493444060171333030557384558094047437549003512698535896499804458852467330758660126612672679083441734591842729171409378101126385516249827456226329736113006816816964592006915111854307460386185361713974620091540781072342680932463016146454609154754732710275480187141087;
            5'd11: xpb[38] = 1024'd1974667477884758603048164611915146492718532654773487298774035067639187167335784066893314118129114133174700152493818430320794585351092757597295963515570359896732439040324215738469034414900665719390360172789983315151570444583578683728412886593821486208085247187067085088243191448320027118222898424390289716164;
            5'd12: xpb[38] = 1024'd47269344770101460802888516814749044444674190941838598554346894642870711577933269494798186752380006075988090859977799536560526398870726766308017460204742589317777451523834132564740851794988801047084101137002614469752389885080593754236442628896252330142209325445570295743576764515959532498831776399925986775572;
            5'd13: xpb[38] = 1024'd92564022062318163002728869017582942396629849228903709809919754218102235988530754922703059386630898018801481567461780642800258212390360775018738956893914818738822464007344049391012669175076936374777842101215245624353209325577608824744472371198683174076333403704073506398910337583599037879440654375461683834980;
            5'd14: xpb[38] = 1024'd13792003670410123803770293815602407603887080390233136937360758728356865061819101440592860806224115652171722867488268314460926185068774449174300328566756007226176801921282748879654247363647865981161385457040636932589667915853727122287523543817884568743637578548459659024137382577309910242930842524371786410057;
            5'd15: xpb[38] = 1024'd59086680962626826003610646018436305555842738677298248192933618303588389472416586868497733440475007594985113574972249420700657998588408457885021825255928236647221814404792665705926064743736001308855126421253268087190487356350742192795553286120315412677761656806962869679470955644949415623539720499907483469465;
            5'd16: xpb[38] = 1024'd104381358254843528203450998221270203507798396964363359448506477878819913883014072296402606074725899537798504282456230526940389812108042466595743321945100466068266826888302582532197882123824136636548867385465899241791306796847757263303583028422746256611885735065466080334804528712588921004148598475443180528873;
            5'd17: xpb[38] = 1024'd25609339862935489004492423019289668715055628125692786575947482389074542956302418814292407494319117171168745582482718198601057784786456140751304693617941654555621164802241282020839460312395066242932410741291290550027765387123875560846634201041947651279189909909852232960031573706299793367638786624353283103950;
            5'd18: xpb[38] = 1024'd70904017155152191204332775222123566667011286412757897831520341964306067366899904242197280128570009113982136289966699304840789598306090149462026190307113883976666177285751198847111277692483201570626151705503921704628584827620890631354663943344378495213313988168355443615365146773939298748247664599888980163358;
            5'd19: xpb[38] = 1024'd116198694447368893404173127424957464618966944699823009087093201539537591777497389670102152762820901056795526997450680411080521411825724158172747686996286113397711189769261115673383095072571336898319892669716552859229404268117905701862693685646809339147438066426858654270698719841578804128856542575424677222766;
            5'd20: xpb[38] = 1024'd37426676055460854205214552222976929826224175861152436214534206049792220850785736187991954182414118690165768297477168082741189384504137832328309058669127301885065527683199815162024673261142266504703436025541944167465862858394023999405744858266010733814742241271244806895925764835289676492346730724334779797843;
            5'd21: xpb[38] = 1024'd82721353347677556405054904425810827778179834148217547470107065625023745261383221615896826816665010632979159004961149188980921198023771841039030555358299531306110540166709731988296490641230401832397176989754575322066682298891039069913774600568441577748866319529748017551259337902929181872955608699870476857251;
            5'd22: xpb[38] = 1024'd3949334955769517206096329223830292985437065309546974597548070135278374334671568133786628236258228266349400304987636860641589170702185515194591927031140719793464878080648431476938068829801331438780720345579966630303140889167157367456825773187642972416170494374134170176486382896640054236445796848780579432328;
            5'd23: xpb[38] = 1024'd49244012247986219405936681426664190937392723596612085853120929710509898745269053561691500870509120209162791012471617966881320984221819523905313423720312949214509890564158348303209886209889466766474461309792597784903960329664172437964855515490073816350294572632637380831819955964279559617054674824316276491736;
            5'd24: xpb[38] = 1024'd94538689540202921605777033629498088889348381883677197108693789285741423155866538989596373504760012151976181719955599073121052797741453532616034920409485178635554903047668265129481703589977602094168202274005228939504779770161187508472885257792504660284418650891140591487153529031919064997663552799851973551144;
            5'd25: xpb[38] = 1024'd15766671148294882406818458427517554096605613045006624236134793795996052229154885507486174924353229785346423019982086744781720770419867206771596292082326367122909240961606964618123281778548531700551745629830620247741238360437305806015936430411706054951722825735526744112380574025629937361153740948762076126221;
            5'd26: xpb[38] = 1024'd61061348440511584606658810630351452048561271332071735491707653371227576639752370935391047558604121728159813727466067851021452583939501215482317788771498596543954253445116881444395099158636667028245486594043251402342057800934320876523966172714136898885846903994029954767714147093269442741762618924297773185629;
            5'd27: xpb[38] = 1024'd106356025732728286806499162833185350000516929619136846747280512946459101050349856363295920192855013670973204434950048957261184397459135224193039285460670825964999265928626798270666916538724802355939227558255882556942877241431335947031995915016567742819970982252533165423047720160908948122371496899833470245037;
            5'd28: xpb[38] = 1024'd27584007340820247607540587631204815207774160780466273874721517456713730123638202881185721612448231304343445734976536628921852370137548898348600657133512014452353603842565497759308494727295731962322770914081273865179335831707454244575047087635769137487275157096919318048274765154619820485861685048743572820114;
            5'd29: xpb[38] = 1024'd72878684633036949807380939834038713159729819067531385130294377031945254534235688309090594246699123247156836442460517735161584183657182907059322153822684243873398616326075414585580312107383867290016511878293905019780155272204469315083076829938199981421399235355422528703608338222259325866470563024279269879522;
            5'd30: xpb[38] = 1024'd118173361925253652007221292036872611111685477354596496385867236607176778944833173736995466880950015189970227149944498841401315997176816915770043650511856473294443628809585331411852129487472002617710252842506536174380974712701484385591106572240630825355523313613925739358941911289898831247079440999814966938930;
            5'd31: xpb[38] = 1024'd39401343533345612808262716834892076318942708515925923513308241117431408018121520254885268300543232823340468449970986513061983969855230589925605022184697661781797966723524030900493707676042932224093796198331927482617433302977602683134157744859832220022827488458311891984168956283609703610569629148725069514007;
        endcase
    end

    always_comb begin
        case(flag[13][5:0])
            6'd0: xpb[39] = 1024'd0;
            6'd1: xpb[39] = 1024'd104381358254843528203450998221270203507798396964363359448506477878819913883014072296402606074725899537798504282456230526940389812108042466595743321945100466068266826888302582532197882123824136636548867385465899241791306796847757263303583028422746256611885735065466080334804528712588921004148598475443180528873;
            6'd2: xpb[39] = 1024'd84696020825562315008103069037725974270898366802991034768881100692662932428719005682790140934794124766153859157454967619301715783374864598636326518873869891202842979207033947726765525056131067551787537162544558637218252743474617753642187487162263063956951566716815102639502529351249208991178507124260766573415;
            6'd3: xpb[39] = 1024'd65010683396281101812755139854181745033998336641618710089255723506505950974423939069177675794862349994509214032453704711663041754641686730676909715802639316337419131525765312921333167988437998467026206939623218032645198690101478243980791945901779871302017398368164124944200529989909496978208415773078352617957;
            6'd4: xpb[39] = 1024'd45325345966999888617407210670637515797098306480246385409630346320348969520128872455565210654930575222864568907452441804024367725908508862717492912731408741471995283844496678115900810920744929382264876716701877428072144636728338734319396404641296678647083230019513147248898530628569784965238324421895938662499;
            6'd5: xpb[39] = 1024'd25640008537718675422059281487093286560198276318874060730004969134191988065833805841952745514998800451219923782451178896385693697175330994758076109660178166606571436163228043310468453853051860297503546493780536823499090583355199224658000863380813485992149061670862169553596531267230072952268233070713524707041;
            6'd6: xpb[39] = 1024'd5954671108437462226711352303549057323298246157501736050379591948035006611538739228340280375067025679575278657449915988747019668442153126798659306588947591741147588481959408505036096785358791212742216270859196218926036529982059714996605322120330293337214893322211191858294531905890360939298141719531110751583;
            6'd7: xpb[39] = 1024'd110336029363280990430162350524819260831096643121865095498886069826854920494552811524742886449792925217373782939906146515687409480550195593394402628534048057809414415370261991037233978909182927849291083656325095460717343326829816978300188350543076549949100628387677272193099060618479281943446740194974291280456;
            6'd8: xpb[39] = 1024'd90650691933999777234814421341275031594196612960492770819260692640697939040257744911130421309861150445729137814904883608048735451817017725434985825462817482943990567688993356231801621841489858764529753433403754856144289273456677468638792809282593357294166460039026294497797061257139569930476648843791877324998;
            6'd9: xpb[39] = 1024'd70965354504718564039466492157730802357296582799120446139635315454540957585962678297517956169929375674084492689903620700410061423083839857475569022391586908078566720007724721426369264773796789679768423210482414251571235220083537958977397268022110164639232291690375316802495061895799857917506557492609463369540;
            6'd10: xpb[39] = 1024'd51280017075437350844118562974186573120396552637748121460009938268383976131667611683905491029997600902439847564902357792771387394350661989516152219320356333213142872326456086620936907706103720595007092987561073646998181166710398449316001726761626971984298123341724339107193062534460145904536466141427049414082;
            6'd11: xpb[39] = 1024'd31594679646156137648770633790642343883496522476375796780384561082226994677372545070293025890065826130795202439901094885132713365617484121556735416249125758347719024645187451815504550638410651510245762764639733042425127113337258939654606185501143779329363954993073361411891063173120433891566374790244635458624;
            6'd12: xpb[39] = 1024'd11909342216874924453422704607098114646596492315003472100759183896070013223077478456680560750134051359150557314899831977494039336884306253597318613177895183482295176963918817010072193570717582425484432541718392437852073059964119429993210644240660586674429786644422383716589063811780721878596283439062221503166;
            6'd13: xpb[39] = 1024'd116290700471718452656873702828368318154394889279366831549265661774889927106091550753083166824859950896949061597356062504434429148992348720193061935122995649550562003852221399542270075694541719062033299927184291679643379856811876693296793672663406843286315521709888464051393592524369642882744881914505402032039;
            6'd14: xpb[39] = 1024'd96605363042437239461525773644824088917494859117994506869640284588732945651796484139470701684928176125304416472354799596795755120259170852233645132051765074685138156170952764736837718626848649977271969704262951075070325803438737183635398131402923650631381353361237486356091593163029930869774790563322988076581;
            6'd15: xpb[39] = 1024'd76920025613156026266177844461279859680594828956622182190014907402575964197501417525858236544996401353659771347353536689157081091525992984274228328980534499819714308489684129931405361559155580892510639481341610470497271750065597673974002590142440457976447185012586508660789593801690218856804699212140574121123;
            6'd16: xpb[39] = 1024'd57234688183874813070829915277735630443694798795249857510389530216418982743206350912245771405064626582015126222352273781518407062792815116314811525909303924954290460808415495125973004491462511807749309258420269865924217696692458164312607048881957265321513016663935530965487594440350506843834607860958160165665;
            6'd17: xpb[39] = 1024'd37549350754593599875481986094191401206794768633877532830764153030262001288911284298633306265132851810370481097351010873879733034059637248355394722838073350088866613127146860320540647423769442722987979035498929261351163643319318654651211507621474072666578848315284553270185595079010794830864516509775746210207;
            6'd18: xpb[39] = 1024'd17864013325312386680134056910647171969894738472505208151138775844105019834616217685020841125201077038725835972349747966241059005326459380395977919766842775223442765445878225515108290356076373638226648812577588656778109589946179144989815966360990880011644679966633575574883595717671082817894425158593332254749;
            6'd19: xpb[39] = 1024'd122245371580155914883585055131917375477693135436868567599645253722924933717630289981423447199926976576524340254805978493181448817434501846991721241711943241291709592334180808047306172479900510274775516198043487898569416386793936408293398994783737136623530415032099655909688124430260003822043023634036512783622;
            6'd20: xpb[39] = 1024'd102560034150874701688237125948373146240793105275496242920019876536767952263335223367810982059995201804879695129804715585542774788701323979032304438640712666426285744652912173241873815412207441190014185975122147293996362333420796898632003453523253943968596246683448678214386125068920291809072932282854098828164;
            6'd21: xpb[39] = 1024'd82874696721593488492889196764828917003893075114123918240394499350610970809040156754198516920063427033235050004803452677904100759968146111072887635569482091560861896971643538436441458344514372105252855752200806689423308280047657388970607912262770751313662078334797700519084125707580579796102840931671684872706;
            6'd22: xpb[39] = 1024'd63189359292312275297541267581284687766993044952751593560769122164453989354745090140586051780131652261590404879802189770265426731234968243113470832498251516695438049290374903631009101276821303020491525529279466084850254226674517879309212371002287558658727909986146722823782126346240867783132749580489270917248;
            6'd23: xpb[39] = 1024'd43504021863031062102193338397740458530093014791379268881143744978297007900450023526973586640199877489945759754800926862626752702501790375154054029427020941830014201609106268825576744209128233935730195306358125480277200173301378369647816829741804366003793741637495745128480126984901155770162658229306856961790;
            6'd24: xpb[39] = 1024'd23818684433749848906845409214196229293192984630006944201518367792140026446154956913361121500268102718301114629799663954988078673768612507194637226355790366964590353927837634020144387141435164850968865083436784875704146119928238859986421288481321173348859573288844767433178127623561443757192566878124443006332;
            6'd25: xpb[39] = 1024'd4133347004468635711497480030652000056292954468634619521892990605983044991859890299748656360336327946656469504798401047349404645035434639235220423284559792099166506246568999214712030073742095766207534860515444271131092066555099350325025747220837980693925404940193789737876128262221731744222475526942029050874;
            6'd26: xpb[39] = 1024'd108514705259312163914948478251922203564091351432997978970399468484802958874873962596151262435062227484454973787254631574289794457143477105830963745229660258167433333134871581746909912197566232402756402245981343512922398863402856613628608775643584237305811140005659870072680656974810652748371074002385209579747;
            6'd27: xpb[39] = 1024'd88829367830030950719600549068377974327191321271625654290774091298645977420578895982538797295130452712810328662253368666651120428410299237871546942158429683302009485453602946941477555129873163317995072023060002908349344810029717103967213234383101044650876971657008892377378657613470940735400982651202795624289;
            6'd28: xpb[39] = 1024'd69144030400749737524252619884833745090291291110253329611148714112488995966283829368926332155198677941165683537252105759012446399677121369912130139087199108436585637772334312136045198062180094233233741800138662303776290756656577594305817693122617851995942803308357914682076658252131228722430891300020381668831;
            6'd29: xpb[39] = 1024'd49458692971468524328904690701289515853391260948881004931523336926332014511988762755313867015266903169521038412250842851373772370943943501952713336015968533571161790091065677330612840994487025148472411577217321699203236703283438084644422151862134659341008634959706936986774658890791516709460799948837967713373;
            6'd30: xpb[39] = 1024'd29773355542187311133556761517745286616491230787508680251897959740175033057693696141701401875335128397876393287249579943735098342210765633993296532944737958705737942409797042525180483926793956063711081354295981094630182649910298574983026610601651466686074466611055959291472659529451804696490708597655553757915;
            6'd31: xpb[39] = 1024'd10088018112906097938208832334201057379591200626136355572272582554018051603398629528088936735403353626231748162248317036096424313477587766033879729873507383840314094728528407719748126859100886978949751131374640490057128596537159065321631069341168274031140298262404981596170660168112092683520617246473139802457;
            6'd32: xpb[39] = 1024'd114469376367749626141659830555471260887389597590499715020779060432837965486412701824491542810129253164030252444704547563036814125585630232629623051818607849908580921616830990251946008982925023615498618516840539731848435393384916328625214097763914530643026033327871061930975188880701013687669215721916320331330;
            6'd33: xpb[39] = 1024'd94784038938468412946311901371927031650489567429127390341153683246680984032117635210879077670197478392385607319703284655398140096852452364670206248747377275043157073935562355446513651915231954530737288293919199127275381340011776818963818556503431337988091864979220084235673189519361301674699124370733906375872;
            6'd34: xpb[39] = 1024'd75098701509187199750963972188382802413589537267755065661528306060524002577822568597266612530265703620740962194702021747759466068119274496710789445676146700177733226254293720641081294847538885445975958070997858522702327286638637309302423015242948145333157696630569106540371190158021589661729033019551492420414;
            6'd35: xpb[39] = 1024'd55413364079905986555616043004838573176689507106382740981902928874367021123527501983654147390333928849096317069700758840120792039386096628751372642604916125312309378573025085835648937779845816361214627848076517918129273233265497799641027473982464952678223528281918128845069190796681877648758941668369078464956;
            6'd36: xpb[39] = 1024'd35728026650624773360268113821294343939789476945010416302277551688210039669232435370041682250402154077451671944699495932482118010652918760791955839533685550446885530891756451030216580712152747276453297625155177313556219179892358289979631932721981760023289359933267151149767191435342165635788850317186664509498;
            6'd37: xpb[39] = 1024'd16042689221343560164920184637750114702889446783638091622652174502053058214937368756429217110470379305807026819698233024843443981919740892832539036462454975581461683210487816224784223644459678191691967402233836708983165126519218780318236391461498567368355191584616173454465192074002453622818758966004250554040;
            6'd38: xpb[39] = 1024'd120424047476187088368371182859020318210687843748001451071158652380872972097951441052831823185196278843605531102154463551783833794027783359428282358407555441649728510098790398756982105768283814828240834787699735950774471923366976043621819419884244823980240926650082253789269720786591374626967357441447431082913;
            6'd39: xpb[39] = 1024'd100738710046905875173023253675476088973787813586629126391533275194715990643656374439219358045264504071960885977153200644145159765294605491468865555336324866784304662417521763951549748700590745743479504564778395346201417869993836533960423878623761631325306758301431276093967721425251662613997266090265017127455;
            6'd40: xpb[39] = 1024'd81053372617624661977675324491931859736887783425256801711907898008559009189361307825606892905332729300316240852151937736506485736561427623509448752265094291918880814736253129146117391632897676658718174341857054741628363816620697024299028337363278438670372589952780298398665722063911950601027174739082603171997;
            6'd41: xpb[39] = 1024'd61368035188343448782327395308387630499987753263884477032282520822402027735066241211994427765400954528671595727150674828867811707828249755550031949193863717053456967054984494340685034565204607573956844118935714137055309763247557514637632796102795246015438421604129320703363722702572238588057083387900189216539;
            6'd42: xpb[39] = 1024'd41682697759062235586979466124843401263087723102512152352657143636245046280771174598381962625469179757026950602149411921229137679095071887590615146122633142188033119373715859535252677497511538489195513896014373532482255709874418004976237254842312053360504253255478343008061723341232526575086992036717775261081;
            6'd43: xpb[39] = 1024'd21997360329781022391631536941299172026187692941139827673031766450088064826476107984769497485537404985382305477148149013590463650361894019631198343051402567322609271692447224729820320429818469404434183673093032927909201656501278495314841713581828860705570084906827365312759723979892814562116900685535361305623;
            6'd44: xpb[39] = 1024'd2312022900499809196283607757754942789287662779767502993406389263931083372181041371157032345605630213737660352146886105951789621628716151671781539980171992457185424011178589924387963362125400319672853450171692323336147603128138985653446172321345668050635916558176387617457724618553102549146809334352947350165;
            6'd45: xpb[39] = 1024'd106693381155343337399734605979025146297086059744130862441912867142750997255195113667559638420331529751536164634603116632892179433736758618267524861925272458525452250899481172456585845485949536956221720835637591565127454399975896248957029200744091924662521651623642467952262253331142023553295407809796127879038;
            6'd46: xpb[39] = 1024'd87008043726062124204386676795480917060186029582758537762287489956594015800900047053947173280399754979891519509601853725253505405003580750308108058854041883660028403218212537651153488418256467871460390612716250960554400346602756739295633659483608732007587483274991490256960253969802311540325316458613713923580;
            6'd47: xpb[39] = 1024'd67322706296780911009038747611936687823285999421386213082662112770437034346604980440334708140467980208246874384600590817614831376270402882348691255782811308794604555536943902845721131350563398786699060389794910355981346293229617229634238118223125539352653314926340512561658254608462599527355225107431299968122;
            6'd48: xpb[39] = 1024'd47637368867499697813690818428392458586385969260013888403036735584280052892309913826722243000536205436602229259599327909976157347537225014389274452711580733929180707855675268040288774282870329701937730166873569751408292239856477719972842576962642346697719146577689534866356255247122887514385133756248886012664;
            6'd49: xpb[39] = 1024'd27952031438218484618342889244848229349485939098641563723411358398123071438014847213109777860604430664957584134598065002337483318804047146429857649640350159063756860174406633234856417215177260617176399943952229146835238186483338210311447035702159154042784978229038557171054255885783175501415042405066472057206;
            6'd50: xpb[39] = 1024'd8266694008937271422994960061304000112585908937269239043785981211966089983719780599497312720672655893312939009596802094698809290070869278470440846569119584198333012493137998429424060147484191532415069721030888542262184133110198700650051494441675961387850809880387579475752256524443463488444951053884058101748;
            6'd51: xpb[39] = 1024'd112648052263780799626445958282574203620384305901632598492292459090786003866733852895899918795398555431111443292053032621639199102178911745066184168514220050266599839381440580961621942271308328168963937106496787784053490929957955963953634522864422217999736544945853659810556785237032384492593549529327238630621;
            6'd52: xpb[39] = 1024'd92962714834499586431098029099029974383484275740260273812667081904629022412438786282287453655466780659466798167051769714000525073445733877106767365442989475401175991700171946156189585203615259084202606883575447179480436876584816454292238981603939025344802376597202682115254785875692672479623458178144824675163;
            6'd53: xpb[39] = 1024'd73277377405218373235750099915485745146584245578887949133041704718472040958143719668674988515535005887822153042050506806361851044712556009147350562371758900535752144018903311350757228135922189999441276660654106574907382823211676944630843440343455832689868208248551704419952786514352960466653366826962410719705;
            6'd54: xpb[39] = 1024'd53592039975937160040402170731941515909684215417515624453416327532315059503848653055062523375603231116177507917049243898723177015979378141187933759300528325670328296337634676545324871068229120914679946437732765970334328769838537434969447899082972640034934039899900726724650787153013248453683275475779996764247;
            6'd55: xpb[39] = 1024'd33906702546655946845054241548397286672784185256143299773790950346158078049553586441450058235671456344532862792047980991084502987246200273228516956229297750804904448656366041739892514000536051829918616214811425365761274716465397925308052357822489447379999871551249749029348787791673536440713184124597582808789;
            6'd56: xpb[39] = 1024'd14221365117374733649706312364853057435884155094770975094165573160001096595258519827837593095739681572888217667046718083445828958513022405269100153158067175939480600975097406934460156932842982745157285991890084761188220663092258415646656816562006254725065703202598771334046788430333824427743092773415168853331;
            6'd57: xpb[39] = 1024'd118602723372218261853157310586123260943682552059134334542672051038821010478272592124240199170465581110686721949502948610386218770621064871864843475103167642007747427863399989466658039056667119381706153377355984002979527459940015678950239844984752511336951438268064851668851317142922745431891691248858349382204;
            6'd58: xpb[39] = 1024'd98917385942937048657809381402579031706782521897762009863046673852664029023977525510627734030533806339042076824501685702747544741887887003905426672031937067142323580182131354661225681988974050296944823154434643398406473406566876169288844303724269318682017269919413873973549317781583033418921599897675935426746;
            6'd59: xpb[39] = 1024'd79232048513655835462461452219034802469882491736389685183421296666507047569682458897015268890602031567397431699500422795108870713154709135946009868960706492276899732500862719855793324921280981212183492931513302793833419353193736659627448762463786126027083101570762896278247318420243321405951508546493521471288;
            6'd60: xpb[39] = 1024'd59546711084374622267113523035490573232982461575017360503795919480350066115387392283402803750670256795752786574499159887470196684421531267986593065889475917411475884819594085050360967853587912127422162708591962189260365299820597149966053221203302933372148933222111918582945319058903609392981417195311107515830;
            6'd61: xpb[39] = 1024'd39861373655093409071765593851946343996082431413645035824170542294193084661092325669790338610738482024108141449497896979831522655688353400027176262818245342546052037138325450244928610785894843042660832485670621584687311246447457640304657679942819740717214764873460940887643319697563897380011325844128693560372;
            6'd62: xpb[39] = 1024'd20176036225812195876417664668402114759182401252272711144545165108036103206797259056177873470806707252463496324496634072192848626955175532067759459747014767680628189457056815439496253718201773957899502262749280980114257193074318130643262138682336548062280596524809963192341320336224185367041234492946279604914;
            6'd63: xpb[39] = 1024'd490698796530982681069735484857885522282371090900386464919787921879121752502192442565408330874932480818851199495371164554174598221997664108342656675784192815204341775788180634063896650508704873138172039827940375541203139701178620981866597421853355407346428176158985497039320974884473354071143141763865649456;
        endcase
    end

    always_comb begin
        case(flag[13][11:6])
            6'd0: xpb[40] = 1024'd0;
            6'd1: xpb[40] = 1024'd104872057051374510884520733706128089030080768055263745913426265800699035635516264738968014405600832018617355481951601691494564410330040130704085978620884658883471168664090763166261778774332841509687039425293839617332509936548935884285449625844599612019232163241625065831843849687473394358219741617207046178329;
            6'd2: xpb[40] = 1024'd85677418418624280370242540007441745315463108984791807698720676536421175933723390567920957596543989727791561556445709948410064979818859926853011832225438276833251662758610308994893318357148477298063881242200439388300659022876974995605920682005969774771644423069133073633581171301018155699320793407788497872327;
            6'd3: xpb[40] = 1024'd66482779785874049855964346308755401600845449914319869484015087272143316231930516396873900787487147436965767630939818205325565549307679723001937685829991894783032156853129854823524857939964113086440723059107039159268808109205014106926391738167339937524056682896641081435318492914562917040421845198369949566325;
            6'd4: xpb[40] = 1024'd47288141153123819341686152610069057886227790843847931269309498007865456530137642225826843978430305146139973705433926462241066118796499519150863539434545512732812650947649400652156397522779748874817564876013638930236957195533053218246862794328710100276468942724149089237055814528107678381522896988951401260323;
            6'd5: xpb[40] = 1024'd28093502520373588827407958911382714171610131773375993054603908743587596828344768054779787169373462855314179779928034719156566688285319315299789393039099130682593145042168946480787937105595384663194406692920238701205106281861092329567333850490080263028881202551657097038793136141652439722623948779532852954321;
            6'd6: xpb[40] = 1024'd8898863887623358313129765212696370456992472702904054839898319479309737126551893883732730360316620564488385854422142976072067257774139111448715246643652748632373639136688492309419476688411020451571248509826838472173255368189131440887804906651450425781293462379165104840530457755197201063725000570114304648319;
            6'd7: xpb[40] = 1024'd113770920938997869197650498918824459487073240758167800753324585280008772762068158622700744765917452583105741336373744667566631668104179242152801225264537407515844807800779255475681255462743861961258287935120678089505765304738067325173254532496050037800525625620790170672374307442670595421944742187321350826648;
            6'd8: xpb[40] = 1024'd94576282306247638683372305220138115772455581687695862538618996015730913060275284451653687956860610292279947410867852924482132237592999038301727078869091025465625301895298801304312795045559497749635129752027277860473914391066106436493725588657420200552937885448298178474111629056215356763045793977902802520646;
            6'd9: xpb[40] = 1024'd75381643673497408169094111521451772057837922617223924323913406751453053358482410280606631147803768001454153485361961181397632807081818834450652932473644643415405795989818347132944334628375133538011971568933877631442063477394145547814196644818790363305350145275806186275848950669760118104146845768484254214644;
            6'd10: xpb[40] = 1024'd56187005040747177654815917822765428343220263546751986109207817487175193656689536109559574338746925710628359559856069438313133376570638630599578786078198261365186290084337892961575874211190769326388813385840477402410212563722184659134667700980160526057762405103314194077586272283304879445247897559065705908642;
            6'd11: xpb[40] = 1024'd36992366407996947140537724124079084628602604476280047894502228222897333954896661938512517529690083419802565634350177695228633946059458426748504639682751879314966784178857438790207413794006405114765655202747077173378361650050223770455138757141530688810174664930822201879323593896849640786348949349647157602640;
            6'd12: xpb[40] = 1024'd17797727775246716626259530425392740913984945405808109679796638958619474253103787767465460720633241128976771708844285952144134515548278222897430493287305497264747278273376984618838953376822040903142497019653676944346510736378262881775609813302900851562586924758330209681060915510394402127450001140228609296638;
            6'd13: xpb[40] = 1024'd122669784826621227510780264131520829944065713461071855593222904759318509888620052506433475126234073147594127190795887643638698925878318353601516471908190156148218446937467747785100732151154882412829536444947516561679020672927198766061059439147500463581819087999955275512904765197867796485669742757435655474967;
            6'd14: xpb[40] = 1024'd103475146193870996996502070432834486229448054390599917378517315495040650186827178335386418317177230856768333265289995900554199495367138149750442325512743774097998941031987293613732271733970518201206378261854116332647169759255237877381530495308870626334231347827463283314642086811412557826770794548017107168965;
            6'd15: xpb[40] = 1024'd84280507561120766482223876734148142514830395320127979163811726230762790485034304164339361508120388565942539339784104157469700064855957945899368179117297392047779435126506839442363811316786153989583220078760716103615318845583276988702001551470240789086643607654971291116379408424957319167871846338598558862963;
            6'd16: xpb[40] = 1024'd65085868928370535967945683035461798800212736249656040949106136966484930783241429993292304699063546275116745414278212414385200634344777742048294032721851009997559929221026385270995350899601789777960061895667315874583467931911316100022472607631610951839055867482479298918116730038502080508972898129180010556961;
            6'd17: xpb[40] = 1024'd45891230295620305453667489336775455085595077179184102734400547702207071081448555822245247890006703984290951488772320671300701203833597538197219886326404627947340423315545931099626890482417425566336903712573915645551617018239355211342943663792981114591468127309987306719854051652046841850073949919761462250959;
            6'd18: xpb[40] = 1024'd26696591662870074939389295638089111370977418108712164519694958437929211379655681651198191080949861693465157563266428928216201773322417334346145739930958245897120917410065476928258430065233061354713745529480515416519766104567394322663414719954351277343880387137495314521591373265591603191175001710342913944957;
            6'd19: xpb[40] = 1024'd7501953030119844425111101939402767656359759038240226304989369173651351677862807480151134271893019402639363637760537185131702342811237130495071593535511863846901411504585022756889969648048697143090587346387115187487915190895433433983885776115721440096292646965003322323328694879136364532276053500924365638955;
            6'd20: xpb[40] = 1024'd112374010081494355309631835645530856686440527093503972218415634974350387313379072219119148677493851421256719119712138876626266753141277261199157572156396522730372580168675785923151748422381538652777626771680954804820425127444369318269335401960321052115524810206628388155172544566609758890495795118131411817284;
            6'd21: xpb[40] = 1024'd93179371448744124795353641946844512971822868023032034003710045710072527611586198048072091868437009130430925194206247133541767322630097057348083425760950140680153074263195331751783288005197174441154468588587554575788574213772408429589806458121691214867937070034136395956909866180154520231596846908712863511282;
            6'd22: xpb[40] = 1024'd73984732815993894281075448248158169257205208952560095789004456445794667909793323877025035059380166839605131268700355390457267892118916853497009279365503758629933568357714877580414827588012810229531310405494154346756723300100447540910277514283061377620349329861644403758647187793699281572697898699294315205280;
            6'd23: xpb[40] = 1024'd54790094183243663766797254549471825542587549882088157574298867181516808208000449705977978250323324548779337343194463647372768461607736649645935132970057376579714062452234423409046367170828446017908152222400754117724872386428486652230748570444431540372761589689152411560384509407244042913798950489875766899278;
            6'd24: xpb[40] = 1024'd35595455550493433252519060850785481827969890811616219359593277917238948506207575534930921441266482257953543417688571904288269031096556445794860986574610994529494556546753969237677906753644081806284994039307353888693021472756525763551219626605801703125173849516660419362121831020788804254900002280457218593276;
            6'd25: xpb[40] = 1024'd16400816917743202738240867152099138113352231741144281144887688652961088804414701363883864632209639967127749492182680161203769600585376241943786840179164612479275050641273515066309446336459717594661835856213953659661170559084564874871690682767171865877586109344168427163859152634333565596001054071038670287274;
            6'd26: xpb[40] = 1024'd121272873969117713622761600858227227143432999796408027058313954453660124439930966102851879037810471985745104974134281852698334010915416372647872818800049271362746219305364278232571225110792559104348875281507793276993680495633500759157140308611771477896818272585793492995703002321806959954220795688245716465603;
            6'd27: xpb[40] = 1024'd102078235336367483108483407159540883428815340725936088843608365189382264738138091931804822228753629694919311048628390109613834580404236168796798672404602889312526713399883824061202764693608194892725717098414393047961829581961539870477611364773141640649230532413301500797440323935351721295321847478827168159601;
            6'd28: xpb[40] = 1024'd82883596703617252594205213460854539714197681655464150628902775925104405036345217760757765419696787404093517123122498366529335149893055964945724526009156507262307207494403369889834304276423830681102558915320992818929978668289578981798082420934511803401642792240809508599177645548896482636422899269408619853599;
            6'd29: xpb[40] = 1024'd63688958070867022079927019762168195999580022584992212414197186660826545334552343589710708610639945113267723197616606623444835719381875761094650379613710125212087701588922915718465843859239466469479400732227592589898127754617618093118553477095881966154055052068317516400914967162441243977523951059990071547597;
            6'd30: xpb[40] = 1024'd44494319438116791565648826063481852284962363514520274199491597396548685632759469418663651801583102822441929272110714880360336288870695557243576233218263743161868195683442461547097383442055102257856242549134192360866276840945657204439024533257252128906467311895825524202652288775986005318625002850571523241595;
            6'd31: xpb[40] = 1024'd25299680805366561051370632364795508570344704444048335984786008132270825930966595247616594992526260531616135346604823137275836858359515353392502086822817361111648689777962007375728923024870738046233084366040792131834425927273696315759495589418622291658879571723333532004389610389530766659726054641152974935593;
            6'd32: xpb[40] = 1024'd6105042172616330537092438666109164855727045373576397770080418867992966229173721076569538183469418240790341421098931394191337427848335149541427940427370979061429183872481553204360462607686373834609926182947391902802575013601735427079966645579992454411291831550841539806126932003075528000827106431734426629591;
            6'd33: xpb[40] = 1024'd110977099223990841421613172372237253885807813428840143683506684668692001864689985815537552589070250259407696903050533085685901838178375280245513919048255637944900352536572316370622241382019215344296965608241231520135084950150671311365416271424592066430523994792466605637970781690548922359046848048941472807920;
            6'd34: xpb[40] = 1024'd91782460591240610907334978673550910171190154358368205468801095404414142162897111644490495780013407968581902977544641342601402407667195076394439772652809255894680846631091862199253780964834851132673807425147831291103234036478710422685887327585962229182936254619974613439708103304093683700147899839522924501918;
            6'd35: xpb[40] = 1024'd72587821958490380393056784974864566456572495287896267254095506140136282461104237473443438970956565677756109052038749599516902977156014872543365626257362873844461340725611408027885320547650486921050649242054431062071383122806749534006358383747332391935348514447482621241445424917638445041248951630104376195916;
            6'd36: xpb[40] = 1024'd53393183325740149878778591276178222741954836217424329039389916875858422759311363302396382161899723386930315126532857856432403546644834668692291479861916491794241834820130953856516860130466122709427491058961030833039532209134788645326829439908702554687760774274990629043182746531183206382350003420685827889914;
            6'd37: xpb[40] = 1024'd34198544692989919364500397577491879027337177146952390824684327611580563057518489131349325352842881096104521201026966113347904116133654464841217333466470109744022328914650499685148399713281758497804332875867630604007681295462827756647300496070072717440173034102498636844920068144727967723451055211267279583912;
            6'd38: xpb[40] = 1024'd15003906060239688850222203878805535312719518076480452609978738347302703355725614960302268543786038805278727275521074370263404685622474260990143187071023727693802823009170045513779939296097394286181174692774230374975830381790866867967771552231442880192585293930006644646657389758272729064552107001848731277910;
            6'd39: xpb[40] = 1024'd119875963111614199734742937584933624342800286131744198523405004148001738991241879699270282949386870823896082757472676061757969095952514391694229165691908386577273991673260808680041718070430235795868214118068069992308340318339802752253221178076042492211817457171631710478501239445746123422771848619055777456239;
            6'd40: xpb[40] = 1024'd100681324478863969220464743886247280628182627061272260308699414883723879289449005528223226140330028533070288831966784318673469665441334187843155019296462004527054485767780354508673257653245871584245055934974669763276489404667841863573692234237412654964229716999139718280238561059290884763872900409637229150237;
            6'd41: xpb[40] = 1024'd81486685846113738706186550187560936913564967990800322093993825619446019587656131357176169331273186242244494906460892575588970234930153983992080872901015622476834979862299900337304797236061507372621897751881269534244638490995880974894163290398782817716641976826647726081975882672835646104973952200218680844235;
            6'd42: xpb[40] = 1024'd62292047213363508191908356488874593198947308920328383879288236355168159885863257186129112522216343951418700980955000832504470804418973780141006726505569240426615473956819446165936336818877143160998739568787869305212787577323920086214634346560152980469054236654155733883713204286380407446075003990800132538233;
            6'd43: xpb[40] = 1024'd43097408580613277677630162790188249484329649849856445664582647090890300184070383015082055713159501660592907055449109089419971373907793576289932580110122858376395968051338991994567876401692778949375581385694469076180936663651959197535105402721523143221466496481663741685450525899925168787176055781381584232231;
            6'd44: xpb[40] = 1024'd23902769947863047163351969091501905769711990779384507449877057826612440482277508844034998904102659369767113129943217346335471943396613372438858433714676476326176462145858537823199415984508414737752423202601068847149085749979998308855576458882893305973878756309171749487187847513469930128277107571963035926229;
            6'd45: xpb[40] = 1024'd4708131315112816649073775392815562055094331708912569235171468562334580780484634672987942095045817078941319204437325603250972512885433168587784287319230094275956956240378083651830955567324050526129265019507668618117234836308037420176047515044263468726291016136679757288925169127014691469378159362544487620227;
            6'd46: xpb[40] = 1024'd109580188366487327533594509098943651085175099764176315148597734363033616416000899411955956500646649097558674686388927294745536923215473299291870265940114753159428124904468846818092734341656892035816304444801508235449744772856973304461497140888863080745523179378304823120769018814488085827597900979751533798556;
            6'd47: xpb[40] = 1024'd90385549733737097019316315400257307370557440693704376933892145098755756714208025240908899691589806806732880760883035551661037492704293095440796119544668371109208618998988392646724273924472527824193146261708108006417893859185012415781968197050233243497935439205812830922506340428032847168698952770332985492554;
            6'd48: xpb[40] = 1024'd71190911100986866505038121701570963655939781623232438719186555834477897012415151069861842882532964515907086835377143808576538062193112891589721973149221989058989113093507938475355813507288163612569988078614707777386042945513051527102439253211603406250347699033320838724243662041577608509800004560914437186552;
            6'd49: xpb[40] = 1024'd51996272468236635990759928002884619941322122552760500504480966570200037310622276898814786073476122225081292909871252065492038631681932687738647826753775607008769607188027484303987353090103799400946829895521307548354192031841090638422910309372973569002759958860828846525980983655122369850901056351495888880550;
            6'd50: xpb[40] = 1024'd32801633835486405476481734304198276226704463482288562289775377305922177608829402727767729264419279934255498984365360322407539201170752483887573680358329224958550101282547030132618892672919435189323671712427907319322341118169129749743381365534343731755172218688336854327718305268667131192002108142077340574548;
            6'd51: xpb[40] = 1024'd13606995202736174962203540605511932512086804411816624075069788041644317907036528556720672455362437643429705058859468579323039770659572280036499533962882842908330595377066575961250432255735070977700513529334507090290490204497168861063852421695713894507584478515844862129455626882211892533103159932658792268546;
            6'd52: xpb[40] = 1024'd118479052254110685846724274311640021542167572467080369988496053842343353542552793295688686860963269662047060540811070270817604180989612410740585512583767501791801764041157339127512211030067912487387552954628346707623000141046104745349302047540313506526816641757469927961299476569685286891322901549865838446875;
            6'd53: xpb[40] = 1024'd99284413621360455332446080612953677827549913396608431773790464578065493840759919124641630051906427371221266615305178527733104750478432206889511366188321119741582258135676884956143750612883548275764394771534946478591149227374143856669773103701683669279228901584977935763036798183230048232423953340447290140873;
            6'd54: xpb[40] = 1024'd80089774988610224818167886914267334112932254326136493559084875313787634138967044953594573242849585080395472689799286784648605319967252003038437219792874737691362752230196430784775290195699184064141236588441546249559298313702182967990244159863053832031641161412485943564774119796774809573525005131028741834871;
            6'd55: xpb[40] = 1024'd60895136355859994303889693215580990398314595255664555344379286049509774437174170782547516433792742789569678764293395041564105889456071799187363073397428355641143246324715976613406829778514819852518078405348146020527447400030222079310715216024423994784053421239993951366511441410319570914626056921610193528869;
            6'd56: xpb[40] = 1024'd41700497723109763789611499516894646683696936185192617129673696785231914735381296611500459624735900498743884838787503298479606458944891595336288927001981973590923740419235522442038369361330455640894920222254745791495596486358261190631186272185794157536465681067501959168248763023864332255727108712191645222867;
            6'd57: xpb[40] = 1024'd22505859090359533275333305818208302969079277114720678914968107520954055033588422440453402815679058207918090913281611555395107028433711391485214780606535591540704234513755068270669908944146091429271762039161345562463745572686300301951657328347164320288877940895009966969986084637409093596828160502773096916865;
            6'd58: xpb[40] = 1024'd3311220457609302761055112119521959254461618044248740700262518256676195331795548269406346006622215917092296987775719812310607597922531187634140634211089209490484728608274614099301448526961727217648603856067945333431894659014339413272128384508534483041290200722517974771723406250953854937929212293354548610863;
            6'd59: xpb[40] = 1024'd108183277508983813645575845825650048284542386099512486613688784057375230967311813008374360412223047935709652469727321503805172008252571318338226612831973868373955897272365377265563227301294568727335643281361784950764404595563275297557578010353134095060522363964143040603567255938427249296148953910561594789192;
            6'd60: xpb[40] = 1024'd88988638876233583131297652126963704569924727029040548398983194793097371265518938837327303603166205644883858544221429760720672577741391114487152466436527486323736391366884923094194766884110204515712485098268384721732553681891314408878049066514504257812934623791651048405304577551972010637250005701143046483190;
            6'd61: xpb[40] = 1024'd69794000243483352617019458428277360855307067958568610184277605528819511563726064666280246794109363354058064618715538017636173147230210910636078320041081104273516885461404468922826306466925840304089326915174984492700702768219353520198520122675874420565346883619159056207041899165516771978351057491724498177188;
            6'd62: xpb[40] = 1024'd50599361610733122102741264729591017140689408888096671969572016264541651861933190495233189985052521063232270693209646274551673716719030706785004173645634722223297379555924014751457846049741476092466168732081584263668851854547392631518991178837244583317759143446667064008779220779061533319452109282305949871186;
            6'd63: xpb[40] = 1024'd31404722977982891588463071030904673426071749817624733754866427000263792160140316324186133175995678772406476767703754531467174286207850502933930027250188340173077873650443560580089385632557111880843010548988184034637000940875431742839462234998614746070171403274175071810516542392606294660553161072887401565184;
        endcase
    end

    always_comb begin
        case(flag[13][16:12])
            5'd0: xpb[41] = 1024'd0;
            5'd1: xpb[41] = 1024'd12210084345232661074184877332218329711454090747152795540160837735985932458347442153139076366938836481580682842197862788382674855696670299082855880854741958122858367744963106408720925215372747669219852365894783805605150027203470854159933291159984908822583663101683079612253864006151056001654212863468853259182;
            5'd2: xpb[41] = 1024'd24420168690465322148369754664436659422908181494305591080321675471971864916694884306278152733877672963161365684395725576765349711393340598165711761709483916245716735489926212817441850430745495338439704731789567611210300054406941708319866582319969817645167326203366159224507728012302112003308425726937706518364;
            5'd3: xpb[41] = 1024'd36630253035697983222554631996654989134362272241458386620482513207957797375042326459417229100816509444742048526593588365148024567090010897248567642564225874368575103234889319226162775646118243007659557097684351416815450081610412562479799873479954726467750989305049238836761592018453168004962638590406559777546;
            5'd4: xpb[41] = 1024'd48840337380930644296739509328873318845816362988611182160643350943943729833389768612556305467755345926322731368791451153530699422786681196331423523418967832491433470979852425634883700861490990676879409463579135222420600108813883416639733164639939635290334652406732318449015456024604224006616851453875413036728;
            5'd5: xpb[41] = 1024'd61050421726163305370924386661091648557270453735763977700804188679929662291737210765695381834694182407903414210989313941913374278483351495414279404273709790614291838724815532043604626076863738346099261829473919028025750136017354270799666455799924544112918315508415398061269320030755280008271064317344266295910;
            5'd6: xpb[41] = 1024'd73260506071395966445109263993309978268724544482916773240965026415915594750084652918834458201633018889484097053187176730296049134180021794497135285128451748737150206469778638452325551292236486015319114195368702833630900163220825124959599746959909452935501978610098477673523184036906336009925277180813119555092;
            5'd7: xpb[41] = 1024'd85470590416628627519294141325528307980178635230069568781125864151901527208432095071973534568571855371064779895385039518678723989876692093579991165983193706860008574214741744861046476507609233684538966561263486639236050190424295979119533038119894361758085641711781557285777048043057392011579490044281972814274;
            5'd8: xpb[41] = 1024'd97680674761861288593479018657746637691632725977222364321286701887887459666779537225112610935510691852645462737582902307061398845573362392662847046837935664982866941959704851269767401722981981353758818927158270444841200217627766833279466329279879270580669304813464636898030912049208448013233702907750826073456;
            5'd9: xpb[41] = 1024'd109890759107093949667663895989964967403086816724375159861447539623873392125126979378251687302449528334226145579780765095444073701270032691745702927692677623105725309704667957678488326938354729022978671293053054250446350244831237687439399620439864179403252967915147716510284776055359504014887915771219679332638;
            5'd10: xpb[41] = 1024'd122100843452326610741848773322183297114540907471527955401608377359859324583474421531390763669388364815806828421978627883826748556966702990828558808547419581228583677449631064087209252153727476692198523658947838056051500272034708541599332911599849088225836631016830796122538640061510560016542128634688532591820;
            5'd11: xpb[41] = 1024'd10244232113434530417234723249587194081296571092945066813637360030868361704512724774514768821669526987944361856718997237630359571822152955356254564385830498417751370625022953158299938177583018640108178416455382015292289449017282622794287633076604547781600390704396817704685975993732983001077651671531791366671;
            5'd12: xpb[41] = 1024'd22454316458667191491419600581805523792750661840097862353798197766854294162860166927653845188608363469525044698916860026013034427518823254439110445240572456540609738369986059567020863392955766309328030782350165820897439476220753476954220924236589456604184053806079897316939839999884039002731864535000644625853;
            5'd13: xpb[41] = 1024'd34664400803899852565604477914023853504204752587250657893959035502840226621207609080792921555547199951105727541114722814395709283215493553521966326095314414663468106114949165975741788608328513978547883148244949626502589503424224331114154215396574365426767716907762976929193704006035095004386077398469497885035;
            5'd14: xpb[41] = 1024'd46874485149132513639789355246242183215658843334403453434119873238826159079555051233931997922486036432686410383312585602778384138912163852604822206950056372786326473859912272384462713823701261647767735514139733432107739530627695185274087506556559274249351380009446056541447568012186151006040290261938351144217;
            5'd15: xpb[41] = 1024'd59084569494365174713974232578460512927112934081556248974280710974812091537902493387071074289424872914267093225510448391161058994608834151687678087804798330909184841604875378793183639039074009316987587880034517237712889557831166039434020797716544183071935043111129136153701432018337207007694503125407204403399;
            5'd16: xpb[41] = 1024'd71294653839597835788159109910678842638567024828709044514441548710798023996249935540210150656363709395847776067708311179543733850305504450770533968659540289032043209349838485201904564254446756986207440245929301043318039585034636893593954088876529091894518706212812215765955296024488263009348715988876057662581;
            5'd17: xpb[41] = 1024'd83504738184830496862343987242897172350021115575861840054602386446783956454597377693349227023302545877428458909906173967926408706002174749853389849514282247154901577094801591610625489469819504655427292611824084848923189612238107747753887380036514000717102369314495295378209160030639319011002928852344910921763;
            5'd18: xpb[41] = 1024'd95714822530063157936528864575115502061475206323014635594763224182769888912944819846488303390241382359009141752104036756309083561698845048936245730369024205277759944839764698019346414685192252324647144977718868654528339639441578601913820671196498909539686032416178374990463024036790375012657141715813764180945;
            5'd19: xpb[41] = 1024'd107924906875295819010713741907333831772929297070167431134924061918755821371292261999627379757180218840589824594301899544691758417395515348019101611223766163400618312584727804428067339900564999993866997343613652460133489666645049456073753962356483818362269695517861454602716888042941431014311354579282617440127;
            5'd20: xpb[41] = 1024'd120134991220528480084898619239552161484383387817320226675084899654741753829639704152766456124119055322170507436499762333074433273092185647101957492078508121523476680329690910836788265115937747663086849709508436265738639693848520310233687253516468727184853358619544534214970752049092487015965567442751470699309;
            5'd21: xpb[41] = 1024'd8278379881636399760284569166956058451139051438737338087113882325750790950678007395890461276400217494308040871240131686878044287947635611629653247916919038712644373505082799907878951139793289610996504467015980224979428870831094391428641974993224186740617118307110555797118087981314910000501090479594729474160;
            5'd22: xpb[41] = 1024'd20488464226869060834469446499174388162593142185890133627274720061736723409025449549029537643339053975888723713437994475260719143644305910712509128771660996835502741250045906316599876355166037280216356832910764030584578898034565245588575266153209095563200781408793635409371951987465966002155303343063582733342;
            5'd23: xpb[41] = 1024'd32698548572101721908654323831392717874047232933042929167435557797722655867372891702168614010277890457469406555635857263643393999340976209795365009626402954958361108995009012725320801570538784949436209198805547836189728925238036099748508557313194004385784444510476715021625815993617022003809516206532435992524;
            5'd24: xpb[41] = 1024'd44908632917334382982839201163611047585501323680195724707596395533708588325720333855307690377216726939050089397833720052026068855037646508878220890481144913081219476739972119134041726785911532618656061564700331641794878952441506953908441848473178913208368107612159794633879679999768078005463729070001289251706;
            5'd25: xpb[41] = 1024'd57118717262567044057024078495829377296955414427348520247757233269694520784067776008446766744155563420630772240031582840408743710734316807961076771335886871204077844484935225542762652001284280287875913930595115447400028979644977808068375139633163822030951770713842874246133544005919134007117941933470142510888;
            5'd26: xpb[41] = 1024'd69328801607799705131208955828047707008409505174501315787918071005680453242415218161585843111094399902211455082229445628791418566430987107043932652190628829326936212229898331951483577216657027957095766296489899253005179006848448662228308430793148730853535433815525953858387408012070190008772154796938995770070;
            5'd27: xpb[41] = 1024'd81538885953032366205393833160266036719863595921654111328078908741666385700762660314724919478033236383792137924427308417174093422127657406126788533045370787449794579974861438360204502432029775626315618662384683058610329034051919516388241721953133639676119096917209033470641272018221246010426367660407849029252;
            5'd28: xpb[41] = 1024'd93748970298265027279578710492484366431317686668806906868239746477652318159110102467863995844972072865372820766625171205556768277824327705209644413900112745572652947719824544768925427647402523295535471028279466864215479061255390370548175013113118548498702760018892113082895136024372302012080580523876702288434;
            5'd29: xpb[41] = 1024'd105959054643497688353763587824702696142771777415959702408400584213638250617457544621003072211910909346953503608823033993939443133520998004292500294754854703695511315464787651177646352862775270964755323394174250669820629088458861224708108304273103457321286423120575192695149000030523358013734793387345555547616;
            5'd30: xpb[41] = 1024'd118169138988730349427948465156921025854225868163112497948561421949624183075804986774142148578849745828534186451020896782322117989217668303375356175609596661818369683209750757586367278078148018633975175760069034475425779115662332078868041595433088366143870086222258272307402864036674414015389006250814408806798;
            5'd31: xpb[41] = 1024'd6312527649838269103334415084324922820981531784529609360590404620633220196843290017266153731130908000671719885761266136125729004073118267903051931448007579007537376385142646657457964102003560581884830517576578434666568292644906160062996316909843825699633845909824293889550199968896836999924529287657667581649;
        endcase
    end

    always_comb begin
        case(flag[14][5:0])
            6'd0: xpb[42] = 1024'd0;
            6'd1: xpb[42] = 1024'd71294653839597835788159109910678842638567024828709044514441548710798023996249935540210150656363709395847776067708311179543733850305504450770533968659540289032043209349838485201904564254446756986207440245929301043318039585034636893593954088876529091894518706212812215765955296024488263009348715988876057662581;
            6'd2: xpb[42] = 1024'd18522611995070930177519292416543252532435622531682404900751242356619152655190732170405230098069744482252402727959128924508403859769788566985907812302749537130395744130105753066178889317376308251104682883471362240271718319848377014222929608069828734522217509011507373501804063975047893001578742151126520840831;
            6'd3: xpb[42] = 1024'd89817265834668765965678402327222095171002647360391449415192791067417176651440667710615380754433453878100178795667440104052137710075293017756441780962289826162438953479944238268083453571823065237312123129400663283589757904883013907816883696946357826416736215224319589267759359999536156010927458140002578503412;
            6'd4: xpb[42] = 1024'd37045223990141860355038584833086505064871245063364809801502484713238305310381464340810460196139488964504805455918257849016807719539577133971815624605499074260791488260211506132357778634752616502209365766942724480543436639696754028445859216139657469044435018023014747003608127950095786003157484302253041681662;
            6'd5: xpb[42] = 1024'd108339877829739696143197694743765347703438269892073854315944033424036329306631399881020610852503198360352581523626569028560541569845081584742349593265039363292834697610049991334262342889199373488416806012872025523861476224731390922039813305016186560938953724235826962769563423974584049012506200291129099344243;
            6'd6: xpb[42] = 1024'd55567835985212790532557877249629757597306867595047214702253727069857457965572196511215690294209233446757208183877386773525211579309365700957723436908248611391187232390317259198536667952128924753314048650414086720815154959545131042668788824209486203566652527034522120505412191925143679004736226453379562522493;
            6'd7: xpb[42] = 1024'd2795794140685884921918059755494167491175465298020575088563420715678586624512993141410769735915268533161834844128204518489881588773649817173097280551457859489539767170584527062810993015058476018211291287956147917768833694358871163297764343402785846194351329833217278241260959875703308996966252615630025700743;
            6'd8: xpb[42] = 1024'd74090447980283720710077169666173010129742490126729619603004969426476610620762928681620920392278977929009610911836515698033615439079154267943631249210998148521582976520423012264715557269505233004418731533885448961086873279393508056891718432279314938088870036046029494007216255900191572006314968604506083363324;
            6'd9: xpb[42] = 1024'd21318406135756815099437352172037420023611087829702979989314663072297739279703725311815999833985013015414237572087333442998285448543438384159005092854207396619935511300690280128989882332434784269315974171427510158040552014207248177520693951472614580716568838844724651743065023850751201998544994766756546541574;
            6'd10: xpb[42] = 1024'd92613059975354650887596462082716262662178112658412024503756211783095763275953660852026150490348722411262013639795644622542019298848942834929539061513747685651978720650528765330894446586881541255523414417356811201358591599241885071114648040349143672611087545057536867509020319875239465007893710755632604204155;
            6'd11: xpb[42] = 1024'd39841018130827745276956644588580672556046710361385384890065905428916891934894457482221229932054757497666640300046462367506689308313226951144912905156956933750331255430796033195168771649811092520420657054898872398312270334055625191743623559542443315238786347856232025244869087825799095000123736917883067382405;
            6'd12: xpb[42] = 1024'd111135671970425581065115754499259515194613735190094429404507454139714915931144393022431380588418466893514416367754773547050423158618731401915446873816497222782374464780634518397073335904257849506628097300828173441630309919090262085337577648418972407133305054069044241010824383850287358009472452906759125044986;
            6'd13: xpb[42] = 1024'd58363630125898675454475937005123925088482332893067789790817147785536044590085189652626460030124501979919043028005591292015093168083015518130820717459706470880726999560901786261347660967187400771525339938370234638583988653904002205966553167612272049761003856867739398746673151800846988001702479069009588223236;
            6'd14: xpb[42] = 1024'd5591588281371769843836119510988334982350930596041150177126841431357173249025986282821539471830537066323669688256409036979763177547299634346194561102915718979079534341169054125621986030116952036422582575912295835537667388717742326595528686805571692388702659666434556482521919751406617993932505231260051401486;
            6'd15: xpb[42] = 1024'd76886242120969605631995229421667177620917955424750194691568390142155197245275921823031690128194246462171445755964720216523497027852804085116728529762456008011122743691007539327526550284563709022630022821841596878855706973752379220189482775682100784283221365879246772248477215775894881003281221220136109064067;
            6'd16: xpb[42] = 1024'd24114200276442700021355411927531587514786553127723555077878083787976325904216718453226769569900281548576072416215537961488167037317088201332102373405665256109475278471274807191800875347493260287527265459383658075809385708566119340818458294875400426910920168677941929984325983726454510995511247382386572242317;
            6'd17: xpb[42] = 1024'd95408854116040535809514521838210430153353577956432599592319632498774349900466653993436920226263990944423848483923849141031900887622592652102636342065205545141518487821113292393705439601940017273734705705312959119127425293600756234412412383751929518805438874890754145750281279750942774004859963371262629904898;
            6'd18: xpb[42] = 1024'd42636812271513630198874704344074840047222175659405959978629326144595478559407450623631999667970026030828475144174666885996570897086876768318010185708414793239871022601380560257979764664869568538631948342855020316081104028414496355041387902945229161433137677689449303486130047701502403997089989533513093083148;
            6'd19: xpb[42] = 1024'd113931466111111465987033814254753682685789200488115004493070874855393502555657386163842150324333735426676251211882978065540304747392381219088544154367955082271914231951219045459884328919316325524839388588784321359399143613449133248635341991821758253327656383902261519252085343725990667006438705522389150745729;
            6'd20: xpb[42] = 1024'd61159424266584560376393996760618092579657798191088364879380568501214631214598182794037229766039770513080877872133795810504974756856665335303917998011164330370266766731486313324158653982245876789736631226326382556352822348262873369264317511015057895955355186700956676987934111676550296998668731684639613923979;
            6'd21: xpb[42] = 1024'd8387382422057654765754179266482502473526395894061725265690262147035759873538979424232309207745805599485504532384613555469644766320949451519291841654373578468619301511753581188432979045175428054633873863868443753306501083076613489893293030208357538583053989499651834723782879627109926990898757846890077102229;
            6'd22: xpb[42] = 1024'd79682036261655490553913289177161345112093420722770769780131810857833783869788914964442459864109514995333280600092924735013378616626453902289825810313913867500662510861592066390337543299622185040841314109797744796624540668111250383487247119084886630477572695712464050489738175651598190000247473835766134764810;
            6'd23: xpb[42] = 1024'd26909994417128584943273471683025755005962018425744130166441504503654912528729711594637539305815550081737907260343742479978048626090738018505199653957123115599015045641859334254611868362551736305738556747339805993578219402924990504116222638278186273105271498511159208225586943602157819992477499998016597943060;
            6'd24: xpb[42] = 1024'd98204648256726420731432581593704597644529043254453174680883053214452936524979647134847689962179259477585683328052053659521782476396242469275733622616663404631058254991697819456516432616998493291945996993269107036896258987959627397710176727154715364999790204723971423991542239626646083001826215986892655605641;
            6'd25: xpb[42] = 1024'd45432606412199515120792764099569007538397640957426535067192746860274065183920443765042769403885294563990309988302871404486452485860526585491107466259872652729410789771965087320790757679928044556843239630811168233849937722773367518339152246348015007627489007522666581727391007577205712994056242149143118783891;
            6'd26: xpb[42] = 1024'd116727260251797350908951874010247850176964665786135579581634295571072089180170379305252920060249003959838086056011182584030186336166031036261641434919412941761453999121803572522695321934374801543050679876740469277167977307808004411933106335224544099522007713735478797493346303601693976003404958138019176446472;
            6'd27: xpb[42] = 1024'd63955218407270445298312056516112260070833263489108939967943989216893217839111175935447999501955039046242712716262000328994856345630315152477015278562622189859806533902070840386969646997304352807947922514282530474121656042621744532562081854417843742149706516534173955229195071552253605995634984300269639624722;
            6'd28: xpb[42] = 1024'd11183176562743539687672239021976669964701861192082300354253682862714346498051972565643078943661074132647339376512818073959526355094599268692389122205831437958159068682338108251243972060233904072845165151824591671075334777435484653191057373611143384777405319332869112965043839502813235987865010462520102802972;
            6'd29: xpb[42] = 1024'd82477830402341375475831348932655512603268886020791344868695231573512370494301908105853229600024783528495115444221129253503260205400103719462923090865371726990202278032176593453148536314680661059052605397753892714393374362470121546785011462487672476671924025545681328730999135527301498997213726451396160465553;
            6'd30: xpb[42] = 1024'd29705788557814469865191531438519922497137483723764705255004925219333499153242704736048309041730818614899742104471946998467930214864387835678296934508580975088554812812443861317422861377610212323949848035295953911347053097283861667413986981680972119299622828344376486466847903477861128989443752613646623643803;
            6'd31: xpb[42] = 1024'd101000442397412305653350641349198765135704508552473749769446473930131523149492640276258459698094528010747518172180258178011664065169892286448830903168121264120598022162282346519327425632056969310157288281225254954665092682318498561007941070557501211194141534557188702232803199502349391998792468602522681306384;
            6'd32: xpb[42] = 1024'd48228400552885400042710823855063175029573106255447110155756167575952651808433436906453539139800563097152144832431075922976334074634176402664204746811330512218950556942549614383601750694986520575054530918767316151618771417132238681636916589750800853821840337355883859968651967452909021991022494764773144484634;
            6'd33: xpb[42] = 1024'd119523054392483235830869933765742017668140131084156154670197716286750675804683372446663689796164272492999920900139387102520067924939680853434738715470870801250993766292388099585506314949433277561261971164696617194936811002166875575230870678627329945716359043568696075734607263477397285000371210753649202147215;
            6'd34: xpb[42] = 1024'd66751012547956330220230116271606427562008728787129515056507409932571804463624169076858769237870307579404547560390204847484737934403964969650112559114080049349346301072655367449780640012362828826159213802238678391890489736980615695859846197820629588344057846367391233470456031427956914992601236915899665325465;
            6'd35: xpb[42] = 1024'd13978970703429424609590298777470837455877326490102875442817103578392933122564965707053848679576342665809174220641022592449407943868249085865486402757289297447698835852922635314054965075292380091056456439780739588844168471794355816488821717013929230971756649166086391206304799378516544984831263078150128503715;
            6'd36: xpb[42] = 1024'd85273624543027260397749408688149680094444351318811919957258652289190957118814901247263999335940052061656950288349333771993141794173753536636020371416829586479742045202761120515959529329739137077263896685710040632162208056828992710082775805890458322866275355378898606972260095403004807994179979067026186166296;
            6'd37: xpb[42] = 1024'd32501582698500354787109591194014089988312949021785280343568345935012085777755697877459078777646087148061576948600151516957811803638037652851394215060038834578094579983028388380233854392668688342161139323252101829115886791642732830711751325083757965493974158177593764708108863353564437986410005229276649344546;
            6'd38: xpb[42] = 1024'd103796236538098190575268701104692932626879973850494324858009894645810109774005633417669229434009796543909353016308462696501545653943542103621928183719579123610137789332866873582138418647115445328368579569181402872433926376677369724305705413960287057388492864390405980474064159378052700995758721218152707007127;
            6'd39: xpb[42] = 1024'd51024194693571284964628883610557342520748571553467685244319588291631238432946430047864308875715831630313979676559280441466215663407826219837302027362788371708490324113134141446412743710044996593265822206723464069387605111491109844934680933153586700016191667189101138209912927328612330987988747380403170185377;
            6'd40: xpb[42] = 1024'd122318848533169120752787993521236185159315596382176729758761137002429262429196365588074459532079541026161755744267591621009949513713330670607835996022328660740533533462972626648317307964491753579473262452652765112705644696525746738528635022030115791910710373401913353975868223353100593997337463369279227847958;
            6'd41: xpb[42] = 1024'd69546806688642215142148176027100595053184194085150090145070830648250391088137162218269538973785576112566382404518409365974619523177614786823209839665537908838886068243239894512591633027421304844370505090194826309659323431339486859157610541223415434538409176200608511711716991303660223989567489531529691026208;
            6'd42: xpb[42] = 1024'd16774764844115309531508358532965004947052791788123450531380524294071519747077958848464618415491611198971009064769227110939289532641898903038583683308747156937238603023507162376865958090350856109267747727736887506613002166153226979786586060416715077166107978999303669447565759254219853981797515693780154204458;
            6'd43: xpb[42] = 1024'd88069418683713145319667468443643847585619816616832495045822073004869543743327894388674769071855320594818785132477538290483023382947403353809117651968287445969281812373345647578770522344797613095475187973666188549931041751187863873380540149293244169060626685212115885213521055278708116991146231682656211867039;
            6'd44: xpb[42] = 1024'd35297376839186239709027650949508257479488414319805855432131766650690672402268691018869848513561355681223411792728356035447693392411687470024491495611496694067634347153612915443044847407727164360372430611208249746884720486001603994009515668486543811688325488010811042949369823229267746983376257844906675045289;
            6'd45: xpb[42] = 1024'd106592030678784075497186760860187100118055439148514899946573315361488696398518626559079999169925065077071187860436667214991427242717191920795025464271036983099677556503451400644949411662173921346579870857137550790202760071036240887603469757363072903582844194223623258715325119253756009992724973833782732707870;
            6'd46: xpb[42] = 1024'd53819988834257169886546943366051510011924036851488260332883009007309825057459423189275078611631100163475814520687484959956097252181476037010399307914246231198030091283718668509223736725103472611477113494679611987156438805849981008232445276556372546210542997022318416451173887204315639984954999996033195886120;
            6'd47: xpb[42] = 1024'd1047946989730264275907125871915919905792634554461620719192702653130953716400219819470158053337135249880441180938302704920767261645760153225773151557455479296382626063985936373498061788033023876374356132221673184110117540663721128861420795749672188838241799821013574187022655154875269977185026158283659064370;
            6'd48: xpb[42] = 1024'd72342600829328100064066235782594762544359659383170665233634251363928977712650155359680308709700844645728217248646613884464501111951264603996307120216995768328425835413824421575402626042479780862581796378150974227428157125698358022455374884626201280732760506033825789952977951179363532986533742147159716726951;
            6'd49: xpb[42] = 1024'd19570558984801194453426418288459172438228257086144025619943945009750106371590951989875388151406879732132843908897431629429171121415548720211680963860205016426778370194091689439676951105409332127479039015693035424381835860512098143084350403819500923360459308832520947688826719129923162978763768309410179905201;
            6'd50: xpb[42] = 1024'd90865212824399030241585528199138015076795281914853070134385493720548130367840887530085538807770589127980619976605742808972904971721053170982214932519745305458821579543930174641581515359856089113686479261622336467699875445546735036678304492696030015254978015045333163454782015154411425988112484298286237567782;
            6'd51: xpb[42] = 1024'd38093170979872124630945710705002424970663879617826430520695187366369259026781684160280618249476624214385246636856560553937574981185337287197588776162954553557174114324197442505855840422785640378583721899164397664653554180360475157307280011889329657882676817844028321190630783104971055980342510460536700746032;
            6'd52: xpb[42] = 1024'd109387824819469960419104820615681267609230904446535475035136736077167283023031619700490768905840333610233022704564871733481308831490841737968122744822494842589217323674035927707760404677232397364791162145093698707971593765395112050901234100765858749777195524056840536956586079129459318989691226449412758408613;
            6'd53: xpb[42] = 1024'd56615782974943054808465003121545677503099502149508835421446429722988411681972416330685848347546368696637649364815689478445978840955125854183496588465704090687569858454303195572034729740161948629688404782635759904925272500208852171530209619959158392404894326855535694692434847080018948981921252611663221586863;
            6'd54: xpb[42] = 1024'd3843741130416149197825185627410087396968099852482195807756123368809540340913212960880927789252403783042276025066507223410648850419409970398870432108913338785922393234570463436309054803091499894585647420177821101878951235022592292159185139152458035032593129654230852428283615030578578974151278773913684765113;
            6'd55: xpb[42] = 1024'd75138394970013984985984295538088930035535124681191240322197672079607564337163148501091078445616113178890052092774818402954382700724914421169404400768453627817965602584408948638213619057538256880793087666107122145196990820057229185753139228028987126927111835867043068194238911055066841983499994762789742427694;
            6'd56: xpb[42] = 1024'd22366353125487079375344478043953339929403722384164600708507365725428692996103945131286157887322148265294678753025636147919052710189198537384778244411662875916318137364676216502487944120467808145690330303649183342150669554870969306382114747222286769554810638665738225930087679005626471975730020925040205605944;
            6'd57: xpb[42] = 1024'd93661006965084915163503587954632182567970747212873645222948914436226716992353880671496308543685857661142454820733947327462786560494702988155312213071203164948361346714514701704392508374914565131897770549578484385468709139905606199976068836098815861449329344878550441696042975030114734985078736913916263268525;
            6'd58: xpb[42] = 1024'd40888965120558009552863770460496592461839344915847005609258608082047845651294677301691387985391892747547081480984765072427456569958987104370686056714412413046713881494781969568666833437844116396795013187120545582422387874719346320605044355292115504077028147677245599431891742980674364977308763076166726446775;
            6'd59: xpb[42] = 1024'd112183618960155845341022880371175435100406369744556050123700156792845869647544612841901538641755602143394857548693076251971190420264491555141220025373952702078757090844620454770571397692290873383002453433049846625740427459753983214198998444168644595971546853890057815197847039005162627986657479065042784109356;
            6'd60: xpb[42] = 1024'd59411577115628939730383062877039844994274967447529410510009850438666998306485409472096618083461637229799484208943893996935860429728775671356593869017161950177109625624887722634845722755220424647899696070591907822694106194567723334827973963361944238599245656688752972933695806955722257978887505227293247287606;
            6'd61: xpb[42] = 1024'd6639535271102034119743245382904254888143565150502770896319544084488126965426206102291697525167672316204110869194711741900530439193059787571967712660371198275462160405154990499120047818149975912796938708133969019647784929381463455456949482555243881226944459487448130669544574906281887971117531389543710465856;
            6'd62: xpb[42] = 1024'd77934189110699869907902355293583097526710589979211815410761092795286150961676141642501848181531381712051886936903022921444264289498564238342501681319911487307505369754993475701024612072596732899004378954063270062965824514416100349050903571431772973121463165700260346435499870930770150980466247378419768128437;
            6'd63: xpb[42] = 1024'd25162147266172964297262537799447507420579187682185175797070786441107279620616938272696927623237416798456513597153840666408934298962848354557875524963120735405857904535260743565298937135526284163901621591605331259919503249229840469679879090625072615749161968498955504171348638881329780972696273540670231306687;
        endcase
    end

    always_comb begin
        case(flag[14][11:6])
            6'd0: xpb[43] = 1024'd0;
            6'd1: xpb[43] = 1024'd96456801105770800085421647710126350059146212510894220311512335151905303616866873812907078279601126194304289664862151845952668149268352805328409493622661024437901113885099228767203501389973041150109061837534632303237542834264477363273833179501601707643680674711767719937303934905818043982044989529546288969268;
            6'd2: xpb[43] = 1024'd68846906527416858772044368015438267373593997896052756494892815238833711896424608715799085344544578079165429922266810257326272457695485276101658862228991007942111553200627240196776763588428876578907926066682024760110724818308057953582687789319973966020541446009418381844501341737707454946971289232466983454205;
            6'd3: xpb[43] = 1024'd41237011949062917458667088320750184688041783281211292678273295325762120175982343618691092409488029964026570179671468668699876766122617746874908230835320991446321992516155251626350025786884712007706790295829417216983906802351638543891542399138346224397402217307069043751698748569596865911897588935387677939142;
            6'd4: xpb[43] = 1024'd13627117370708976145289808626062102002489568666369828861653775412690528455540078521583099474431481848887710437076127080073481074549750217648157599441650974950532431831683263055923287985340547436505654524976809673857088786395219134200397008956718482774262988604719705658896155401486276876823888638308372424079;
            6'd5: xpb[43] = 1024'd110083918476479776230711456336188452061635781177264049173166110564595832072406952334490177754032608043192000101938278926026149223818103022976567093064311999388433545716782491823126789375313588586614716362511441977094631620659696497474230188458320190417943663316487425596200090307304320858868878167854661393347;
            6'd6: xpb[43] = 1024'd82474023898125834917334176641500369376083566562422585356546590651524240351964687237382184818976059928053140359342937337399753532245235493749816461670641982892643985032310503252700051573769424015413580591658834433967813604703277087783084798276692448794804434614138087503397497139193731823795177870775355878284;
            6'd7: xpb[43] = 1024'd54864129319771893603956896946812286690531351947581121539927070738452648631522422140274191883919511812914280616747595748773357840672367964523065830276971966396854424347838514682273313772225259444212444820806226890840995588746857678091939408095064707171665205911788749410594903971083142788721477573696050363221;
            6'd8: xpb[43] = 1024'd27254234741417952290579617252124204004979137332739657723307550825381056911080157043166198948862963697775420874152254160146962149099500435296315198883301949901064863663366526111846575970681094873011309049953619347714177572790438268400794017913436965548525977209439411317792310802972553753647777276616744848158;
            6'd9: xpb[43] = 1024'd123711035847188752376001264962250554064125349843633878034819885977286360527947030856073277228464089892079710539014406006099630298367853240624724692505962974338965977548465754879050077360654136023120370887488251650951720407054915631674627197415038673192206651921207131255096245708790597735692766806163033817426;
            6'd10: xpb[43] = 1024'd96101141268834811062623985267562471378573135228792414218200366064214768807504765758965284293407541776940850796419064417473234606794985711397974061112292957843176416863993766308623339559109971451919235116635644107824902391098496221983481807233410931569067423218857793162293652540680008700619066509083728302363;
            6'd11: xpb[43] = 1024'd68491246690480869749246705572874388693020920613950950401580846151143177087062500661857291358350993661801991053823722828846838915222118182171223429718622941347386856179521777738196601757565806880718099345783036564698084375142076812292336417051783189945928194516508455069491059372569419665545366212004422787300;
            6'd12: xpb[43] = 1024'd40881352112126928435869425878186306007468705999109486584961326238071585366620235564749298423294445546663131311228381240220443223649250652944472798324952924851597295495049789167769863956021642309516963574930429021571266359185657402601191026870155448322788965814159116976688466204458830630471665914925117272237;
            6'd13: xpb[43] = 1024'd13271457533772987122492146183498223321916491384268022768341806324999993646177970467641305488237897431524271568633039651594047532076383123717722166931282908355807734810577800597343126154477477738315827804077821478444448343229237992910045636688527706699649737111809778883885873036348241595397965617845811757174;
            6'd14: xpb[43] = 1024'd109728258639543787207913793893624573381062703895162243079854141476905297263044844280548383767839023625828561233495191497546715681344735929046131660553943932793708848695677029364546627544450518888424889641612453781681991177493715356183878816190129414343330411823577498821189807942166285577442955147392100726442;
            6'd15: xpb[43] = 1024'd82118364061189845894536514198936490695510489280320779263234621563833705542602579183440390832782475510689701490899849908920319989771868399819381029160273916297919288011205040794119889742906354317223753870759846238555173161537295946492733426008501672720191183121228160728387214774055696542369254850312795211379;
            6'd16: xpb[43] = 1024'd54508469482835904581159234504248408009958274665479315446615101650762113822160314086332397897725927395550841748304508320293924298199000870592630397766603899802129727326733052223693151941362189746022618099907238695428355145580876536801588035826873931097051954418878822635584621605945107507295554553233489696316;
            6'd17: xpb[43] = 1024'd26898574904481963267781954809560325324406060050637851629995581737690522101718048989224404962669379280411982005709166731667528606626133341365879766372933883306340166642261063653266414139818025174821482329054631152301537129624457127110442645645246189473912725716529484542782028437834518472221854256154184181253;
            6'd18: xpb[43] = 1024'd123355376010252763353203602519686675383552272561532071941507916889595825718584922802131483242270505474716271670571318577620196755894486146694289259995594907744241280527360292420469915529791066324930544166589263455539079963888934490384275825146847897117593400428297204480085963343652562454266843785700473150521;
            6'd19: xpb[43] = 1024'd95745481431898822039826322824998592698000057946690608124888396976524233998142657705023490307213957359577411927975976988993801064321618617467538628601924891248451719842888303850043177728246901753729408395736655912412261947932515080693130434965220155494454171725947866387283370175541973419193143488621167635458;
            6'd20: xpb[43] = 1024'd68135586853544880726449043130310510012447843331849144308268877063452642277700392607915497372157409244438552185380635400367405372748751088240787997208254874752662159158416315279616439926702737182528272624884048369285443931976095671001985044783592413871314943023598528294480777007431384384119443191541862120395;
            6'd21: xpb[43] = 1024'd40525692275190939413071763435622427326895628717007680491649357150381050557258127510807504437100861129299692442785293811741009681175883559014037365814584858256872598473944326709189702125158572611327136854031440826158625916019676261310839654601964672248175714321249190201678183839320795349045742894462556605332;
            6'd22: xpb[43] = 1024'd12915797696836998099694483740934344641343414102166216675029837237309458836815862413699511502044313014160832700189952223114613989603016029787286734420914841761083037789472338138762964323614408040126001083178833283031807900063256851619694264420336930625036485618899852108875590671210206313972042597383251090269;
            6'd23: xpb[43] = 1024'd109372598802607798185116131451060694700489626613060436986542172389214762453682736226606589781645439208465122365052104069067282138871368835115696228043575866198984151674571566905966465713587449190235062920713465586269350734327734214893527443921938638268717160330667572046179525577028250296017032126929540059537;
            6'd24: xpb[43] = 1024'd81762704224253856871738851756372612014937411998218973169922652476143170733240471129498596846588891093326262622456762480440886447298501305888945596649905849703194590990099578335539727912043284619033927149860858043142532718371314805202382053740310896645577931628318233953376932408917661260943331829850234544474;
            6'd25: xpb[43] = 1024'd54152809645899915558361572061684529329385197383377509353303132563071579012798206032390603911532342978187402879861420891814490755725633776662194965256235833207405030305627589765112990110499120047832791379008250500015714702414895395511236663558683155022438702925968895860574339240807072225869631532770929029411;
            6'd26: xpb[43] = 1024'd26542915067545974244984292366996446643832982768536045536683612649999987292355940935282610976475794863048543137266079303188095064152766247435444333862565816711615469621155601194686252308954955476631655608155642956888896686458475985820091273377055413399299474223619557767771746072696483190795931235691623514348;
            6'd27: xpb[43] = 1024'd122999716173316774330405940077122796702979195279430265848195947801905290909222814748189689256076921057352832802128231149140763213421119052763853827485226841149516583506254829961889753698927996626740717445690275260126439520722953349093924452878657121042980148935387277705075680978514527172840920765237912483616;
            6'd28: xpb[43] = 1024'd95389821594962833017028660382434714017426980664588802031576427888833699188780549651081696321020372942213973059532889560514367521848251523537103196091556824653727022821782841391463015897383832055539581674837667716999621504766533939402779062697029379419840920233037939612273087810403938137767220468158606968553;
            6'd29: xpb[43] = 1024'd67779927016608891703651380687746631331874766049747338214956907975762107468338284553973703385963824827075113316937547971887971830275383994310352564697886808157937462137310852821036278095839667484338445903985060173872803488810114529711633672515401637796701691530688601519470494642293349102693520171079301453490;
            6'd30: xpb[43] = 1024'd40170032438254950390274100993058548646322551434905874398337388062690515747896019456865710450907276711936253574342206383261576138702516465083601933304216791662147901452838864250609540294295502913137310133132452630745985472853695120020488282333773896173562462828339263426667901474182760067619819873999995938427;
            6'd31: xpb[43] = 1024'd12560137859901009076896821298370465960770336820064410581717868149618924027453754359757717515850728596797393831746864794635180447129648935856851301910546775166358340768366875680182802492751338341936174362279845087619167456897275710329342892152146154550423234125989925333865308306072171032546119576920690423364;
            6'd32: xpb[43] = 1024'd109016938965671809162318469008496816019916549330958630893230203301524227644320628172664795795451854791101683496609016640587848596398001741185260795533207799604259454653466104447386303882724379492045236199814477390856710291161753073603176071653747862194103908837757645271169243211890215014591109106466979392632;
            6'd33: xpb[43] = 1024'd81407044387317867848941189313808733334364334716117167076610683388452635923878363075556802860395306675962823754013675051961452904825134211958510164139537783108469893968994115876959566081180214920844100428961869847729892275205333663912030681472120120570964680135408307178366650043779625979517408809387673877569;
            6'd34: xpb[43] = 1024'd53797149808963926535563909619120650648812120101275703259991163475381044203436097978448809925338758560823964011418333463335057213252266682731759532745867766612680333284522127306532828279636050349642964658109262304603074259248914254220885291290492378947825451433058969085564056875669036944443708512308368362506;
            6'd35: xpb[43] = 1024'd26187255230609985222186629924432567963259905486434239443371643562309452482993832881340816990282210445685104268822991874708661521679399153505008901352197750116890772600050138736106090478091885778441828887256654761476256243292494844529739901108864637324686222730709630992761463707558447909370008215229062847443;
            6'd36: xpb[43] = 1024'd122644056336380785307608277634558918022406117997328459754883978714214756099860706694247895269883336639989393933685143720661329670947751958833418394974858774554791886485149367503309591868064926928550890724791287064713799077556972207803573080610466344968366897442477350930065398613376491891414997744775351816711;
            6'd37: xpb[43] = 1024'd95034161758026843994230997939870835336853903382486995938264458801143164379418441597139902334826788524850534191089802132034933979374884429606667763581188758059002325800677378932882854066520762357349754953938679521586981061600552798112427690428838603345227668740128012837262805445265902856341297447696046301648;
            6'd38: xpb[43] = 1024'd67424267179672902680853718245182752651301688767645532121644938888071572658976176500031909399770240409711674448494460543408538287802016900379917132187518741563212765116205390362456116264976597786148619183086071978460163045644133388421282300247210861722088440037778674744460212277155313821267597150616740786585;
            6'd39: xpb[43] = 1024'd39814372601318961367476438550494669965749474152804068305025418974999980938533911402923916464713692294572814705899118954782142596229149371153166500793848725067423204431733401792029378463432433214947483412233464435333345029687713978730136910065583120098949211335429336651657619109044724786193896853537435271522;
            6'd40: xpb[43] = 1024'd12204478022965020054099158855806587280197259537962604488405899061928389218091646305815923529657144179433954963303777366155746904656281841926415869400178708571633643747261413221602640661888268643746347641380856892206527013731294569038991519883955378475809982633079998558855025940934135751120196556458129756459;
            6'd41: xpb[43] = 1024'd108661279128735820139520806565932937339343472048856824799918234213833692834958520118723001809258270373738244628165929212108415053924634647254825363022839733009534757632360641988806142051861309793855409478915489195444069847995771932312824699385557086119490657344847718496158960846752179733165186086004418725727;
            6'd42: xpb[43] = 1024'd81051384550381878826143526871244854653791257434015360983298714300762101114516255021615008874201722258599384885570587623482019362351767118028074731629169716513745196947888653418379404250317145222654273708062881652317251832039352522621679309203929344496351428642498380403356367678641590698091485788925113210664;
            6'd43: xpb[43] = 1024'd53441489972027937512766247176556771968239042819173897166679194387690509394073989924507015939145174143460525142975246034855623670778899588801324100235499700017955636263416664847952666448772980651453137937210274109190433816082933112930533919022301602873212199940149042310553774510531001663017785491845807695601;
            6'd44: xpb[43] = 1024'd25831595393673996199388967481868689282686828204332433350059674474618917673631724827399023004088626028321665400379904446229227979206032059574573468841829683522166075578944676277525928647228816080252002166357666566063615800126513703239388528840673861250072971237799704217751181342420412627944085194766502180538;
            6'd45: xpb[43] = 1024'd122288396499444796284810615191995039341833040715226653661572009626524221290498598640306101283689752222625955065242056292181896128474384864902982962464490707960067189464043905044729430037201857230361064003892298869301158634390991066513221708342275568893753645949567424155055116248238456609989074724312791149806;
            6'd46: xpb[43] = 1024'd94678501921090854971433335497306956656280826100385189844952489713452629570056333543198108348633204107487095322646714703555500436901517335676232331070820691464277628779571916474302692235657692659159928233039691326174340618434571656822076318160647827270614417247218086062252523080127867574915374427233485634743;
            6'd47: xpb[43] = 1024'd67068607342736913658056055802618873970728611485543726028332969800381037849614068446090115413576655992348235580051373114929104745328649806449481699677150674968488068095099927903875954434113528087958792462187083783047522602478152247130930927979020085647475188544868747969449929912017278539841674130154180119680;
            6'd48: xpb[43] = 1024'd39458712764382972344678776107930791285176396870702262211713449887309446129171803348982122478520107877209375837456031526302709053755782277222731068283480658472698507410627939333449216632569363516757656691334476239920704586521732837439785537797392344024335959842519409876647336743906689504767973833074874604617;
            6'd49: xpb[43] = 1024'd11848818186029031031301496413242708599624182255860798395093929974237854408729538251874129543463559762070516094860689937676313362182914747995980436889810641976908946726155950763022478831025198945556520920481868696793886570565313427748640147615764602401196731140170071783844743575796100469694273535995569089554;
            6'd50: xpb[43] = 1024'd108305619291799831116723144123369058658770394766755018706606265126143158025596412064781207823064685956374805759722841783628981511451267553324389930512471666414810060611255179530225980220998240095665582758016501000031429404829790791022473327117366310044877405851937791721148678481614144451739263065541858058822;
            6'd51: xpb[43] = 1024'd80695724713445889803345864428680975973218180151913554889986745213071566305154146967673214888008137841235946017127500195002585819878400024097639299118801649919020499926783190959799242419454075524464446987163893456904611388873371381331327936935738568421738177149588453628346085313503555416665562768462552543759;
            6'd52: xpb[43] = 1024'd53085830135091948489968584733992893287665965537072091073367225299999974584711881870565221952951589726097086274532158606376190128305532494870888667725131633423230939242311202389372504617909910953263311216311285913777793372916951971640182546754110826798598948447239115535543492145392966381591862471383247028696;
            6'd53: xpb[43] = 1024'd25475935556738007176591305039304810602113750922230627256747705386928382864269616773457229017895041610958226531936817017749794436732664965644138036331461616927441378557839213818945766816365746382062175445458678370650975356960532561949037156572483085175459719744889777442740898977282377346518162174303941513633;
            6'd54: xpb[43] = 1024'd121932736662508807262012952749431160661259963433124847568260040538833686481136490586364307297496167805262516196798968863702462586001017770972547529954122641365342492442938442586149268206338787532171237282993310673888518191225009925222870336074084792819140394456657497380044833883100421328563151703850230482901;
            6'd55: xpb[43] = 1024'd94322842084154865948635673054743077975707748818283383751640520625762094760694225489256314362439619690123656454203627275076066894428150241745796898560452624869552931758466454015722530404794622960970101512140703130761700175268590515531724945892457051196001165754308159287242240714989832293489451406770924967838;
            6'd56: xpb[43] = 1024'd66712947505800924635258393360054995290155534203441919935021000712690503040251960392148321427383071574984796711608285686449671202855282712519046267166782608373763371073994465445295792603250458389768965741288095587634882159312171105840579555710829309572861937051958821194439647546879243258415751109691619452775;
            6'd57: xpb[43] = 1024'd39103052927446983321881113665366912604603319588600456118401480799618911319809695295040328492326523459845936969012944097823275511282415183292295635773112591877973810389522476874869054801706293818567829970435488044508064143355751696149434165529201567949722708349609483101637054378768654223342050812612313937712;
            6'd58: xpb[43] = 1024'd11493158349093042008503833970678829919051104973758992301781960886547319599367430197932335557269975344707077226417602509196879819709547654065545004379442575382184249705050488304442317000162129247366694199582880501381246127399332286458288775347573826326583479647260145008834461210658065188268350515533008422649;
            6'd59: xpb[43] = 1024'd107949959454863842093925481680805179978197317484653212613294296038452623216234304010839413836871101539011366891279754355149547968977900459393954498002103599820085363590149717071645818390135170397475756037117512804618788961663809649732121954849175533970264154359027864946138396116476109170313340045079297391917;
            6'd60: xpb[43] = 1024'd80340064876509900780548201986117097292645102869811748796674776125381031495792038913731420901814553423872507148684412766523152277405032930167203866608433583324295802905677728501219080588591005826274620266264905261491970945707390240040976564667547792347124925656678526853335802948365520135239639747999991876854;
            6'd61: xpb[43] = 1024'd52730170298155959467170922291429014607092888254970284980055256212309439775349773816623427966758005308733647406089071177896756585832165400940453235214763566828506242221205739930792342787046841255073484495412297718365152929750970830349831174485920050723985696954329188760533209780254931100165939450920686361791;
            6'd62: xpb[43] = 1024'd25120275719802018153793642596740931921540673640128821163435736299237848054907508719515435031701457193594787663493729589270360894259297871713702603821093550332716681536733751360365604985502676683872348724559690175238334913794551420658685784304292309100846468251979850667730616612144342065092239153841380846728;
            6'd63: xpb[43] = 1024'd121577076825572818239215290306867281980686886151023041474948071451143151671774382532422513311302583387899077328355881435223029043527650677042112097443754574770617795421832980127569106375475717833981410562094322478475877748059028783932518963805894016744527142963747570605034551517962386047137228683387669815996;
        endcase
    end

    always_comb begin
        case(flag[14][16:12])
            5'd0: xpb[44] = 1024'd0;
            5'd1: xpb[44] = 1024'd93967182247218876925838010612179199295134671536181577658328551538071559951332117435314520376246035272760217585760539846596633351954783147815361466050084558274828234737360991557142368573931553262780274791241714935349059732102609374241373573624266275121387914261398232512231958349851797012063528386308364300933;
            5'd2: xpb[44] = 1024'd63867668810313012452877093819543965845570915946627471188525248011166224565355095960613969537834396236077285764063586258614202863068345961075562807083838075615965794905150765776654497956345900804250351974096190024333758613984321975517768577565303100975955925108679406994357388625774961007008366945991134117535;
            5'd3: xpb[44] = 1024'd33768155373407147979916177026908732396007160357073364718721944484260889179378074485913418699422757199394353942366632670631772374181908774335764148117591592957103355072940539996166627338760248345720429156950665113318457495866034576794163581506339926830523935955960581476482818901698125001953205505673903934137;
            5'd4: xpb[44] = 1024'd3668641936501283506955260234273498946443404767519258248918640957355553793401053011212867861011118162711422120669679082649341885295471587595965489151345110298240915240730314215678756721174595887190506339805140202303156377747747178070558585447376752685091946803241755958608249177621288996898044065356673750739;
            5'd5: xpb[44] = 1024'd97635824183720160432793270846452698241578076303700835907247192495427113744733170446527388237257153435471639706430218929245975237250254735411326955201429668573069149978091305772821125295106149149970781131046855137652216109850356552311932159071643027806479861064639988470840207527473086008961572451665038051672;
            5'd6: xpb[44] = 1024'd67536310746814295959832354053817464792014320714146729437443888968521778358756148971826837398845514398788707884733265341263544748363817548671528296235183185914206710145881079992333254677520496691440858313901330226636914991732069153588327163012679853661047871911921162952965637803396250003906411011347807868274;
            5'd7: xpb[44] = 1024'd37436797309908431486871437261182231342450565124592622967640585441616442972779127497126286560433875362105776063036311753281114259477380361931729637268936703255344270313670854211845384059934844232910935496755805315621613873613781754864722166953716679515615882759202337435091068079319413998851249571030577684876;
            5'd8: xpb[44] = 1024'd7337283873002567013910520468546997892886809535038516497837281914711107586802106022425735722022236325422844241339358165298683770590943175191930978302690220596481830481460628431357513442349191774381012679610280404606312755495494356141117170894753505370183893606483511917216498355242577993796088130713347501478;
            5'd9: xpb[44] = 1024'd101304466120221443939748531080726197188021481071220094156165833452782667538134223457740256098268271598183061827099898011895317122545726323007292444352774778871310065218821619988499882016280745037161287470851995339955372487598103730382490744519019780491571807867881744429448456705094375005859616517021711802411;
            5'd10: xpb[44] = 1024'd71204952683315579466787614288090963738457725481665987686362529925877332152157201983039705259856632561500130005402944423912886633659289136267493785386528296212447625386611394208012011398695092578631364653706470428940071369479816331658885748460056606346139818715162918911573886981017539000804455076704481619013;
            5'd11: xpb[44] = 1024'd41105439246409714993826697495455730288893969892111881216559226398971996766180180508339154421444993524817198183705990835930456144772851949527695126420281813553585185554401168427524140781109440120101441836560945517924770251361528932935280752401093432200707829562444093393699317256940702995749293636387251435615;
            5'd12: xpb[44] = 1024'd11005925809503850520865780702820496839330214302557774746755922872066661380203159033638603583033354488134266362009037247948025655886414762787896467454035330894722745722190942647036270163523787661571519019415420606909469133243241534211675756342130258055275840409725267875824747532863866990694132196070021252217;
            5'd13: xpb[44] = 1024'd104973108056722727446703791314999696134464885838739352405084474410138221331535276468953123959279389760894483947769577094544659007841197910603257933504119889169550980459551934204178638737455340924351793810657135542258528865345850908453049329966396533176663754671123500388056705882715664002757660582378385553150;
            5'd14: xpb[44] = 1024'd74873594619816862973742874522364462684901130249185245935281170883232885945558254994252573120867750724211552126072623506562228518954760723863459274537873406510688540627341708423690768119869688465821870993511610631243227747227563509729444333907433359031231765518404674870182136158638827997702499142061155369752;
            5'd15: xpb[44] = 1024'd44774081182910998500781957729729229235337374659631139465477867356327550559581233519552022282456111687528620304375669918579798030068323537123660615571626923851826100795131482643202897502284036007291948176366085720227926629109276111005839337848470184885799776365685849352307566434561991992647337701743925186354;
            5'd16: xpb[44] = 1024'd14674567746005134027821040937093995785773619070077032995674563829422215173604212044851471444044472650845688482678716330597367541181886350383861956605380441192963660962921256862715026884698383548762025359220560809212625510990988712282234341789507010740367787212967023834432996710485155987592176261426695002956;
            5'd17: xpb[44] = 1024'd108641749993224010953659051549273195080908290606258610654003115367493775124936329480165991820290507923605906068439256177194000893136669498199223422655464999467791895700282248419857395458629936811542300150462275744561685243093598086523607915413773285861755701474365256346664955060336952999655704647735059303889;
            5'd18: xpb[44] = 1024'd78542236556318146480698134756637961631344535016704504184199811840588439738959308005465440981878868886922974246742302589211570404250232311459424763689218516808929455868072022639369524841044284353012377333316750833546384124975310687800002919354810111716323712321646430828790385336260116994600543207417829120491;
            5'd19: xpb[44] = 1024'd48442723119412282007737217964002728181780779427150397714396508313683104352982286530764890143467229850240042425045349001229139915363795124719626104722972034150067016035861796858881654223458631894482454516171225922531083006857023289076397923295846937570891723168927605310915815612183280989545381767100598937093;
            5'd20: xpb[44] = 1024'd18343209682506417534776301171367494732217023837596291244593204786777768967005265056064339305055590813557110603348395413246709426477357937979827445756725551491204576203651571078393783605872979435952531699025701011515781888738735890352792927236883763425459734016208779793041245888106444984490220326783368753695;
            5'd21: xpb[44] = 1024'd112310391929725294460614311783546694027351695373777868902921756324849328918337382491378859681301626086317328189108935259843342778432141085795188911806810109766032810941012562635536152179804532698732806490267415946864841620841345264594166500861150038546847648277607012305273204237958241996553748713091733054628;
            5'd22: xpb[44] = 1024'd82210878492819429987653394990911460577787939784223762433118452797943993532360361016678308842889987049634396367411981671860912289545703899055390252840563627107170371108802336855048281562218880240202883673121891035849540502723057865870561504802186864401415659124888186787398634513881405991498587272774502871230;
            5'd23: xpb[44] = 1024'd52111365055913565514692478198276227128224184194669655963315149271038658146383339541977758004478348012951464545715028083878481800659266712315591593874317144448307931276592111074560410944633227781672960855976366124834239384604770467146956508743223690255983669972169361269524064789804569986443425832457272687832;
            5'd24: xpb[44] = 1024'd22011851619007701041731561405640993678660428605115549493511845744133322760406318067277207166066708976268532724018074495896051311772829525575792934908070661789445491444381885294072540327047575323143038038830841213818938266486483068423351512684260516110551680819450535751649495065727733981388264392140042504434;
            5'd25: xpb[44] = 1024'd115979033866226577967569572017820192973795100141297127151840397282204882711738435502591727542312744249028750309778614342492684663727612673391154400958155220064273726181742876851214908900979128585923312830072556149167997998589092442664725086308526791231939595080848768263881453415579530993451792778448406805367;
            5'd26: xpb[44] = 1024'd85879520429320713494608655225184959524231344551743020682037093755299547325761414027891176703901105212345818488081660754510254174841175486651355741991908737405411286349532651070727038283393476127393390012927031238152696880470805043941120090249563617086507605928129942746006883691502694988396631338131176621969;
            5'd27: xpb[44] = 1024'd55780006992414849021647738432549726074667588962188914212233790228394211939784392553190625865489466175662886666384707166527823685954738299911557083025662254746548846517322425290239167665807823668863467195781506327137395762352517645217515094190600442941075616775411117228132313967425858983341469897813946438571;
            5'd28: xpb[44] = 1024'd25680493555508984548686821639914492625103833372634807742430486701488876553807371078490075027077827138979954844687753578545393197068301113171758424059415772087686406685112199509751297048222171210333544378635981416122094644234230246493910098131637268795643627622692291710257744243349022978286308457496716255173;
            5'd29: xpb[44] = 1024'd119647675802727861474524832252093691920238504908816385400759038239560436505139488513804595403323862411740172430448293425142026549023084260987119890109500330362514641422473191066893665622153724473113819169877696351471154376336839620735283671755903543917031541884090524222489702593200819990349836843805080556106;
            5'd30: xpb[44] = 1024'd89548162365821997001563915459458458470674749319262278930955734712655101119162467039104044564912223375057240608751339837159596060136647074247321231143253847703652201590262965286405795004568072014583896352732171440455853258218552222011678675696940369771599552731371698704615132869123983985294675403487850372708;
            5'd31: xpb[44] = 1024'd59448648928916132528602998666823225021110993729708172461152431185749765733185445564403493726500584338374308787054386249177165571250209887507522572177007365044789761758052739505917924386982419556053973535586646529440552140100264823288073679637977195626167563578652873186740563145047147980239513963170620189310;
        endcase
    end

    always_comb begin
        case(flag[15][5:0])
            6'd0: xpb[45] = 1024'd0;
            6'd1: xpb[45] = 1024'd14674567746005134027821040937093995785773619070077032995674563829422215173604212044851471444044472650845688482678716330597367541181886350383861956605380441192963660962921256862715026884698383548762025359220560809212625510990988712282234341789507010740367787212967023834432996710485155987592176261426695002956;
            6'd2: xpb[45] = 1024'd29349135492010268055642081874187991571547238140154065991349127658844430347208424089702942888088945301691376965357432661194735082363772700767723913210760882385927321925842513725430053769396767097524050718441121618425251021981977424564468683579014021480735574425934047668865993420970311975184352522853390005912;
            6'd3: xpb[45] = 1024'd44023703238015402083463122811281987357320857210231098987023691488266645520812636134554414332133417952537065448036148991792102623545659051151585869816141323578890982888763770588145080654095150646286076077661682427637876532972966136846703025368521032221103361638901071503298990131455467962776528784280085008868;
            6'd4: xpb[45] = 1024'd58698270984020536111284163748375983143094476280308131982698255317688860694416848179405885776177890603382753930714865322389470164727545401535447826421521764771854643851685027450860107538793534195048101436882243236850502043963954849128937367158028042961471148851868095337731986841940623950368705045706780011824;
            6'd5: xpb[45] = 1024'd73372838730025670139105204685469978928868095350385164978372819147111075868021060224257357220222363254228442413393581652986837705909431751919309783026902205964818304814606284313575134423491917743810126796102804046063127554954943561411171708947535053701838936064835119172164983552425779937960881307133475014780;
            6'd6: xpb[45] = 1024'd88047406476030804166926245622563974714641714420462197974047382976533291041625272269108828664266835905074130896072297983584205247091318102303171739632282647157781965777527541176290161308190301292572152155323364855275753065945932273693406050737042064442206723277802143006597980262910935925553057568560170017736;
            6'd7: xpb[45] = 1024'd102721974222035938194747286559657970500415333490539230969721946805955506215229484313960300108311308555919819378751014314181572788273204452687033696237663088350745626740448798039005188192888684841334177514543925664488378576936920985975640392526549075182574510490769166841030976973396091913145233829986865020692;
            6'd8: xpb[45] = 1024'd117396541968041072222568327496751966286188952560616263965396510635377721388833696358811771552355781206765507861429730644778940329455090803070895652843043529543709287703370054901720215077587068390096202873764486473701004087927909698257874734316056085922942297703736190675463973683881247900737410091413560023648;
            6'd9: xpb[45] = 1024'd8004414029921464851590441029031529327264144504957612832939219399823041225128769493648171781742579548168046936650953540797244029795756818899597484432092929802982274096720094426805002770768246217548030624597807436549268748698001637575130506422333647396490181502586156479790442320437770871210896526214660542273;
            6'd10: xpb[45] = 1024'd22678981775926598879411481966125525113037763575034645828613783229245256398732981538499643225787052199013735419329669871394611570977643169283459441037473370995945935059641351289520029655466629766310055983818368245761894259688990349857364848211840658136857968715553180314223439030922926858803072787641355545229;
            6'd11: xpb[45] = 1024'd37353549521931732907232522903219520898811382645111678824288347058667471572337193583351114669831524849859423902008386201991979112159529519667321397642853812188909596022562608152235056540165013315072081343038929054974519770679979062139599190001347668877225755928520204148656435741408082846395249049068050548185;
            6'd12: xpb[45] = 1024'd52028117267936866935053563840313516684585001715188711819962910888089686745941405628202586113875997500705112384687102532589346653341415870051183354248234253381873256985483865014950083424863396863834106702259489864187145281670967774421833531790854679617593543141487227983089432451893238833987425310494745551141;
            6'd13: xpb[45] = 1024'd66702685013942000962874604777407512470358620785265744815637474717511901919545617673054057557920470151550800867365818863186714194523302220435045310853614694574836917948405121877665110309561780412596132061480050673399770792661956486704067873580361690357961330354454251817522429162378394821579601571921440554097;
            6'd14: xpb[45] = 1024'd81377252759947134990695645714501508256132239855342777811312038546934117093149829717905529001964942802396489350044535193784081735705188570818907267458995135767800578911326378740380137194260163961358157420700611482612396303652945198986302215369868701098329117567421275651955425872863550809171777833348135557053;
            6'd15: xpb[45] = 1024'd96051820505952269018516686651595504041905858925419810806986602376356332266754041762757000446009415453242177832723251524381449276887074921202769224064375576960764239874247635603095164078958547510120182779921172291825021814643933911268536557159375711838696904780388299486388422583348706796763954094774830560009;
            6'd16: xpb[45] = 1024'd110726388251957403046337727588689499827679477995496843802661166205778547440358253807608471890053888104087866315401967854978816818068961271586631180669756018153727900837168892465810190963656931058882208139141733101037647325634922623550770898948882722579064691993355323320821419293833862784356130356201525562965;
            6'd17: xpb[45] = 1024'd1334260313837795675359841120969062868754669939838192670203874970223867276653326942444872119440686445490405390623190750997120518409627287415333012258805418413000887230518931990894978656838108886334035889975054063885911986405014562868026671055160284052612575792205289125147887930390385754829616791002626081590;
            6'd18: xpb[45] = 1024'd16008828059842929703180882058063058654528289009915225665878438799646082450257538987296343563485159096336093873301907081594488059591513637799194968864185859605964548193440188853610005541536492435096061249195614873098537497396003275150261012844667294792980363005172312959580884640875541742421793052429321084546;
            6'd19: xpb[45] = 1024'd30683395805848063731001922995157054440301908079992258661553002629068297623861751032147815007529631747181782355980623412191855600773399988183056925469566300798928209156361445716325032426234875983858086608416175682311163008386991987432495354634174305533348150218139336794013881351360697730013969313856016087502;
            6'd20: xpb[45] = 1024'd45357963551853197758822963932251050226075527150069291657227566458490512797465963076999286451574104398027470838659339742789223141955286338566918882074946741991891870119282702579040059310933259532620111967636736491523788519377980699714729696423681316273715937431106360628446878061845853717606145575282711090458;
            6'd21: xpb[45] = 1024'd60032531297858331786644004869345046011849146220146324652902130287912727971070175121850757895618577048873159321338056073386590683137172688950780838680327183184855531082203959441755086195631643081382137326857297300736414030368969411996964038213188327014083724644073384462879874772331009705198321836709406093414;
            6'd22: xpb[45] = 1024'd74707099043863465814465045806439041797622765290223357648576694117334943144674387166702229339663049699718847804016772403983958224319059039334642795285707624377819192045125216304470113080330026630144162686077858109949039541359958124279198380002695337754451511857040408297312871482816165692790498098136101096370;
            6'd23: xpb[45] = 1024'd89381666789868599842286086743533037583396384360300390644251257946757158318278599211553700783707522350564536286695488734581325765500945389718504751891088065570782853008046473167185139965028410178906188045298418919161665052350946836561432721792202348494819299070007432131745868193301321680382674359562796099326;
            6'd24: xpb[45] = 1024'd104056234535873733870107127680627033369170003430377423639925821776179373491882811256405172227751995001410224769374205065178693306682831740102366708496468506763746513970967730029900166849726793727668213404518979728374290563341935548843667063581709359235187086282974455966178864903786477667974850620989491102282;
            6'd25: xpb[45] = 1024'd118730802281878867897928168617721029154943622500454456635600385605601588665487023301256643671796467652255913252052921395776060847864718090486228665101848947956710174933888986892615193734425177276430238763739540537586916074332924261125901405371216369975554873495941479800611861614271633655567026882416186105238;
            6'd26: xpb[45] = 1024'd9338674343759260526950282150000592196018814444795805503143094370046908501782096436093043901183265993658452327274144291794364548205384106314930496690898348215983161327239026417699981427606355103882066514572861500435180735103016200443157177477493931449102757294791445604938330250828156626040513317217286623863;
            6'd27: xpb[45] = 1024'd24013242089764394554771323087094587981792433514872838498817658199469123675386308480944515345227738644504140809952860622391732089387270456698792453296278789408946822290160283280415008312304738652644091873793422309647806246094004912725391519267000942189470544507758469439371326961313312613632689578643981626819;
            6'd28: xpb[45] = 1024'd38687809835769528582592364024188583767566052584949871494492222028891338848990520525795986789272211295349829292631576952989099630569156807082654409901659230601910483253081540143130035197003122201406117233013983118860431757084993625007625861056507952929838331720725493273804323671798468601224865840070676629775;
            6'd29: xpb[45] = 1024'd53362377581774662610413404961282579553339671655026904490166785858313554022594732570647458233316683946195517775310293283586467171751043157466516366507039671794874144216002797005845062081701505750168142592234543928073057268075982337289860202846014963670206118933692517108237320382283624588817042101497371632731;
            6'd30: xpb[45] = 1024'd68036945327779796638234445898376575339113290725103937485841349687735769196198944615498929677361156597041206257989009614183834712932929507850378323112420112987837805178924053868560088966399889298930167951455104737285682779066971049572094544635521974410573906146659540942670317092768780576409218362924066635687;
            6'd31: xpb[45] = 1024'd82711513073784930666055486835470571124886909795180970481515913517157984369803156660350401121405629247886894740667725944781202254114815858234240279717800554180801466141845310731275115851098272847692193310675665546498308290057959761854328886425028985150941693359626564777103313803253936564001394624350761638643;
            6'd32: xpb[45] = 1024'd97386080819790064693876527772564566910660528865258003477190477346580199543407368705201872565450101898732583223346442275378569795296702208618102236323180995373765127104766567593990142735796656396454218669896226355710933801048948474136563228214535995891309480572593588611536310513739092551593570885777456641599;
            6'd33: xpb[45] = 1024'd112060648565795198721697568709658562696434147935335036472865041176002414717011580750053344009494574549578271706025158605975937336478588559001964192928561436566728788067687824456705169620495039945216244029116787164923559312039937186418797570004043006631677267785560612445969307224224248539185747147204151644555;
            6'd34: xpb[45] = 1024'd2668520627675591350719682241938125737509339879676385340407749940447734553306653884889744238881372890980810781246381501994241036819254574830666024517610836826001774461037863981789957313676217772668071779950108127771823972810029125736053342110320568105225151584410578250295775860780771509659233582005252163180;
            6'd35: xpb[45] = 1024'd17343088373680725378540723179032121523282958949753418336082313769869949726910865929741215682925845541826499263925097832591608578001140925214527981122991278018965435423959120844504984198374601321430097139170668936984449483801017838018287683899827578845592938797377602084728772571265927497251409843431947166136;
            6'd36: xpb[45] = 1024'd32017656119685859406361764116126117309056578019830451331756877599292164900515077974592687126970318192672187746603814163188976119183027275598389937728371719211929096386880377707220011083072984870192122498391229746197074994792006550300522025689334589585960726010344625919161769281751083484843586104858642169092;
            6'd37: xpb[45] = 1024'd46692223865690993434182805053220113094830197089907484327431441428714380074119290019444158571014790843517876229282530493786343660364913625982251894333752160404892757349801634569935037967771368418954147857611790555409700505782995262582756367478841600326328513223311649753594765992236239472435762366285337172048;
            6'd38: xpb[45] = 1024'd61366791611696127462003845990314108880603816159984517323106005258136595247723502064295630015059263494363564711961246824383711201546799976366113850939132601597856418312722891432650064852469751967716173216832351364622326016773983974864990709268348611066696300436278673588027762702721395460027938627712032175004;
            6'd39: xpb[45] = 1024'd76041359357701261489824886927408104666377435230061550318780569087558810421327714109147101459103736145209253194639963154981078742728686326749975807544513042790820079275644148295365091737168135516478198576052912173834951527764972687147225051057855621807064087649245697422460759413206551447620114889138727177960;
            6'd40: xpb[45] = 1024'd90715927103706395517645927864502100452151054300138583314455132916981025594931926153998572903148208796054941677318679485578446283910572677133837764149893483983783740238565405158080118621866519065240223935273472983047577038755961399429459392847362632547431874862212721256893756123691707435212291150565422180916;
            6'd41: xpb[45] = 1024'd105390494849711529545466968801596096237924673370215616310129696746403240768536138198850044347192681446900630159997395816175813825092459027517699720755273925176747401201486662020795145506564902614002249294494033792260202549746950111711693734636869643287799662075179745091326752834176863422804467411992117183872;
            6'd42: xpb[45] = 1024'd120065062595716663573288009738690092023698292440292649305804260575825455942140350243701515791237154097746318642676112146773181366274345377901561677360654366369711062164407918883510172391263286162764274653714594601472828060737938823993928076426376654028167449288146768925759749544662019410396643673418812186828;
            6'd43: xpb[45] = 1024'd10672934657597056202310123270969655064773484384633998173346969340270775778435423378537916020623952439148857717897335042791485066615011393730263508949703766628984048557757958408594960084444463990216102404547915564321092721508030763311183848532654215501715333086996734730086218181218542380870130108219912705453;
            6'd44: xpb[45] = 1024'd25347502403602190230131164208063650850547103454711031169021533169692990952039635423389387464668425089994546200576051373388852607796897744114125465555084207821947709520679215271309986969142847538978127763768476373533718232499019475593418190322161226242083120299963758564519214891703698368462306369646607708409;
            6'd45: xpb[45] = 1024'd40022070149607324257952205145157646636320722524788064164696096999115206125643847468240858908712897740840234683254767703986220148978784094497987422160464649014911370483600472134025013853841231087740153122989037182746343743490008187875652532111668236982450907512930782398952211602188854356054482631073302711365;
            6'd46: xpb[45] = 1024'd54696637895612458285773246082251642422094341594865097160370660828537421299248059513092330352757370391685923165933484034583587690160670444881849378765845090207875031446521728996740040738539614636502178482209597991958969254480996900157886873901175247722818694725897806233385208312674010343646658892499997714321;
            6'd47: xpb[45] = 1024'd69371205641617592313594287019345638207867960664942130156045224657959636472852271557943801796801843042531611648612200365180955231342556795265711335371225531400838692409442985859455067623237998185264203841430158801171594765471985612440121215690682258463186481938864830067818205023159166331238835153926692717277;
            6'd48: xpb[45] = 1024'd84045773387622726341415327956439633993641579735019163151719788487381851646456483602795273240846315693377300131290916695778322772524443145649573291976605972593802353372364242722170094507936381734026229200650719610384220276462974324722355557480189269203554269151831853902251201733644322318831011415353387720233;
            6'd49: xpb[45] = 1024'd98720341133627860369236368893533629779415198805096196147394352316804066820060695647646744684890788344222988613969633026375690313706329496033435248581986413786766014335285499584885121392634765282788254559871280419596845787453963037004589899269696279943922056364798877736684198444129478306423187676780082723189;
            6'd50: xpb[45] = 1024'd113394908879632994397057409830627625565188817875173229143068916146226281993664907692498216128935260995068677096648349356973057854888215846417297205187366854979729675298206756447600148277333148831550279919091841228809471298444951749286824241059203290684289843577765901571117195154614634294015363938206777726145;
            6'd51: xpb[45] = 1024'd4002780941513387026079523362907188606264009819514578010611624910671601829959980827334616358322059336471216171869572252991361555228881862245999036776416255239002661691556795972684935970514326659002107669925162191657735959215043688604080013165480852157837727376615867375443663791171157264488850373007878244770;
            6'd52: xpb[45] = 1024'd18677348687518521053900564300001184392037628889591611006286188740093817003564192872186087802366531987316904654548288583588729096410768212629860993381796696431966322654478052835399962855212710207764133029145723000870361470206032400886314354954987862898205514589582891209876660501656313252081026634434573247726;
            6'd53: xpb[45] = 1024'd33351916433523655081721605237095180177811247959668644001960752569516032177168404917037559246411004638162593137227004914186096637592654563013722949987177137624929983617399309698114989739911093756526158388366283810082986981197021113168548696744494873638573301802549915044309657212141469239673202895861268250682;
            6'd54: xpb[45] = 1024'd48026484179528789109542646174189175963584867029745676997635316398938247350772616961889030690455477289008281619905721244783464178774540913397584906592557578817893644580320566560830016624609477305288183747586844619295612492188009825450783038534001884378941089015516938878742653922626625227265379157287963253638;
            6'd55: xpb[45] = 1024'd62701051925533923137363687111283171749358486099822709993309880228360462524376829006740502134499949939853970102584437575380831719956427263781446863197938020010857305543241823423545043509307860854050209106807405428508238003178998537733017380323508895119308876228483962713175650633111781214857555418714658256594;
            6'd56: xpb[45] = 1024'd77375619671539057165184728048377167535132105169899742988984444057782677697981041051591973578544422590699658585263153905978199261138313614165308819803318461203820966506163080286260070394006244402812234466027966237720863514169987250015251722113015905859676663441450986547608647343596937202449731680141353259550;
            6'd57: xpb[45] = 1024'd92050187417544191193005768985471163320905724239976775984659007887204892871585253096443445022588895241545347067941870236575566802320199964549170776408698902396784627469084337148975097278704627951574259825248527046933489025160975962297486063902522916600044450654418010382041644054082093190041907941568048262506;
            6'd58: xpb[45] = 1024'd106724755163549325220826809922565159106679343310053808980333571716627108045189465141294916466633367892391035550620586567172934343502086314933032733014079343589748288432005594011690124163403011500336285184469087856146114536151964674579720405692029927340412237867385034216474640764567249177634084202994743265462;
            6'd59: xpb[45] = 1024'd121399322909554459248647850859659154892452962380130841976008135546049323218793677186146387910677840543236724033299302897770301884683972665316894689619459784782711949394926850874405151048101395049098310543689648665358740047142953386861954747481536938080780025080352058050907637475052405165226260464421438268418;
            6'd60: xpb[45] = 1024'd12007194971434851877669964391938717933528154324472190843550844310494643055088750320982788140064638884639263108520525793788605585024638681145596521208509185041984935788276890399489938741282572876550138294522969628207004707913045326179210519587814499554327908879202023855234106111608928135699746899222538787043;
            6'd61: xpb[45] = 1024'd26681762717439985905491005329032713719301773394549223839225408139916858228692962365834259584109111535484951591199242124385973126206525031529458477813889626234948596751198147262204965625980956425312163653743530437419630218904034038461444861377321510294695696092169047689667102822094084123291923160649233789999;
            6'd62: xpb[45] = 1024'd41356330463445119933312046266126709505075392464626256834899971969339073402297174410685731028153584186330640073877958454983340667388411381913320434419270067427912257714119404124919992510679339974074189012964091246632255729895022750743679203166828521035063483305136071524100099532579240110884099422075928792955;
            6'd63: xpb[45] = 1024'd56030898209450253961133087203220705290849011534703289830574535798761288575901386455537202472198056837176328556556674785580708208570297732297182391024650508620875918677040660987635019395377723522836214372184652055844881240886011463025913544956335531775431270518103095358533096243064396098476275683502623795911;
        endcase
    end

    always_comb begin
        case(flag[15][11:6])
            6'd0: xpb[46] = 1024'd0;
            6'd1: xpb[46] = 1024'd70705465955455387988954128140314701076622630604780322826249099628183503749505598500388673916242529488022017039235391116178075749752184082681044347630030949813839579639961917850350046280076107071598239731405212865057506751877000175308147886745842542515799057731070119192966092953549552086068451944929318798867;
            6'd2: xpb[46] = 1024'd17344236226786034579109328875814969408546834083824961524366344191390112161702058090762276617827384666600884671013288797777087658663147830806928570243730858693988484710352618363069853368635008421886281854423185883750652653533103577651317203808455635764778212048023180355825657833170471155018214063233043113403;
            6'd3: xpb[46] = 1024'd88049702182241422568063457016129670485169464688605284350615443819573615911207656591150950534069914154622901710248679913955163408415331913487972917873761808507828064350314536213419899648711115493484521585828398748808159405410103752959465090554298178280577269779093299548791750786720023241086666008162361912270;
            6'd4: xpb[46] = 1024'd34688472453572069158218657751629938817093668167649923048732688382780224323404116181524553235654769333201769342026577595554175317326295661613857140487461717387976969420705236726139706737270016843772563708846371767501305307066207155302634407616911271529556424096046360711651315666340942310036428126466086226806;
            6'd5: xpb[46] = 1024'd105393938409027457147172785891944639893716298772430245874981788010963728072909714681913227151897298821223786381261968711732251067078479744294901488117492667201816549060667154576489753017346123915370803440251584632558812058943207330610782294362753814045355481827116479904617408619890494396104880071395405025673;
            6'd6: xpb[46] = 1024'd52032708680358103737327986627444908225640502251474884573099032574170336485106174272286829853482153999802654013039866393331262975989443492420785710731192576081965454131057855089209560105905025265658845563269557651251957960599310732953951611425366907294334636144069541067476973499511413465054642189699129340209;
            6'd7: xpb[46] = 1024'd122738174635813491726282114767759609302263132856255207399348132202353840234611772772675503769724683487824671052275257509509338725741627575101830058361223525895805033771019772939559606385981132337257085294674770516309464712476310908262099498171209449810133693875139660260443066453060965551123094134628448139076;
            6'd8: xpb[46] = 1024'd69376944907144138316437315503259877634187336335299846097465376765560448646808232363049106471309538666403538684053155191108350634652591323227714280974923434775953938841410473452279413474540033687545127417692743535002610614132414310605268815233822543059112848192092721423302631332681884620072856252932172453612;
            6'd9: xpb[46] = 1024'd16015715178474784906592516238760145966111539814344484795582621328767057059004691953422709172894393844982406315831052872707362543563555071353598503588623343656102843911801173964999220563098935037833169540710716553695756515788517712948438132296435636308092002509045782586162196212302803689022618371235896768148;
            6'd10: xpb[46] = 1024'd86721181133930172895546644379074847042734170419124807621831720956950560808510290453811383089136923333004423355066443988885438293315739154034642851218654293469942423551763091815349266843175042109431409272115929418753263267665517888256586019042278178823891060240115901779128289165852355775091070316165215567015;
            6'd11: xpb[46] = 1024'd33359951405260819485701845114575115374658373898169446319948965520157169220706750044184985790721778511583290986844341670484450202226702902160527073832354202350091328622153792328069073931733943459719451395133902437446409169321621290599755336104891272072870214557068962941987854045473274844040832434468939881551;
            6'd12: xpb[46] = 1024'd104065417360716207474655973254889816451281004502949769146198065148340672970212348544573659706964307999605308026079732786662525951978886984841571421462385152163930908262115710178419120211810050531317691126539115302503915921198621465907903222850733814588669272288139082134953946999022826930109284379398258680418;
            6'd13: xpb[46] = 1024'd50704187632046854064811173990390084783205207981994407844315309711547281382408808134947262408549163178184175657857630468261537860889850732967455644076085061044079813332506410691138927300368951881605733249557088321197061822854724868251072539913346907837648426605092143297813511878643745999059046497701982994954;
            6'd14: xpb[46] = 1024'd121409653587502242053765302130704785859827838586774730670564409339730785131914406635335936324791692666206192697093021584439613610642034815648499991706116010857919392972468328541488973580445058953203972980962301186254568574731725043559220426659189450353447484336162262490779604832193298085127498442631301793821;
            6'd15: xpb[46] = 1024'd68048423858832888643920502866205054191752042065819369368681653902937393544110866225709539026376547844785060328870919266038625519552998563774384214319815919738068298042859029054208780669003960303492015103980274204947714476387828445902389743721802543602426638653115323653639169711814217154077260560935026108357;
            6'd16: xpb[46] = 1024'd14687194130163535234075703601705322523676245544864008066798898466144001956307325816083141727961403023363927960648816947637637428463962311900268436933515828618217203113249729566928587757562861653780057226998247223640860378043931848245559060784415636851405792970068384816498734591435136223027022679238750422893;
            6'd17: xpb[46] = 1024'd85392660085618923223029831742020023600298876149644330893047998094327505705812924316471815644203932511385944999884208063815713178216146394581312784563546778432056782753211647417278634037638968725378296958403460088698367129920932023553706947530258179367204850701138504009464827544984688309095474624168069221760;
            6'd18: xpb[46] = 1024'd32031430356949569813185032477520291932223079628688969591165242657534114118009383906845418345788787689964812631662105745414725087127110142707197007177246687312205687823602347929998441126197870075666339081421433107391513031577035425896876264592871272616184005018091565172324392424605607378045236742471793536296;
            6'd19: xpb[46] = 1024'd102736896312404957802139160617834993008845710233469292417414342285717617867514982407234092262031317177986829670897496861592800836879294225388241354807277637126045267463564265780348487406273977147264578812826645972449019783454035601205024151338713815131983062749161684365290485378155159464113688687401112335163;
            6'd20: xpb[46] = 1024'd49375666583735604392294361353335261340769913712513931115531586848924226279711441997607694963616172356565697302675394543191812745790257973514125577420977546006194172533954966293068294494832878497552620935844618991142165685110139003548193468401326908380962217066114745528150050257776078533063450805704836649699;
            6'd21: xpb[46] = 1024'd120081132539190992381248489493649962417392544317294253941780686477107730029217040497996368879858701844587714341910785659369888495542442056195169925051008495820033752173916884143418340774908985569150860667249831856199672436987139178856341355147169450896761274797184864721116143211325630619131902750634155448566;
            6'd22: xpb[46] = 1024'd66719902810521638971403690229150230749316747796338892639897931040314338441413500088369971581443557023166581973688683340968900404453405804321054147664708404700182657244307584656138147863467886919438902790267804874892818338643242581199510672209782544145740429114137925883975708090946549688081664868937879763102;
            6'd23: xpb[46] = 1024'd13358673081852285561558890964650499081240951275383531338015175603520946853609959678743574283028412201745449605466581022567912313364369552446938370278408313580331562314698285168857954952026788269726944913285777893585964240299345983542679989272395637394719583431090987046835272970567468757031426987241604077638;
            6'd24: xpb[46] = 1024'd84064139037307673550513019104965200157863581880163854164264275231704450603115558179132248199270941689767466644701972138745988063116553635127982717908439263394171141954660203019208001232102895341325184644690990758643470992176346158850827876018238179910518641162161106239801365924117020843099878932170922876505;
            6'd25: xpb[46] = 1024'd30702909308638320140668219840465468489787785359208492862381519794911059015312017769505850900855796868346334276479869820344999972027517383253866940522139172274320047025050903531927808320661796691613226767708963777336616893832449561193997193080851273159497795479114167402660930803737939912049641050474647191041;
            6'd26: xpb[46] = 1024'd101408375264093708129622347980780169566410415963988815688630619423094562764817616269894524817098326356368351315715260936523075721779701465934911288152170122088159626665012821382277854600737903763211466499114176642394123645709449736502145079826693815675296853210184286595627023757287491998118092995403965989908;
            6'd27: xpb[46] = 1024'd48047145535424354719777548716280437898334619443033454386747863986301171177014075860268127518683181534947218947493158618122087630690665214060795510765870030968308531735403521894997661689296805113499508622132149661087269547365553138845314396889306908924276007527137347758486588636908411067067855113707690304444;
            6'd28: xpb[46] = 1024'd118752611490879742708731676856595138974957250047813777212996963614484674926519674360656801434925711022969235986728549734300163380442849296741839858395900980782148111375365439745347707969372912185097748353537362526144776299242553314153462283635149451440075065258207466951452681590457963153136307058637009103311;
            6'd29: xpb[46] = 1024'd65391381762210389298886877592095407306881453526858415911114208177691283338716133951030404136510566201548103618506447415899175289353813044867724081009600889662297016445756140258067515057931813535385790476555335544837922200898656716496631600697762544689054219575160528114312246470078882222086069176940733417847;
            6'd30: xpb[46] = 1024'd12030152033541035889042078327595675638805657005903054609231452740897891750912593541404006838095421380126971250284345097498187198264776792993608303623300798542445921516146840770787322146490714885673832599573308563531068102554760118839800917760375637938033373892113589277171811349699801291035831295244457732383;
            6'd31: xpb[46] = 1024'd82735617988996423877996206467910376715428287610683377435480552369081395500418192041792680754337950868148988289519736213676262948016960875674652651253331748356285501156108758621137368426566821957272072330978521428588574854431760294147948804506218180453832431623183708470137904303249353377104283240173776531250;
            6'd32: xpb[46] = 1024'd29374388260327070468151407203410645047352491089728016133597796932288003912614651632166283455922806046727855921297633895275274856927924623800536873867031657236434406226499459133857175515125723307560114453996494447281720756087863696491118121568831273702811585940136769632997469182870272446054045358477500845786;
            6'd33: xpb[46] = 1024'd100079854215782458457105535343725346123975121694508338959846896560471507662120250132554957372165335534749872960533025011453350606680108706481581221497062607050273985866461376984207221795201830379158354185401707312339227507964863871799266008314673816218610643671206888825963562136419824532122497303406819644653;
            6'd34: xpb[46] = 1024'd46718624487113105047260736079225614455899325173552977657964141123678116074316709722928560073750190713328740592310922693052362515591072454607465444110762515930422890936852077496927028883760731729446396308419680331032373409620967274142435325377286909467589797988159949988823127016040743601072259421710543959189;
            6'd35: xpb[46] = 1024'd117424090442568493036214864219540315532521955778333300484213240751861619823822308223317233989992720201350757631546313809230438265343256537288509791740793465744262470576813995347277075163836838801044636039824893196089880161497967449450583212123129451983388855719230069181789219969590295687140711366639862758056;
            6'd36: xpb[46] = 1024'd64062860713899139626370064955040583864446159257377939182330485315068228236018767813690836691577575379929625263324211490829450174254220285414394014354493374624411375647204695859996882252395740151332678162842866214783026063154070851793752529185742545232368010036183130344648784849211214756090473484943587072592;
            6'd37: xpb[46] = 1024'd10701630985229786216525265690540852196370362736422577880447729878274836648215227404064439393162430558508492895102109172428462083165184033540278236968193283504560280717595396372716689340954641501620720285860839233476171964810174254136921846248355638481347164353136191507508349728832133825040235603247311387128;
            6'd38: xpb[46] = 1024'd81407096940685174205479393830855553272992993341202900706696829506458340397720825904453113309404960046530509934337500288606537832917368116221322584598224233318399860357557314223066735621030748573218960017266052098533678716687174429445069732994198180997146222084206310700474442682381685911108687548176630185995;
            6'd39: xpb[46] = 1024'd28045867212015820795634594566355821604917196820247539404814074069664948809917285494826716010989815225109377566115397970205549741828331864347206807211924142198548765427948014735786542709589649923507002140284025117226824618343277831788239050056811274246125376401159371863334007562002604980058449666480354500531;
            6'd40: xpb[46] = 1024'd98751333167471208784588722706670522681539827425027862231063173697848452559422883995215389927232344713131394605350789086383625491580515947028251154841955092012388345067909932586136588989665756995105241871689237982284331370220278007096386936802653816761924434132229491056300100515552157066126901611409673299398;
            6'd41: xpb[46] = 1024'd45390103438801855374743923442170791013464030904072500929180418261055060971619343585588992628817199891710262237128686767982637400491479695154135377455655000892537250138300633098856396078224658345393283994707211000977477271876381409439556253865266910010903588449182552219159665395173076135076663729713397613934;
            6'd42: xpb[46] = 1024'd116095569394257243363698051582485492090086661508852823755429517889238564721124942085977666545059729379732279276364077884160713150243663777835179725085685950706376829778262550949206442358300765416991523726112423866034984023753381584747704140611109452526702646180252671412125758348722628221145115674642716412801;
            6'd43: xpb[46] = 1024'd62734339665587889953853252317985760422010864987897462453546762452445173133321401676351269246644584558311146908141975565759725059154627525961063947699385859586525734848653251461926249446859666767279565849130396884728129925409484987090873457673722545775681800497205732574985323228343547290094877792946440727337;
            6'd44: xpb[46] = 1024'd9373109936918536544008453053486028753935068466942101151664007015651781545517861266724871948229439736890014539919873247358736968065591274086948170313085768466674639919043951974646056535418568117567607972148369903421275827065588389434042774736335639024660954814158793737844888107964466359044639911250165041873;
            6'd45: xpb[46] = 1024'd80078575892373924532962581193800729830557699071722423977913106643835285295023459767113545864471969224912031579155264363536812717817775356767992517943116718280514219559005869824996102815494675189165847703553582768478782578942588564742190661482178181540460012545228912930810981061514018445113091856179483840740;
            6'd46: xpb[46] = 1024'd26717346163704571123117781929300998162481902550767062676030351207041893707219919357487148566056824403490899210933162045135824626728739104893876740556816627160663124629396570337715909904053576539453889826571555787171928480598691967085359978544791274789439166862181974093670545941134937514062853974483208155276;
            6'd47: xpb[46] = 1024'd97422812119159959112071910069615699239104533155547385502279450835225397456725517857875822482299353891512916250168553161313900376480923187574921088186847576974502704269358488188065956184129683611052129557976768652229435232475692142393507865290633817305238224593252093286636638894684489600131305919412526954143;
            6'd48: xpb[46] = 1024'd44061582390490605702227110805115967571028736634592024200396695398432005868921977448249425183884209070091783881946450842912912285391886935700805310800547485854651609339749188700785763272688584961340171680994741670922581134131795544736677182353246910554217378910205154449496203774305408669081068037716251268679;
            6'd49: xpb[46] = 1024'd114767048345945993691181238945430668647651367239372347026645795026615509618427575948638099100126738558113800921181841959090988035144071018381849658430578435668491188979711106551135809552764692032938411412399954535980087886008795720044825069099089453070016436641275273642462296727854960755149519982645570067546;
            6'd50: xpb[46] = 1024'd61405818617276640281336439680930936979575570718416985724763039589822118030624035539011701801711593736692668552959739640689999944055034766507733881044278344548640094050101807063855616641323593383226453535417927554673233787664899122387994386161702546318995590958228334805321861607475879824099282100949294382082;
            6'd51: xpb[46] = 1024'd8044588888607286871491640416431205311499774197461624422880284153028726442820495129385304503296448915271536184737637322289011852965998514633618103657978253428788999120492507576575423729882494733514495658435900573366379689321002524731163703224315639567974745275181395968181426487096798893049044219253018696618;
            6'd52: xpb[46] = 1024'd78750054844062674860445768556745906388122404802241947249129383781212230192326093629773978419538978403293553223973028438467087602718182597314662451288009203242628578760454425426925470009958601805112735389841113438423886441198002700039311589970158182083773803006251515161147519440646350979117496164182337495485;
            6'd53: xpb[46] = 1024'd25388825115393321450600969292246174720046608281286585947246628344418838604522553220147581121123833581872420855750926120066099511629146345440546673901709112122777483830845125939645277098517503155400777512859086457117032342854106102382480907032771275332752957323204576324007084320267270048067258282486061810021;
            6'd54: xpb[46] = 1024'd96094291070848709439555097432560875796669238886066908773495727972602342354028151720536255037366363069894437894986317236244175261381330428121591021531740061936617063470807043789995323378593610226999017244264299322174539094731106277690628793778613817848552015054274695516973177273816822134135710227415380608888;
            6'd55: xpb[46] = 1024'd42733061342179356029710298168061144128593442365111547471612972535808950766224611310909857738951218248473305526764214917843187170292294176247475244145439970816765968541197744302715130467152511577287059367282272340867684996387209680033798110841226911097531169371227756679832742153437741203085472345719104923424;
            6'd56: xpb[46] = 1024'd113438527297634744018664426308375845205216072969891870297862072163992454515730209811298531655193747736495322565999606034021262920044478258928519591775470920630605548181159662153065176747228618648885299098687485205925191748264209855341945997587069453613330227102297875872798835106987293289153924290648423722291;
            6'd57: xpb[46] = 1024'd60077297568965390608819627043876113537140276448936508995979316727199062927926669401672134356778602915074190197777503715620274828955442007054403814389170829510754453251550362665784983835787519999173341221705458224618337649920313257685115314649682546862309381419250937035658399986608212358103686408952148036827;
            6'd58: xpb[46] = 1024'd6716067840296037198974827779376381869064479927981147694096561290405671340123128992045737058363458093653057829555401397219286737866405755180288037002870738390903358321941063178504790924346421349461383344723431243311483551576416660028284631712295640111288535736203998198517964866229131427053448527255872351363;
            6'd59: xpb[46] = 1024'd77421533795751425187928955919691082945687110532761470520345660918589175089628727492434410974605987581675074868790792513397362487618589837861332384632901688204742937961902981028854837204422528421059623076128644108368990303453416835336432518458138182627087593467274117391484057819778683513121900472185191150230;
            6'd60: xpb[46] = 1024'd24060304067082071778084156655191351277611314011806109218462905481795783501825187082808013676190842760253942500568690194996374396529553585987216607246601597084891843032293681541574644292981429771347665199146617127062136205109520237679601835520751275876066747784227178554343622699399602582071662590488915464766;
            6'd61: xpb[46] = 1024'd94765770022537459767038284795506052354233944616586432044712005109979287251330785583196687592433372248275959539804081311174450146281737668668260954876632546898731422672255599391924690573057536842945904930551829992119642956986520412987749722266593818391865805515297297747309715652949154668140114535418234263633;
            6'd62: xpb[46] = 1024'd41404540293868106357193485531006320686158148095631070742829249673185895663527245173570290294018227426854827171581978992773462055192701416794145177490332455778880327742646299904644497661616438193233947053569803010812788858642623815330919039329206911640844959832250358910169280532570073737089876653721958578169;
            6'd63: xpb[46] = 1024'd112110006249323494346147613671321021762780778700411393569078349301369399413032843673958964210260756914876844210817370108951537804944885499475189525120363405592719907382608217754994543941692545264832186784975015875870295610519623990639066926075049454156644017563320478103135373486119625823158328598651277377036;
        endcase
    end

    always_comb begin
        case(flag[15][16:12])
            5'd0: xpb[47] = 1024'd0;
            5'd1: xpb[47] = 1024'd58748776520654140936302814406821290094704982179456032267195593864576007825229303264332566911845612093455711842595267790550549713855849247601073747734063314472868812452998918267714351030251446615120228907992988894563441512175727392982236243137662547405623171880273539265994938365740544892108090716955001691572;
            5'd2: xpb[47] = 1024'd117497553041308281872605628813642580189409964358912064534391187729152015650458606528665133823691224186911423685190535581101099427711698495202147495468126628945737624905997836535428702060502893230240457815985977789126883024351454785964472486275325094811246343760547078531989876731481089784216181433910003383144;
            5'd3: xpb[47] = 1024'd52179633877837681410109515815649437539416519412632412673454926528751128138378770882982629520879161970923986120328309937072585300726327408248061118185858902484915762789425537465512813899237134124050489115591726837325963686306285405981730159729758192950049612226703559767878287023293001659205582324239410590385;
            5'd4: xpb[47] = 1024'd110928410398491822346412330222470727634121501592088444940650520393327135963608074147315196432724774064379697962923577727623135014582176655849134865919922216957784575242424455733227164929488580739170718023584715731889405198482012798963966402867420740355672784106977099033873225389033546551313673041194412281957;
            5'd5: xpb[47] = 1024'd45610491235021221883916217224477584984128056645808793079714259192926248451528238501632692129912711848392260398061352083594620887596805568895048488637654490496962713125852156663311276768222821632980749323190464780088485860436843418981224076321853838494476052573133580269761635680845458426303073931523819489198;
            5'd6: xpb[47] = 1024'd104359267755675362820219031631298875078833038825264825346909853057502256276757541765965259041758323941847972240656619874145170601452654816496122236371717804969831525578851074931025627798474268248100978231183453674651927372612570811963460319459516385900099224453407119535756574046586003318411164648478821180770;
            5'd7: xpb[47] = 1024'd39041348592204762357722918633305732428839593878985173485973591857101368764677706120282754738946261725860534675794394230116656474467283729542035859089450078509009663462278775861109739637208509141911009530789202722851008034567401431980717992913949484038902492919563600771644984338397915193400565538808228388011;
            5'd8: xpb[47] = 1024'd97790125112858903294025733040127022523544576058441205753169185721677376589907009384615321650791873819316246518389662020667206188323132977143109606823513392981878475915277694128824090667459955757031238438782191617414449546743128824962954236051612031444525664799837140037639922704138460085508656255763230079583;
            5'd9: xpb[47] = 1024'd32472205949388302831529620042133879873551131112161553892232924521276489077827173738932817347979811603328808953527436376638692061337761890189023229541245666521056613798705395058908202506194196650841269738387940665613530208697959444980211909506045129583328933265993621273528332995950371960498057146092637286824;
            5'd10: xpb[47] = 1024'd91220982470042443767832434448955169968256113291617586159428518385852496903056477003265384259825423696784520796122704167189241775193611137790096977275308980993925426251704313326622553536445643265961498646380929560176971720873686837962448152643707676988952105146267160539523271361690916852606147863047638978396;
            5'd11: xpb[47] = 1024'd25903063306571843305336321450962027318262668345337934298492257185451609390976641357582879957013361480797083231260478523160727648208240050836010599993041254533103564135132014256706665375179884159771529945986678608376052382828517457979705826098140775127755373612423641775411681653502828727595548753377046185637;
            5'd12: xpb[47] = 1024'd84651839827225984241639135857783317412967650524793966565687851050027617216205944621915446868858973574252795073855746313711277362064089298437084347727104569005972376588130932524421016405431330774891758853979667502939493895004244850961942069235803322533378545492697181041406620019243373619703639470332047877209;
            5'd13: xpb[47] = 1024'd19333920663755383779143022859790174762974205578514314704751589849626729704126108976232942566046911358265357508993520669682763235078718211482997970444836842545150514471558633454505128244165571668701790153585416551138574556959075470979199742690236420672181813958853662277295030311055285494693040360661455084450;
            5'd14: xpb[47] = 1024'd78082697184409524715445837266611464857679187757970346971947183714202737529355412240565509477892523451721069351588788460233312948934567459084071718178900157018019326924557551722219479274417018283822019061578405445702016069134802863961435985827898968077804985839127201543289968676795830386801131077616456776022;
            5'd15: xpb[47] = 1024'd12764778020938924252949724268618322207685742811690695111010922513801850017275576594883005175080461235733631786726562816204798821949196372129985340896632430557197464807985252652303591113151259177632050361184154493901096731089633483978693659282332066216608254305283682779178378968607742261790531967945863983263;
            5'd16: xpb[47] = 1024'd71513554541593065189252538675439612302390724991146727378206516378377857842504879859215572086926073329189343629321830606755348535805045619731059088630695745030066277260984170920017942143402705792752279269177143388464538243265360876960929902419994613622231426185557222045173317334348287153898622684900865674835;
            5'd17: xpb[47] = 1024'd6195635378122464726756425677446469652397280044867075517270255177976970330425044213533067784114011113201906064459604962726834408819674532776972711348428018569244415144411871850102053982136946686562310568782892436663618905220191496978187575874427711761034694651713703281061727626160199028888023575230272882076;
            5'd18: xpb[47] = 1024'd64944411898776605663059240084267759747102262224323107784465849042552978155654347477865634695959623206657617907054872753277384122675523780378046459082491333042113227597410790117816405012388393301682539476775881331227060417395918889960423819012090259166657866531987242547056665991900743920996114292185274573648;
            5'd19: xpb[47] = 1024'd123693188419430746599362054491089049841807244403779140051661442907128985980883650742198201607805235300113329749650140543827933836531373027979120206816554647514982040050409708385530756042639839916802768384768870225790501929571646282942660062149752806572281038412260781813051604357641288813104205009140276265220;
            5'd20: xpb[47] = 1024'd58375269255960146136865941493095907191813799457499488190725181706728098468803815096515697304993173084125892184787914899799419709546001941025033829534286921054160177933837409315614867881374080810612799684374619273989582591526476902959917735604185904711084306878417263048940014649453200688093605899469683472461;
            5'd21: xpb[47] = 1024'd117124045776614287073168755899917197286518781636955520457920775571304106294033118360848264216838785177581604027383182690349969423401851188626107577268350235527028990386836327583329218911625527425733028592367608168553024103702204295942153978741848452116707478758690802314934953015193745580201696616424685164033;
            5'd22: xpb[47] = 1024'd51806126613143686610672642901924054636525336690675868596984514370903218781953282715165759914026722961594166462520957046321455296416480101672021199986082509066207128270264028513413330750359768319543059891973357216752104765657034915959411652196281550255510747224847283550823363307005657455191097506754092371274;
            5'd23: xpb[47] = 1024'd110554903133797827546975457308745344731230318870131900864180108235479226607182585979498326825872335055049878305116224836872005010272329349273094947720145823539075940723262946781127681780611214934663288799966346111315546277832762308941647895333944097661133919105120822816818301672746202347299188223709094062846;
            5'd24: xpb[47] = 1024'd45236983970327227084479344310752202081236873923852249003243847035078339095102750333815822523060272839062440740253999192843490883286958262319008570437878097078254078606690647711211793619345455828473320099572095159514626939787592928958905568788377195799937187571277304052706711964558114222288589114038501270087;
            5'd25: xpb[47] = 1024'd103985760490981368020782158717573492175941856103308281270439440899654346920332053598148389434905884932518152582849266983394040597142807509920082318171941411551122891059689565978926144649596902443593549007565084054078068451963320321941141811926039743205560359451550843318701650330298659114396679830993502961659;
            5'd26: xpb[47] = 1024'd38667841327510767558286045719580349525948411157028629409503179699253459408252217952465885132093822716530715017987041339365526470157436422965995940889673685090301028943117266909010256488331143337403580307170833102277149113918150941958399485380472841344363627917707324554590060622110570989386080721322910168900;
            5'd27: xpb[47] = 1024'd97416617848164908494588860126401639620653393336484661676698773563829467233481521216798452043939434809986426860582309129916076184013285670567069688623736999563169841396116185176724607518582589952523809215163821996840590626093878334940635728518135388749986799797980863820584998987851115881494171438277911860472;
            5'd28: xpb[47] = 1024'd32098698684694308032092747128408496970659948390205009815762512363428579721401685571115947741127372593998989295720083485887562057027914583612983311341469273102347979279543886106808719357316830846333840514769571045039671288048708954957893401972568486888790068264137345056473409279663027756483572328607319067713;
            5'd29: xpb[47] = 1024'd90847475205348448968395561535229787065364930569661042082958106228004587546630988835448514652972984687454701138315351276438111770883763831214057059075532587575216791732542804374523070387568277461454069422762559939603112800224436347940129645110231034294413240144410884322468347645403572648591663045562320759285;
            5'd30: xpb[47] = 1024'd25529556041877848505899448537236644415371485623381390222021845027603700034551153189766010350160922471467263573453125632409597643898392744259970681793264861114394929615970505304607182226302518355264100722368308987802193462179266967957387318564664132433216508610567365558356757937215484523581063935891727966526;
            5'd31: xpb[47] = 1024'd84278332562531989442202262944057934510076467802837422489217438892179707859780456454098577262006534564922975416048393422960147357754241991861044429527328175587263742068969423572321533256553964970384329630361297882365634974354994360939623561702326679838839680490840904824351696302956029415689154652846729658098;
        endcase
    end

    always_comb begin
        case(flag[16][5:0])
            6'd0: xpb[48] = 1024'd0;
            6'd1: xpb[48] = 1024'd71513554541593065189252538675439612302390724991146727378206516378377857842504879859215572086926073329189343629321830606755348535805045619731059088630695745030066277260984170920017942143402705792752279269177143388464538243265360876960929902419994613622231426185557222045173317334348287153898622684900865674835;
            6'd2: xpb[48] = 1024'd18960413399061388979706149946064791860083022856557770628281177691778820347700620808416072959194472348935537851186167778931633230768870904906958052245060449126441879952397124502405645095288205864194360929967046930564715636309824980956881235156759777977642948956997386060240106594767941290678555543176136865339;
            6'd3: xpb[48] = 1024'd90473967940654454168958688621504404162473747847704498006487694070156678190205500667631645046120545678124881480507998385686981766573916524638017140875756194156508157213381295422423587238690911656946640199144190319029253879575185857917811137576754391599874375142554608105413423929116228444577178228077002540174;
            6'd4: xpb[48] = 1024'd37920826798122777959412299892129583720166045713115541256562355383557640695401241616832145918388944697871075702372335557863266461537741809813916104490120898252883759904794249004811290190576411728388721859934093861129431272619649961913762470313519555955285897913994772120480213189535882581357111086352273730678;
            6'd5: xpb[48] = 1024'd109434381339715843148664838567569196022556770704262268634768871761935498537906121476047718005315018027060419331694166164618614997342787429544975193120816643282950037165778419924829232333979117521141001129111237249593969515885010838874692372733514169577517324099551994165653530523884169735255733771253139405513;
            6'd6: xpb[48] = 1024'd56881240197184166939118449838194375580249068569673311884843533075336461043101862425248218877583417046806613553558503336794899692306612714720874156735181347379325639857191373507216935285864617592583082789901140791694146908929474942870643705470279333932928846870992158180720319784303823872035666629528410596017;
            6'd7: xpb[48] = 1024'd4328099054652490729572061108819555137941366435084355134918194388737423548297603374448719749851816066552807775422840508971184387270437999896773120349546051475701242548604327089604638237750117664025164450691044333794324301973939046866595038207044498288340369642432322195787109044723478008815599487803681786521;
            6'd8: xpb[48] = 1024'd75841653596245555918824599784259167440332091426231082513124710767115281390802483233664291836777889395742151404744671115726532923075483619627832208980241796505767519809588498009622580381152823456777443719868187722258862545239299923827524940627039111910571795827989544240960426379071765162714222172704547461356;
            6'd9: xpb[48] = 1024'd23288512453713879709278211054884346998024389291642125763199372080516243895998224182864792709046288415488345626609008287902817618039308904803731172594606500602143122501001451592010283333038323528219525380658091264359039938283764027823476273363804276265983318599429708256027215639491419299494155030979818651860;
            6'd10: xpb[48] = 1024'd94802066995306944898530749730323959300415114282788853141405888458894101738503104042080364795972361744677689255930838894658166153844354524534790261225302245632209399761985622512028225476441029320971804649835234652823578181549124904784406175783798889888214744784986930301200532973839706453392777715880684326695;
            6'd11: xpb[48] = 1024'd42248925852775268688984361000949138858107412148199896391480549772295064243698844991280865668240760764423883477795176066834450848808179809710689224839666949728585002453398576094415928428326529392413886310625138194923755574593589008780357508520564054243626267556427094316267322234259360590172710574155955517199;
            6'd12: xpb[48] = 1024'd113762480394368333878236899676388751160498137139346623769687066150672922086203724850496437755166834093613227107117006673589799384613225429441748313470362694758651279714382747014433870571729235185166165579802281583388293817858949885741287410940558667865857693741984316361440639568607647744071333259056821192034;
            6'd13: xpb[48] = 1024'd61209339251836657668690510947013930718190435004757667019761727464073884591399465799696938627435233113359421328981343845766084079577050714617647277084727398855026882405795700596821573523614735256608247240592185125488471210903413989737238743677323832221269216513424480376507428829027301880851266117332092382538;
            6'd14: xpb[48] = 1024'd8656198109304981459144122217639110275882732870168710269836388777474847096595206748897439499703632133105615550845681017942368774540875999793546240699092102951402485097208654179209276475500235328050328901382088667588648603947878093733190076414088996576680739284864644391574218089446956017631198975607363573042;
            6'd15: xpb[48] = 1024'd80169752650898046648396660893078722578273457861315437648042905155852704939100086608113011586629705462294959180167511624697717310345921619524605329329787847981468762358192825099227218618902941120802608170559232056053186847213238970694119978834083610198912165470421866436747535423795243171529821660508229247877;
            6'd16: xpb[48] = 1024'd27616611508366370438850272163703902135965755726726480898117566469253667444295827557313512458898104482041153402031848796874002005309746904700504292944152552077844365049605778681614921570788441192244689831349135598153364240257703074690071311570848774554323688241862030451814324684214897308309754518783500438381;
            6'd17: xpb[48] = 1024'd99130166049959435628102810839143514438356480717873208276324082847631525286800707416529084545824177811230497031353679403629350541114792524431563381574848297107910642310589949601632863714191146984996969100526278986617902483523063951651001213990843388176555114427419252496987642018563184462208377203684366113216;
            6'd18: xpb[48] = 1024'd46577024907427759418556422109768693996048778583284251526398744161032487791996448365729585418092576830976691253218016575805635236078617809607462345189213001204286245002002903184020566666076647056439050761316182528718079876567528055646952546727608552531966637198859416512054431278982838598988310061959637303720;
            6'd19: xpb[48] = 1024'd118090579449020824607808960785208306298439503574430978904605260539410345634501328224945157505018650160166034882539847182560983771883663429338521433819908746234352522262987074104038508809479352849191330030493325917182618119832888932607882449147603166154198063384416638557227748613331125752886932746860502978555;
            6'd20: xpb[48] = 1024'd65537438306489148398262572055833485856131801439842022154679921852811308139697069174145658377287049179912229104404184354737268466847488714514420397434273450330728124954400027686426211761364852920633411691283229459282795512877353036603833781884368330509609586155856802572294537873750779889666865605135774169059;
            6'd21: xpb[48] = 1024'd12984297163957472188716183326458665413824099305253065404754583166212270644892810123346159249555448199658423326268521526913553161811313999690319361048638154427103727645812981268813914713250352992075493352073133001382972905921817140599785114621133494865021108927296966587361327134170434026446798463411045359563;
            6'd22: xpb[48] = 1024'd84497851705550537377968722001898277716214824296399792782961099544590128487397689982561731336481521528847766955590352133668901697616359619421378449679333899457170004906797152188831856856653058784827772621250276389847511149187178017560715017041128108487252535112854188632534644468518721180345421148311911034398;
            6'd23: xpb[48] = 1024'd31944710563018861168422333272523457273907122161810836033035760857991090992593430931762232208749920548593961177454689305845186392580184904597277413293698603553545607598210105771219559808538558856269854282040179931947688542231642121556666349777893272842664057884294352647601433728938375317125354006587182224902;
            6'd24: xpb[48] = 1024'd103458265104611926357674871947963069576297847152957563411242277236368948835098310790977804295675993877783304806776519912600534928385230524328336501924394348583611884859194276691237501951941264649022133551217323320412226785497002998517596252197887886464895484069851574692774751063286662471023976691488047899737;
            6'd25: xpb[48] = 1024'd50905123962080250148128483218588249133990145018368606661316938549769911340294051740178305167944392897529499028640857084776819623349055809504235465538759052679987487550607230273625204903826764720464215212007226862512404178541467102513547584934653050820307006841291738707841540323706316607803909549763319090241;
            6'd26: xpb[48] = 1024'd122418678503673315337381021894027861436380870009515334039523454928147769182798931599393877254870466226718842657962687691532168159154101429235294554169454797710053764811591401193643147047229470513216494481184370250976942421806827979474477487354647664442538433026848960753014857658054603761702532234664184765076;
            6'd27: xpb[48] = 1024'd69865537361141639127834633164653040994073167874926377289598116241548731687994672548594378127138865246465036879827024863708452854117926714411193517783819501806429367503004354776030849999114970584658576141974273793077119814851292083470428820091412828797949955798289124768081646918474257898482465092939455955580;
            6'd28: xpb[48] = 1024'd17312396218609962918288244435278220551765465740337420539672777554949694193190413497794878999407264266211231101691362035884737549081751999587092481398184205902804970194417308358418552951000470656100657802764177335177297207895756187466380152828177993153361478569729288783148436178893912035262397951214727146084;
            6'd29: xpb[48] = 1024'd88825950760203028107540783110717832854156190731484147917879293933327552035695293357010451086333337595400574731013192642640086084886797619318151570028879950932871247455401479278436495094403176448852937071941320723641835451161117064427310055248172606775592904755286510828321753513242199189161020636115592820919;
            6'd30: xpb[48] = 1024'd36272809617671351897994394381343012411848488596895191167953955246728514540891034306210951958601736615146768952877529814816370779850622904494050533643244655029246850146814432860824198046288676520295018732731224265742012844205581168423261387984937771131004427526726674843388542773661853325940953494390864011423;
            6'd31: xpb[48] = 1024'd107786364159264417087246933056782624714239213588041918546160471625106372383395914165426524045527809944336112582199360421571719315655668524225109622273940400059313127407798603780842140189691382313047298001908367654206551087470942045384191290404932384753235853712283896888561860108010140479839576179291729686258;
            6'd32: xpb[48] = 1024'd55233223016732740877700544327407804271931511453452961796235132938507334888591655114627024917796208964082306804063697593748004010619493809401008585888305104155688730099211557363229843141576882384489379662698271196306728480515406149380142623141697549108647376483724060903628649368429794616619509037567000876762;
            6'd33: xpb[48] = 1024'd2680081874201064668154155598032983829623809318864005046309794251908297393787396063827525790064607983828501025928034765924288705583319094576907549502669808252064332790624510945617546093462382455931461323488174738406905873559870253376093955878462713464058899255164224918695438628849448753399441895842272067266;
            6'd34: xpb[48] = 1024'd74193636415794129857406694273472596132014534310010732424516310630286155236292275923043097876990681313017844655249865372679637241388364714307966638133365553282130610051608681865635488236865088248683740592665318126871444116825231130337023858298457327086290325440721446963868755963197735907298064580743137742101;
            6'd35: xpb[48] = 1024'd21640495273262453647860305544097775689706832175421775674590971943687117741488016872243598749259080332764038877114202544855921936352189999483865601747730257378506212743021635448023191188750588320125822253455221668971621509869695234332975191035222491441701848212161610978935545223617390044077997439018408932605;
            6'd36: xpb[48] = 1024'd93154049814855518837112844219537387992097557166568503052797488322064975583992896731459170836185153661953382506436033151611270472157235619214924690378426002408572490004005806368041133332153294112878101522632365057436159753135056111293905093455217105063933274397718833024108862557965677197976620123919274607440;
            6'd37: xpb[48] = 1024'd40600908672323842627566455490162567549789855031979546302872149635465938089188637680659671708453552681699576728300370323787555167121060904390823653992790706504948092695418759950428836284038794184320183183422268599536337146179520215289856426191982269419344797169158997039175651818385331334756552982194545797944;
            6'd38: xpb[48] = 1024'd112114463213916907816818994165602179852180580023126273681078666013843795931693517539875243795379626010888920357622200930542903702926106524121882742623486451535014369956402930870446778427441499977072462452599411988000875389444881092250786328611976883041576223354716219084348969152733618488655175667095411472779;
            6'd39: xpb[48] = 1024'd59561322071385231607272605436227359409872877888537316931153327327244758436889258489075744667648025030635114579486538102719188397889931809297781706237851155631389972647815884452834481379327000048514544113389315530101052782489345196246737661348742047396987746126156383099415758413153272625435108525370682663283;
            6'd40: xpb[48] = 1024'd7008180928853555397726216706852538967565175753948360181227988640645720942084999438276245539916424050381308801350875274895473092853757094473680669852215859727765575339228838035222184331212500119956625774179219072201230175533809300242688994085507211752399268897596547114482547673572926762215041383645953853787;
            6'd41: xpb[48] = 1024'd78521735470446620586978755382292151269955900745095087559434505019023578784589879297491817626842497379570652430672705881650821628658802714204739758482911604757831852600213008955240126474615205912708905043356362460665768418799170177203618896505501825374630695083153769159655865007921213916113664068546819528622;
            6'd42: xpb[48] = 1024'd25968594327914944377432366652917330827648198610506130809509166332424541289785620246692318499110896399316846652537043053827106323622627999380638722097276308854207455291625962537627829426500705984150986704146266002765945811843634281199570229242266989730042217854593933174722654268340868052893596926822090719126;
            6'd43: xpb[48] = 1024'd97482148869508009566684905328356943130038923601652858187715682710802399132290500105907890586036969728506190281858873660582454859427673619111697810727972053884273732552610133457645771569903411776903265973323409391230484055108995158160500131662261603352273644040151155219895971602689155206792219611722956393961;
            6'd44: xpb[48] = 1024'd44929007726976333357138516598982122687731221467063901437790344024203361637486241055108391458305368748252384503723210832758739554391498904287596774342336757980649335244023087040033474521788911848345347634113312933330661448153459262156451464399026767707685166811591319234962760863108809343572152469998227584465;
            6'd45: xpb[48] = 1024'd116442562268569398546391055274421734990121946458210628815996860402581219479991120914323963545231442077441728133045041439514088090196544524018655862973032503010715612505007257960051416665191617641097626903290456321795199691418820139117381366819021381329916592997148541280136078197457096497470775154899093259300;
            6'd46: xpb[48] = 1024'd63889421126037722336844666545046914547814244323621672066071521715982181985186861863524464417499841097187922354909378611690372785160369809194554826587397207107091215196420211542439119617077117712539708564080359863895377084463284243113332699555786545685328115768588705295202867457876750634250708013174364449804;
            6'd47: xpb[48] = 1024'd11336279983506046127298277815672094105506542189032715316146183029383144490382602812724965289768240116934116576773715783866657480124195094370453790201761911203466817887833165124826822568962617783981790224870263405995554477507748347109284032292551710040739638540028869310269656718296404771030640871449635640308;
            6'd48: xpb[48] = 1024'd82849834525099111316550816491111706407897267180179442694352699407761002332887482671940537376694313446123460206095546390622006015929240714101512878832457656233533095148817336044844764712365323576734069494047406794460092720773109224070213934712546323662971064725586091355442974052644691924929263556350501315143;
            6'd49: xpb[48] = 1024'd30296693382567435107004427761736885965589565045590485944427360721161964838083223621141038248962712465869654427959883562798290710893065999277411842446822360329908697840230289627232467664250823648176151154837310336560270113817573328066165267449311488018382587497026255370509763313064346061709196414625772505647;
            6'd50: xpb[48] = 1024'd101810247924160500296256966437176498267980290036737213322633877099539822680588103480356610335888785795058998057281714169553639246698111619008470931077518105359974975101214460547250409807653529440928430424014453725024808357082934205027095169869306101640614013682583477415683080647412633215607819099526638180482;
            6'd51: xpb[48] = 1024'd49257106781628824086710577707801677825672587902148256572708538412940785185783844429557111208157184814805192279146051341729923941661936904184369894691882809456350577792627414129638112759539029512370512084804357267124985750127398309023046502606071265996025536454023641430749869907832287352387751957801909370986;
            6'd52: xpb[48] = 1024'd120770661323221889275963116383241290128063312893294983950915054791318643028288724288772683295083258143994535908467881948485272477466982523915428983322578554486416855053611585049656054902941735305122791353981500655589523993392759185983976405026065879618256962639580863475923187242180574506286374642702775045821;
            6'd53: xpb[48] = 1024'd68217520180690213066416727653866469685755610758706027200989716104719605533484465237973184167351657163740730130332219120661557172430807809091327946936943258582792457745024538632043757854827235376564873014771404197689701386437223289979927737762831043973668485411021027490989976502600228643066307500978046236325;
            6'd54: xpb[48] = 1024'd15664379038158536856870338924491649243447908624117070451064377418120568038680206187173685039620056183486924352196556292837841867394633094267226910551307962679168060436437492214431460806712735448006954675561307739789878779481687393975879070499596208329080008182461191506056765763019882779846240359253317426829;
            6'd55: xpb[48] = 1024'd87177933579751602046122877599931261545838633615263797829270893796498425881185086046389257126546129512676267981518386899593190403199678713998285999182003707709234337697421663134449402950115441240759233944738451128254417022747048270936808972919590821951311434368018413551230083097368169933744863044154183101664;
            6'd56: xpb[48] = 1024'd34624792437219925836576488870556441103530931480674841079345555109899388386380826995589757998814528532422462203382724071769475098163503999174184962796368411805609940388834616716837105902000941312201315605528354670354594415791512374932760305656355986306722957139458577566296872357787824070524795902429454292168;
            6'd57: xpb[48] = 1024'd106138346978812991025829027545996053405921656471821568457552071488277246228885706854805330085740601861611805832704554678524823633968549618905244051427064156835676217649818787636855048045403647104953594874705498058819132659056873251893690208076350599928954383325015799611470189692136111224423418587330319967003;
            6'd58: xpb[48] = 1024'd53585205836281314816282638816621232963613954337232611707626732801678208734081447804005830958009000881358000054568891850701108328932374904081143015041428860932051820341231741219242750997289147176395676535495401600919310052101337355889641540813115764284365906096455963626536978952555765361203351445605591157507;
            6'd59: xpb[48] = 1024'd1032064693749638606736250087246412521306252202643654957701394115079171239277188753206331830277399901104194276433229022877393023896200189257041978655793565028427423032644694801630453949174647247837758196285305143019487445145801459885592873549880928639777428867896127641603768212975419497983284303880862348011;
            6'd60: xpb[48] = 1024'd72545619235342703795988788762686024823696977193790382335907910493457029081782068612421903917203473230293537905755059629632741559701245808988101067286489310058493700293628865721648396092577353040590037465462448531484025688411162336846522775969875542262008855053453349686777085547323706651881906988781728022846;
            6'd61: xpb[48] = 1024'd19992478092811027586442400033311204381389275059201425585982571806857991586977809561622404789471872250039732127619396801809026254665071094164000030900854014154869302985041819304036099044462853112032119126252352073584203081455626440842474108706640706617420377824893513701843874807743360788661839847056999213350;
            6'd62: xpb[48] = 1024'd91506032634404092775694938708750816683780000050348152964189088185235849429482689420837976876397945579229075756941227408564374790470116713895059119531549759184935580246025990224054041187865558904784398395429495462048741324720987317803404011126635320239651804010450735747017192142091647942560462531957864888185;
            6'd63: xpb[48] = 1024'd38952891491872416566148549979375996241472297915759196214263749498636811934678430370038477748666344598975269978805564580740659485433941999070958083145914463281311182937438943806441744139751058976226480056219399004148918717765451421799355343863400484595063326781890899762083981402511302079340395390233136078689;
        endcase
    end

    always_comb begin
        case(flag[16][11:6])
            6'd0: xpb[49] = 1024'd0;
            6'd1: xpb[49] = 1024'd110466446033465481755401088654815608543863022906905923592470265877014669777183310229254049835592417928164613608127395187496008021238987618802017171776610208311377460198423114726459686283153764768978759325396542392613456961030812298760285246283395098217294752967448121807257298736859589233239018075134001753524;
            6'd2: xpb[49] = 1024'd96866196382806222112003249904816784343027618688076163056808676689052444217057481548493028456527161546886077808797296940412952201636754903048874218536889375689064245827275012115289133374790323816647321042405844938862553071840727824555591922883560747167769602520779185584408069399790545449359346323642409022717;
            6'd3: xpb[49] = 1024'd83265946732146962468605411154817960142192214469246402521147087501090218656931652867732007077461905165607542009467198693329896382034522187295731265297168543066751031456126909504118580466426882864315882759415147485111649182650643350350898599483726396118244452074110249361558840062721501665479674572150816291910;
            6'd4: xpb[49] = 1024'd69665697081487702825207572404819135941356810250416641985485498313127993096805824186970985698396648784329006210137100446246840562432289471542588312057447710444437817084978806892948027558063441911984444476424450031360745293460558876146205276083892045068719301627441313138709610725652457881600002820659223561103;
            6'd5: xpb[49] = 1024'd56065447430828443181809733654820311740521406031586881449823909125165767536679995506209964319331392403050470410807002199163784742830056755789445358817726877822124602713830704281777474649700000959653006193433752577609841404270474401941511952684057694019194151180772376915860381388583414097720331069167630830296;
            6'd6: xpb[49] = 1024'd42465197780169183538411894904821487539686001812757120914162319937203541976554166825448942940266136021771934611476903952080728923227824040036302405578006045199811388342682601670606921741336560007321567910443055123858937515080389927736818629284223342969669000734103440693011152051514370313840659317676038099489;
            6'd7: xpb[49] = 1024'd28864948129509923895014056154822663338850597593927360378500730749241316416428338144687921561200879640493398812146805704997673103625591324283159452338285212577498173971534499059436368832973119054990129627452357670108033625890305453532125305884388991920143850287434504470161922714445326529960987566184445368682;
            6'd8: xpb[49] = 1024'd15264698478850664251616217404823839138015193375097599842839141561279090856302509463926900182135623259214863012816707457914617284023358608530016499098564379955184959600386396448265815924609678102658691344461660216357129736700220979327431982484554640870618699840765568247312693377376282746081315814692852637875;
            6'd9: xpb[49] = 1024'd1664448828191404608218378654825014937179789156267839307177552373316865296176680783165878803070366877936327213486609210831561464421125892776873545858843547332871745229238293837095263016246237150327253061470962762606225847510136505122738659084720289821093549394096632024463464040307238962201644063201259907068;
            6'd10: xpb[49] = 1024'd112130894861656886363619467309640623481042812063173762899647818250331535073359991012419928638662784806100940821614004398327569485660113511578890717635453755644249205427661408563554949299400001919306012386867505155219682808540948803883023905368115388038388302361544753831720762777166828195440662138335261660592;
            6'd11: xpb[49] = 1024'd98530645210997626720221628559641799280207407844344002363986229062369309513234162331658907259597528424822405022283906151244513666057880795825747764395732923021935991056513305952384396391036560966974574103876807701468778919350864329678330581968281036988863151914875817608871533440097784411560990386843668929785;
            6'd12: xpb[49] = 1024'd84930395560338367076823789809642975079372003625514241828324639874407083953108333650897885880532272043543869222953807904161457846455648080072604811156012090399622776685365203341213843482673120014643135820886110247717875030160779855473637258568446685939338001468206881386022304103028740627681318635352076198978;
            6'd13: xpb[49] = 1024'd71330145909679107433425951059644150878536599406684481292663050686444858392982504970136864501467015662265333423623709657078402026853415364319461857916291257777309562314217100730043290574309679062311697537895412793966971140970695381268943935168612334889812851021537945163173074765959696843801646883860483468171;
            6'd14: xpb[49] = 1024'd57729896259019847790028112309645326677701195187854720757001461498482632832856676289375843122401759280986797624293611409995346207251182648566318904676570425154996347943068998118872737665946238109980259254904715340216067251780610907064250611768777983840287700574869008940323845428890653059921975132368890737364;
            6'd15: xpb[49] = 1024'd44129646608360588146630273559646502476865790969024960221339872310520407272730847608614821743336502899708261824963513162912290387648949932813175951436849592532683133571920895507702184757582797157648820971914017886465163362590526432859557288368943632790762550128200072717474616091821609276042303380877298006557;
            6'd16: xpb[49] = 1024'd30529396957701328503232434809647678276030386750195199685678283122558181712605018927853800364271246518429726025633414915829234568046717217060032998197128759910369919200772792896531631849219356205317382688923320432714259473400441958654863964969109281741237399681531136494625386754752565492162631629385705275750;
            6'd17: xpb[49] = 1024'd16929147307042068859834596059648854075194982531365439150016693934595956152479190247092778985205990137151190226303316668746178748444484501306890044957407927288056704829624690285361078940855915252985944405932622978963355584210357484450170641569274930691712249234862200271776157417683521708282959877894112544943;
            6'd18: xpb[49] = 1024'd3328897656382809216436757309650029874359578312535678614355104746633730592353361566331757606140733755872654426973218421663122928842251785553747091717687094665743490458476587674190526032492474300654506122941925525212451695020273010245477318169440579642187098788193264048926928080614477924403288126402519814136;
            6'd19: xpb[49] = 1024'd113795343689848290971837845964465638418222601219441602206825370623648400369536671795585807441733151684037268035100613609159130950081239404355764263494297302977120950656899702400650212315646239069633265448338467917825908656051085309005762564452835677859481851755641385856184226817474067157642306201536521567660;
            6'd20: xpb[49] = 1024'd100195094039189031328440007214466814217387197000611841671163781435686174809410843114824786062667895302758732235770515362076075130479006688602621310254576470354807736285751599789479659407282798117301827165347770464075004766861000834801069241053001326809956701308972449633334997480405023373762634450044928836853;
            6'd21: xpb[49] = 1024'd86594844388529771685042168464467990016551792781782081135502192247723949249285014434063764683602638921480196436440417114993019310876773972849478357014855637732494521914603497178309106498919357164970388882357073010324100877670916360596375917653166975760431550862303513410485768143335979589882962698553336106046;
            6'd22: xpb[49] = 1024'd72994594737870512041644329714469165815716388562952320599840603059761723689159185753302743304537382540201660637110318867909963491274541257096335403775134805110181307543455394567138553590555916212638950599366375556573196988480831886391682594253332624710906400415634577187636538806266935806003290947061743375239;
            6'd23: xpb[49] = 1024'd59394345087211252398246490964470341614880984344122560064179013871799498129033357072541721925472126158923124837780220620826907671672308541343192450535413972487868093172307291955968000682192475260307512316375678102822293099290747412186989270853498273661381249968965640964787309469197892022123619195570150644432;
            6'd24: xpb[49] = 1024'd45794095436551992754848652214471517414045580125292799528517424683837272568907528391780700546406869777644589038450122373743851852070075825590049497295693139865554878801159189344797447773829034307976074033384980649071389210100662937982295947453663922611856099522296704741938080132128848238243947444078557913625;
            6'd25: xpb[49] = 1024'd32193845785892733111450813464472693213210175906463038992855835495875047008781699711019679167341613396366053239120024126660796032467843109836906544055972307243241664430011086733626894865465593355644635750394283195320485320910578463777602624053829571562330949075627768519088850795059804454364275692586965182818;
            6'd26: xpb[49] = 1024'd18593596135233473468052974714473869012374771687633278457194246307912821448655871030258657788276357015087517439789925879577740212865610394083763590816251474620928450058862984122456341957102152403313197467403585741569581431720493989572909300653995220512805798628958832296239621457990760670484603941095372452011;
            6'd27: xpb[49] = 1024'd4993346484574213824655135964475044811539367468803517921532657119950595888530042349497636409211100633808981640459827632494684393263377678330620637576530641998615235687714881511285789048738711450981759184412888287818677542530409515368215977254160869463280648182289896073390392120921716886604932189603779721204;
            6'd28: xpb[49] = 1024'd115459792518039695580056224619290653355402390375709441514002922996965265665713352578751686244803518561973595248587222819990692414502365297132637809353140850309992695886137996237745475331892476219960518509809430680432134503561221814128501223537555967680575401149738017880647690857781306119843950264737781474728;
            6'd29: xpb[49] = 1024'd101859542867380435936658385869291829154566986156879680978341333809003040105587523897990664865738262180695059449257124572907636594900132581379494856113420017687679481514989893626574922423529035267629080226818733226681230614371137339923807900137721616631050250703069081657798461520712262335964278513246188743921;
            6'd30: xpb[49] = 1024'd88259293216721176293260547119293004953731581938049920442679744621040814545461695217229643486673005799416523649927026325824580775297899865626351902873699185065366267143841791015404369515165594315297641943828035772930326725181052865719114576737887265581525100256400145434949232183643218552084606761754596013114;
            6'd31: xpb[49] = 1024'd74659043566061916649862708369294180752896177719220159907018155433078588985335866536468622107607749418137987850596928078741524955695667149873208949633978352443053052772693688404233816606802153362966203660837338319179422835990968391514421253338052914531999949809731209212100002846574174768204935010263003282307;
            6'd32: xpb[49] = 1024'd61058793915402657006464869619295356552060773500390399371356566245116363425210037855707600728542493036859452051266829831658469136093434434120065996394257519820739838401545585793063263698438712410634765377846640865428518946800883917309727929938218563482474799363062272989250773509505130984325263258771410551500;
            6'd33: xpb[49] = 1024'd47458544264743397363067030869296532351225369281560638835694977057154137865084209174946579349477236655580916251936731584575413316491201718366923043154536687198426624030397483181892710790075271458303327094855943411677615057610799443105034606538384212432949648916393336766401544172436087200445591507279817820693;
            6'd34: xpb[49] = 1024'd33858294614084137719669192119297708150389965062730878300033387869191912304958380494185557970411980274302380452606633337492357496888969002613780089914815854576113409659249380570722157881711830505971888811865245957926711168420714968900341283138549861383424498469724400543552314835367043416565919755788225089886;
            6'd35: xpb[49] = 1024'd20258044963424878076271353369298883949554560843901117764371798681229686744832551813424536591346723893023844653276535090409301677286736286860637136675095021953800195288101277959551604973348389553640450528874548504175807279230630494695647959738715510333899348023055464320703085498297999632686248004296632359079;
            6'd36: xpb[49] = 1024'd6657795312765618432873514619300059748719156625071357228710209493267461184706723132663515212281467511745308853946436843326245857684503571107494183435374189331486980916953175348381052064984948601309012245883851050424903390040546020490954636338881159284374197576386528097853856161228955848806576252805039628272;
            6'd37: xpb[49] = 1024'd117124241346231100188274603274115668292582179531977280821180475370282130961890033361917565047873885439909922462073832030822253878923491189909511355211984397642864441115376290074840738348138713370287771571280393443038360351071358319251239882622276257501668950543834649905111154898088545082045594327939041381796;
            6'd38: xpb[49] = 1024'd103523991695571840544876764524116844091746775313147520285518886182319905401764204681156543668808629058631386662743733783739198059321258474156368401972263565020551226744228187463670185439775272417956333288289695989287456461881273845046546559222441906452143800097165713682261925561019501298165922576447448650989;
            6'd39: xpb[49] = 1024'd89923742044912580901478925774118019890911371094317759749857296994357679841638376000395522289743372677352850863413635536656142239719025758403225448732542732398238012373080084852499632531411831465624895005298998535536552572691189370841853235822607555402618649650496777459412696223950457514286250824955855920182;
            6'd40: xpb[49] = 1024'd76323492394253321258081087024119195690075966875487999214195707806395454281512547319634500910678116296074315064083537289573086420116793042650082495492821899775924798001931982241329079623048390513293456722308301081785648683501104896637159912422773204353093499203827841236563466886881413730406579073464263189375;
            6'd41: xpb[49] = 1024'd62723242743594061614683248274120371489240562656658238678534118618433228721386718638873479531612859914795779264753439042490030600514560326896939542253101067153611583630783879630158526714684949560962018439317603628034744794311020422432466589022938853303568348757158905013714237549812369946526907321972670458568;
            6'd42: xpb[49] = 1024'd49122993092934801971285409524121547288405158437828478142872529430471003161260889958112458152547603533517243465423340795406974780912327611143796589013380234531298369259635777018987973806321508608630580156326906174283840905120935948227773265623104502254043198310489968790865008212743326162647235570481077727761;
            6'd43: xpb[49] = 1024'd35522743442275542327887570774122723087569754218998717607210940242508777601135061277351436773482347152238707666093242548323918961310094895390653635773659401908985154888487674407817420897958067656299141873336208720532937015930851474023079942223270151204518047863821032568015778875674282378767563818989484996954;
            6'd44: xpb[49] = 1024'd21922493791616282684489732024123898886734350000168957071549351054546552041009232596590415394417090770960171866763144301240863141707862179637510682533938569286671940517339571796646867989594626703967703590345511266782033126740766999818386618823435800154992897417152096345166549538605238594887892067497892266147;
            6'd45: xpb[49] = 1024'd8322244140957023041091893274125074685898945781339196535887761866584326480883403915829394015351834389681636067433046054157807322105629463884367729294217736664358726146191469185476315081231185751636265307354813813031129237550682525613693295423601449105467746970483160122317320201536194811008220316006299535340;
            6'd46: xpb[49] = 1024'd118788690174422504796492981928940683229761968688245120128358027743598996258066714145083443850944252317846249675560441241653815343344617082686384901070827944975736186344614583911936001364384950520615024632751356205644586198581494824373978541706996547322762499937931281929574618938395784044247238391140301288864;
            6'd47: xpb[49] = 1024'd105188440523763245153095143178941859028926564469415359592696438555636770697940885464322422471878995936567713876230342994570759523742384366933241947831107112353422971973466481300765448456021509568283586349760658751893682309391410350169285218307162196273237349491262345706725389601326740260367566639648708558057;
            6'd48: xpb[49] = 1024'd91588190873103985509697304428943034828091160250585599057034849367674545137815056783561401092813739555289178076900244747487703704140151651180098994591386279731109757602318378689594895547658068615952148066769961298142778420201325875964591894907327845223712199044593409483876160264257696476487894888157115827250;
            6'd49: xpb[49] = 1024'd77987941222444725866299465678944210627255756031755838521373260179712319577689228102800379713748483174010642277570146500404647884537918935426956041351665447108796543231170276078424342639294627663620709783779263844391874531011241401759898571507493494174187048597924473261026930927188652692608223136665523096443;
            6'd50: xpb[49] = 1024'd64387691571785466222901626928945386426420351812926077985711670991750094017563399422039358334683226792732106478240048253321592064935686219673813088111944614486483328860022173467253789730931186711289271500788566390640970641821156927555205248107659143124661898151255537038177701590119608908728551385173930365636;
            6'd51: xpb[49] = 1024'd50787441921126206579503788178946562225584947594096317450050081803787868457437570741278336955617970411453570678909950006238536245333453503920670134872223781864170114488874070856083236822567745758957833217797868936890066752631072453350511924707824792075136747704586600815328472253050565124848879633682337634829;
            6'd52: xpb[49] = 1024'd37187192270466946936105949428947738024749543375266556914388492615825642897311742060517315576552714030175034879579851759155480425731220788167527181632502949241856900117725968244912683914204304806626394934807171483139162863440987979145818601307990441025611597257917664592479242915981521340969207882190744904022;
            6'd53: xpb[49] = 1024'd23586942619807687292708110678948913823914139156436796378726903427863417337185913379756294197487457648896499080249753512072424606128988072414384228392782116619543685746577865633742131005840863854294956651816474029388258974250903504941125277908156089976086446811248728369630013578912477557089536130699152173215;
            6'd54: xpb[49] = 1024'd9986692969148427649310271928950089623078734937607035843065314239901191777060084698995272818422201267617963280919655264989368786526755356661241275153061283997230471375429763022571578097477422901963518368825776575637355085060819030736431954508321738926561296364579792146780784241843433773209864379207559442408;
            6'd55: xpb[49] = 1024'd120453139002613909404711360583765698166941757844512959435535580116915861554243394928249322654014619195782576889047050452485376807765742975463258446929671492308607931573852877749031264380631187670942277694222318968250812046091631329496717200791716837143856049332027913954038082978703023006448882454341561195932;
            6'd56: xpb[49] = 1024'd106852889351954649761313521833766873966106353625683198899873990928953635994117566247488301274949362814504041089716952205402320988163510259710115493689950659686294717202704775137860711472267746718610839411231621514499908156901546855292023877391882486094330898885358977731188853641633979222569210702849968465125;
            6'd57: xpb[49] = 1024'd93252639701295390117915683083768049765270949406853438364212401740991410433991737566727279895884106433225505290386853958319265168561277543956972540450229827063981502831556672526690158563904305766279401128240924060749004267711462381087330553992048135044805748438690041508339624304564935438689538951358375734318;
            6'd58: xpb[49] = 1024'd79652390050636130474517844333769225564435545188023677828550812553029184873865908885966258516818850051946969491056755711236209348959044828203829587210508994441668288460408569915519605655540864813947962845250226606998100378521377906882637230592213783995280597992021105285490394967495891654809867199866783003511;
            6'd59: xpb[49] = 1024'd66052140399976870831120005583770401363600140969193917292889223365066959313740080205205237137753593670668433691726657464153153529356812112450686633970788161819355074089260467304349052747177423861616524562259529153247196489331293432677943907192379432945755447545352169062641165630426847870930195448375190272704;
            6'd60: xpb[49] = 1024'd52451890749317611187722166833771577162764736750364156757227634177104733753614251524444215758688337289389897892396559217070097709754579396697543680731067329197041859718112364693178499838813982909285086279268831699496292600141208958473250583792545081896230297098683232839791936293357804087050523696883597541897;
            6'd61: xpb[49] = 1024'd38851641098658351544324328083772752961929332531534396221566044989142508193488422843683194379623080908111362093066460969987041890152346680944400727491346496574728645346964262082007946930450541956953647996278134245745388710951124484268557260392710730846705146652014296616942706956288760303170851945392004811090;
            6'd62: xpb[49] = 1024'd25251391447999091900926489333773928761093928312704635685904455801180282633362594162922173000557824526832826293736362722903986070550113965191257774251625663952415430975816159470837394022087101004622209713287436791994484821761040010063863936992876379797179996205345360394093477619219716519291180193900412080283;
            6'd63: xpb[49] = 1024'd11651141797339832257528650583775104560258524093874875150242866613218057073236765482161151621492568145554290494406264475820930250947881249438114821011904831330102216604668056859666841113723660052290771430296739338243580932570955535859170613593042028747654845758676424171244248282150672735411508442408819349476;
        endcase
    end

    always_comb begin
        case(flag[16][16:12])
            5'd0: xpb[50] = 1024'd0;
            5'd1: xpb[50] = 1024'd122117587830805314012929739238590713104121547000780798742713132490232726850420075711415201457084986073718904102533659663316938272186868868240131992788515039641479676803091171586126527396877424821269530755693281730857037893601767834619455859876437126964949598726124545978501547019010261968650526517542821103000;
            5'd2: xpb[50] = 1024'd120168479977485886627060551072366993463544666875825913357294409915488558363531012512815331699512297837994658797609825892054812703532517401925103860560699038349268679036611125834622815602237643921228863902999323615349714936982638896273933150069644804663079294038132033926896565964091890920182363208460047721669;
            5'd3: xpb[50] = 1024'd118219372124166459241191362906143273822967786750871027971875687340744389876641949314215461941939609602270413492685992120792687134878165935610075728332883037057057681270131080083119103807597863021188197050305365499842391980363509957928410440262852482361208989350139521875291584909173519871714199899377274340338;
            5'd4: xpb[50] = 1024'd116270264270847031855322174739919554182390906625916142586456964766000221389752886115615592184366921366546168187762158349530561566223814469295047596105067035764846683503651034331615392012958082121147530197611407384335069023744381019582887730456060160059338684662147009823686603854255148823246036590294500959007;
            5'd5: xpb[50] = 1024'd114321156417527604469452986573695834541814026500961257201038242191256052902863822917015722426794233130821922882838324578268435997569463002980019463877251034472635685737170988580111680218318301221106863344917449268827746067125252081237365020649267837757468379974154497772081622799336777774777873281211727577676;
            5'd6: xpb[50] = 1024'd112372048564208177083583798407472114901237146376006371815619519616511884415974759718415852669221544895097677577914490807006310428915111536664991331649435033180424687970690942828607968423678520321066196492223491153320423110506123142891842310842475515455598075286161985720476641744418406726309709972128954196345;
            5'd7: xpb[50] = 1024'd110422940710888749697714610241248395260660266251051486430200797041767715929085696519815982911648856659373432272990657035744184860260760070349963199421619031888213690204210897077104256629038739421025529639529533037813100153886994204546319601035683193153727770598169473668871660689500035677841546663046180815014;
            5'd8: xpb[50] = 1024'd108473832857569322311845422075024675620083386126096601044782074467023547442196633321216113154076168423649186968066823264482059291606408604034935067193803030596002692437730851325600544834398958520984862786835574922305777197267865266200796891228890870851857465910176961617266679634581664629373383353963407433683;
            5'd9: xpb[50] = 1024'd106524725004249894925976233908800955979506506001141715659363351892279378955307570122616243396503480187924941663142989493219933722952057137719906934965987029303791694671250805574096833039759177620944195934141616806798454240648736327855274181422098548549987161222184449565661698579663293580905220044880634052352;
            5'd10: xpb[50] = 1024'd104575617150930467540107045742577236338929625876186830273944629317535210468418506924016373638930791952200696358219155721957808154297705671404878802738171028011580696904770759822593121245119396720903529081447658691291131284029607389509751471615306226248116856534191937514056717524744922532437056735797860671021;
            5'd11: xpb[50] = 1024'd102626509297611040154237857576353516698352745751231944888525906742791041981529443725416503881358103716476451053295321950695682585643354205089850670510355026719369699138290714071089409450479615820862862228753700575783808327410478451164228761808513903946246551846199425462451736469826551483968893426715087289690;
            5'd12: xpb[50] = 1024'd100677401444291612768368669410129797057775865626277059503107184168046873494640380526816634123785415480752205748371488179433557016989002738774822538282539025427158701371810668319585697655839834920822195376059742460276485370791349512818706052001721581644376247158206913410846755414908180435500730117632313908359;
            5'd13: xpb[50] = 1024'd98728293590972185382499481243906077417198985501322174117688461593302705007751317328216764366212727245027960443447654408171431448334651272459794406054723024134947703605330622568081985861200054020781528523365784344769162414172220574473183342194929259342505942470214401359241774359989809387032566808549540527028;
            5'd14: xpb[50] = 1024'd96779185737652757996630293077682357776622105376367288732269739018558536520862254129616894608640039009303715138523820636909305879680299806144766273826907022842736705838850576816578274066560273120740861670671826229261839457553091636127660632388136937040635637782221889307636793305071438338564403499466767145697;
            5'd15: xpb[50] = 1024'd94830077884333330610761104911458638136045225251412403346851016443814368033973190931017024851067350773579469833599986865647180311025948339829738141599091021550525708072370531065074562271920492220700194817977868113754516500933962697782137922581344614738765333094229377256031812250153067290096240190383993764366;
            5'd16: xpb[50] = 1024'd92880970031013903224891916745234918495468345126457517961432293869070199547084127732417155093494662537855224528676153094385054742371596873514710009371275020258314710305890485313570850477280711320659527965283909998247193544314833759436615212774552292436895028406236865204426831195234696241628076881301220383035;
            5'd17: xpb[50] = 1024'd90931862177694475839022728579011198854891465001502632576013571294326031060195064533817285335921974302130979223752319323122929173717245407199681877143459018966103712539410439562067138682640930420618861112589951882739870587695704821091092502967759970135024723718244353152821850140316325193159913572218447001704;
            5'd18: xpb[50] = 1024'd88982754324375048453153540412787479214314584876547747190594848719581862573306001335217415578349286066406733918828485551860803605062893940884653744915643017673892714772930393810563426888001149520578194259895993767232547631076575882745569793160967647833154419030251841101216869085397954144691750263135673620373;
            5'd19: xpb[50] = 1024'd87033646471055621067284352246563759573737704751592861805176126144837694086416938136617545820776597830682488613904651780598678036408542474569625612687827016381681717006450348059059715093361368620537527407202035651725224674457446944400047083354175325531284114342259329049611888030479583096223586954052900239042;
            5'd20: xpb[50] = 1024'd85084538617736193681415164080340039933160824626637976419757403570093525599527874938017676063203909594958243308980818009336552467754191008254597480460011015089470719239970302307556003298721587720496860554508077536217901717838318006054524373547383003229413809654266816998006906975561212047755423644970126857711;
            5'd21: xpb[50] = 1024'd83135430764416766295545975914116320292583944501683091034338680995349357112638811739417806305631221359233998004056984238074426899099839541939569348232195013797259721473490256556052291504081806820456193701814119420710578761219189067709001663740590680927543504966274304946401925920642840999287260335887353476380;
            5'd22: xpb[50] = 1024'd81186322911097338909676787747892600652007064376728205648919958420605188625749748540817936548058533123509752699133150466812301330445488075624541216004379012505048723707010210804548579709442025920415526849120161305203255804600060129363478953933798358625673200278281792894796944865724469950819097026804580095049;
            5'd23: xpb[50] = 1024'd79237215057777911523807599581668881011430184251773320263501235845861020138860685342218066790485844887785507394209316695550175761791136609309513083776563011212837725940530165053044867914802245020374859996426203189695932847980931191017956244127006036323802895590289280843191963810806098902350933717721806713718;
            5'd24: xpb[50] = 1024'd77288107204458484137938411415445161370853304126818434878082513271116851651971622143618197032913156652061262089285482924288050193136785142994484951548747009920626728174050119301541156120162464120334193143732245074188609891361802252672433534320213714021932590902296768791586982755887727853882770408639033332387;
            5'd25: xpb[50] = 1024'd75338999351139056752069223249221441730276424001863549492663790696372683165082558945018327275340468416337016784361649153025924624482433676679456819320931008628415730407570073550037444325522683220293526291038286958681286934742673314326910824513421391720062286214304256739982001700969356805414607099556259951056;
            5'd26: xpb[50] = 1024'd73389891497819629366200035082997722089699543876908664107245068121628514678193495746418457517767780180612771479437815381763799055828082210364428687093115007336204732641090027798533732530882902320252859438344328843173963978123544375981388114706629069418191981526311744688377020646050985756946443790473486569725;
            5'd27: xpb[50] = 1024'd71440783644500201980330846916774002449122663751953778721826345546884346191304432547818587760195091944888526174513981610501673487173730744049400554865299006043993734874609982047030020736243121420212192585650370727666641021504415437635865404899836747116321676838319232636772039591132614708478280481390713188394;
            5'd28: xpb[50] = 1024'd69491675791180774594461658750550282808545783626998893336407622972140177704415369349218718002622403709164280869590147839239547918519379277734372422637483004751782737108129936295526308941603340520171525732956412612159318064885286499290342695093044424814451372150326720585167058536214243660010117172307939807063;
            5'd29: xpb[50] = 1024'd67542567937861347208592470584326563167968903502044007950988900397396009217526306150618848245049715473440035564666314067977422349865027811419344290409667003459571739341649890544022597146963559620130858880262454496651995108266157560944819985286252102512581067462334208533562077481295872611541953863225166425732;
            5'd30: xpb[50] = 1024'd65593460084541919822723282418102843527392023377089122565570177822651840730637242952018978487477027237715790259742480296715296781210676345104316158181851002167360741575169844792518885352323778720090192027568496381144672151647028622599297275479459780210710762774341696481957096426377501563073790554142393044401;
            5'd31: xpb[50] = 1024'd63644352231222492436854094251879123886815143252134237180151455247907672243748179753419108729904339001991544954818646525453171212556324878789288025954035000875149743808689799041015173557683997820049525174874538265637349195027899684253774565672667457908840458086349184430352115371459130514605627245059619663070;
        endcase
    end

    always_comb begin
        case(flag[17][5:0])
            6'd0: xpb[51] = 1024'd0;
            6'd1: xpb[51] = 1024'd92880970031013903224891916745234918495468345126457517961432293869070199547084127732417155093494662537855224528676153094385054742371596873514710009371275020258314710305890485313570850477280711320659527965283909998247193544314833759436615212774552292436895028406236865204426831195234696241628076881301220383035;
            6'd2: xpb[51] = 1024'd61695244377903065050984906085655404246238263127179351794732732673163503756859116554819238972331650766267299649894812754191045643901973412474259893726218999582938746042209753289511461763044216920008858322180580150130026238408770745908251855865875135606970153398356672378747134316540759466137463935976846281739;
            6'd3: xpb[51] = 1024'd30509518724792226877077895426075889997008181127901185628033171477256807966634105377221322851168638994679374771113472413997036545432349951433809778081162978907562781778529021265452073048807722519358188679077250302012858932502707732379888498957197978777045278390476479553067437437846822690646850990652472180443;
            6'd4: xpb[51] = 1024'd123390488755806130101969812171310808492476526254358703589465465346327007513718233109638477944663301532534599299789625508382091287803946824948519787452437999165877492084419506579022923526088433840017716644361160300260052476817541491816503711731750271213940306796713344757494268633081518932274927871953692563478;
            6'd5: xpb[51] = 1024'd92204763102695291928062801511731294243246444255080537422765904150420311723493221932040561823500289760946674421008285168188082189334323363908069671807381978490501527820738774554963534811851939439367047001257830452142885170911478478288140354823073114384015431788833151931814571754387582156784314926629318462182;
            6'd6: xpb[51] = 1024'd61019037449584453754155790852151779994016362255802371256066342954513615933268210754442645702337277989358749542226944827994073090864699902867619556162325957815125563557058042530904146097615445038716377358154500604025717865005415464759776997914395957554090556780952959106134874875693645381293701981304944360886;
            6'd7: xpb[51] = 1024'd29833311796473615580248780192572265744786280256524205089366781758606920143043199576844729581174266217770824663445604487800063992395076441827169440517269937139749599293377310506844757383378950638065707715051170755908550559099352451231413641005718800724165681773072766280455177996999708605803089035980570259590;
            6'd8: xpb[51] = 1024'd122714281827487518805140696937807184240254625382981723050799075627677119690127327309261884674668928755626049192121757582185118734766673315341879449888544957398064309599267795820415607860659661958725235680335080754155744103414186210668028853780271093161060710179309631484882009192234404847431165917281790642625;
            6'd9: xpb[51] = 1024'd91528556174376680631233686278227669991024543383703556884099514431770423899902316131663968553505916984038124313340417241991109636297049854301429334243488936722688345335587063796356219146423167558074566037231750906038576797508123197139665496871593936331135835171429438659202312313540468071940552971957416541329;
            6'd10: xpb[51] = 1024'd60342830521265842457326675618648155741794461384425390717399953235863728109677304954066052432342905212450199434559076901797100537827426393260979218598432916047312381071906331772296830432186673157423896394128421057921409491602060183611302139962916779501210960163549245833522615434846531296449940026633042440033;
            6'd11: xpb[51] = 1024'd29157104868155004283419664959068641492564379385147224550700392039957032319452293776468136311179893440862274555777736561603091439357802932220529102953376895371936416808225599748237441717950178756773226751025091209804242185695997170082938783054239622671286085155669053007842918556152594520959327081308668338737;
            6'd12: xpb[51] = 1024'd122038074899168907508311581704303559988032724511604742512132685909027231866536421508885291404674555978717499084453889655988146181729399805735239112324651915630251127114116085061808292195230890077432754716309001208051435730010830929519553995828791915108181113561905918212269749751387290762587403962609888721772;
            6'd13: xpb[51] = 1024'd90852349246058069334404571044724045738802642512326576345433124713120536076311410331287375283511544207129574205672549315794137083259776344694788996679595894954875162850435353037748903480994395676782085073205671359934268424104767915991190638920114758278256238554025725386590052872693353987096791017285514620476;
            6'd14: xpb[51] = 1024'd59666623592947231160497560385144531489572560513048410178733563517213840286086399153689459162348532435541649326891208975600127984790152883654338881034539874279499198586754621013689514766757901276131415430102341511817101118198704902462827282011437601448331363546145532560910355993999417211606178071961140519180;
            6'd15: xpb[51] = 1024'd28480897939836392986590549725565017240342478513770244012034002321307144495861387976091543041185520663953724448109868635406118886320529422613888765389483853604123234323073888989630126052521406875480745786999011663699933812292641888934463925102760444618406488538265339735230659115305480436115565126636766417884;
            6'd16: xpb[51] = 1024'd121361867970850296211482466470799935735810823640227761973466296190377344042945515708508698134680183201808948976786021729791173628692126296128598774760758873862437944628964374303200976529802118196140273752282921661947127356607475648371079137877312737055301516944502204939657490310540176677743642007937986800919;
            6'd17: xpb[51] = 1024'd90176142317739458037575455811220421486580741640949595806766734994470648252720504530910782013517171430221024098004681389597164530222502835088148659115702853187061980365283642279141587815565623795489604109179591813829960050701412634842715780968635580225376641936622012113977793431846239902253029062613612699623;
            6'd18: xpb[51] = 1024'd58990416664628619863668445151640907237350659641671429640067173798563952462495493353312865892354159658633099219223341049403155431752879374047698543470646832511686016101602910255082199101329129394838934466076261965712792744795349621314352424059958423395451766928741819288298096553152303126762416117289238598327;
            6'd19: xpb[51] = 1024'd27804691011517781689761434492061392988120577642393263473367612602657256672270482175714949771191147887045174340442000709209146333283255913007248427825590811836310051837922178231022810387092634994188264822972932117595625438889286607785989067151281266565526891920861626462618399674458366351271803171964864497031;
            6'd20: xpb[51] = 1024'd120685661042531684914653351237296311483588922768850781434799906471727456219354609908132104864685810424900398869118153803594201075654852786521958437196865832094624762143812663544593660864373346314847792788256842115842818983204120367222604279925833559002421920327098491667045230869693062592899880053266084880066;
            6'd21: xpb[51] = 1024'd89499935389420846740746340577716797234358840769572615268100345275820760429129598730534188743522798653312473990336813463400191977185229325481508321551809811419248797880131931520534272150136851914197123145153512267725651677298057353694240923017156402172497045319218298841365533990999125817409267107941710778770;
            6'd22: xpb[51] = 1024'd58314209736310008566839329918137282985128758770294449101400784079914064638904587552936272622359786881724549111555473123206182878715605864441058205906753790743872833616451199496474883435900357513546453502050182419608484371391994340165877566108479245342572170311338106015685837112305189041918654162617336677474;
            6'd23: xpb[51] = 1024'd27128484083199170392932319258557768735898676771016282934701222884007368848679576375338356501196775110136624232774132783012173780245982403400608090261697770068496869352770467472415494721663863112895783858946852571491317065485931326637514209199802088512647295303457913190006140233611252266428041217292962576178;
            6'd24: xpb[51] = 1024'd120009454114213073617824236003792687231367021897473800896133516753077568395763704107755511594691437647991848761450285877397228522617579276915318099632972790326811579658660952785986345198944574433555311824230762569738510609800765086074129421974354380949542323709694778394432971428845948508056118098594182959213;
            6'd25: xpb[51] = 1024'd88823728461102235443917225344213172982136939898195634729433955557170872605538692930157595473528425876403923882668945537203219424147955815874867983987916769651435615394980220761926956484708080032904642181127432721621343303894702072545766065065677224119617448701814585568753274550152011732565505153269808857917;
            6'd26: xpb[51] = 1024'd57638002807991397270010214684633658732906857898917468562734394361264176815313681752559679352365414104815999003887605197009210325678332354834417868342860748976059651131299488737867567770471585632253972538024102873504175997988639059017402708157000067289692573693934392743073577671458074957074892207945434756621;
            6'd27: xpb[51] = 1024'd26452277154880559096103204025054144483676775899639302396034833165357481025088670574961763231202402333228074125106264856815201227208708893793967752697804728300683686867618756713808179056235091231603302894920773025387008692082576045489039351248322910459767698686054199917393880792764138181584279262621060655325;
            6'd28: xpb[51] = 1024'd119333247185894462320995120770289062979145121026096820357467127034427680572172798307378918324697064871083298653782417951200255969580305767308677762069079748558998397173509242027379029533515802552262830860204683023634202236397409804925654564022875202896662727092291065121820711987998834423212356143922281038360;
            6'd29: xpb[51] = 1024'd88147521532783624147088110110709548729915039026818654190767565838520984781947787129781002203534053099495373775001077611006246871110682306268227646424023727883622432909828510003319640819279308151612161217101353175517034930491346791397291207114198046066737852084410872296141015109304897647721743198597906937064;
            6'd30: xpb[51] = 1024'd56961795879672785973181099451130034480684957027540488024068004642614288991722775952183086082371041327907448896219737270812237772641058845227777530778967707208246468646147777979260252105042813750961491573998023327399867624585283777868927850205520889236812977076530679470461318230610960872231130253273532835768;
            6'd31: xpb[51] = 1024'd25776070226561947799274088791550520231454875028262321857368443446707593201497764774585169961208029556319524017438396930618228674171435384187327415133911686532870504382467045955200863390806319350310821930894693479282700318679220764340564493296843732406888102068650486644781621351917024096740517307949158734472;
            6'd32: xpb[51] = 1024'd118657040257575851024166005536785438726923220154719839818800737315777792748581892507002325054702692094174748546114550025003283416543032257702037424505186706791185214688357531268771713868087030670970349896178603477529893862994054523777179706071396024843783130474887351849208452547151720338368594189250379117507;
            6'd33: xpb[51] = 1024'd87471314604465012850258994877205924477693138155441673652101176119871096958356881329404408933539680322586823667333209684809274318073408796661587308860130686115809250424676799244712325153850536270319680253075273629412726557087991510248816349162718868013858255467007159023528755668457783562877981243926005016211;
            6'd34: xpb[51] = 1024'd56285588951354174676351984217626410228463056156163507485401614923964401168131870151806492812376668550998898788551869344615265219603785335621137193215074665440433286160996067220652936439614041869669010609971943781295559251181928496720452992254041711183933380459126966197849058789763846787387368298601630914915;
            6'd35: xpb[51] = 1024'd25099863298243336502444973558046895979232974156885341318702053728057705377906858974208576691213656779410973909770529004421256121134161874580687077570018644765057321897315335196593547725377547469018340966868613933178391945275865483192089635345364554354008505451246773372169361911069910011896755353277256813619;
            6'd36: xpb[51] = 1024'd117980833329257239727336890303281814474701319283342859280134347597127904924990986706625731784708319317266198438446682098806310863505758748095397086941293665023372032203205820510164398202658258789677868932152523931425585489590699242628704848119916846790903533857483638576596193106304606253524832234578477196654;
            6'd37: xpb[51] = 1024'd86795107676146401553429879643702300225471237284064693113434786401221209134765975529027815663545307545678273559665341758612301765036135287054946971296237644347996067939525088486105009488421764389027199289049194083308418183684636229100341491211239689960978658849603445750916496227610669478034219289254103095358;
            6'd38: xpb[51] = 1024'd55609382023035563379522868984122785976241155284786526946735225205314513344540964351429899542382295774090348680884001418418292666566511826014496855651181623672620103675844356462045620774185269988376529645945864235191250877778573215571978134302562533131053783841723252925236799348916732702543606343929728994062;
            6'd39: xpb[51] = 1024'd24423656369924725205615858324543271727011073285508360780035664009407817554315953173831983421219284002502423802102661078224283568096888364974046740006125602997244139412163624437986232059948775587725860002842534387074083571872510202043614777393885376301128908833843060099557102470222795927052993398605354892766;
            6'd40: xpb[51] = 1024'd117304626400938628430507775069778190222479418411965878741467957878478017101400080906249138514713946540357648330778814172609338310468485238488756749377400623255558849718054109751557082537229486908385387968126444385321277116187343961480229990168437668738023937240079925303983933665457492168681070279906575275801;
            6'd41: xpb[51] = 1024'd86118900747827790256600764410198675973249336412687712574768396682571321311175069728651222393550934768769723451997473832415329211998861777448306633732344602580182885454373377727497693822992992507734718325023114537204109810281280947951866633259760511908099062232199732478304236786763555393190457334582201174505;
            6'd42: xpb[51] = 1024'd54933175094716952082693753750619161724019254413409546408068835486664625520950058551053306272387922997181798573216133492221320113529238316407856518087288581904806921190692645703438305108756498107084048681919784689086942504375217934423503276351083355078174187224319539652624539908069618617699844389257827073209;
            6'd43: xpb[51] = 1024'd23747449441606113908786743091039647474789172414131380241369274290757929730725047373455390151224911225593873694434793152027311015059614855367406402442232561229430956927011913679378916394520003706433379038816454840969775198469154920895139919442406198248249312216439346826944843029375681842209231443933452971913;
            6'd44: xpb[51] = 1024'd116628419472620017133678659836274565970257517540588898202801568159828129277809175105872545244719573763449098223110946246412365757431211728882116411813507581487745667232902398992949766871800715027092907004100364839216968742783988680331755132216958490685144340622676212031371674224610378083837308325234673354948;
            6'd45: xpb[51] = 1024'd85442693819509178959771649176695051721027435541310732036102006963921433487584163928274629123556561991861173344329605906218356658961588267841666296168451560812369702969221666968890378157564220626442237360997034991099801436877925666803391775308281333855219465614796019205691977345916441308346695379910299253652;
            6'd46: xpb[51] = 1024'd54256968166398340785864638517115537471797353542032565869402445768014737697359152750676713002393550220273248465548265566024347560491964806801216180523395540136993738705540934944830989443327726225791567717893705142982634130971862653275028418399604177025294590606915826380012280467222504532856082434585925152356;
            6'd47: xpb[51] = 1024'd23071242513287502611957627857536023222567271542754399702702884572108041907134141573078796881230538448685323586766925225830338462022341345760766064878339519461617774441860202920771600729091231825140898074790375294865466825065799639746665061490927020195369715599035633554332583588528567757365469489261551051060;
            6'd48: xpb[51] = 1024'd115952212544301405836849544602770941718035616669211917664135178441178241454218269305495951974725200986540548115443078320215393204393938219275476074249614539719932484747750688234342451206371943145800426040074285293112660369380633399183280274265479312632264744005272498758759414783763263998993546370562771434095;
            6'd49: xpb[51] = 1024'd84766486891190567662942533943191427468805534669933751497435617245271545663993258127898035853562189214952623236661737980021384105924314758235025958604558519044556520484069956210283062492135448745149756396970955444995493063474570385654916917356802155802339868997392305933079717905069327223502933425238397332799;
            6'd50: xpb[51] = 1024'd53580761238079729489035523283611913219575452670655585330736056049364849873768246950300119732399177443364698357880397639827375007454691297194575842959502498369180556220389224186223673777898954344499086753867625596878325757568507372126553560448124998972414993989512113107400021026375390448012320479914023231503;
            6'd51: xpb[51] = 1024'd22395035584968891315128512624032398970345370671377419164036494853458154083543235772702203611236165671776773479099057299633365908985067836154125727314446477693804591956708492162164285063662459943848417110764295748761158451662444358598190203539447842142490118981631920281720324147681453672521707534589649130207;
            6'd52: xpb[51] = 1024'd115276005615982794540020429369267317465813715797834937125468788722528353630627363505119358704730828209631998007775210394018420651356664709668835736685721497952119302262598977475735135540943171264507945076048205747008351995977278118034805416314000134579385147387868785486147155342916149914149784415890869513242;
            6'd53: xpb[51] = 1024'd84090279962871956366113418709687803216583633798556770958769227526621657840402352327521442583567816438044073128993870053824411552887041248628385621040665477276743337998918245451675746826706676863857275432944875898891184690071215104506442059405322977749460272379988592660467458464222213138659171470566495411946;
            6'd54: xpb[51] = 1024'd52904554309761118192206408050108288967353551799278604792069666330714962050177341149923526462404804666456148250212529713630402454417417787587935505395609456601367373735237513427616358112470182463206605789841546050774017384165152090978078702496645820919535397372108399834787761585528276363168558525242121310650;
            6'd55: xpb[51] = 1024'd21718828656650280018299397390528774718123469800000438625370105134808266259952329972325610341241792894868223371431189373436393355947794326547485389750553435925991409471556781403556969398233688062555936146738216202656850078259089077449715345587968664089610522364228207009108064706834339587677945579917747209354;
            6'd56: xpb[51] = 1024'd114599798687664183243191314135763693213591814926457956586802399003878465807036457704742765434736455432723447900107342467821448098319391200062195399121828456184306119777447266717127819875514399383215464112022126200904043622573922836886330558362520956526505550770465072213534895902069035829306022461218967592389;
            6'd57: xpb[51] = 1024'd83414073034553345069284303476184178964361732927179790420102837807971770016811446527144849313573443661135523021326002127627438999849767739021745283476772435508930155513766534693068431161277904982564794468918796352786876316667859823357967201453843799696580675762584879387855199023375099053815409515894593491093;
            6'd58: xpb[51] = 1024'd52228347381442506895377292816604664715131650927901624253403276612065074226586435349546933192410431889547598142544661787433429901380144277981295167831716414833554191250085802669009042447041410581914124825815466504669709010761796809829603844545166642866655800754704686562175502144681162278324796570570219389797;
            6'd59: xpb[51] = 1024'd21042621728331668721470282157025150465901568928623458086703715416158378436361424171949017071247420117959673263763321447239420802910520816940845052186660394158178226986405070644949653732804916181263455182712136656552541704855733796301240487636489486036730925746824493736495805265987225502834183625245845288501;
            6'd60: xpb[51] = 1024'd113923591759345571946362198902260068961369914055080976048136009285228577983445551904366172164742082655814897792439474541624475545282117690455555061557935414416492937292295555958520504210085627501922983147996046654799735249170567555737855700411041778473625954153061358940922636461221921744462260506547065671536;
            6'd61: xpb[51] = 1024'd82737866106234733772455188242680554712139832055802809881436448089321882193220540726768256043579070884226972913658134201430466446812494229415104945912879393741116973028614823934461115495849133101272313504892716806682567943264504542209492343502364621643701079145181166115242939582527984968971647561222691570240;
            6'd62: xpb[51] = 1024'd51552140453123895598548177583101040462909750056524643714736886893415186402995529549170339922416059112639048034876793861236457348342870768374654830267823373065741008764934091910401726781612638700621643861789386958565400637358441528681128986593687464813776204137300973289563242703834048193481034615898317468944;
            6'd63: xpb[51] = 1024'd20366414800013057424641166923521526213679668057246477548037325697508490612770518371572423801253047341051123156095453521042448249873247307334204714622767352390365044501253359886342338067376144299970974218686057110448233331452378515152765629685010307983851329129420780463883545825140111417990421670573943367648;
        endcase
    end

    always_comb begin
        case(flag[17][11:6])
            6'd0: xpb[52] = 1024'd0;
            6'd1: xpb[52] = 1024'd113247384831026960649533083668756444709148013183703995509469619566578690159854646103989578894747709878906347684771606615427502992244844180848914723994042372648679754807143845199913188544656855620630502183969967108695426875767212274589380842459562600420746357535657645668310377020374807659618498551875163750683;
            6'd2: xpb[52] = 1024'd102428073977929179900267239932698456673597599241672306890807384068180484982400153297964086574837745448369545962085719796275942143648468027142669322971753704363668835044716473062196137897796505519950806759552694371026492901313527776213783115235895751574672811657198233306514225966820982302118307277124733017035;
            6'd3: xpb[52] = 1024'd91608763124831399151001396196640468638047185299640618272145148569782279804945660491938594254927781017832744239399832977124381295052091873436423921949465036078657915282289100924479087250936155419271111335135421633357558926859843277838185388012228902728599265778738820944718074913267156944618116002374302283387;
            6'd4: xpb[52] = 1024'd80789452271733618401735552460582480602496771357608929653482913071384074627491167685913101935017816587295942516713946157972820446455715719730178520927176367793646995519861728786762036604075805318591415910718148895688624952406158779462587660788562053882525719900279408582921923859713331587117924727623871549739;
            6'd5: xpb[52] = 1024'd69970141418635837652469708724524492566946357415577241034820677572985869450036674879887609615107852156759140794028059338821259597859339566023933119904887699508636075757434356649044985957215455217911720486300876158019690977952474281086989933564895205036452174021819996221125772806159506229617733452873440816091;
            6'd6: xpb[52] = 1024'd59150830565538056903203864988466504531395943473545552416158442074587664272582182073862117295197887726222339071342172519669698749262963412317687718882599031223625155995006984511327935310355105117232025061883603420350757003498789782711392206341228356190378628143360583859329621752605680872117542178123010082443;
            6'd7: xpb[52] = 1024'd48331519712440276153938021252408516495845529531513863797496206576189459095127689267836624975287923295685537348656285700518137900666587258611442317860310362938614236232579612373610884663494755016552329637466330682681823029045105284335794479117561507344305082264901171497533470699051855514617350903372579348795;
            6'd8: xpb[52] = 1024'd37512208859342495404672177516350528460295115589482175178833971077791253917673196461811132655377958865148735625970398881366577052070211104905196916838021694653603316470152240235893834016634404915872634213049057945012889054591420785960196751893894658498231536386441759135737319645498030157117159628622148615147;
            6'd9: xpb[52] = 1024'd26692898006244714655406333780292540424744701647450486560171735579393048740218703655785640335467994434611933903284512062215016203473834951198951515815733026368592396707724868098176783369774054815192938788631785207343955080137736287584599024670227809652157990507982346773941168591944204799616968353871717881499;
            6'd10: xpb[52] = 1024'd15873587153146933906140490044234552389194287705418797941509500080994843562764210849760148015558030004075132180598625243063455354877458797492706114793444358083581476945297495960459732722913704714513243364214512469675021105684051789209001297446560960806084444629522934412145017538390379442116777079121287147851;
            6'd11: xpb[52] = 1024'd5054276300049153156874646308176564353643873763387109322847264582596638385309718043734655695648065573538330457912738423911894506281082643786460713771155689798570557182870123822742682076053354613833547939797239732006087131230367290833403570222894111960010898751063522050348866484836554084616585804370856414203;
            6'd12: xpb[52] = 1024'd118301661131076113806407729976933009062791886947091104832316884149175328545164364147724234590395775452444678142684345039339397498525926824635375437765198062447250311990013969022655870620710210234464050123767206840701514006997579565422784412682456712380757256286721167718659243505211361744235084356246020164886;
            6'd13: xpb[52] = 1024'd107482350277978333057141886240875021027241473005059416213654648650777123367709871341698742270485811021907876419998458220187836649929550670929130036742909394162239392227586596884938819973849860133784354699349934103032580032543895067047186685458789863534683710408261755356863092451657536386734893081495589431238;
            6'd14: xpb[52] = 1024'd96663039424880552307876042504817032991691059063027727594992413152378918190255378535673249950575846591371074697312571401036275801333174517222884635720620725877228472465159224747221769326989510033104659274932661365363646058090210568671588958235123014688610164529802342995066941398103711029234701806745158697590;
            6'd15: xpb[52] = 1024'd85843728571782771558610198768759044956140645120996038976330177653980713012800885729647757630665882160834272974626684581884714952736798363516639234698332057592217552702731852609504718680129159932424963850515388627694712083636526070295991231011456165842536618651342930633270790344549885671734510531994727963942;
            6'd16: xpb[52] = 1024'd75024417718684990809344355032701056920590231178964350357667942155582507835346392923622265310755917730297471251940797762733154104140422209810393833676043389307206632940304480471787668033268809831745268426098115890025778109182841571920393503787789316996463072772883518271474639290996060314234319257244297230294;
            6'd17: xpb[52] = 1024'd64205106865587210060078511296643068885039817236932661739005706657184302657891900117596772990845953299760669529254910943581593255544046056104148432653754721022195713177877108334070617386408459731065573001680843152356844134729157073544795776564122468150389526894424105909678488237442234956734127982493866496646;
            6'd18: xpb[52] = 1024'd53385796012489429310812667560585080849489403294900973120343471158786097480437407311571280670935988869223867806569024124430032406947669902397903031631466052737184793415449736196353566739548109630385877577263570414687910160275472575169198049340455619304315981015964693547882337183888409599233936707743435762998;
            6'd19: xpb[52] = 1024'd42566485159391648561546823824527092813938989352869284501681235660387892302982914505545788351026024438687066083883137305278471558351293748691657630609177384452173873653022364058636516092687759529706182152846297677018976185821788076793600322116788770458242435137505281186086186130334584241733745432993005029350;
            6'd20: xpb[52] = 1024'd31747174306293867812280980088469104778388575410837595883019000161989687125528421699520296031116060008150264361197250486126910709754917594985412229586888716167162953890594991920919465445827409429026486728429024939350042211368103578418002594893121921612168889259045868824290035076780758884233554158242574295702;
            6'd21: xpb[52] = 1024'd20927863453196087063015136352411116742838161468805907264356764663591481948073928893494803711206095577613462638511363666975349861158541441279166828564600047882152034128167619783202414798967059328346791304011752201681108236914419080042404867669455072766095343380586456462493884023226933526733362883492143562054;
            6'd22: xpb[52] = 1024'd10108552600098306313749292616353128707287747526774218645694529165193276770619436087469311391296131147076660915825476847823789012562165287572921427542311379597141114365740247645485364152106709227667095879594479464012174262460734581666807140445788223920021797502127044100697732969673108169233171608741712828406;
            6'd23: xpb[52] = 1024'd123355937431125266963282376285109573416435760710478214155164148731771966930474082191458890286043841025983008600597083463251292004807009468421836151536353752245820869172884092845398552696763564848297598063564446572707601138227946856256187982905350824340768155037784689769008109990047915828851670160616876579089;
            6'd24: xpb[52] = 1024'd112536626578027486214016532549051585380885346768446525536501913233373761753019589385433397966133876595446206877911196644099731156210633314715590750514065083960809949410456720707681502049903214747617902639147173835038667163774262357880590255681683975494694609159325277407211958936494090471351478885866445845441;
            6'd25: xpb[52] = 1024'd101717315724929705464750688812993597345334932826414836917839677734975556575565096579407905646223912164909405155225309824948170307614257161009345349491776415675799029648029348569964451403042864646938207214729901097369733189320577859504992528458017126648621063280865865045415807882940265113851287611116015111793;
            6'd26: xpb[52] = 1024'd90898004871831924715484845076935609309784518884383148299177442236577351398110603773382413326313947734372603432539423005796609459017881007303099948469487747390788109885601976432247400756182514546258511790312628359700799214866893361129394801234350277802547517402406452683619656829386439756351096336365584378145;
            6'd27: xpb[52] = 1024'd80078694018734143966219001340877621274234104942351459680515206738179146220656110967356921006403983303835801709853536186645048610421504853596854547447199079105777190123174604294530350109322164445578816365895355622031865240413208862753797074010683428956473971523947040321823505775832614398850905061615153644497;
            6'd28: xpb[52] = 1024'd69259383165636363216953157604819633238683691000319771061852971239780941043201618161331428686494018873298999987167649367493487761825128699890609146424910410820766270360747232156813299462461814344899120941478082884362931265959524364378199346787016580110400425645487627960027354722278789041350713786864722910849;
            6'd29: xpb[52] = 1024'd58440072312538582467687313868761645203133277058288082443190735741382735865747125355305936366584054442762198264481762548341926913228752546184363745402621742535755350598319860019096248815601464244219425517060810146693997291505839866002601619563349731264326879767028215598231203668724963683850522512114292177201;
            6'd30: xpb[52] = 1024'd47620761459440801718421470132703657167582863116256393824528500242984530688292632549280444046674090012225396541795875729190366064632376392478118344380333074250744430835892487881379198168741114143539730092643537409025063317052155367627003892339682882418253333888568803236435052615171138326350331237363861443553;
            6'd31: xpb[52] = 1024'd36801450606343020969155626396645669132032449174224705205866264744586325510838139743254951726764125581688594819109988910038805216036000238771872943358044405965733511073465115743662147521880764042860034668226264671356129342598470869251406165116016033572179788010109390874638901561617312968850139962613430709905;
            6'd32: xpb[52] = 1024'd25982139753245240219889782660587681096482035232193016587204029246188120333383646937229459406854161151151793096424102090887244367439624085065627542335755737680722591311037743605945096875020413942180339243808991933687195368144786370875808437892349184726106242131649978512842750508063487611349948687862999976257;
            6'd33: xpb[52] = 1024'd15162828900147459470623938924529693060931621290161327968541793747789915155929154131203967086944196720614991373738215271735683518843247931359382141313467069395711671548610371468228046228160063841500643819391719196018261393691101872500210710668682335880032696253190566151046599454509662253849757413112569242609;
            6'd34: xpb[52] = 1024'd4343518047049678721358095188471705025381207348129639349879558249391709978474661325178474767034232290078189651052328452584122670246871777653136740291178401110700751786182999330510995581299713740820948394974446458349327419237417374124612983445015487033959150374731153789250448400955836896349566138362138508961;
            6'd35: xpb[52] = 1024'd117590902878076639370891178857228149734529220531833634859349177815970400138329307429168053661781942168984537335823935068011625662491715958502051464285220773759380506593326844530424184125956569361451450578944413567044754295004629648713993825904578087454705507910388799457560825421330644555968064690237302259644;
            6'd36: xpb[52] = 1024'd106771592024978858621625335121170161698978806589801946240686942317572194960874814623142561341871977738447735613138048248860064813895339804795806063262932105474369586830899472392707133479096219260771755154527140829375820320550945150338396098680911238608631962031929387095764674367776819198467873415486871525996;
            6'd37: xpb[52] = 1024'd95952281171881077872359491385112173663428392647770257622024706819173989783420321817117069021962013307910933890452161429708503965298963651089560662240643437189358667068472100254990082832235869160092059730109868091706886346097260651962798371457244389762558416153469974733968523314222993840967682140736440792348;
            6'd38: xpb[52] = 1024'd85132970318783297123093647649054185627877978705738569003362471320775784605965829011091576702052048877374132167766274610556943116702587497383315261218354768904347747306044728117273032185375519059412364305692595354037952371643576153587200644233577540916484870275010562372172372260669168483467490865986010058700;
            6'd39: xpb[52] = 1024'd74313659465685516373827803912996197592327564763706880384700235822377579428511336205066084382142084446837330445080387791405382268106211343677069860196066100619336827543617355979555981538515168958732668881275322616369018397189891655211602917009910692070411324396551150010376221207115343125967299591235579325052;
            6'd40: xpb[52] = 1024'd63494348612587735624561960176938209556777150821675191766038000323979374251056843399040592062232120016300528722394500972253821419509835189970824459173777432334325907781189983841838930891654818858052973456858049878700084422736207156836005189786243843224337778518091737648580070153561517768467108316485148591404;
            6'd41: xpb[52] = 1024'd52675037759489954875296116440880221521226736879643503147375764825581169073602350593015099742322155585763726999708614153102260570913459036264579058151488764049314988018762611704121880244794468757373278032440777141031150448282522658460407462562576994378264232639632325286783919100007692410966917041734717857756;
            6'd42: xpb[52] = 1024'd41855726906392174126030272704822233485676322937611814528713529327182963896147857786989607422412191155226925277022727333950699722317082882558333657129200095764304068256335239566404829597934118656693582608023504403362216473828838160084809735338910145532190686761172912924987768046453867053466725766984287124108;
            6'd43: xpb[52] = 1024'd31036416053294393376764428968764245450125908995580125910051293828784758718693364980964115102502226724690123554336840514799138873720706728852088256106911427479293148493907867428687778951073768556013887183606231665693282499375153661709212008115243296686117140882713500563191616992900041695966534492233856390460;
            6'd44: xpb[52] = 1024'd20217105200196612627498585232706257414575495053548437291389058330386553541238872174938622782592262294153321831650953695647578025124330575145842855084622759194282228731480495290970728304213418455334191759188958928024348524921469163333614280891576447840043595004254088201395465939346216338466343217483425656812;
            6'd45: xpb[52] = 1024'd9397794347098831878232741496648269379025081111516748672726822831988348363784379368913130462682297863616520108965066876496017176527954421439597454062334090909271308969053123153253677657353068354654496334771686190355414550467784664958016553667909598993970049125794675839599314885792390980966151942732994923164;
            6'd46: xpb[52] = 1024'd122645179178125792527765825165404714088173094295220744182196442398567038523639025472902709357430007742522867793736673491923520168772798602288512178056376463557951063776196968353166866202009923975284998518741653299050841426234996939547397396127472199414716406661452321507909691906167198640584650494608158673847;
            6'd47: xpb[52] = 1024'd111825868325028011778499981429346726052622680353189055563534206900168833346184532666877217037520043311986066071050786672771959320176422448582266777034087795272940144013769596215449815555149573874605303094324380561381907451781312441171799668903805350568642860782992909146113540852613373283084459219857727940199;
            6'd48: xpb[52] = 1024'd101006557471930231029234137693288738017072266411157366944871971401770628168730039860851724717610078881449264348364899853620398471580046294876021376011799126987929224251342224077732764908289223773925607669907107823712973477327627942796201941680138501722569314904533496784317389799059547925584267945107297206551;
            6'd49: xpb[52] = 1024'd90187246618832450279968293957230749981521852469125678326209735903372422991275547054826232397700114450912462625679013034468837622983670141169775974989510458702918304488914851940015714261428873673245912245489835086044039502873943444420604214456471652876495769026074084422521238745505722568084076670356866472903;
            6'd50: xpb[52] = 1024'd79367935765734669530702450221172761945971438527093989707547500404974217813821054248800740077790150020375660902993126215317276774387293987463530573967221790417907384726487479802298663614568523572566216821072562348375105528420258946045006487232804804030422223147614672060725087691951897210583885395606435739255;
            6'd51: xpb[52] = 1024'd68548624912636888781436606485114773910421024585062301088885264906576012636366561442775247757880185589838859180307239396165715925790917833757285172944933122132896464964060107664581612967708173471886521396655289610706171553966574447669408760009137955184348677269155259698928936638398071853083694120856005005607;
            6'd52: xpb[52] = 1024'd57729314059539108032170762749056785874870610643030612470223029408177807458912068636749755437970221159302057457621352577014155077194541680051039771922644453847885545201632735526864562320847823371206825972238016873037237579512889949293811032785471106338275131390695847337132785584844246495583502846105574271959;
            6'd53: xpb[52] = 1024'd46910003206441327282904919012998797839320196700998923851560793909779602281457575830724263118060256728765255734935465757862594228598165526344794370900355785562874625439205363389147511673987473270527130547820744135368303605059205450918213305561804257492201585512236434975336634531290421138083311571355143538311;
            6'd54: xpb[52] = 1024'd36090692353343546533639075276940809803769782758967235232898558411381397104003083024698770798150292298228454012249578938711033380001789372638548969878067117277863705676777991251430461027127123169847435123403471397699369630605520952542615578338137408646128039633777022613540483477736595780583120296604712804663;
            6'd55: xpb[52] = 1024'd25271381500245765784373231540882821768219368816935546614236322912983191926548590218673278478240327867691652289563692119559472531405413218932303568855778448992852785914350619113713410380266773069167739698986198660030435656151836454167017851114470559800054493755317610251744332424182770423082929021854282071015;
            6'd56: xpb[52] = 1024'd14452070647147985035107387804824833732668954874903857995574087414584986749094097412647786158330363437154850566877805300407911682809037065226058167833489780707841866151923246975996359733406422968488044274568925922361501681698151955791420123890803710953980947876858197889948181370628945065582737747103851337367;
            6'd57: xpb[52] = 1024'd3632759794050204285841544068766845697118540932872169376911851916186781571639604606622293838420399006618048844191918481256350834212660911519812766811201112422830946389495874838279309086546072867808348850151653184692567707244467457415822396667136862107907401998398785528152030317075119708082546472353420603719;
            6'd58: xpb[52] = 1024'd116880144625077164935374627737523290406266554116576164886381471482765471731494250710611872733168108885524396528963525096683853826457505092368727490805243485071510701196639720038192497631202928488438851034121620293387994583011679732005203239126699462528653759534056431196462407337449927367701045024228584354402;
            6'd59: xpb[52] = 1024'd106060833771979384186108784001465302370716140174544476267719235984367266554039757904586380413258144454987594806277638277532292977861128938662482089782954816786499781434212347900475446984342578387759155609704347555719060608557995233629605511903032613682580213655597018834666256283896102010200853749478153620754;
            6'd60: xpb[52] = 1024'd95241522918881603436842940265407314335165726232512787649057000485969061376585265098560888093348180024450793083591751458380732129264752784956236688760666148501488861671784975762758396337482228287079460185287074818050126634104310735254007784679365764836506667777137606472870105230342276652700662474727722887106;
            6'd61: xpb[52] = 1024'd84422212065783822687577096529349326299615312290481099030394764987570856199130772292535395773438215593913991360905864639229171280668376631249991287738377480216477941909357603625041345690621878186399764760869802080381192659650626236878410057455698915990433121898678194111073954176788451295200471199977292153458;
            6'd62: xpb[52] = 1024'd73602901212686041938311252793291338264064898348449410411732529489172651021676279486509903453528251163377189638219977820077610432072000477543745886716088811931467022146930231487324295043761528085720069336452529342712258685196941738502812330232032067144359576020218781749277803123234625937700279925226861419810;
            6'd63: xpb[52] = 1024'd62783590359588261189045409057233350228514484406417721793070293990774445844221786680484411133618286732840387915534091000926049583475624323837500485693800143646456102384502859349607244396901177985040373912035256605043324710743257240127214603008365218298286030141759369387481652069680800580200088650476430686162;
        endcase
    end

    always_comb begin
        case(flag[17][16:12])
            5'd0: xpb[53] = 1024'd0;
            5'd1: xpb[53] = 1024'd51964279506490480439779565321175362192964070464386033174408058492376240666767293874458918813708322302303586192848204181774488734879248170131255084671511475361445182622075487211890193750040827884360678487617983867374390736289572741751616875784698369452212484263299957025685501016126975222699897375725999952514;
            5'd2: xpb[53] = 1024'd103928559012980960879559130642350724385928140928772066348816116984752481333534587748917837627416644604607172385696408363548977469758496340262510169343022950722890365244150974423780387500081655768721356975235967734748781472579145483503233751569396738904424968526599914051371002032253950445399794751451999905028;
            5'd3: xpb[53] = 1024'd31826142835346699920539768558711653834193784267422415395092320412151826662992742713361685226467292597467609171087119110744402363796524175838605128998203385150644873296655244298040342058605277931771837854466711755758811358647821452289872057670865659089817549375782813046949974974452292650981002300552405373211;
            5'd4: xpb[53] = 1024'd83790422341837180360319333879887016027157854731808448569500378904528067329760036587820604040175614899771195363935323292518891098675772345969860213669714860512090055918730731509930535808646105816132516342084695623133202094937394194041488933455564028542030033639082770072635475990579267873680899676278405325725;
            5'd5: xpb[53] = 1024'd11688006164202919401299971796247945475423498070458797615776582331927412659218191552264451639226262892631632149326034039714315992713800181545955173324895294939844563971235001384190490367169727979182997221315439644143231981006070162828127239557032948727422614488265669068214448932777610079262107225378810793908;
            5'd6: xpb[53] = 1024'd63652285670693399841079537117423307668387568534844830790184640824303653325985485426723370452934585194935218342174238221488804727593048351677210257996406770301289746593310488596080684117210555863543675708933423511517622717295642904579744115341731318179635098751565626093899949948904585301962004601104810746422;
            5'd7: xpb[53] = 1024'd115616565177183880280859102438598669861351638999230863964592699316679893992752779301182289266642907497238804535022442403263293462472296521808465342667918245662734929215385975807970877867251383747904354196551407378892013453585215646331360991126429687631847583014865583119585450965031560524661901976830810698936;
            5'd8: xpb[53] = 1024'd43514148999549619321839740354959599309617282337881213010868902744079239322210934265626136865693555490099241320413153150458718356510324357384560302323098680090489437267890245682230832425775005910954835075782151399902043339653891615117999297227898607817240163864048482115164423907229902730243109525931216167119;
            5'd9: xpb[53] = 1024'd95478428506040099761619305676134961502581352802267246185276961236455479988978228140085055679401877792402827513261357332233207091389572527515815386994610155451934619889965732894121026175815833795315513563400135267276434075943464356869616173012596977269452648127348439140849924923356877952943006901657216119633;
            5'd10: xpb[53] = 1024'd23376012328405838802599943592495890950846996140917595231553164663854825318436383104528903278452525785263264298652068079428631985427600363091910346649790589879689127942470002768380980734339455958365994442630879288286463962012140325656254479114065897454845228976531338136428897865555220158524214450757621587816;
            5'd11: xpb[53] = 1024'd75340291834896319242379508913671253143811066605303628405961223156231065985203676978987822092160848087566850491500272261203120720306848533223165431321302065241134310564545489980271174484380283842726672930248863155660854698301713067407871354898764266907057713239831295162114398881682195381224111826483621540330;
            5'd12: xpb[53] = 1024'd3237875657262058283360146830032182592076709943953977452237426583630411314661831943431669691211496080427287276890983008398545614344876368799260390976482499668888818617049759854531129042903906005777153809479607176670884584370389036194509661000233187092450294089014194157693371823880537586805319375584027008513;
            5'd13: xpb[53] = 1024'd55202155163752538723139712151207544785040780408340010626645485076006651981429125817890588504919818382730873469739187190173034349224124538930515475647993975030334001239125247066421322792944733890137832297097591044045275320659961777946126536784931556544662778352314151183378872840007512809505216751310026961027;
            5'd14: xpb[53] = 1024'd107166434670243019162919277472382906978004850872726043801053543568382892648196419692349507318628140685034459662587391371947523084103372709061770560319505450391779183861200734278311516542985561774498510784715574911419666056949534519697743412569629925996875262615614108209064373856134488032205114127036026913541;
            5'd15: xpb[53] = 1024'd35064018492608758203899915388743836426270494211376392847329746995782237977654574656793354917678788677894896447978102119142947978141400544637865519974685884819533691913705004152571471101509183937548991663946318932429695943018210488484381718671098846182267843464797007204643346798332830237786321676136432381724;
            5'd16: xpb[53] = 1024'd87028297999099238643679480709919198619234564675762426021737805488158478644421868531252273731387110980198482640826306300917436713020648714769120604646197360180978874535780491364461664851550011821909670151564302799804086679307783230235998594455797215634480327728096964230328847814459805460486219051862432334238;
            5'd17: xpb[53] = 1024'd14925881821464977684660118626280128067500208014412775068014008915557823973880023495696121330437758973058919426217017048112861607058676550345215564301377794608733382588284761238721619410073633984960151030795046820814116565376459199022636900557266135819872908577279863225907820756658147666067426600962837802421;
            5'd18: xpb[53] = 1024'd66890161327955458124439683947455490260464278478798808242422067407934064640647317370155040144146081275362505619065221229887350341937924720476470648972889269970178565210360248450611813160114461869320829518413030688188507301666031940774253776341964505272085392840579820251593321772785122888767323976688837754935;
            5'd19: xpb[53] = 1024'd118854440834445938564219249268630852453428348943184841416830125900310305307414611244613958957854403577666091811913425411661839076817172890607725733644400745331623747832435735662502006910155289753681508006031014555562898037955604682525870652126662874724297877103879777277278822788912098111467221352414837707449;
            5'd20: xpb[53] = 1024'd46752024656811677605199887184991781901693992281835190463106329327709650636872766209057806556905051570526528597304136158857263970855200726183820693299581179759378255884940005536761961468678911916731988885261758576572927924024280651312508958228131794909690457953062676272857795731110440317048428901515243175632;
            5'd21: xpb[53] = 1024'd98716304163302158044979452506167144094658062746221223637514387820085891303640060083516725370613373872830114790152340340631752705734448896315075777971092655120823438507015492748652155218719739801092667372879742443947318660313853393064125834012830164361902942216362633298543296747237415539748326277241243128146;
            5'd22: xpb[53] = 1024'd26613887985667897085960090422528073542923706084871572683790591247485236633098215047960572969664021865690551575543051087827177599772476731891170737626273089548577946559519762622912109777243361964143148252110486464957348546382529361850764140114299084547295523065545532294122269689435757745329533826341648596329;
            5'd23: xpb[53] = 1024'd78578167492158377525739655743703435735887776549257605858198649739861477299865508922419491783372344167994137768391255269601666334651724902022425822297784564910023129181595249834802303527284189848503826739728470332331739282672102103602381015898997453999508007328845489319807770705562732968029431202067648548843;
            5'd24: xpb[53] = 1024'd6475751314524116566720293660064365184153419887907954904474853167260822629323663886863339382422992160854574553781966016797091228689752737598520781952964999337777637234099519709062258085807812011554307618959214353341769168740778072389019322000466374184900588178028388315386743647761075173610638751168054017026;
            5'd25: xpb[53] = 1024'd58440030821014597006499858981239727377117490352293988078882911659637063296090957761322258196131314463158160746630170198571579963569000907729775866624476474699222819856175006920952451835848639895914986106577198220716159905030350814140636197785164743637113072441328345341072244663888050396310536126894053969540;
            5'd26: xpb[53] = 1024'd110404310327505077446279424302415089570081560816680021253290970152013303962858251635781177009839636765461746939478374380346068698448249077861030951295987950060668002478250494132842645585889467780275664594195182088090550641319923555892253073569863113089325556704628302366757745680015025619010433502620053922054;
            5'd27: xpb[53] = 1024'd38301894149870816487260062218776019018347204155330370299567173579412649292316406600225024608890284758322183724869085127541493592486276913437125910951168384488422510530754764007102600144413089943326145473425926109100580527388599524678891379671332033274718137553811201362336718622213367824591641051720459390237;
            5'd28: xpb[53] = 1024'd90266173656361296927039627539951381211311274619716403473975232071788889959083700474683943422598607060625769917717289309315982327365525083568380995622679859849867693152830251218992793894453917827686823961043909976474971263678172266430508255456030402726930621817111158388022219638340343047291538427446459342751;
            5'd29: xpb[53] = 1024'd18163757478727035968020265456312310659576917958366752520251435499188235288541855439127791021649255053486206703108000056511407221403552919144475955277860294277622201205334521093252748452977539990737304840274653997485001149746848235217146561557499322912323202666294057383601192580538685252872745976546864810934;
            5'd30: xpb[53] = 1024'd70128036985217516407799830777487672852540988422752785694659493991564475955309149313586709835357577355789792895956204238285895956282801089275731039949371769639067383827410008305142942203018367875097983327892637864859391886036420976968763437342197692364535686929594014409286693596665660475572643352272864763448;
            5'd31: xpb[53] = 1024'd122092316491707996847579396098663035045505058887138818869067552483940716622076443188045628649065899658093379088804408420060384691162049259406986124620883245000512566449485495517033135953059195759458661815510621732233782622325993718720380313126896061816748171192893971434972194612792635698272540727998864715962;
        endcase
    end

    always_comb begin
        case(flag[18][5:0])
            6'd0: xpb[54] = 1024'd0;
            6'd1: xpb[54] = 1024'd87028297999099238643679480709919198619234564675762426021737805488158478644421868531252273731387110980198482640826306300917436713020648714769120604646197360180978874535780491364461664851550011821909670151564302799804086679307783230235998594455797215634480327728096964230328847814459805460486219051862432334238;
            6'd2: xpb[54] = 1024'd49989900314073735888560034015023964493770702225789167915343755911340061951534598152489476248116547650953815874195119167255809585200077094983081084276063679428267074501989765391293090511582817922509142694741365753243812508394669687507018619228364982002140752042076870430551167554990977903853748277099270184145;
            6'd3: xpb[54] = 1024'd12951502629048233133440587320128730368306839775815909808949706334521645258647327773726678764845984321709149107563932033594182457379505475197041563905929998675555274468199039418124516171615624023108615237918428706683538337481556144778038644000932748369801176356056776630773487295522150347221277502336108034052;
            6'd4: xpb[54] = 1024'd99979800628147471777120068030047928987541404451578335830687511822680123903069196304978952496233095301907631748390238334511619170400154189966162168552127358856534149003979530782586181023165635845018285389482731506487625016789339375014037238456729964004281504084153740861102335109981955807707496554198540368290;
            6'd5: xpb[54] = 1024'd62941402943121969022000621335152694862077542001605077724293462245861707210181925926216155012962531972662964981759051200849992042579582570180122648181993678103822348970188804809417606683198441945617757932659794459927350845876225832285057263229297730371941928398133647061324654850513128251075025779435378218197;
            6'd6: xpb[54] = 1024'd25903005258096466266881174640257460736613679551631819617899412669043290517294655547453357529691968643418298215127864067188364914759010950394083127811859997351110548936398078836249032343231248046217230475836857413367076674963112289556077288001865496739602352712113553261546974591044300694442555004672216068104;
            6'd7: xpb[54] = 1024'd112931303257195704910560655350176659355848244227394245639637218157201769161716524078705631261079079623616780855954170368105801627779659665163203732458057357532089423472178570200710697194781259868126900627401160213171163354270895519792075882457662712374082680440210517491875822405504106154928774056534648402342;
            6'd8: xpb[54] = 1024'd75892905572170202155441208655281425230384381777420987533243168580383352468829253699942833777808516294372114089322983234444174499959088045377164212087923676779377623438387844227542122854814065968726373170578223166610889183357781977063095907230230478741743104754190423692098142146035278598296303281771486252249;
            6'd9: xpb[54] = 1024'd38854507887144699400321761960386191104920519327447729426849119003564935775941983321180036294537952965127447322691796100782547372138516425591124691717789996026665823404597118254373548514846872069325845713755286120050615012444668434334115932002798245109403529068170329892320461886566451041663832507008324102156;
            6'd10: xpb[54] = 1024'd1816110202119196645202315265490956979456656877474471320455069426746519083054712942417238811267389635882780556060608967120920244317944805805085171347656315273954023370806392281204974174879678169925318256932349073490340841531554891605135956775366011477063953382150236092542781627097623485031361732245161952063;
            6'd11: xpb[54] = 1024'd88844408201218435288881795975410155598691221553236897342192874914904997727476581473669512542654500616081263196886915268038356957338593520574205775993853675454932897906586883645666639026429689991834988408496651873294427520839338121841134551231163227111544281110247200322871629441557428945517580784107594286301;
            6'd12: xpb[54] = 1024'd51806010516192932533762349280514921473227359103263639235798825338086581034589311094906715059383937286836596430255728134376729829518021900788166255623719994702221097872796157672498064686462496092434460951673714826734153349926224579112154576003730993479204705424227106523093949182088601388885110009344432136208;
            6'd13: xpb[54] = 1024'd14767612831167429778642902585619687347763496653290381129404775761268164341702040716143917576113373957591929663624541000715102701697450281002126735253586313949509297839005431699329490346495302193033933494850777780173879179013111036383174600776298759846865129738207012723316268922619773832252639234581269986115;
            6'd14: xpb[54] = 1024'd101795910830266668422322383295538885966998061329052807151142581249426642986123909247396191307500484937790412304450847301632539414718098995771247339899783674130488172374785923063791155198045314014943603646415080579977965858320894266619173195232095975481345457466303976953645116737079579292738858286443702320353;
            6'd15: xpb[54] = 1024'd64757513145241165667202936600643651841534198879079549044748531672608226293236638868633393824229921608545745537819660167970912286897527375985207819529649993377776372340995197090622580858078120115543076189592143533417691687407780723890193220004663741849005881780283883153867436477610751736106387511680540170260;
            6'd16: xpb[54] = 1024'd27719115460215662912083489905748417716070336429106290938354482095789809600349368489870596340959358279301078771188473034309285159076955756199168299159516312625064572307204471117454006518110926216142548732769206486857417516494667181161213244777231508216666306094263789354089756218141924179473916736917378020167;
            6'd17: xpb[54] = 1024'd114747413459314901555762970615667616335304901104868716960092287583948288244771237021122870072346469259499561412014779335226721872097604470968288903805713672806043446842984962481915671369660938038052218884333509286661504195802450411397211839233028723851146633822360753584418604032601729639960135788779810354405;
            6'd18: xpb[54] = 1024'd77709015774289398800643523920772382209841038654895458853698238007129871551883966642360072589075905930254894645383592201565094744277032851182249383435579992053331646809194236508747097029693744138651691427510572240101230024889336868668231864005596490218807058136340659784640923773132902083327665014016648204312;
            6'd19: xpb[54] = 1024'd40670618089263896045524077225877148084377176204922200747304188430311454858996696263597275105805342601010227878752405067903467616456461231396209863065446311300619846775403510535578522689726550239251163970687635193540955853976223325939251888778164256586467482450320565984863243513664074526695194239253486054219;
            6'd20: xpb[54] = 1024'd3632220404238393290404630530981913958913313754948942640910138853493038166109425884834477622534779271765561112121217934241840488635889611610170342695312630547908046741612784562409948349759356339850636513864698146980681683063109783210271913550732022954127906764300472185085563254195246970062723464490323904126;
            6'd21: xpb[54] = 1024'd90660518403337631934084111240901112578147878430711368662647944341651516810531294416086751353921890251964043752947524235159277201656538326379290947341509990728886921277393275926871613201309368161760306665429000946784768362370893013446270508006529238588608234492397436415414411068655052430548942516352756238364;
            6'd22: xpb[54] = 1024'd53622120718312129178964664546005878452684015980738110556253894764833100117644024037323953870651326922719376986316337101497650073835966706593251426971376309976175121243602549953703038861342174262359779208606063900224494191457779470717290532779097004956268658806377342615636730809186224873916471741589594088271;
            6'd23: xpb[54] = 1024'd16583723033286626423845217851110644327220153530764852449859845188014683424756753658561156387380763593474710219685149967836022946015395086807211906601242629223463321209811823980534464521374980362959251751783126853664220020544665927988310557551664771323929083120357248815859050549717397317284000966826431938178;
            6'd24: xpb[54] = 1024'd103612021032385865067524698561029842946454718206527278471597650676173162069178622189813430118767874573673192860511456268753459659036043801576332511247439989404442195745592315344996129372924992184868921903347429653468306699852449158224309152007461986958409410848454213046187898364177202777770220018688864272416;
            6'd25: xpb[54] = 1024'd66573623347360362312405251866134608820990855756554020365203601099354745376291351811050632635497311244428526093880269135091832531215472181790292990877306308651730395711801589371827555032957798285468394446524492606908032528939335615495329176780029753326069835162434119246410218104708375221137749243925702122323;
            6'd26: xpb[54] = 1024'd29535225662334859557285805171239374695526993306580762258809551522536328683404081432287835152226747915183859327249082001430205403394900562004253470507172627899018595678010863398658980692990604386067866989701555560347758358026222072766349201552597519693730259476414025446632537845239547664505278469162539972230;
            6'd27: xpb[54] = 1024'd116563523661434098200965285881158573314761557982343188280547357010694807327825949963540108883613858895382341968075388302347642116415549276773374075153369988079997470213791354763120645544540616207977537141265858360151845037334005303002347796008394735328210587204510989676961385659699353124991497521024972306468;
            6'd28: xpb[54] = 1024'd79525125976408595445845839186263339189297695532369930174153307433876390634938679584777311400343295566137675201444201168686014988594977656987334554783236307327285670180000628789952071204573422308577009684442921313591570866420891760273367820780962501695871011518490895877183705400230525568359026746261810156375;
            6'd29: xpb[54] = 1024'd42486728291383092690726392491368105063833833082396672067759257857057973942051409206014513917072732236893008434813014035024387860774406037201295034413102626574573870146209902816783496864606228409176482227619984267031296695507778217544387845553530268063531435832470802077406025140761698011726555971498648006282;
            6'd30: xpb[54] = 1024'd5448330606357589935606945796472870938369970632423413961365208280239557249164138827251716433802168907648341668181826901362760732953834417415255514042968945821862070112419176843614922524639034509775954770797047220471022524594664674815407870326098034431191860146450708277628344881292870455094085196735485856189;
            6'd31: xpb[54] = 1024'd92476628605456828579286426506392069557604535308185839983103013768398035893586007358503990165189279887846824309008133202280197445974483132184376118689166306002840944648199668208076587376189046331685624922361350020275109203902447905051406464781895250065672187874547672507957192695752675915580304248597918190427;
            6'd32: xpb[54] = 1024'd55438230920431325824166979811496835432140672858212581876708964191579619200698736979741192681918716558602157542376946068618570318153911512398336598319032625250129144614408942234908013036221852432285097465538412973714835032989334362322426489554463016433332612188527578708179512436283848358947833473834756040334;
            6'd33: xpb[54] = 1024'd18399833235405823069047533116601601306676810408239323770314914614761202507811466600978395198648153229357490775745758934956943190333339892612297077948898944497417344580618216261739438696254658532884570008715475927154560862076220819593446514327030782800993036502507484908401832176815020802315362699071593890241;
            6'd34: xpb[54] = 1024'd105428131234505061712727013826520799925911375084001749792052720102919681152233335132230668930035264209555973416572065235874379903353988607381417682595096304678396219116398707626201103547804670354794240160279778726958647541384004049829445108782827998435473364230604449138730679991274826262801581750934026224479;
            6'd35: xpb[54] = 1024'd68389733549479558957607567131625565800447512634028491685658670526101264459346064753467871446764700880311306649940878102212752775533416987595378162224962623925684419082607981653032529207837476455393712703456841680398373370470890507100465133555395764803133788544584355338952999731805998706169110976170864074386;
            6'd36: xpb[54] = 1024'd31351335864454056202488120436730331674983650184055233579264620949282847766458794374705073963494137551066639883309690968551125647712845367809338641854828943172972619048817255679863954867870282555993185246633904633838099199557776964371485158327963531170794212858564261539175319472337171149536640201407701924293;
            6'd37: xpb[54] = 1024'd118379633863553294846167601146649530294218214859817659601002426437441326410880662905957347694881248531265122524135997269468562360733494082578459246501026303353951493584597747044325619719420294377902855398198207433642185878865560194607483752783760746805274540586661225769504167286796976610022859253270134258531;
            6'd38: xpb[54] = 1024'd81341236178527792091048154451754296168754352409844401494608376860622909717993392527194550211610685202020455757504810135806935232912922462792419726130892622601239693550807021071157045379453100478502327941375270387081911707952446651878503777556328513172934964900641131969726487027328149053390388478506972108438;
            6'd39: xpb[54] = 1024'd44302838493502289335928707756859062043290489959871143388214327283804493025106122148431752728340121872775788990873623002145308105092350843006380205760758941848527893517016295097988471039485906579101800484552333340521637537039333109149523802328896279540595389214621038169948806767859321496757917703743809958345;
            6'd40: xpb[54] = 1024'd7264440808476786580809261061963827917826627509897885281820277706986076332218851769668955245069558543531122224242435868483680977271779223220340685390625261095816093483225569124819896699518712679701273027729396293961363366126219566420543827101464045908255813528600944370171126508390493940125446928980647808252;
            6'd41: xpb[54] = 1024'd94292738807576025224488741771883026537061192185660311303558083195144554976640720300921228976456669523729604865068742169401117690292427937989461290036822621276794968019006060489281561551068724501610943179293699093765450045434002796656542421557261261542736141256697908600499974322850299400611665980843080142490;
            6'd42: xpb[54] = 1024'd57254341122550522469369295076987792411597329735687053197164033618326138283753449922158431493186106194484938098437555035739490562471856318203421769666688940524083167985215334516112987211101530602210415722470762047205175874520889253927562446329829027910396565570677814800722294063381471843979195206079917992397;
            6'd43: xpb[54] = 1024'd20215943437525019714249848382092558286133467285713795090769984041507721590866179543395634009915542865240271331806367902077863434651284698417382249296555259771371367951424608542944412871134336702809888265647825000644901703607775711198582471102396794278056989884657721000944613803912644287346724431316755842304;
            6'd44: xpb[54] = 1024'd107244241436624258357929329092011756905368031961476221112507789529666200235288048074647907741302653845438753972632674202995300147671933413186502853942752619952350242487205099907406077722684348524719558417212127800448988382915558941434581065558194009912537317612754685231273461618372449747832943483179188176542;
            6'd45: xpb[54] = 1024'd70205843751598755602809882397116522779904169511502963006113739952847783542400777695885110258032090516194087206001487069333673019851361793400463333572618939199638442453414373934237503382717154625319030960389190753888714212002445398705601090330761776280197741926734591431495781358903622191200472708416026026449;
            6'd46: xpb[54] = 1024'd33167446066573252847690435702221288654440307061529704899719690376029366849513507317122312774761527186949420439370299935672045892030790173614423813202485258446926642419623647961068929042749960725918503503566253707328440041089331855976621115103329542647858166240714497631718101099434794634568001933652863876356;
            6'd47: xpb[54] = 1024'd120195744065672491491369916412140487273674871737292130921457495864187845493935375848374586506148638167147903080196606236589482605051438888383544417848682618627905516955404139325530593894299972547828173655130556507132526720397115086212619709559126758282338493968811461862046948913894600095054220985515296210594;
            6'd48: xpb[54] = 1024'd83157346380646988736250469717245253148211009287318872815063446287369428801048105469611789022878074837903236313565419102927855477230867268597504897478548937875193716921613413352362019554332778648427646198307619460572252549484001543483639734331694524649998918282791368062269268654425772538421750210752134060501;
            6'd49: xpb[54] = 1024'd46118948695621485981131023022350019022747146837345614708669396710551012108160835090848991539607511508658569546934231969266228349410295648811465377108415257122481916887822687379193445214365584749027118741484682414011978378570888000754659759104262291017659342596771274262491588394956944981789279435988971910408;
            6'd50: xpb[54] = 1024'd9080551010595983226011576327454784897283284387372356602275347133732595415273564712086194056336948179413902780303044835604601221589724029025425856738281576369770116854031961406024870874398390849626591284661745367451704207657774458025679783876830057385319766910751180462713908135488117425156808661225809760315;
            6'd51: xpb[54] = 1024'd96108849009695221869691057037373983516517849063134782624013152621891074059695433243338467787724059159612385421129351136522037934610372743794546461384478936550748991389812452770486535725948402671536261436226048167255790886965557688261678378332627273019800094638848144693042755949947922885643027713088242094553;
            6'd52: xpb[54] = 1024'd59070451324669719114571610342478749391053986613161524517619103045072657366808162864575670304453495830367718654498164002860410806789801124008506941014345255798037191356021726797317961385981208772135733979403111120695516716052444145532698403105195039387460518952828050893265075690479095329010556938325079944460;
            6'd53: xpb[54] = 1024'd22032053639644216359452163647583515265590124163188266411225053468254240673920892485812872821182932501123051887866976869198783678969229504222467420644211575045325391322231000824149387046014014872735206522580174074135242545139330602803718427877762805755120943266807957093487395431010267772378086163561917794367;
            6'd54: xpb[54] = 1024'd109060351638743455003131644357502713884824688838950692432962858956412719318342761017065146552570043481321534528693283170116220391989878218991588025290408935226304265858011492188611051897564026694644876674144476873939329224447113833039717022333560021389601270994904921323816243245470073232864305215424350128605;
            6'd55: xpb[54] = 1024'd72021953953717952248012197662607479759360826388977434326568809379594302625455490638302349069299480152076867762062096036454593264169306599205548504920275254473592465824220766215442477557596832795244349217321539827379055053534000290310737047106127787757261695308884827524038562986001245676231834440661187978512;
            6'd56: xpb[54] = 1024'd34983556268692449492892750967712245633896963939004176220174759802775885932568220259539551586028916822832200995430908902792966136348734979419508984550141573720880665790430040242273903217629638895843821760498602780818780882620886747581757071878695554124922119622864733724260882726532418119599363665898025828419;
            6'd57: xpb[54] = 1024'd122011854267791688136572231677631444253131528614766602241912565290934364576990088790791825317416027803030683636257215203710402849369383694188629589196338933901859540326210531606735568069179650717753491912062905580622867561928669977817755666334492769759402447350961697954589730540992223580085582717760458162657;
            6'd58: xpb[54] = 1024'd84973456582766185381452784982736210127667666164793344135518515714115947884102818412029027834145464473786016869626028070048775721548812074402590068826205253149147740292419805633566993729212456818352964455239968534062593391015556435088775691107060536127062871664941604154812050281523396023453111942997296012564;
            6'd59: xpb[54] = 1024'd47935058897740682626333338287840976002203803714820086029124466137297531191215548033266230350874901144541350102994840936387148593728240454616550548456071572396435940258629079660398419389245262918952436998417031487502319220102442892359795715879628302494723295978921510355034370022054568466820641168234133862471;
            6'd60: xpb[54] = 1024'd10896661212715179871213891592945741876739941264846827922730416560479114498328277654503432867604337815296683336363653802725521465907668834830511028085937891643724140224838353687229845049278069019551909541594094440942045049189329349630815740652196068862383720292901416555256689762585740910188170393470971712378;
            6'd61: xpb[54] = 1024'd97924959211814418514893372302864940495974505940609253944468222048637593142750146185755706598991448795495165977189960103642958178928317549599631632732135251824703014760618845051691509900828080841461579693158397240746131728497112579866814335107993284496864048020998380785585537577045546370674389445333404046616;
            6'd62: xpb[54] = 1024'd60886561526788915759773925607969706370510643490635995838074172471819176449862875806992909115720885466250499210558772969981331051107745929813592112362001571071991214726828119078522935560860886942061052236335460194185857557583999037137834359880561050864524472334978286985807857317576718814041918670570241896523;
            6'd63: xpb[54] = 1024'd23848163841763413004654478913074472245046781040662737731680122895000759756975605428230111632450322137005832443927585836319703923287174310027552591991867890319279414693037393105354361220893693042660524779512523147625583386670885494408854384653128817232184896648958193186030177058107891257409447895807079746430;
        endcase
    end

    always_comb begin
        case(flag[18][11:6])
            6'd0: xpb[55] = 1024'd0;
            6'd1: xpb[55] = 1024'd110876461840862651648333959622993670864281345716425163753417928383159238401397473959482385363837433117204315084753892137237140636307823024796673196638065250500258289228817884469816026072443704864570194931076825947429670065978668724644852979108926032866665224377055157416359024872567696717895666947669512080668;
            6'd2: xpb[55] = 1024'd97686227997600561897868991841172908983864264307114643378704001701341581465485809008949699513017191924965480762050290839895217431774425715038186268259799460066825903888064551602001812953370204007830192253766412048494979281736440676324727388534622616466510545339993256802611521671206760418672644068713429677005;
            6'd3: xpb[55] = 1024'd84495994154338472147404024059352147103447182897804123003990075019523924529574144058417013662196950732726646439346689542553294227241028405279699339881533669633393518547311218734187599834296703151090189576455998149560288497494212628004601797960319200066355866302931356188864018469845824119449621189757347273342;
            6'd4: xpb[55] = 1024'd71305760311076382396939056277531385223030101488493602629276148337706267593662479107884327811376709540487812116643088245211371022707631095521212411503267879199961133206557885866373386715223202294350186899145584250625597713251984579684476207386015783666201187265869455575116515268484887820226598310801264869679;
            6'd5: xpb[55] = 1024'd58115526467814292646474088495710623342613020079183082254562221655888610657750814157351641960556468348248977793939486947869447818174233785762725483125002088766528747865804552998559173596149701437610184221835170351690906929009756531364350616811712367266046508228807554961369012067123951521003575431845182466016;
            6'd6: xpb[55] = 1024'd44925292624552202896009120713889861462195938669872561879848294974070953721839149206818956109736227156010143471235885650527524613640836476004238554746736298333096362525051220130744960477076200580870181544524756452756216144767528483044225026237408950865891829191745654347621508865763015221780552552889100062353;
            6'd7: xpb[55] = 1024'd31735058781290113145544152932069099581778857260562041505134368292253296785927484256286270258915985963771309148532284353185601409107439166245751626368470507899663977184297887262930747358002699724130178867214342553821525360525300434724099435663105534465737150154683753733874005664402078922557529673933017658690;
            6'd8: xpb[55] = 1024'd18544824938028023395079185150248337701361775851251521130420441610435639850015819305753584408095744771532474825828683055843678204574041856487264697990204717466231591843544554395116534238929198867390176189903928654886834576283072386403973845088802118065582471117621853120126502463041142623334506794976935255027;
            6'd9: xpb[55] = 1024'd5354591094765933644614217368427575820944694441941000755706514928617982914104154355220898557275503579293640503125081758501755000040644546728777769611938927032799206502791221527302321119855698010650173512593514755952143792040844338083848254514498701665427792080559952506378999261680206324111483916020852851364;
            6'd10: xpb[55] = 1024'd116231052935628585292948176991421246685226040158366164509124443311777221315501628314703283921112936696497955587878973895738895636348467571525450966250004177533057495731609105997118347192299402875220368443670340703381813858019513062728701233623424734532093016457615109922738024134247903042007150863690364932032;
            6'd11: xpb[55] = 1024'd103040819092366495542483209209600484804808958749055644134410516629959564379589963364170598070292695504259121265175372598396972431815070261766964037871738387099625110390855773129304134073225902018480365766359926804447123073777285014408575643049121318131938337420553209308990520932886966742784127984734282528369;
            6'd12: xpb[55] = 1024'd89850585249104405792018241427779722924391877339745123759696589948141907443678298413637912219472454312020286942471771301055049227281672952008477109493472596666192725050102440261489920954152401161740363089049512905512432289535056966088450052474817901731783658383491308695243017731526030443561105105778200124706;
            6'd13: xpb[55] = 1024'd76660351405842316041553273645958961043974795930434603384982663266324250507766633463105226368652213119781452619768170003713126022748275642249990181115206806232760339709349107393675707835078900305000360411739099006577741505292828917768324461900514485331628979346429408081495514530165094144338082226822117721043;
            6'd14: xpb[55] = 1024'd63470117562580226291088305864138199163557714521124083010268736584506593571854968512572540517831971927542618297064568706371202818214878332491503252736941015799327954368595774525861494716005399448260357734428685107643050721050600869448198871326211068931474300309367507467748011328804157845115059347866035317380;
            6'd15: xpb[55] = 1024'd50279883719318136540623338082317437283140633111813562635554809902688936635943303562039854667011730735303783974360967409029279613681481022733016324358675225365895569027842441658047281596931898591520355057118271208708359936808372821128073280751907652531319621272305606854000508127443221545892036468909952913717;
            6'd16: xpb[55] = 1024'd37089649876056046790158370300496675402723551702503042260840883220871279700031638611507168816191489543064949651657366111687356409148083712974529395980409434932463183687089108790233068477858397734780352379807857309773669152566144772807947690177604236131164942235243706240253004926082285246669013589953870510054;
            6'd17: xpb[55] = 1024'd23899416032793957039693402518675913522306470293192521886126956539053622764119973660974482965371248350826115328953764814345433204614686403216042467602143644499030798346335775922418855358784896878040349702497443410838978368323916724487822099603300819731010263198181805626505501724721348947445990710997788106391;
            6'd18: xpb[55] = 1024'd10709182189531867289228434736855151641889388883882001511413029857235965828208308710441797114551007158587281006250163517003510000081289093457555539223877854065598413005582443054604642239711396021300347025187029511904287584081688676167696509028997403330855584161119905012757998523360412648222967832041705702728;
            6'd19: xpb[55] = 1024'd121585644030394518937562394359848822506170734600307165264830958240395204229605782669924182478388440275791596091004055654240650636389112118254228735861943104565856702234400327524420668312155100885870541956263855459333957650060357400812549488137923436197520808538175062429117023395928109366118634779711217783396;
            6'd20: xpb[55] = 1024'd108395410187132429187097426578028060625753653190996644890117031558577547293694117719391496627568199083552761768300454356898727431855714808495741807483677314132424316893646994656606455193081600029130539278953441560399266865818129352492423897563620019797366129501113161815369520194567173066895611900755135379733;
            6'd21: xpb[55] = 1024'd95205176343870339436632458796207298745336571781686124515403104876759890357782452768858810776747957891313927445596853059556804227322317498737254879105411523698991931552893661788792242074008099172390536601643027661464576081575901304172298306989316603397211450464051261201622016993206236767672589021799052976070;
            6'd22: xpb[55] = 1024'd82014942500608249686167491014386536864919490372375604140689178194942233421870787818326124925927716699075093122893251762214881022788920188978767950727145733265559546212140328920978028954934598315650533924332613762529885297333673255852172716415013186997056771426989360587874513791845300468449566142842970572407;
            6'd23: xpb[55] = 1024'd68824708657346159935702523232565774984502408963065083765975251513124576485959122867793439075107475506836258800189650464872957818255522879220281022348879942832127160871386996053163815835861097458910531247022199863595194513091445207532047125840709770596902092389927459974127010590484364169226543263886888168744;
            6'd24: xpb[55] = 1024'd55634474814084070185237555450745013104085327553754563391261324831306919550047457917260753224287234314597424477486049167531034613722125569461794093970614152398694775530633663185349602716787596602170528569711785964660503728849217159211921535266406354196747413352865559360379507389123427870003520384930805765081;
            6'd25: xpb[55] = 1024'd42444240970821980434772587668924251223668246144444043016547398149489262614135792966728067373466993122358590154782447870189111409188728259703307165592348361965262390189880330317535389597714095745430525892401372065725812944606989110891795944692102937796592734315803658746632004187762491570780497505974723361418;
            6'd26: xpb[55] = 1024'd29254007127559890684307619887103489343251164735133522641833471467671605678224128016195381522646751930119755832078846572847188204655330949944820237214082571531830004849126997449721176478640594888690523215090958166791122160364761062571670354117799521396438055278741758132884500986401555271557474627018640957755;
            6'd27: xpb[55] = 1024'd16063773284297800933842652105282727462834083325823002267119544785853948742312463065662695671826510737880921509375245275505265000121933640186333308835816781098397619508373664581906963359567094031950520537780544267856431376122533014251544763543496104996283376241679857519136997785040618972334451748062558554092;
            6'd28: xpb[55] = 1024'd2873539441035711183377684323461965582417001916512481892405618104036291806400798115130009821006269545642087186671643978163341795588536330427846380457550990664965234167620331714092750240493593175210517860470130368921740591880304965931419172969192688596128697204617956905389494583679682673111428869106476150429;
            6'd29: xpb[55] = 1024'd113750001281898362831711643946455636446698347632937645645823546487195530207798272074612395184843702662846402271425536115400482431896359355224519577095616241165223523396438216183908776312937298039780712791546956316351410657858973690576272152078118721462793921581673114321748519456247379391007095816775988231097;
            6'd30: xpb[55] = 1024'd100559767438636273081246676164634874566281266223627125271109619805377873271886607124079709334023461470607567948721934818058559227362962045466032648717350450731791138055684883316094563193863797183040710114236542417416719873616745642256146561503815305062639242544611213708001016254886443091784072937819905827434;
            6'd31: xpb[55] = 1024'd87369533595374183330781708382814112685864184814316604896395693123560216335974942173547023483203220278368733626018333520716636022829564735707545720339084660298358752714931550448280350074790296326300707436926128518482029089374517593936020970929511888662484563507549313094253513053525506792561050058863823423771;
            6'd32: xpb[55] = 1024'd74179299752112093580316740600993350805447103405006084521681766441742559400063277223014337632382979086129899303314732223374712818296167425949058791960818869864926367374178217580466136955716795469560704759615714619547338305132289545615895380355208472262329884470487412480506009852164570493338027179907741020108;
            6'd33: xpb[55] = 1024'd60989065908850003829851772819172588925030021995695564146967839759924902464151612272481651781562737893891064980611130926032789613762770116190571863582553079431493982033424884712651923836643294612820702082305300720612647520890061497295769789780905055862175205433425511866758506650803634194115004300951658616445;
            6'd34: xpb[55] = 1024'd47798832065587914079386805037351827044612940586385043772253913078107245528239947321948965930742496701652230657907529628690866409229372806432084935204287288998061596692671551844837710717569793756080699404994886821677956736647833448975644199206601639462020526396363611253011003449442697894891981421995576212782;
            6'd35: xpb[55] = 1024'd34608598222325824328921837255531065164195859177074523397539986396289588592328282371416280079922255509413396335203928331348943204695975496673598006826021498564629211351918218977023497598496292899340696727684472922743265952405605400655518608632298223061865847359301710639263500248081761595668958543039493809119;
            6'd36: xpb[55] = 1024'd21418364379063734578456869473710303283778777767764003022826059714471931656416617420883594229102014317174562012500327034007020000162578186915111078447755708131196826011164886109209284479422792042600694050374059023808575168163377352335393018057994806661711168322239810025515997046720825296445935664083411405456;
            6'd37: xpb[55] = 1024'd8228130535801644827991901691889541403361696358453482648112133032654274720504952470350908378281773124935727689796725736665096795629180877156624150069489917697764440670411553241395071360349291185860691373063645124873884383921149304015267427483691390261556489285177909411768493845359888997222912785127329001793;
            6'd38: xpb[55] = 1024'd119104592376664296476325861314883212267643042074878646401530061415813513121902426429833293742119206242140042774550617873902237431937003901953297346707555168198022729899229437711211097432792996050430886304140471072303554449899818028660120406592617423128221713662233066828127518717927585715118579732796841082461;
            6'd39: xpb[55] = 1024'd105914358533402206725860893533062450387225960665568126026816134733995856185990761479300607891298965049901208451847016576560314227403606592194810418329289377764590344558476104843396884313719495193690883626830057173368863665657589980339994816018314006728067034625171166214380015516566649415895556853840758678798;
            6'd40: xpb[55] = 1024'd92724124690140116975395925751241688506808879256257605652102208052178199250079096528767922040478723857662374129143415279218391022870209282436323489951023587331157959217722771975582671194645994336950880949519643274434172881415361932019869225444010590327912355588109265600632512315205713116672533974884676275135;
            6'd41: xpb[55] = 1024'd79533890846878027224930957969420926626391797846947085277388281370360542314167431578235236189658482665423539806439813981876467818336811972677836561572757796897725573876969439107768458075572493480210878272209229375499482097173133883699743634869707173927757676551047364986885009113844776817449511095928593871472;
            6'd42: xpb[55] = 1024'd66343657003615937474465990187600164745974716437636564902674354688542885378255766627702550338838241473184705483736212684534544613803414662919349633194492006464293188536216106239954244956498992623470875594898815476564791312930905835379618044295403757527602997513985464373137505912483840518226488216972511467809;
            6'd43: xpb[55] = 1024'd53153423160353847724001022405779402865557635028326044527960428006725228442344101677169864488018000280945871161032611387192621409270017353160862704816226216030860803195462773372140031837425491766730872917588401577630100528688677787059492453721100341127448318476923563759390002711122904219003465338016429064146;
            6'd44: xpb[55] = 1024'd39963189317091757973536054623958640985140553619015524153246501324907571506432436726637178637197759088707036838329010089850698204736620043402375776437960425597428417854709440504325818718351990909990870240277987678695409744446449738739366863146796924727293639439861663145642499509761967919780442459060346660483;
            6'd45: xpb[55] = 1024'd26772955473829668223071086842137879104723472209705003778532574643089914570520771776104492786377517896468202515625408792508775000203222733643888848059694635163996032513956107636511605599278490053250867562967573779760718960204221690419241272572493508327138960402799762531894996308401031620557419580104264256820;
            6'd46: xpb[55] = 1024'd13582721630567578472606119060317117224306390800394483403818647961272257634609106825571806935557276704229368192921807495166851795669825423885401919681428844730563647173202774768697392480204989196510864885657159880826028175961993642099115681998190091926984281365737861918147493107040095321334396701148181853157;
            6'd47: xpb[55] = 1024'd392487787305488722141151278496355343889309391083963029104721279454600698697441875039121084737035511990533870218206197824928591136428114126914991303163054297131261832449441900883179361131488339770862208346745981891337391719765593778990091423886675526829602328675961304399989905679159022111373822192099449494;
            6'd48: xpb[55] = 1024'd111268949628168140370475110901490026208170655107509126782522649662613839100094915834521506448574468629194848954972098335062069227444251138923588187941228304797389551061267326370699205433575193204341057139423571929321007457698434318423843070532812708393494826705731118720759014778246855740007040769861611530162;
            6'd49: xpb[55] = 1024'd98078715784906050620010143119669264327753573698198606407808722980796182164183250883988820597754227436956014632268497037720146022910853829165101259562962514363957165720513993502884992314501692347601054462113158030386316673456206270103717479958509291993340147668669218107011511576885919440784017890905529126499;
            6'd50: xpb[55] = 1024'd84888481941643960869545175337848502447336492288888086033094796298978525228271585933456134746933986244717180309564895740378222818377456519406614331184696723930524780379760660635070779195428191490861051784802744131451625889213978221783591889384205875593185468631607317493264008375524983141560995011949446722836;
            6'd51: xpb[55] = 1024'd71698248098381871119080207556027740566919410879577565658380869617160868292359920982923448896113745052478345986861294443036299613844059209648127402806430933497092395039007327767256566076354690634121049107492330232516935104971750173463466298809902459193030789594545416879516505174164046842337972132993364319173;
            6'd52: xpb[55] = 1024'd58508014255119781368615239774206978686502329470267045283666942935343211356448256032390763045293503860239511664157693145694376409310661899889640474428165143063660009698253994899442352957281189777381046430181916333582244320729522125143340708235599042792876110557483516265769001972803110543114949254037281915510;
            6'd53: xpb[55] = 1024'd45317780411857691618150271992386216806085248060956524908953016253525554420536591081858077194473262668000677341454091848352453204777264590131153546049899352630227624357500662031628139838207688920641043752871502434647553536487294076823215117661295626392721431520421615652021498771442174243891926375081199511847;
            6'd54: xpb[55] = 1024'd32127546568595601867685304210565454925668166651646004534239089571707897484624926131325391343653021475761843018750490551010530000243867280372666617671633562196795239016747329163813926719134188063901041075561088535712862752245066028503089527086992209992566752483359715038273995570081237944668903496125117108184;
            6'd55: xpb[55] = 1024'd18937312725333512117220336428744693045251085242335484159525162889890240548713261180792705492832780283523008696046889253668606795710469970614179689293367771763362853675993996295999713600060687207161038398250674636778171968002837980182963936512688793592412073446297814424526492368720301645445880617169034704521;
            6'd56: xpb[55] = 1024'd5747078882071422366755368646923931164834003833024963784811236208072583612801596230260019642012539091284174373343287956326683591177072660855692760915101981329930468335240663428185500480987186350421035720940260737843481183760609931862838345938385377192257394409235913810778989167359365346222857738212952300858;
            6'd57: xpb[55] = 1024'd116623540722934074015089328269917602029115349549450127538229164591231822014199070189742405005849972208488489458097180093563824227484895685652365957553167231830188757564058547898001526553430891214991230652017086685273151249739278656507691325047311410058922618786291071227138014039927062064118524685882464381526;
            6'd58: xpb[55] = 1024'd103433306879671984264624360488096840148698268140139607163515237909414165078287405239209719155029731016249655135393578796221901022951498375893879029174901441396756372223305215030187313434357390358251227974706672786338460465497050608187565734473007993658767939749229170613390510838566125764895501806926381977863;
            6'd59: xpb[55] = 1024'd90243073036409894514159392706276078268281186730829086788801311227596508142375740288677033304209489824010820812689977498879977818418101066135392100796635650963323986882551882162373100315283889501511225297396258887403769681254822559867440143898704577258613260712167269999643007637205189465672478927970299574200;
            6'd60: xpb[55] = 1024'd77052839193147804763694424924455316387864105321518566414087384545778851206464075338144347453389248631771986489986376201538054613884703756376905172418369860529891601541798549294558887196210388644771222620085844988469078897012594511547314553324401160858458581675105369385895504435844253166449456049014217170537;
            6'd61: xpb[55] = 1024'd63862605349885715013229457142634554507447023912208046039373457863961194270552410387611661602569007439533152167282774904196131409351306446618418244040104070096459216201045216426744674077136887788031219942775431089534388112770366463227188962750097744458303902638043468772148001234483316867226433170058134766874;
            6'd62: xpb[55] = 1024'd50672371506623625262764489360813792627029942502897525664659531182143537334640745437078975751748766247294317844579173606854208204817909136859931315661838279663026830860291883558930460958063386931291217265465017190599697328528138414907063372175794328058149223600981568158400498033122380568003410291102052363211;
            6'd63: xpb[55] = 1024'd37482137663361535512299521578993030746612861093587005289945604500325880398729080486546289900928525055055483521875572309512285000284511827101444387283572489229594445519538550691116247838989886074551214588154603291665006544285910366586937781601490911657994544563919667544652994831761444268780387412145969959548;
        endcase
    end

    always_comb begin
        case(flag[18][16:12])
            5'd0: xpb[56] = 1024'd0;
            5'd1: xpb[56] = 1024'd24291903820099445761834553797172268866195779684276484915231677818508223462817415536013604050108283862816649199171971012170361795751114517342957458905306698796162060178785217823302034719916385217811211910844189392730315760043682318266812191027187495257839865526857766930905491630400507969557364533189887555885;
            5'd2: xpb[56] = 1024'd48583807640198891523669107594344537732391559368552969830463355637016446925634831072027208100216567725633298398343942024340723591502229034685914917810613397592324120357570435646604069439832770435622423821688378785460631520087364636533624382054374990515679731053715533861810983260801015939114729066379775111770;
            5'd3: xpb[56] = 1024'd72875711460298337285503661391516806598587339052829454745695033455524670388452246608040812150324851588449947597515913036511085387253343552028872376715920096388486180536355653469906104159749155653433635732532568178190947280131046954800436573081562485773519596580573300792716474891201523908672093599569662667655;
            5'd4: xpb[56] = 1024'd97167615280397783047338215188689075464783118737105939660926711274032893851269662144054416200433135451266596796687884048681447183004458069371829835621226795184648240715140871293208138879665540871244847643376757570921263040174729273067248764108749981031359462107431067723621966521602031878229458132759550223540;
            5'd5: xpb[56] = 1024'd121459519100497228809172768985861344330978898421382424576158389092541117314087077680068020250541419314083245995859855060851808978755572586714787294526533493980810300893926089116510173599581926089056059554220946963651578800218411591334060955135937476289199327634288834654527458152002539847786822665949437779425;
            5'd6: xpb[56] = 1024'd21684727236471933172208395378219180452476250979923225363258211846072445439595354306066553085992028867456745787574332638443106933665466769502584628415509151843281686503140089602181969127981105585557073856677896510017533710041197136635894576479895522280219289747029543555326421708474414800225497372513730850979;
            5'd7: xpb[56] = 1024'd45976631056571378934042949175391449318672030664199710278489889664580668902412769842080157136100312730273394986746303650613468729416581286845542087320815850639443746681925307425484003847897490803368285767522085902747849470084879454902706767507083017538059155273887310486231913338874922769782861905703618406864;
            5'd8: xpb[56] = 1024'd70268534876670824695877502972563718184867810348476195193721567483088892365230185378093761186208596593090044185918274662783830525167695804188499546226122549435605806860710525248786038567813876021179497678366275295478165230128561773169518958534270512795899020800745077417137404969275430739340226438893505962749;
            5'd9: xpb[56] = 1024'd94560438696770270457712056769735987051063590032752680108953245301597115828047600914107365236316880455906693385090245674954192320918810321531457005131429248231767867039495743072088073287730261238990709589210464688208480990172244091436331149561458008053738886327602844348042896599675938708897590972083393518634;
            5'd10: xpb[56] = 1024'd118852342516869716219546610566908255917259369717029165024184923120105339290865016450120969286425164318723342584262216687124554116669924838874414464036735947027929927218280960895390108007646646456801921500054654080938796750215926409703143340588645503311578751854460611278948388230076446678454955505273281074519;
            5'd11: xpb[56] = 1024'd19077550652844420582582236959266092038756722275569965811284745873636667416373293076119502121875773872096842375976694264715852071579819021662211797925711604890401312827494961381061903536045825953302935802511603627304751660038711955004976961932603549302598713967201320179747351786548321630893630211837574146073;
            5'd12: xpb[56] = 1024'd43369454472943866344416790756438360904952501959846450726516423692144890879190708612133106171984057734913491575148665276886213867330933539005169256831018303686563373006280179204363938255962211171114147713355793020035067420082394273271789152959791044560438579494059087110652843416948829600450994745027461701958;
            5'd13: xpb[56] = 1024'd67661358293043312106251344553610629771148281644122935641748101510653114342008124148146710222092341597730140774320636289056575663082048056348126715736325002482725433185065397027665972975878596388925359624199982412765383180126076591538601343986978539818278445020916854041558335047349337570008359278217349257843;
            5'd14: xpb[56] = 1024'd91953262113142757868085898350782898637344061328399420556979779329161337804825539684160314272200625460546789973492607301226937458833162573691084174641631701278887493363850614850968007695794981606736571535044171805495698940169758909805413535014166035076118310547774620972463826677749845539565723811407236813728;
            5'd15: xpb[56] = 1024'd116245165933242203629920452147955167503539841012675905472211457147669561267642955220173918322308909323363439172664578313397299254584277091034041633546938400075049553542635832674270042415711366824547783445888361198226014700213441228072225726041353530333958176074632387903369318308150353509123088344597124369613;
            5'd16: xpb[56] = 1024'd16470374069216907992956078540313003625037193571216706259311279901200889393151231846172451157759518876736938964379055890988597209494171273821838967435914057937520939151849833159941837944110546321048797748345310744591969610036226773374059347385311576324978138187373096804168281864622228461561763051161417441167;
            5'd17: xpb[56] = 1024'd40762277889316353754790632337485272491232973255493191174542957719709112855968647382186055207867802739553588163551026903158959005245285791164796426341220756733682999330635050983243872664026931538860009659189500137322285370079909091640871538412499071582818003714230863735073773495022736431119127584351304997052;
            5'd18: xpb[56] = 1024'd65054181709415799516625186134657541357428752939769676089774635538217336318786062918199659257976086602370237362722997915329320800996400308507753885246527455529845059509420268806545907383943316756671221570033689530052601130123591409907683729439686566840657869241088630665979265125423244400676492117541192552937;
            5'd19: xpb[56] = 1024'd89346085529515245278459739931829810223624532624046161005006313356725559781603478454213263308084370465186886561894968927499682596747514825850711344151834154326007119688205486629847942103859701974482433480877878922782916890167273728174495920466874062098497734767946397596884756755823752370233856650731080108822;
            5'd20: xpb[56] = 1024'd113637989349614691040294293729002079089820312308322645920237991175233783244420893990226867358192654328003535761066939939670044392498629343193668803057140853122169179866990704453149976823776087192293645391722068315513232650210956046441308111494061557356337600294804164527790248386224260339791221183920967664707;
            5'd21: xpb[56] = 1024'd13863197485589395403329920121359915211317664866863446707337813928765111369929170616225400193643263881377035552781417517261342347408523525981466136946116510984640565476204704938821772352175266688794659694179017861879187560033741591743141732838019603347357562407544873428589211942696135292229895890485260736261;
            5'd22: xpb[56] = 1024'd38155101305688841165164473918532184077513444551139931622569491747273334832746586152239004243751547744193684751953388529431704143159638043324423595851423209780802625654989922762123807072091651906605871605023207254609503320077423910009953923865207098605197427934402640359494703573096643261787260423675148292146;
            5'd23: xpb[56] = 1024'd62447005125788286926999027715704452943709224235416416537801169565781558295564001688252608293859831607010333951125359541602065938910752560667381054756729908576964685833775140585425841792008037124417083515867396647339819080121106228276766114892394593863037293461260407290400195203497151231344624956865035848031;
            5'd24: xpb[56] = 1024'd86738908945887732688833581512876721809905003919692901453032847384289781758381417224266212343968115469826983150297330553772427734661867078010338513662036607373126746012560358408727876511924422342228295426711586040070134840164788546543578305919582089120877158988118174221305686833897659200901989490054923403916;
            5'd25: xpb[56] = 1024'd111030812765987178450668135310048990676100783603969386368264525202798005221198832760279816394076399332643632349469301565942789530412981595353295972567343306169288806191345576232029911231840807560039507337555775432800450600208470864810390496946769584378717024514975941152211178464298167170459354023244810959801;
            5'd26: xpb[56] = 1024'd11256020901961882813703761702406826797598136162510187155364347956329333346707109386278349229527008886017132141183779143534087485322875778141093306456318964031760191800559576717701706760239987056540521640012724979166405510031256410112224118290727630369736986627716650053010142020770042122898028729809104031355;
            5'd27: xpb[56] = 1024'd35547924722061328575538315499579095663793915846786672070596025774837556809524524922291953279635292748833781340355750155704449281073990295484050765361625662827922251979344794541003741480156372274351733550856914371896721270074938728379036309317915125627576852154574416983915633651170550092455393262998991587240;
            5'd28: xpb[56] = 1024'd59839828542160774337372869296751364529989695531063156985827703593345780272341940458305557329743576611650430539527721167874811076825104812827008224266932361624084312158130012364305776200072757492162945461701103764627037030118621046645848500345102620885416717681432183914821125281571058062012757796188879143125;
            5'd29: xpb[56] = 1024'd84131732362260220099207423093923633396185475215339641901059381411854003735159355994319161379851860474467079738699692180045172872576219330169965683172239060420246372336915230187607810919989142709974157372545293157357352790162303364912660691372290116143256583208289950845726616911971566031570122329378766699010;
            5'd30: xpb[56] = 1024'd108423636182359665861041976891095902262381254899616126816291059230362227197976771530332765429960144337283728937871663192215534668327333847512923142077545759216408432515700448010909845639905527927785369283389482550087668550205985683179472882399477611401096448735147717776632108542372074001127486862568654254895;
            5'd31: xpb[56] = 1024'd8648844318334370224077603283453738383878607458156927603390881983893555323485048156331298265410753890657228729586140769806832623237228030300720475966521417078879818124914448496581641168304707424286383585846432096453623460028771228481306503743435657392116410847888426677431072098843948953566161569132947326449;
        endcase
    end

    always_comb begin
        case(flag[19][5:0])
            6'd0: xpb[57] = 1024'd0;
            6'd1: xpb[57] = 1024'd16470374069216907992956078540313003625037193571216706259311279901200889393151231846172451157759518876736938964379055890988597209494171273821838967435914057937520939151849833159941837944110546321048797748345310744591969610036226773374059347385311576324978138187373096804168281864622228461561763051161417441167;
            6'd2: xpb[57] = 1024'd32940748138433815985912157080626007250074387142433412518622559802401778786302463692344902315519037753473877928758111781977194418988342547643677934871828115875041878303699666319883675888221092642097595496690621489183939220072453546748118694770623152649956276374746193608336563729244456923123526102322834882334;
            6'd3: xpb[57] = 1024'd49411122207650723978868235620939010875111580713650118777933839703602668179453695538517353473278556630210816893137167672965791628482513821465516902307742173812562817455549499479825513832331638963146393245035932233775908830108680320122178042155934728974934414562119290412504845593866685384685289153484252323501;
            6'd4: xpb[57] = 1024'd65881496276867631971824314161252014500148774284866825037245119604803557572604927384689804631038075506947755857516223563954388837976685095287355869743656231750083756607399332639767351776442185284195190993381242978367878440144907093496237389541246305299912552749492387216673127458488913846247052204645669764668;
            6'd5: xpb[57] = 1024'd82351870346084539964780392701565018125185967856083531296556399506004446965756159230862255788797594383684694821895279454942986047470856369109194837179570289687604695759249165799709189720552731605243988741726553722959848050181133866870296736926557881624890690936865484020841409323111142307808815255807087205835;
            6'd6: xpb[57] = 1024'd98822244415301447957736471241878021750223161427300237555867679407205336358907391077034706946557113260421633786274335345931583256965027642931033804615484347625125634911098998959651027664663277926292786490071864467551817660217360640244356084311869457949868829124238580825009691187733370769370578306968504647002;
            6'd7: xpb[57] = 1024'd115292618484518355950692549782191025375260354998516943815178959308406225752058622923207158104316632137158572750653391236920180466459198916752872772051398405562646574062948832119592865608773824247341584238417175212143787270253587413618415431697181034274846967311611677629177973052355599230932341358129922088169;
            6'd8: xpb[57] = 1024'd7696296869610522544849700917689596255599121443997965946358384144630219807900715859364538047418476704452362307574953693329713835112149856019551614470981422566476838645227447941904464361367164847080184378375246110371396030068917414027496209399263161333005202084867716403239726843049194675375414582665745045005;
            6'd9: xpb[57] = 1024'd24166670938827430537805779458002599880636315015214672205669664045831109201051947705536989205177995581189301271954009584318311044606321129841390581906895480503997777797077281101846302305477711168128982126720556854963365640105144187401555556784574737657983340272240813207408008707671423136937177633827162486172;
            6'd10: xpb[57] = 1024'd40637045008044338530761857998315603505673508586431378464980943947031998594203179551709440362937514457926240236333065475306908254100492403663229549342809538441518716948927114261788140249588257489177779875065867599555335250141370960775614904169886313982961478459613910011576290572293651598498940684988579927339;
            6'd11: xpb[57] = 1024'd57107419077261246523717936538628607130710702157648084724292223848232887987354411397881891520697033334663179200712121366295505463594663677485068516778723596379039656100776947421729978193698803810226577623411178344147304860177597734149674251555197890307939616646987006815744572436915880060060703736149997368506;
            6'd12: xpb[57] = 1024'd73577793146478154516674015078941610755747895728864790983603503749433777380505643244054342678456552211400118165091177257284102673088834951306907484214637654316560595252626780581671816137809350131275375371756489088739274470213824507523733598940509466632917754834360103619912854301538108521622466787311414809673;
            6'd13: xpb[57] = 1024'd90048167215695062509630093619254614380785089300081497242914783650634666773656875090226793836216071088137057129470233148272699882583006225128746451650551712254081534404476613741613654081919896452324173120101799833331244080250051280897792946325821042957895893021733200424081136166160336983184229838472832250840;
            6'd14: xpb[57] = 1024'd106518541284911970502586172159567618005822282871298203502226063551835556166808106936399244993975589964873996093849289039261297092077177498950585419086465770191602473556326446901555492026030442773372970868447110577923213690286278054271852293711132619282874031209106297228249418030782565444745992889634249692007;
            6'd15: xpb[57] = 1024'd122988915354128878495542250699880621630859476442514909761537343453036445559959338782571696151735108841610935058228344930249894301571348772772424386522379828129123412708176280061497329970140989094421768616792421322515183300322504827645911641096444195607852169396479394032417699895404793906307755940795667133174;
            6'd16: xpb[57] = 1024'd15392593739221045089699401835379192511198242887995931892716768289260439615801431718729076094836953408904724615149907386659427670224299712039103228941962845132953677290454895883808928722734329694160368756750492220742792060137834828054992418798526322666010404169735432806479453686098389350750829165331490090010;
            6'd17: xpb[57] = 1024'd31862967808437953082655480375692196136235436459212638152028048190461329008952663564901527252596472285641663579528963277648024879718470985860942196377876903070474616442304729043750766666844876015209166505095802965334761670174061601429051766183837898990988542357108529610647735550720617812312592216492907531177;
            6'd18: xpb[57] = 1024'd48333341877654861075611558916005199761272630030429344411339328091662218402103895411073978410355991162378602543908019168636622089212642259682781163813790961007995555594154562203692604610955422336257964253441113709926731280210288374803111113569149475315966680544481626414816017415342846273874355267654324972344;
            6'd19: xpb[57] = 1024'd64803715946871769068567637456318203386309823601646050670650607992863107795255127257246429568115510039115541508287075059625219298706813533504620131249705018945516494746004395363634442555065968657306762001786424454518700890246515148177170460954461051640944818731854723218984299279965074735436118318815742413511;
            6'd20: xpb[57] = 1024'd81274090016088677061523715996631207011347017172862756929961887894063997188406359103418880725875028915852480472666130950613816508200984807326459098685619076883037433897854228523576280499176514978355559750131735199110670500282741921551229808339772627965922956919227820023152581144587303196997881369977159854678;
            6'd21: xpb[57] = 1024'd97744464085305585054479794536944210636384210744079463189273167795264886581557590949591331883634547792589419437045186841602413717695156081148298066121533134820558373049704061683518118443287061299404357498477045943702640110318968694925289155725084204290901095106600916827320863009209531658559644421138577295845;
            6'd22: xpb[57] = 1024'd114214838154522493047435873077257214261421404315296169448584447696465775974708822795763783041394066669326358401424242732591010927189327354970137033557447192758079312201553894843459956387397607620453155246822356688294609720355195468299348503110395780615879233293974013631489144873831760120121407472299994737012;
            6'd23: xpb[57] = 1024'd6618516539614659641593024212755785141760170760777191579763872532689770030550915731921162984495911236620147958345805189000544295842278294236815875977030209761909576783832510665771555139990948220191755386780427586522218480170525468708429280812477907674037468067230052405550898664525355564564480696835817693848;
            6'd24: xpb[57] = 1024'd23088890608831567634549102753068788766797364331993897839075152433890659423702147578093614142255430113357086922724861079989141505336449568058654843412944267699430515935682343825713393084101494541240553135125738331114188090206752242082488628197789483999015606254603149209719180529147584026126243747997235135015;
            6'd25: xpb[57] = 1024'd39559264678048475627505181293381792391834557903210604098386432335091548816853379424266065300014948990094025887103916970977738714830620841880493810848858325636951455087532176985655231028212040862289350883471049075706157700242979015456547975583101060323993744441976246013887462393769812487688006799158652576182;
            6'd26: xpb[57] = 1024'd56029638747265383620461259833694796016871751474427310357697712236292438210004611270438516457774467866830964851482972861966335924324792115702332778284772383574472394239382010145597068972322587183338148631816359820298127310279205788830607322968412636648971882629349342818055744258392040949249769850320070017349;
            6'd27: xpb[57] = 1024'd72500012816482291613417338374007799641908945045644016617008992137493327603155843116610967615533986743567903815862028752954933133818963389524171745720686441511993333391231843305538906916433133504386946380161670564890096920315432562204666670353724212973950020816722439622224026123014269410811532901481487458516;
            6'd28: xpb[57] = 1024'd88970386885699199606373416914320803266946138616860722876320272038694216996307074962783418773293505620304842780241084643943530343313134663346010713156600499449514272543081676465480744860543679825435744128506981309482066530351659335578726017739035789298928159004095536426392307987636497872373295952642904899683;
            6'd29: xpb[57] = 1024'd105440760954916107599329495454633806891983332188077429135631551939895106389458306808955869931053024497041781744620140534932127552807305937167849680592514557387035211694931509625422582804654226146484541876852292054074036140387886108952785365124347365623906297191468633230560589852258726333935059003804322340850;
            6'd30: xpb[57] = 1024'd121911135024133015592285573994946810517020525759294135394942831841095995782609538655128321088812543373778720708999196425920724762301477210989688648028428615324556150846781342785364420748764772467533339625197602798666005750424112882326844712509658941948884435378841730034728871716880954795496822054965739782017;
            6'd31: xpb[57] = 1024'd14314813409225182186442725130445381397359292204775157526122256677319989838451631591285701031914387941072510265920758882330258130954428150256367490448011632328386415429059958607676019501358113067271939765155673696893614510239442882735925490211741069007042670152097768808790625507574550239939895279501562738853;
            6'd32: xpb[57] = 1024'd30785187478442090179398803670758385022396485775991863785433536578520879231602863437458152189673906817809449230299814773318855340448599424078206457883925690265907354580909791767617857445468659388320737513500984441485584120275669656109984837597052645332020808339470865612958907372196778701501658330662980180020;
            6'd33: xpb[57] = 1024'd47255561547658998172354882211071388647433679347208570044744816479721768624754095283630603347433425694546388194678870664307452549942770697900045425319839748203428293732759624927559695389579205709369535261846295186077553730311896429484044184982364221656998946526843962417127189236819007163063421381824397621187;
            6'd34: xpb[57] = 1024'd63725935616875906165310960751384392272470872918425276304056096380922658017905327129803054505192944571283327159057926555296049759436941971721884392755753806140949232884609458087501533333689752030418333010191605930669523340348123202858103532367675797981977084714217059221295471101441235624625184432985815062354;
            6'd35: xpb[57] = 1024'd80196309686092814158267039291697395897508066489641982563367376282123547411056558975975505662952463448020266123436982446284646968931113245543723360191667864078470172036459291247443371277800298351467130758536916675261492950384349976232162879752987374306955222901590156025463752966063464086186947484147232503521;
            6'd36: xpb[57] = 1024'd96666683755309722151223117832010399522545260060858688822678656183324436804207790822147956820711982324757205087816038337273244178425284519365562327627581922015991111188309124407385209221910844672515928506882227419853462560420576749606222227138298950631933361088963252829632034830685692547748710535308649944688;
            6'd37: xpb[57] = 1024'd113137057824526630144179196372323403147582453632075395081989936084525326197359022668320407978471501201494144052195094228261841387919455793187401295063495979953512050340158957567327047166021390993564726255227538164445432170456803522980281574523610526956911499276336349633800316695307921009310473586470067385855;
            6'd38: xpb[57] = 1024'd5540736209618796738336347507821974027921220077556417213169360920749320253201115604477787921573345768787933609116656684671374756572406732454080137483078996957342314922437573389638645918614731593303326395185609062673040930272133523389362352225692654015069734049592388407862070486001516453753546811005890342691;
            6'd39: xpb[57] = 1024'd22011110278835704731292426048134977652958413648773123472480640821950209646352347450650239079332864645524872573495712575659971966066578006275919104918993054894863254074287406549580483862725277914352124143530919807265010540308360296763421699611004230340047872236965485212030352350623744915315309862167307783858;
            6'd40: xpb[57] = 1024'd38481484348052612724248504588447981277995607219989829731791920723151099039503579296822690237092383522261811537874768466648569175560749280097758072354907112832384193226137239709522321806835824235400921891876230551856980150344587070137481046996315806665026010424338582016198634215245973376877072913328725225025;
            6'd41: xpb[57] = 1024'd54951858417269520717204583128760984903032800791206535991103200624351988432654811142995141394851902398998750502253824357637166385054920553919597039790821170769905132377987072869464159750946370556449719640221541296448949760380813843511540394381627382990004148611711678820366916079868201838438835964490142666192;
            6'd42: xpb[57] = 1024'd71422232486486428710160661669073988528069994362423242250414480525552877825806042989167592552611421275735689466632880248625763594549091827741436007226735228707426071529836906029405997695056916877498517388566852041040919370417040616885599741766938959314982286799084775624535197944490430300000599015651560107359;
            6'd43: xpb[57] = 1024'd87892606555703336703116740209386992153107187933639948509725760426753767218957274835340043710370940152472628431011936139614360804043263101563274974662649286644947010681686739189347835639167463198547315136912162785632888980453267390259659089152250535639960424986457872428703479809112658761562362066812977548526;
            6'd44: xpb[57] = 1024'd104362980624920244696072818749699995778144381504856654769037040327954656612108506681512494868130459029209567395390992030602958013537434375385113942098563344582467949833536572349289673583278009519596112885257473530224858590489494163633718436537562111964938563173830969232871761673734887223124125117974394989693;
            6'd45: xpb[57] = 1024'd120833354694137152689028897290012999403181575076073361028348320229155546005259738527684946025889977905946506359770047921591555223031605649206952909534477402519988888985386405509231511527388555840644910633602784274816828200525720937007777783922873688289916701361204066037040043538357115684685888169135812430860;
            6'd46: xpb[57] = 1024'd13237033079229319283186048425511570283520341521554383159527745065379540061101831463842325968991822473240295916691610378001088591684556588473631751954060419523819153567665021331543110279981896440383510773560855173044436960341050937416858561624955815348074936134460104811101797329050711129128961393671635387696;
            6'd47: xpb[57] = 1024'd29707407148446227276142126965824573908557535092771089418839024966580429454253063310014777126751341349977234881070666268989685801178727862295470719389974477461340092719514854491484948224092442761432308521906165917636406570377277710790917909010267391673053074321833201615270079193672939590690724444833052828863;
            6'd48: xpb[57] = 1024'd46177781217663135269098205506137577533594728663987795678150304867781318847404295156187228284510860226714173845449722159978283010672899136117309686825888535398861031871364687651426786168202989082481106270251476662228376180413504484164977256395578967998031212509206298419438361058295168052252487495994470270030;
            6'd49: xpb[57] = 1024'd62648155286880043262054284046450581158631922235204501937461584768982208240555527002359679442270379103451112809828778050966880220167070409939148654261802593336381971023214520811368624112313535403529904018596787406820345790449731257539036603780890544323009350696579395223606642922917396513814250547155887711197;
            6'd50: xpb[57] = 1024'd79118529356096951255010362586763584783669115806421208196772864670183097633706758848532130600029897980188051774207833941955477429661241683760987621697716651273902910175064353971310462056424081724578701766942098151412315400485958030913095951166202120647987488883952492027774924787539624975376013598317305152364;
            6'd51: xpb[57] = 1024'd95588903425313859247966441127076588408706309377637914456084144571383987026857990694704581757789416856924990738586889832944074639155412957582826589133630709211423849326914187131252300000534628045627499515287408896004285010522184804287155298551513696972965627071325588831943206652161853436937776649478722593531;
            6'd52: xpb[57] = 1024'd112059277494530767240922519667389592033743502948854620715395424472584876420009222540877032915548935733661929702965945723932671848649584231404665556569544767148944788478764020291194137944645174366676297263632719640596254620558411577661214645936825273297943765258698685636111488516784081898499539700640140034698;
            6'd53: xpb[57] = 1024'd4462955879622933835079670802888162914082269394335642846574849308808870475851315477034412858650780300955719259887508180342205217302535170671344398989127784152775053061042636113505736697238514966414897403590790538823863380373741578070295423638907400356102000031954724410173242307477677342942612925175962991534;
            6'd54: xpb[57] = 1024'd20933329948839841828035749343201166539119462965552349105886129210009759869002547323206864016410299177692658224266564071330802426796706444493183366425041842090295992212892469273447574641349061287463695151936101283415832990409968351444354771024218976681080138219327821214341524172099905804504375976337380432701;
            6'd55: xpb[57] = 1024'd37403704018056749820991827883514170164156656536769055365197409111210649262153779169379315174169818054429597188645619962319399636290877718315022333860955900027816931364742302433389412585459607608512492900281412028007802600446195124818414118409530553006058276406700918018509806036722134266066139027498797873868;
            6'd56: xpb[57] = 1024'd53874078087273657813947906423827173789193850107985761624508689012411538655305011015551766331929336931166536153024675853307996845785048992136861301296869957965337870516592135593331250529570153929561290648626722772599772210482421898192473465794842129331036414594074014822678087901344362727627902078660215315035;
            6'd57: xpb[57] = 1024'd70344452156490565806903984964140177414231043679202467883819968913612428048456242861724217489688855807903475117403731744296594055279220265958700268732784015902858809668441968753273088473680700250610088396972033517191741820518648671566532813180153705656014552781447111626846369765966591189189665129821632756202;
            6'd58: xpb[57] = 1024'd86814826225707473799860063504453181039268237250419174143131248814813317441607474707896668647448374684640414081782787635285191264773391539780539236168698073840379748820291801913214926417791246571658886145317344261783711430554875444940592160565465281980992690968820208431014651630588819650751428180983050197369;
            6'd59: xpb[57] = 1024'd103285200294924381792816142044766184664305430821635880402442528716014206834758706554069119805207893561377353046161843526273788474267562813602378203604612131777900687972141635073156764361901792892707683893662655006375681040591102218314651507950776858305970829156193305235182933495211048112313191232144467638536;
            6'd60: xpb[57] = 1024'd119755574364141289785772220585079188289342624392852586661753808617215096227909938400241570962967412438114292010540899417262385683761734087424217171040526189715421627123991468233098602306012339213756481642007965750967650650627328991688710855336088434630948967343566402039351215359833276573874954283305885079703;
            6'd61: xpb[57] = 1024'd12159252749233456379929371720577759169681390838333608792933233453439090283752031336398950906069257005408081567462461873671919052414685026690896013460109206719251891706270084055410201058605679813495081781966036649195259410442658992097791633038170561689107202116822440813412969150526872018318027507841708036539;
            6'd62: xpb[57] = 1024'd28629626818450364372885450260890762794718584409550315052244513354639979676903263182571402063828775882145020531841517764660516261908856300512734980896023264656772830858119917215352039002716226134543879530311347393787229020478885765471850980423482138014085340304195537617581251015149100479879790559003125477706;
            6'd63: xpb[57] = 1024'd45100000887667272365841528801203766419755777980767021311555793255840869070054495028743853221588294758881959496220573655649113471403027574334573948331937322594293770009969750375293876946826772455592677278656658138379198630515112538845910327808793714339063478491568634421749532879771328941441553610164542918873;
        endcase
    end

    always_comb begin
        case(flag[19][11:6])
            6'd0: xpb[58] = 1024'd0;
            6'd1: xpb[58] = 1024'd61570374956884180358797607341516770044792971551983727570867073157041758463205726874916304379347813635618898460599629546637710680897198848156412915767851380531814709161819583535235714890937318776641475027001968882971168240551339312219969675194105290664041616678941731225917814744393557403003316661325960360040;
            6'd2: xpb[58] = 1024'd123140749913768360717595214683033540089585943103967455141734146314083516926411453749832608758695627271237796921199259093275421361794397696312825831535702761063629418323639167070471429781874637553282950054003937765942336481102678624439939350388210581328083233357883462451835629488787114806006633322651920720080;
            6'd3: xpb[58] = 1024'd60644429186527799677593894619735877389680487530215498584469364406148380052308041714733841923385766597413545974341395205334068201850376209914078622287223100661753452915887533268076905481294750608614227472618666802549143871433121163694930455899086422725304946622708135647646916159252039191891260157352286595789;
            6'd4: xpb[58] = 1024'd122214804143411980036391501961252647434473459082199226155336437563190138515513768589650146302733580233032444434941024751971778882747575058070491538055074481193568162077707116803312620372232069385255702499620635685520312111984460475914900131093191713389346563301649866873564730903645596594894576818678246955829;
            6'd5: xpb[58] = 1024'd59718483416171418996390181897954984734568003508447269598071655655255001641410356554551379467423719559208193488083160864030425722803553571671744328806594820791692196669955483000918096071652182440586979918235364722127119502314903015169891236604067554786568276566474540069376017574110520980779203653378612831538;
            6'd6: xpb[58] = 1024'd121288858373055599355187789239471754779360975060430997168938728812296760104616083429467683846771533194827091948682790410668136403700752419828157244574446201323506905831775066536153810962589501217228454945237333605098287742866242327389860911798172845450609893245416271295293832318504078383782520314704573191578;
            6'd7: xpb[58] = 1024'd58792537645815038315186469176174092079455519486679040611673946904361623230512671394368917011461672521002841001824926522726783243756730933429410035325966540921630940424023432733759286662009614272559732363852062641705095133196684866644852017309048686847831606510240944491105118988969002769667147149404939067287;
            6'd8: xpb[58] = 1024'd120362912602699218673984076517690862124248491038662768182541020061403381693718398269285221390809486156621739462424556069364493924653929781585822951093817921453445649585843016268995001552946933049201207390854031524676263373748024178864821692503153977511873223189182675717022933733362560172670463810730899427327;
            6'd9: xpb[58] = 1024'd57866591875458657633982756454393199424343035464910811625276238153468244819614986234186454555499625482797488515566692181423140764709908295187075741845338261051569684178091382466600477252367046104532484809468760561283070764078466718119812798014029818909094936454007348912834220403827484558555090645431265303036;
            6'd10: xpb[58] = 1024'd119436966832342837992780363795909969469136007016894539196143311310510003282820713109102758934847439118416386976166321728060851445607107143343488657613189641583384393339910966001836192143304364881173959836470729444254239004629806030339782473208135109573136553132949080138752035148221041961558407306757225663076;
            6'd11: xpb[58] = 1024'd56940646105102276952779043732612306769230551443142582638878529402574866408717301074003992099537578444592136029308457840119498285663085656944741448364709981181508427932159332199441667842724477936505237255085458480861046394960248569594773578719010950970358266397773753334563321818685966347443034141457591538785;
            6'd12: xpb[58] = 1024'd118511021061986457311576651074129076814023522995126310209745602559616624871923027948920296478885392080211034489908087386757208966560284505101154364132561361713323137093978915734677382733661796713146712282087427363832214635511587881814743253913116241634399883076715484560481136563079523750446350802783551898825;
            6'd13: xpb[58] = 1024'd56014700334745896271575331010831414114118067421374353652480820651681487997819615913821529643575531406386783543050223498815855806616263018702407154884081701311447171686227281932282858433081909768477989700702156400439022025842030421069734359423992083031621596341540157756292423233544448136330977637483917774534;
            6'd14: xpb[58] = 1024'd117585075291630076630372938352348184158911038973358081223347893808723246461025342788737834022923345042005682003649853045453566487513461866858820070651933081843261880848046865467518573324019228545119464727704125283410190266393369733289704034618097373695663213020481888982210237977938005539334294298809878134574;
            6'd15: xpb[58] = 1024'd55088754564389515590371618289050521459005583399606124666083111900788109586921930753639067187613484368181431056791989157512213327569440380460072861403453421441385915440295231665124049023439341600450742146318854320016997656723812272544695140128973215092884926285306562178021524648402929925218921133510244010283;
            6'd16: xpb[58] = 1024'd116659129521273695949169225630567291503798554951589852236950185057829868050127657628555371566961298003800329517391618704149924008466639228616485777171304801973200624602114815200359763914376660377092217173320823202988165897275151584764664815323078505756926542964248293403939339392796487328222237794836204370323;
            6'd17: xpb[58] = 1024'd54162808794033134909167905567269628803893099377837895679685403149894731176024245593456604731651437329976078570533754816208570848522617742217738567922825141571324659194363181397965239613796773432423494591935552239594973287605594124019655920833954347154148256229072966599750626063261411714106864629536570246032;
            6'd18: xpb[58] = 1024'd115733183750917315267965512908786398848686070929821623250552476306936489639229972468372909110999250965594977031133384362846281529419816590374151483690676522103139368356182764933200954504734092209064969618937521122566141528156933436239625596028059637818189872908014697825668440807654969117110181290862530606072;
            6'd19: xpb[58] = 1024'd53236863023676754227964192845488736148780615356069666693287694399001352765126560433274142275689390291770726084275520474904928369475795103975404274442196861701263402948431131130806430204154205264396247037552250159172948918487375975494616701538935479215411586172839371021479727478119893502994808125562896481781;
            6'd20: xpb[58] = 1024'd114807237980560934586761800187005506193573586908053394264154767556043111228332287308190446655037203927389624544875150021542639050372993952131817190210048242233078112110250714666042145095091524041037722064554219042144117159038715287714586376733040769879453202851781102247397542222513450905998124786888856841821;
            6'd21: xpb[58] = 1024'd52310917253320373546760480123707843493668131334301437706889985648107974354228875273091679819727343253565373598017286133601285890428972465733069980961568581831202146702499080863647620794511637096368999483168948078750924549369157826969577482243916611276674916116605775443208828892978375291882751621589222717530;
            6'd22: xpb[58] = 1024'd113881292210204553905558087465224613538461102886285165277757058805149732817434602148007984199075156889184272058616915680238996571326171313889482896729419962363016855864318664398883335685448955873010474510170916961722092789920497139189547157438021901940716532795547506669126643637371932694886068282915183077570;
            6'd23: xpb[58] = 1024'd51384971482963992865556767401926950838555647312533208720492276897214595943331190112909217363765296215360021111759051792297643411382149827490735687480940301961140890456567030596488811384869068928341751928785645998328900180250939678444538262948897743337938246060372179864937930307836857080770695117615548953279;
            6'd24: xpb[58] = 1024'd112955346439848173224354374743443720883348618864516936291359350054256354406536916987825521743113109850978919572358681338935354092279348675647148603248791682492955599618386614131724526275806387704983226955787614881300068420802278990664507938143003034001979862739313911090855745052230414483774011778941509313319;
            6'd25: xpb[58] = 1024'd50459025712607612184353054680146058183443163290764979734094568146321217532433504952726754907803249177154668625500817450994000932335327189248401394000312022091079634210634980329330001975226500760314504374402343917906875811132721529919499043653878875399201576004138584286667031722695338869658638613641875189028;
            6'd26: xpb[58] = 1024'd112029400669491792543150662021662828228236134842748707304961641303362975995639231827643059287151062812773567086100446997631711613232526037404814309768163402622894343372454563864565716866163819536955979401404312800878044051684060842139468718847984166063243192683080315512584846467088896272661955274967835549068;
            6'd27: xpb[58] = 1024'd49533079942251231503149341958365165528330679268996750747696859395427839121535819792544292451841202138949316139242583109690358453288504551006067100519683742221018377964702930062171192565583932592287256820019041837484851442014503381394459824358860007460464905947904988708396133137553820658546582109668201424777;
            6'd28: xpb[58] = 1024'd111103454899135411861946949299881935573123650820980478318563932552469597584741546667460596831189015774568214599842212656328069134185703399162480016287535122752833087126522513597406907456521251368928731847021010720456019682565842693614429499552965298124506522626846719934313947881947378061549898770994161784817;
            6'd29: xpb[58] = 1024'd48607134171894850821945629236584272873218195247228521761299150644534460710638134632361829995879155100743963652984348768386715974241681912763732807039055462350957121718770879795012383155941364424260009265635739757062827072896285232869420605063841139521728235891671393130125234552412302447434525605694527660526;
            6'd30: xpb[58] = 1024'd110177509128779031180743236578101042918011166799212249332166223801576219173843861507278134375226968736362862113583978315024426655138880760920145722806906842882771830880590463330248098046878683200901484292637708640033995313447624545089390280257946430185769852570613124356043049296805859850437842267020488020566;
            6'd31: xpb[58] = 1024'd47681188401538470140741916514803380218105711225460292774901441893641082299740449472179367539917108062538611166726114427083073495194859274521398513558427182480895865472838829527853573746298796256232761711252437676640802703778067084344381385768822271582991565835437797551854335967270784236322469101720853896275;
            6'd32: xpb[58] = 1024'd109251563358422650499539523856320150262898682777444020345768515050682840762946176347095671919264921698157509627325743973720784176092058122677811429326278563012710574634658413063089288637236115032874236738254406559611970944329406396564351060962927562247033182514379528777772150711664341639325785763046814256315;
            6'd33: xpb[58] = 1024'd46755242631182089459538203793022487562993227203692063788503733142747703888842764311996905083955061024333258680467880085779431016148036636279064220077798902610834609226906779260694764336656228088205514156869135596218778334659848935819342166473803403644254895779204201973583437382129266025210412597747180132024;
            6'd34: xpb[58] = 1024'd108325617588066269818335811134539257607786198755675791359370806299789462352048491186913209463302874659952157141067509632417141697045235484435477135845650283142649318388726362795930479227593546864846989183871104479189946575211188248039311841667908694308296512458145933199501252126522823428213729259073140492064;
            6'd35: xpb[58] = 1024'd45829296860825708778334491071241594907880743181923834802106024391854325477945079151814442627993013986127906194209645744475788537101213998036729926597170622740773352980974728993535954927013659920178266602485833515796753965541630787294302947178784535705518225722970606395312538796987747814098356093773506367773;
            6'd36: xpb[58] = 1024'd107399671817709889137132098412758364952673714733907562372973097548896083941150806026730747007340827621746804654809275291113499217998412846193142842365022003272588062142794312528771669817950978696819741629487802398767922206092970099514272622372889826369559842401912337621230353541381305217101672755099466727813;
            6'd37: xpb[58] = 1024'd44903351090469328097130778349460702252768259160155605815708315640960947067047393991631980172030966947922553707951411403172146058054391359794395633116542342870712096735042678726377145517371091752151019048102531435374729596423412638769263727883765667766781555666737010817041640211846229602986299589799832603522;
            6'd38: xpb[58] = 1024'd106473726047353508455928385690977472297561230712139333386575388798002705530253120866548284551378780583541452168551040949809856738951590207950808548884393723402526805896862262261612860408308410528792494075104500318345897836974751950989233403077870958430823172345678742042959454956239787005989616251125792963562;
            6'd39: xpb[58] = 1024'd43977405320112947415927065627679809597655775138387376829310606890067568656149708831449517716068919909717201221693177061868503579007568721552061339635914063000650840489110628459218336107728523584123771493719229354952705227305194490244224508588746799828044885610503415238770741626704711391874243085826158839271;
            6'd40: xpb[58] = 1024'd105547780276997127774724672969196579642448746690371104400177680047109327119355435706365822095416733545336099682292806608506214259904767569708474255403765443532465549650930211994454050998665842360765246520721198237923873467856533802464194183782852090492086502289445146464688556371098268794877559747152119199311;
            6'd41: xpb[58] = 1024'd43051459549756566734723352905898916942543291116619147842912898139174190245252023671267055260106872871511848735434942720564861099960746083309727046155285783130589584243178578192059526698085955416096523939335927274530680858186976341719185289293727931889308215554269819660499843041563193180762186581852485075020;
            6'd42: xpb[58] = 1024'd104621834506640747093520960247415686987336262668602875413779971296215948708457750546183359639454686507130747196034572267202571780857944931466139961923137163662404293404998161727295241589023274192737998966337896157501849098738315653939154964487833222553349832233211550886417657785956750583765503243178445435060;
            6'd43: xpb[58] = 1024'd42125513779400186053519640184118024287430807094850918856515189388280811834354338511084592804144825833306496249176708379261218620913923445067392752674657503260528327997246527924900717288443387248069276384952625194108656489068758193194146069998709063950571545498036224082228944456421674969650130077878811310769;
            6'd44: xpb[58] = 1024'd103695888736284366412317247525634794332223778646834646427382262545322570297560065386000897183492639468925394709776337925898929301811122293223805668442508883792343037159066111460136432179380706024710751411954594077079824729620097505414115745192814354614613162176977955308146759200815232372653446739204771670809;
            6'd45: xpb[58] = 1024'd41199568009043805372315927462337131632318323073082689870117480637387433423456653350902130348182778795101143762918474037957576141867100806825058459194029223390467071751314477657741907878800819080042028830569323113686632119950540044669106850703690196011834875441802628503958045871280156758538073573905137546518;
            6'd46: xpb[58] = 1024'd102769942965927985731113534803853901677111294625066417440984553794429191886662380225818434727530592430720042223518103584595286822764299654981471374961880603922281780913134061192977622769738137856683503857571291996657800360501879356889076525897795486675876492120744359729875860615673714161541390235231097906558;
            6'd47: xpb[58] = 1024'd40273622238687424691112214740556238977205839051314460883719771886494055012558968190719667892220731756895791276660239696653933662820278168582724165713400943520405815505382427390583098469158250912014781276186021033264607750832321896144067631408671328073098205385569032925687147286138638547426017069931463782267;
            6'd48: xpb[58] = 1024'd101843997195571605049909822082073009021998810603298188454586845043535813475764695065635972271568545392514689737259869243291644343717477016739137081481252324052220524667202010925818813360095569688656256303187989916235775991383661208364037306602776618737139822064510764151604962030532195950429333731257424142307;
            6'd49: xpb[58] = 1024'd39347676468331044009908502018775346322093355029546231897322063135600676601661283030537205436258684718690438790402005355350291183773455530340389872232772663650344559259450377123424289059515682743987533721802718952842583381714103747619028412113652460134361535329335437347416248700997120336313960565957790018016;
            6'd50: xpb[58] = 1024'd100918051425215224368706109360292116366886326581529959468189136292642435064867009905453509815606498354309337251001634901988001864670654378496802788000624044182159268421269960658660003950453001520629008748804687835813751622265443059838998087307757750798403152008277168573334063445390677739317277227283750378056;
            6'd51: xpb[58] = 1024'd38421730697974663328704789296994453666980871007778002910924354384707298190763597870354742980296637680485086304143771014046648704726632892098055578752144383780283303013518326856265479649873114575960286167419416872420559012595885599093989192818633592195624865273101841769145350115855602125201904061984116253765;
            6'd52: xpb[58] = 1024'd99992105654858843687502396638511223711773842559761730481791427541749056653969324745271047359644451316103984764743400560684359385623831740254468494519995764312098012175337910391501194540810433352601761194421385755391727253147224911313958868012738882859666481952043572995063164860249159528205220723310076613805;
            6'd53: xpb[58] = 1024'd37495784927618282647501076575213561011868386986009773924526645633813919779865912710172280524334590642279733817885536672743006225679810253855721285271516103910222046767586276589106670240230546407933038613036114791998534643477667450568949973523614724256888195216868246190874451530714083914089847558010442489514;
            6'd54: xpb[58] = 1024'd99066159884502463006298683916730331056661358537993501495393718790855678243071639585088584903682404277898632278485166219380716906577009102012134201039367484442036755929405860124342385131167865184574513640038083674969702884029006762788919648717720014920929811895809977416792266275107641317093164219336402849554;
            6'd55: xpb[58] = 1024'd36569839157261901966297363853432668356755902964241544938128936882920541368968227549989818068372543604074381331627302331439363746632987615613386991790887824040160790521654226321947860830587978239905791058652812711576510274359449302043910754228595856318151525160634650612603552945572565702977791054036768725263;
            6'd56: xpb[58] = 1024'd98140214114146082325094971194949438401548874516225272508996010039962299832173954424906122447720357239693279792226931878077074427530186463769799907558739204571975499683473809857183575721525297016547266085654781594547678514910788614263880429422701146982193141839576381838521367689966123105981107715362729085303;
            6'd57: xpb[58] = 1024'd35643893386905521285093651131651775701643418942473315951731228132027162958070542389807355612410496565869028845369067990135721267586164977371052698310259544170099534275722176054789051420945410071878543504269510631154485905241231153518871534933576988379414855104401055034332654360431047491865734550063094961012;
            6'd58: xpb[58] = 1024'd97214268343789701643891258473168545746436390494457043522598301289068921421276269264723659991758310201487927305968697536773431948483363825527465614078110924701914243437541759590024766311882728848520018531271479514125654145792570465738841210127682279043456471783342786260250469104824604894869051211389055321052;
            6'd59: xpb[58] = 1024'd34717947616549140603889938409870883046530934920705086965333519381133784547172857229624893156448449527663676359110833648832078788539342339128718404829631264300038278029790125787630242011302841903851295949886208550732461536123013004993832315638558120440678185048167459456061755775289529280753678046089421196761;
            6'd60: xpb[58] = 1024'd96288322573433320962687545751387653091323906472688814536200592538175543010378584104541197535796263163282574819710463195469789469436541187285131320597482644831852987191609709322865956902240160680492770976888177433703629776674352317213801990832663411104719801727109190681979570519683086683756994707415381556801;
            6'd61: xpb[58] = 1024'd33792001846192759922686225688089990391418450898936857978935810630240406136275172069442430700486402489458323872852599307528436309492519700886384111349002984429977021783858075520471432601660273735824048395502906470310437167004794856468793096343539252501941514991933863877790857190148011069641621542115747432510;
            6'd62: xpb[58] = 1024'd95362376803076940281483833029606760436211422450920585549802883787282164599480898944358735079834216125077222333452228854166146990389718549042797027116854364961791730945677659055707147492597592512465523422504875353281605407556134168688762771537644543165983131670875595103708671934541568472644938203441707792550;
            6'd63: xpb[58] = 1024'd32866056075836379241482512966309097736305966877168628992538101879347027725377486909259968244524355451252971386594364966224793830445697062644049817868374704559915765537926025253312623192017705567796800841119604389888412797886576707943753877048520384563204844935700268299519958605006492858529565038142073668259;
        endcase
    end

    always_comb begin
        case(flag[19][16:12])
            5'd0: xpb[59] = 1024'd0;
            5'd1: xpb[59] = 1024'd94436431032720559600280120307825867781098938429152356563405175036388786188583213784176272623872169086871869847193994512862504511342895910800462733636226085091730474699745608788548338082955024344438275868121573272859581038437916020163723552242625675227246461614641999525437773349400050261532881699468034028299;
            5'd2: xpb[59] = 1024'd64806166381316377801761313210837302817499449732569028998678495007800677039857288658337474033086663864300590286930495591145945181844571487045765342256121129249770274829920000239466436974392842967566354127855906699354801226654935267362468534802021901187673019815166941020769018624871467505947073572310473572267;
            5'd3: xpb[59] = 1024'd35175901729912196003242506113848737853899961035985701433951814979212567891131363532498675442301158641729310726666996669429385852346247063291067950876016173407810074960094391690384535865830661590694432387590240125850021414871954514561213517361418127148099578015691882516100263900342884750361265445152913116235;
            5'd4: xpb[59] = 1024'd5545637078508014204723699016860172890300472339402373869225134950624458742405438406659876851515653419158031166403497747712826522847922639536370559495911217565849875090268783141302634757268480213822510647324573552345241603088973761759958499920814353108526136216216824011431509175814301994775457317995352660203;
            5'd5: xpb[59] = 1024'd99982068111228573805003819324686040671399410768554730432630309987013244930988652190836149475387822506029901013597492260575331034190818550336833293132137302657580349790014391929850972840223504558260786515446146825204822641526889781923682052163440028335772597830858823536869282525214352256308339017463386688502;
            5'd6: xpb[59] = 1024'd70351803459824392006485012227697475707799922071971402867903629958425135782262727064997350884602317283458621453333993338858771704692494126582135901752032346815620149920188783380769071731661323181388864775180480251700042829743909029122427034722836254296199156031383765032200527800685769500722530890305826232470;
            5'd7: xpb[59] = 1024'd40721538808420210207966205130708910744200433375388075303176949929837026633536801939158552293816812060887341893070494417142212375194169702827438510371927390973659950050363174831687170623099141804516943034914813678195263017960928276321172017282232480256625714231908706527531773076157186745136722763148265776438;
            5'd8: xpb[59] = 1024'd11091274157016028409447398033720345780600944678804747738450269901248917484810876813319753703031306838316062332806995495425653045695845279072741118991822435131699750180537566282605269514536960427645021294649147104690483206177947523519916999841628706217052272432433648022863018351628603989550914635990705320406;
            5'd9: xpb[59] = 1024'd105527705189736588009727518341546213561699883107957104301855444937637703673394090597496026326903475925187932180000990008288157557038741189873203852628048520223430224880283175071153607597491984772083297162770720377550064244615863543683640552084254381444298734047075647548300791701028654251083796335458739348705;
            5'd10: xpb[59] = 1024'd75897440538332406211208711244557648598100394411373776737128764909049594524668165471657227736117970702616652619737491086571598227540416766118506461247943564381470025010457566522071706488929803395211375422505053804045284432832882790882385534643650607404725292247600589043632036976500071495497988208301178892673;
            5'd11: xpb[59] = 1024'd46267175886928224412689904147569083634500905714790449172402084880461485375942240345818429145332465480045373059473992164855038898042092342363809069867838608539509825140631957972989805380367622018339453682239387230540504621049902038081130517203046833365151850448125530538963282251971488739912180081143618436641;
            5'd12: xpb[59] = 1024'd16636911235524042614171097050580518670901417018207121607675404851873376227216315219979630554546960257474093499210493243138479568543767918609111678487733652697549625270806349423907904271805440641467531941973720657035724809266921285279875499762443059325578408648650472034294527527442905984326371953986057980609;
            5'd13: xpb[59] = 1024'd111073342268244602214451217358406386452000355447359478171080579888262162415799529004155903178419129344345963346404487756000984079886663829409574412123959737789280099970551958212456242354760464985905807810095293929895305847704837305443599052005068734552824870263292471559732300876842956245859253653454092008908;
            5'd14: xpb[59] = 1024'd81443077616840420415932410261417821488400866750776150606353899859674053267073603878317104587633624121774683786140988834284424750388339405654877020743854781947319900100726349663374341246198283609033886069829627356390526035921856552642344034564464960513251428463817413055063546152314373490273445526296531552876;
            5'd15: xpb[59] = 1024'd51812812965436238617413603164429256524801378054192823041627219831085944118347678752478305996848118899203404225877489912567865420890014981900179629363749826105359700230900741114292440137636102232161964329563960782885746224138875799841089017123861186473677986664342354550394791427785790734687637399138971096844;
            5'd16: xpb[59] = 1024'd22182548314032056818894796067440691561201889357609495476900539802497834969621753626639507406062613676632124665613990990851306091391690558145482237983644870263399500361075132565210539029073920855290042589298294209380966412355895047039833999683257412434104544864867296045726036703257207979101829271981410640812;
            5'd17: xpb[59] = 1024'd116618979346752616419174916375266559342300827786761852040305714838886621158204967410815780029934782763503994512807985503713810602734586468945944971619870955355129975060820741353758877112028945199728318457419867482240547450793811067203557551925883087661351006479509295571163810052657258240634710971449444669111;
            5'd18: xpb[59] = 1024'd86988714695348434620656109278277994378701339090178524475579034810298512009479042284976981439149277540932714952544486581997251273236262045191247580239765999513169775190995132804676976003466763822856396717154200908735767639010830314402302534485279313621777564680034237066495055328128675485048902844291884213079;
            5'd19: xpb[59] = 1024'd57358450043944252822137302181289429415101850393595196910852354781710402860753117159138182848363772318361435392280987660280691943737937621436550188859661043671209575321169524255595074894904582445984474976888534335230987827227849561601047517044675539582204122880559178561826300603600092729463094717134323757047;
            5'd20: xpb[59] = 1024'd27728185392540071023618495084300864451502361697011869346125674753122293712027192033299384257578267095790155832017488738564132614239613197681852797479556087829249375451343915706513173786342401069112553236622867761726208015444868808799792499604071765542630681081084120057157545879071509973877286589976763301015;
            5'd21: xpb[59] = 1024'd122164616425260630623898615392126732232601300126164225909530849789511079900610405817475656881450436182662025679211483251426637125582509108482315531115782172920979850151089524495061511869297425413550829104744441034585789053882784828963516051846697440769877142695726119582595319228471560235410168289444797329314;
            5'd22: xpb[59] = 1024'd92534351773856448825379808295138167269001811429580898344804169760922970751884480691636858290664930960090746118947984329710077796084184684727618139735677217079019650281263915945979610760735244036678907364478774461081009242099804076162261034406093666730303700896251061077926564503942977479824360162287236873282;
            5'd23: xpb[59] = 1024'd62904087122452267026861001198149602305402322732997570780077489732334861603158555565798059699879425737519466558684485407993518466585860260972920748355572261237059450411438307396897709652173062659806985624213107887576229430316823323361006016965489892690730259096776002573257809779414394724238552035129676417250;
            5'd24: xpb[59] = 1024'd33273822471048085228342194101161037341802834036414243215350809703746752454432630439959261109093920514948186998420986486276959137087535837218223356975467305395099250541612698847815808543610881282935063883947441314071449618533842570559750999524886118651156817297300944068589055054885811968652743907972115961218;
            5'd25: xpb[59] = 1024'd3643557819643903429823387004172472378203345339830915650624129675158643305706705314120462518308415292376907438157487564560399807589211413463525965595362349553139050671787090298733907435048699906063142143681774740566669806750861817758495982084282344611583375497825885563920300330357229213066935780814555505186;
            5'd26: xpb[59] = 1024'd98079988852364463030103507311998340159302283768983272214029304711547429494289919098296735142180584379248777285351482077422904318932107324263988699231588434644869525371532699087282245518003724250501418011803348013426250845188777837922219534326908019838829837112467885089358073679757279474599817480282589533485;
            5'd27: xpb[59] = 1024'd68449724200960281231584700215009775195702795072399944649302624682959320345563993972457936551395079156677497725087983155706344989433782900509291307851483478802909325501707090538200344409441542873629496271537681439921471033405797085120964516886304245799256395312992826584689318955228696719014009353125029077453;
            5'd28: xpb[59] = 1024'd38819459549556099433065893118021210232103306375816617084575944654371211196838068846619137960609573934106218164824484233989785659935458476754593916471378522960949125631881481989118443300879361496757574531272014866416691221622816332319709499445700471759682953513517768080020564230700113963428201225967468621421;
            5'd29: xpb[59] = 1024'd9189194898151917634547086021032645268503817679233289519849264625783102048112143720780339369824068711534938604560985312273226330437134052999896525091273567118988925762055873440036542192317180119885652791006348292911911409839835579518454482005096697720109511714042709575351809506171531207842393098809908165389;
            5'd30: xpb[59] = 1024'd103625625930872477234827206328858513049602756108385646083254439662171888236695357504956611993696237798406808451754979825135730841780029963800359258727499652210719400461801482228584880275272204464323928659127921565771492448277751599682178034247722372947355973328684709100789582855571581469375274798277942193688;
            5'd31: xpb[59] = 1024'd73995361279468295436308399231869948086003267411802318518527759633583779087969432379117813402910732575835528891491480903419171512281705540045661867347394696368759200591975873679502979166710023087452006918862254992266712636494770846880923016807118598907782531529209650596120828131042998713789466671120381737656;
        endcase
    end

    always_comb begin
        case(flag[20][5:0])
            6'd0: xpb[60] = 1024'd0;
            6'd1: xpb[60] = 1024'd22182548314032056818894796067440691561201889357609495476900539802497834969621753626639507406062613676632124665613990990851306091391690558145482237983644870263399500361075132565210539029073920855290042589298294209380966412355895047039833999683257412434104544864867296045726036703257207979101829271981410640812;
            6'd2: xpb[60] = 1024'd44365096628064113637789592134881383122403778715218990953801079604995669939243507253279014812125227353264249331227981981702612182783381116290964475967289740526799000722150265130421078058147841710580085178596588418761932824711790094079667999366514824868209089729734592091452073406514415958203658543962821281624;
            6'd3: xpb[60] = 1024'd66547644942096170456684388202322074683605668072828486430701619407493504908865260879918522218187841029896373996841972972553918274175071674436446713950934610790198501083225397695631617087221762565870127767894882628142899237067685141119501999049772237302313634594601888137178110109771623937305487815944231922436;
            6'd4: xpb[60] = 1024'd88730193256128227275579184269762766244807557430437981907602159209991339878487014506558029624250454706528498662455963963405224365566762232581928951934579481053598001444300530260842156116295683421160170357193176837523865649423580188159335998733029649736418179459469184182904146813028831916407317087925642563248;
            6'd5: xpb[60] = 1024'd110912741570160284094473980337203457806009446788047477384502699012489174848108768133197537030313068383160623328069954954256530456958452790727411189918224351316997501805375662826052695145369604276450212946491471046904832061779475235199169998416287062170522724324336480228630183516286039895509146359907053204060;
            6'd6: xpb[60] = 1024'd9028594200067599514569848999829716622512909019921288733271383750010114480421382849821973221718007750349598586226452510528772707508923014317733302885538180646706327596879578053632994982926319410430057927402525409921437623914473509274025428416315025337807365775086718244249692145614614857492285805262869360541;
            6'd7: xpb[60] = 1024'd31211142514099656333464645067270408183714798377530784210171923552507949450043136476461480627780621426981723251840443501380078798900613572463215540869183050910105827957954710618843534012000240265720100516700819619302404036270368556313859428099572437771911910639954014289975728848871822836594115077244280001353;
            6'd8: xpb[60] = 1024'd53393690828131713152359441134711099744916687735140279687072463355005784419664890103100988033843235103613847917454434492231384890292304130608697778852827921173505328319029843184054073041074161121010143105999113828683370448626263603353693427782829850206016455504821310335701765552129030815695944349225690642165;
            6'd9: xpb[60] = 1024'd75576239142163769971254237202151791306118577092749775163973003157503619389286643729740495439905848780245972583068425483082690981683994688754180016836472791436904828680104975749264612070148081976300185695297408038064336860982158650393527427466087262640121000369688606381427802255386238794797773621207101282977;
            6'd10: xpb[60] = 1024'd97758787456195826790149033269592482867320466450359270640873542960001454358908397356380002845968462456878097248682416473933997073075685246899662254820117661700304329041180108314475151099222002831590228284595702247445303273338053697433361427149344675074225545234555902427153838958643446773899602893188511923789;
            6'd11: xpb[60] = 1024'd119941335770227883609043829337033174428522355807968766117774082762499289328530150983019510252031076133510221914296407464785303164467375805045144492803762531963703829402255240879685690128295923686880270873893996456826269685693948744473195426832602087508330090099423198472879875661900654753001432165169922564601;
            6'd12: xpb[60] = 1024'd18057188400135199029139697999659433245025818039842577466542767500020228960842765699643946443436015500699197172452905021057545415017846028635466605771076361293412655193759156107265989965852638820860115854805050819842875247828947018548050856832630050675614731550173436488499384291229229714984571610525738721082;
            6'd13: xpb[60] = 1024'd40239736714167255848034494067100124806227707397452072943443307302518063930464519326283453849498629177331321838066896011908851506409536586780948843754721231556812155554834288672476528994926559676150158444103345029223841660184842065587884856515887463109719276415040732534225420994486437694086400882507149361894;
            6'd14: xpb[60] = 1024'd62422285028199312666929290134540816367429596755061568420343847105015898900086272952922961255561242853963446503680887002760157597801227144926431081738366101820211655915909421237687068024000480531440201033401639238604808072540737112627718856199144875543823821279908028579951457697743645673188230154488560002706;
            6'd15: xpb[60] = 1024'd84604833342231369485824086201981507928631486112671063897244386907513733869708026579562468661623856530595571169294877993611463689192917703071913319722010972083611156276984553802897607053074401386730243622699933447985774484896632159667552855882402287977928366144775324625677494401000853652290059426469970643518;
            6'd16: xpb[60] = 1024'd106787381656263426304718882269422199489833375470280559374144926710011568839329780206201976067686470207227695834908868984462769780584608261217395557705655842347010656638059686368108146082148322242020286211998227657366740897252527206707386855565659700412032911009642620671403531104258061631391888698451381284330;
            6'd17: xpb[60] = 1024'd4903234286170741724814750932048458306336837702154370722913611447532508471642394922826412259091409574416671093065366540735012031135078484807717670672969671676719482429563601595688445919705037376000131192909282020383346459387525480782242285565687663579317552460392858687023039733586636593375028143807197440811;
            6'd18: xpb[60] = 1024'd27085782600202798543709546999489149867538727059763866199814151250030343441264148549465919665154023251048795758679357531586318122526769042953199908656614541940118982790638734160898984948778958231290173782207576229764312871743420527822076285248945076013422097325260154732749076436843844572476857415788608081623;
            6'd19: xpb[60] = 1024'd49268330914234855362604343066929841428740616417373361676714691052528178410885902176105427071216636927680920424293348522437624213918459601098682146640259412203518483151713866726109523977852879086580216371505870439145279284099315574861910284932202488447526642190127450778475113140101052551578686687770018722435;
            6'd20: xpb[60] = 1024'd71450879228266912181499139134370532989942505774982857153615230855026013380507655802744934477279250604313045089907339513288930305310150159244164384623904282466917983512788999291320063006926799941870258960804164648526245696455210621901744284615459900881631187054994746824201149843358260530680515959751429363247;
            6'd21: xpb[60] = 1024'd93633427542298969000393935201811224551144395132592352630515770657523848350129409429384441883341864280945169755521330504140236396701840717389646622607549152730317483873864131856530602036000720797160301550102458857907212108811105668941578284298717313315735731919862042869927186546615468509782345231732840004059;
            6'd22: xpb[60] = 1024'd115815975856331025819288731269251916112346284490201848107416310460021683319751163056023949289404477957577294421135321494991542488093531275535128860591194022993716984234939264421741141065074641652450344139400753067288178521167000715981412283981974725749840276784729338915653223249872676488884174503714250644871;
            6'd23: xpb[60] = 1024'd13931828486238341239384599931878174928849746722075659456184995197542622952063777772648385480809417324766269679291819051263784738644001499125450973558507852323425810026443179649321440902631356786430189120311807430304784083301998990056267713982002688917124918235479576931272731879201251450867313949070066801352;
            6'd24: xpb[60] = 1024'd36114376800270398058279395999318866490051636079685154933085535000040457921685531399287892886872031001398394344905810042115090830035692057270933211542152722586825310387518312214531979931705277641720231709610101639685750495657894037096101713665260101351229463100346872976998768582458459429969143221051477442164;
            6'd25: xpb[60] = 1024'd58296925114302454877174192066759558051253525437294650409986074802538292891307285025927400292934644678030519010519801032966396921427382615416415449525797592850224810748593444779742518960779198497010274298908395849066716908013789084135935713348517513785334007965214169022724805285715667409070972493032888082976;
            6'd26: xpb[60] = 1024'd80479473428334511696068988134200249612455414794904145886886614605036127860929038652566907698997258354662643676133792023817703012819073173561897687509442463113624311109668577344953057989853119352300316888206690058447683320369684131175769713031774926219438552830081465068450841988972875388172801765014298723788;
            6'd27: xpb[60] = 1024'd102662021742366568514963784201640941173657304152513641363787154407533962830550792279206415105059872031294768341747783014669009104210763731707379925493087333377023811470743709910163597018927040207590359477504984267828649732725579178215603712715032338653543097694948761114176878692230083367274631036995709364600;
            6'd28: xpb[60] = 1024'd777874372273883935059652864267199990160766384387452712555839145054902462863406995830851296464811398483743599904280570941251354761233955297702038460401162706732637262247625137743896856483755341570204458416038630845255294860577452290459142715060301820827739145698999129796387321558658329257770482351525521081;
            6'd29: xpb[60] = 1024'd22960422686305940753954448931707891551362655741996948189456378947552737432485160622470358702527425075115868265518271561792557446152924513443184276444046032970132137623322757702954435885557676196860247047714332840226221707216472499330293142398317714254932284010566295175522424024815866308359599754332936161893;
            6'd30: xpb[60] = 1024'd45142971000337997572849244999148583112564545099606443666356918750050572402106914249109866108590038751747992931132262552643863537544615071588666514427690903233531637984397890268164974914631597052150289637012627049607188119572367546370127142081575126689036828875433591221248460728073074287461429026314346802705;
            6'd31: xpb[60] = 1024'd67325519314370054391744041066589274673766434457215939143257458552548407371728667875749373514652652428380117596746253543495169628936305629734148752411335773496931138345473022833375513943705517907440332226310921258988154531928262593409961141764832539123141373740300887266974497431330282266563258298295757443517;
            6'd32: xpb[60] = 1024'd89508067628402111210638837134029966234968323814825434620157998355046242341350421502388880920715266105012242262360244534346475720327996187879630990394980643760330638706548155398586052972779438762730374815609215468369120944284157640449795141448089951557245918605168183312700534134587490245665087570277168084329;
            6'd33: xpb[60] = 1024'd111690615942434168029533633201470657796170213172434930097058538157544077310972175129028388326777879781644366927974235525197781811719686746025113228378625514023730139067623287963796592001853359618020417404907509677750087356640052687489629141131347363991350463470035479358426570837844698224766916842258578725141;
            6'd34: xpb[60] = 1024'd9806468572341483449629501864096916612673675404308741445827222895065016943284789845652824518182819148833342186130733081470024062270156969615435341345939343353438964859127203191376891839410074752000262385818564040766692918775050961564484571131375327158635104920785717374046079467173273186750056287614394881622;
            6'd35: xpb[60] = 1024'd31989016886373540268524297931537608173875564761918236922727762697562851912906543472292331924245432825465466851744724072321330153661847527760917579329584213616838465220202335756587430868483995607290304975116858250147659331130946008604318570814632739592739649785653013419772116170430481165851885559595805522434;
            6'd36: xpb[60] = 1024'd54171565200405597087419093998978299735077454119527732399628302500060686882528297098931839330308046502097591517358715063172636245053538085906399817313229083880237965581277468321797969897557916462580347564415152459528625743486841055644152570497890152026844194650520309465498152873687689144953714831577216163246;
            6'd37: xpb[60] = 1024'd76354113514437653906313890066418991296279343477137227876528842302558521852150050725571346736370660178729716182972706054023942336445228644051882055296873954143637465942352600887008508926631837317870390153713446668909592155842736102683986570181147564460948739515387605511224189576944897124055544103558626804058;
            6'd38: xpb[60] = 1024'd98536661828469710725208686133859682857481232834746723353429382105056356821771804352210854142433273855361840848586697044875248427836919202197364293280518824407036966303427733452219047955705758173160432743011740878290558568198631149723820569864404976895053284380254901556950226280202105103157373375540037444870;
            6'd39: xpb[60] = 1024'd120719210142501767544103482201300374418683122192356218830329921907554191791393557978850361548495887531993965514200688035726554519228609760342846531264163694670436466664502866017429586984779679028450475332310035087671524980554526196763654569547662389329157829245122197602676262983459313082259202647521448085682;
            6'd40: xpb[60] = 1024'd18835062772409082964199350863926633235186584424230030179098606645075131423706172695474797739900826899182940772357185591998796769779079983933168644231477524000145292456006781245009886822336394162430320313221089450688130542689524470838509999547690352496442470695872435618295771612787888044242342092877264242163;
            6'd41: xpb[60] = 1024'd41017611086441139783094146931367324796388473781839525655999146447572966393327926322114305145963440575815065437971176582850102861170770542078650882215122394263544792817081913810220425851410315017720362902519383660069096955045419517878343999230947764930547015560739731664021808316045096023344171364858674882975;
            6'd42: xpb[60] = 1024'd63200159400473196601988942998808016357590363139449021132899686250070801362949679948753812552026054252447190103585167573701408952562461100224133120198767264526944293178157046375430964880484235873010405491817677869450063367401314564918177998914205177364651560425607027709747845019302304002446000636840085523787;
            6'd43: xpb[60] = 1024'd85382707714505253420883739066248707918792252497058516609800226052568636332571433575393319958088667929079314769199158564552715043954151658369615358182412134790343793539232178940641503909558156728300448081115972078831029779757209611958011998597462589798756105290474323755473881722559511981547829908821496164599;
            6'd44: xpb[60] = 1024'd107565256028537310239778535133689399479994141854668012086700765855066471302193187202032827364151281605711439434813149555404021135345842216515097596166057005053743293900307311505852042938632077583590490670414266288211996192113104658997845998280720002232860650155341619801199918425816719960649659180802906805411;
            6'd45: xpb[60] = 1024'd5681108658444625659874403796315658296497604086541823435469450592587410934505801918657263555556220972900414692969647111676263385896312440105419709133370834383452119691811226733432342776188792717570335651325320651228601754248102933072701428280747965400145291606091857816819427055145294922632798626158722961892;
            6'd46: xpb[60] = 1024'd27863656972476682478769199863756349857699493444151318912369990395085245904127555545296770961618834649532539358583638102527569477288002998250901947117015704646851620052886359298642881805262713572860378240623614860609568166603997980112535427964005377834249836470959153862545463758402502901734627898140133602704;
            6'd47: xpb[60] = 1024'd50046205286508739297663995931197041418901382801760814389270530197583080873749309171936278367681448326164664024197629093378875568679693556396384185100660574910251120413961491863853420834336634428150420829921909069990534578959893027152369427647262790268354381335826449908271500461659710880836457170121544243516;
            6'd48: xpb[60] = 1024'd72228753600540796116558791998637732980103272159370309866171070000080915843371062798575785773744062002796788689811620084230181660071384114541866423084305445173650620775036624429063959863410555283440463419220203279371500991315788074192203427330520202702458926200693745953997537164916918859938286442102954884328;
            6'd49: xpb[60] = 1024'd94411301914572852935453588066078424541305161516979805343071609802578750812992816425215293179806675679428913355425611075081487751463074672687348661067950315437050121136111756994274498892484476138730506008518497488752467403671683121232037427013777615136563471065561041999723573868174126839040115714084365525140;
            6'd50: xpb[60] = 1024'd116593850228604909754348384133519116102507050874589300819972149605076585782614570051854800585869289356061038021039602065932793842854765230832830899051595185700449621497186889559485037921558396994020548597816791698133433816027578168271871426697035027570668015930428338045449610571431334818141944986065776165952;
            6'd51: xpb[60] = 1024'd14709702858512225174444252796145374919010513106463112168740834342597525414927184768479236777274228723250013279196099622205036093405235454423153012018909015030158447288690804787065337759115112128000393578727846061150039378162576442346726856697062990737952657381178576061069119200759909780125084431421592322433;
            6'd52: xpb[60] = 1024'd36892251172544281993339048863586066480212402464072607645641374145095360384548938395118744183336842399882137944810090613056342184796926012568635250002553885293557947649765937352275876788189032983290436168026140270531005790518471489386560856380320403172057202246045872106795155904017117759226913703403002963245;
            6'd53: xpb[60] = 1024'd59074799486576338812233844931026758041414291821682103122541913947593195354170692021758251589399456076514262610424081603907648276188616570714117487986198755556957448010841069917486415817262953838580478757324434479911972202874366536426394856063577815606161747110913168152521192607274325738328742975384413604057;
            6'd54: xpb[60] = 1024'd81257347800608395631128640998467449602616181179291598599442453750091030323792445648397758995462069753146387276038072594758954367580307128859599725969843625820356948371916202482696954846336874693870521346622728689292938615230261583466228855746835228040266291975780464198247229310531533717430572247365824244869;
            6'd55: xpb[60] = 1024'd103439896114640452450023437065908141163818070536901094076342993552588865293414199275037266401524683429778511941652063585610260458971997687005081963953488496083756448732991335047907493875410795549160563935921022898673905027586156630506062855430092640474370836840647760243973266013788741696532401519347234885681;
            6'd56: xpb[60] = 1024'd1555748744547767870119305728534399980321532768774905425111678290109804925726813991661702592929622796967487199808561141882502709522467910595404076920802325413465274524495250275487793712967510683140408916832077261690510589721154904580918285430120603641655478291397998259592774643117316658515540964703051042162;
            6'd57: xpb[60] = 1024'd23738297058579824689014101795975091541523422126384400902012218092607639895348567618301209998992236473599611865422552132733808800914158468740886314904447195676864774885570382840698332742041431538430451506130371471071477002077049951620752285113378016075760023156265294305318811346374524637617370236684461682974;
            6'd58: xpb[60] = 1024'd45920845372611881507908897863415783102725311483993896378912757895105474864970321244940717405054850150231736531036543123585114892305849026886368552888092065940264275246645515405908871771115352393720494095428665680452443414432944998660586284796635428509864568021132590351044848049631732616719199508665872323786;
            6'd59: xpb[60] = 1024'd68103393686643938326803693930856474663927200841603391855813297697603309834592074871580224811117463826863861196650534114436420983697539585031850790871736936203663775607720647971119410800189273249010536684726959889833409826788840045700420284479892840943969112885999886396770884752888940595821028780647282964598;
            6'd60: xpb[60] = 1024'd90285942000675995145698489998297166225129090199212887332713837500101144804213828498219732217180077503495985862264525105287727075089230143177333028855381806467063275968795780536329949829263194104300579274025254099214376239144735092740254284163150253378073657750867182442496921456146148574922858052628693605410;
            6'd61: xpb[60] = 1024'd112468490314708051964593286065737857786330979556822382809614377302598979773835582124859239623242691180128110527878516096139033166480920701322815266839026676730462776329870913101540488858337114959590621863323548308595342651500630139780088283846407665812178202615734478488222958159403356554024687324610104246222;
            6'd62: xpb[60] = 1024'd10584342944615367384689154728364116602834441788696194158383062040119919406148196841483675814647630547317085786035013652411275417031390924913137379806340506060171602121374828329120788695893830093570466844234602671611948213635628413854943713846435628979462844066484716503842466788731931516007826769965920402703;
            6'd63: xpb[60] = 1024'd32766891258647424203583950795804808164036331146305689635283601842617754375769950468123183220710244223949210451649004643262581508423081483058619617789985376323571102482449960894331327724967750948860509433532896880992914625991523460894777713529693041413567388931352012549568503491989139495109656041947331043515;
        endcase
    end

    always_comb begin
        case(flag[20][11:6])
            6'd0: xpb[61] = 1024'd0;
            6'd1: xpb[61] = 1024'd54949439572679481022478746863245499725238220503915185112184141645115589345391704094762690626772857900581335117262995634113887599814772041204101855773630246586970602843525093459541866754041671804150552022831191090373881038347418507934611713212950453847671933796219308595294540195246347474211485313928741684327;
            6'd2: xpb[61] = 1024'd109898879145358962044957493726490999450476441007830370224368283290231178690783408189525381253545715801162670234525991268227775199629544082408203711547260493173941205687050186919083733508083343608301104045662382180747762076694837015869223426425900907695343867592438617190589080390492694948422970627857483368654;
            6'd3: xpb[61] = 1024'd40781623033913701668637313184922066431016234386009871208420569870369872698865973374273000665660899392300855944331493467762598958603095789057145442304559698827221133961004063040995361070607809691141458460106333424757282264821358750838856569955621912276195897974540867755777092511810409405515766115160630568650;
            6'd4: xpb[61] = 1024'd95731062606593182691116060048167566156254454889925056320604711515485462044257677469035691292433757292882191061594489101876486558417867830261247298078189945414191736804529156500537227824649481495292010482937524515131163303168777258773468283168572366123867831770760176351071632707056756879727251429089372252977;
            6'd5: xpb[61] = 1024'd26613806495147922314795879506598633136794248268104557304656998095624156052340242653783310704548940884020376771399991301411310317391419536910189028835489151067471665078483032622448855387173947578132364897381475759140683491295298993743101426698293370704719862152862426916259644828374471336820046916392519452973;
            6'd6: xpb[61] = 1024'd81563246067827403337274626369844132862032468772019742416841139740739745397731946748546001331321798784601711888662986935525197917206191578114290884609119397654442267922008126081990722141215619382282916920212666849514564529642717501677713139911243824552391795949081735511554185023620818811031532230321261137300;
            6'd7: xpb[61] = 1024'd12445989956382142960954445828275199842572262150199243400893426320878439405814511933293620743436982375739897598468489135060021676179743284763232615366418603307722196195962002203902349703740085465123271334656618093524084717769239236647346283440964829133243826331183986076742197144938533268124327717624408337296;
            6'd8: xpb[61] = 1024'd67395429529061623983433192691520699567810482654114428513077567965994028751206216028056311370209840276321232715731484769173909275994515325967334471140048849894692799039487095663444216457781757269273823357487809183897965756116657744581957996653915282980915760127403294672036737340184880742335813031553150021623;
            6'd9: xpb[61] = 1024'd122344869101741105005911939554766199293048703158029613625261709611109618096597920122819001996982698176902567832994480403287796875809287367171436326913679096481663401883012189122986083211823429073424375380319000274271846794464076252516569709866865736828587693923622603267331277535431228216547298345481891705950;
            6'd10: xpb[61] = 1024'd53227612990295844629591759013197266273588496536209114609313996191248312104680485307566621409097881768040753542799982602822620634782839073820378057670978302134943330156966065244897710774347895156264729794762951518281366982590597987486202853396586741409439724305724853832519289656748942673640093832785038905946;
            6'd11: xpb[61] = 1024'd108177052562975325652070505876442765998826717040124299721498137836363901450072189402329312035870739668622088660062978236936508234597611115024479913444608548721913933000491158704439577528389566960415281817594142608655248020938016495420814566609537195257111658101944162427813829851995290147851579146713780590273;
            6'd12: xpb[61] = 1024'd39059796451530065275750325334873832979366510418303800705550424416502595458154754587076931447985923259760274369868480436471331993571162821673421644201907754375193861274445034826351205090914033043255636232038093852664768209064538230390447710139258199837963688484046412993001841973313004604944374634016927790269;
            6'd13: xpb[61] = 1024'd94009236024209546298229072198119332704604730922218985817734566061618184803546458681839622074758781160341609487131476070585219593385934862877523499975538000962164464117970128285893071844955704847406188254869284943038649247411956738325059423352208653685635622280265721588296382168559352079155859947945669474596;
            6'd14: xpb[61] = 1024'd24891979912764285921908891656550399685144524300398486801786852641756878811629023866587241486873964751479795196936978270120043352359486569526465230732837206615444392391924004407804699407480170930246542669313236187048169435538478473294692566881929658266487652662367972153484394289877066536248655435248816674592;
            6'd15: xpb[61] = 1024'd79841419485443766944387638519795899410382744804313671913970994286872468157020727961349932113646822652061130314199973904233930952174258610730567086506467453202414995235449097867346566161521842734397094692144427277422050473885896981229304280094880112114159586458587280748778934485123414010460140749177558358919;
            6'd16: xpb[61] = 1024'd10724163373998506568067457978226966390922538182493172898023280867011162165103293146097551525762006243199316024005476103768754711147810317379508817263766658855694923509402973989258193724046308817237449106588378521431570662012418716198937423624601116695011616840689531313966946606441128467552936236480705558915;
            6'd17: xpb[61] = 1024'd65673602946677987590546204841472466116160758686408358010207422512126751510494997240860242152534864143780651141268471737882642310962582358583610673037396905442665526352928067448800060478087980621388001129419569611805451700359837224133549136837551570542683550636908839909261486801687475941764421550409447243242;
            6'd18: xpb[61] = 1024'd120623042519357468613024951704717965841398979190323543122391564157242340855886701335622932779307722044361986258531467371996529910777354399787712528811027152029636129196453160908341927232129652425538553152250760702179332738707255732068160850050502024390355484433128148504556026996933823415975906864338188927569;
            6'd19: xpb[61] = 1024'd51505786407912208236704771163149032821938772568503044106443850737381034863969266520370552191422905635500171968336969571531353669750906106436654259568326357682916057470407037030253554794654118508378907566694711946188852926833777467037793993580223028971207514815230399069744039118251537873068702351641336127565;
            6'd20: xpb[61] = 1024'd106455225980591689259183518026394532547176993072418229218627992382496624209360970615133242818195763536081507085599965205645241269565678147640756115341956604269886660313932130489795421548695790312529459589525903036562733965181195974972405706793173482818879448611449707665038579313497885347280187665570077811892;
            6'd21: xpb[61] = 1024'd37337969869146428882863337484825599527716786450597730202680278962635318217443535799880862230310947127219692795405467405180065028539229854289697846099255809923166588587886006611707049111220256395369814003969854280572254153307717709942038850322894487399731478993551958230226591434815599804372983152873225011888;
            6'd22: xpb[61] = 1024'd92287409441825909905342084348071099252955006954512915314864420607750907562835239894643552857083805027801027912668463039293952628354001895493799701872886056510137191431411100071248915865261928199520366026801045370946135191655136217876650563535844941247403412789771266825521131630061947278584468466801966696215;
            6'd23: xpb[61] = 1024'd23170153330380649529021903806502166233494800332692416298916707187889601570917805079391172269198988618939213622473965238828776387327553602142741432630185262163417119705364976193160543427786394282360720441244996614955655379781657952846283707065565945828255443171873517390709143751379661735677263954105113896211;
            6'd24: xpb[61] = 1024'd78119592903060130551500650669747665958733020836607601411100848833005190916309509174153862895971846519520548739736960872942663987142325643346843288403815508750387722548890069652702410181828066086511272464076187705329536418129076460780895420278516399675927376968092825986003683946626009209888749268033855580538;
            6'd25: xpb[61] = 1024'd9002336791614870175180470128178732939272814214787102395153135413143884924392074358901482308087030110658734449542463072477487746115877349995785019161114714403667650822843945774614037744352532169351626878520138949339056606255598195750528563808237404256779407350195076551191696067943723666981544755337002780534;
            6'd26: xpb[61] = 1024'd63951776364294351197659216991424232664511034718702287507337277058259474269783778453664172934859888011240069566805458706591375345930649391199886874934744960990638253666369039234155904498394203973502178901351330039712937644603016703685140277021187858104451341146414385146486236263190071141193030069265744464861;
            6'd27: xpb[61] = 1024'd118901215936973832220137963854669732389749255222617472619521418703375063615175482548426863561632745911821404684068454340705262945745421432403988730708375207577608856509894132693697771252435875777652730924182521130086818682950435211619751990234138311952123274942633693741780776458436418615404515383194486149188;
            6'd28: xpb[61] = 1024'd49783959825528571843817783313100799370289048600796973603573705283513757623258047733174482973747929502959590393873956540240086704718973139052930461465674413230888784783848008815609398814960341860493085338626472374096338871076956946589385133763859316532975305324735944306968788579754133072497310870497633349184;
            6'd29: xpb[61] = 1024'd104733399398208052866296530176346299095527269104712158715757846928629346968649751827937173600520787403540925511136952174353974304533745180257032317239304659817859387627373102275151265569002013664643637361457663464470219909424375454523996846976809770380647239120955252902263328775000480546708796184426375033511;
            6'd30: xpb[61] = 1024'd35616143286762792489976349634777366076067062482891659699810133508768040976732317012684793012635970994679111220942454373888798063507296886905974047996603865471139315901326978397062893131526479747483991775901614708479740097550897189493629990506530774961499269503057503467451340896318195003801591671729522233507;
            6'd31: xpb[61] = 1024'd90565582859442273512455096498022865801305282986806844811994275153883630322124021107447483639408828895260446338205450008002685663322068928110075903770234112058109918744852071856604759885568151551634543798732805798853621135898315697428241703719481228809171203299276812062745881091564542478013076985658263917834;
            6'd32: xpb[61] = 1024'd21448326747997013136134915956453932781845076364986345796046561734022324330206586292195103051524012486398632048010952207537509422295620634759017634527533317711389847018805947978516387448092617634474898213176757042863141324024837432397874847249202233390023233681379062627933893212882256935105872472961411117830;
            6'd33: xpb[61] = 1024'd76397766320676494158613662819699432507083296868901530908230703379137913675598290386957793678296870386979967165273947841651397022110392675963119490301163564298360449862331041438058254202134289438625450236007948133237022362372255940332486560462152687237695167477598371223228433408128604409317357786890152802157;
            6'd34: xpb[61] = 1024'd7280510209231233782293482278130499487623090247081031892282989959276607683680855571705413090412053978118152875079450041186220781083944382612061221058462769951640378136284917559969881764658755521465804650451899377246542550498777675302119703991873691818547197859700621788416445529446318866410153274193300002153;
            6'd35: xpb[61] = 1024'd62229949781910714804772229141375999212861310750996217004467131604392197029072559666468103717184911878699487992342445675300108380898716423816163076832093016538610980979810011019511748518700427325616356673283090467620423588846196183236731417204824145666219131655919930383710985724692666340621638588122041686480;
            6'd36: xpb[61] = 1024'd117179389354590195827250976004621498938099531254911402116651273249507786374464263761230794343957769779280823109605441309413995980713488465020264932605723263125581583823335104479053615272742099129766908696114281557994304627193614691171343130417774599513891065452139238979005525919939013814833123902050783370807;
            6'd37: xpb[61] = 1024'd48062133243144935450930795463052565918639324633090903100703559829646480382546828945978413756072953370419008819410943508948819739687040171669206663363022468778861512097288980600965242835266565212607263110558232802003824815320136426140976273947495604094743095834241489544193538041256728271925919389353930570803;
            6'd38: xpb[61] = 1024'd103011572815824416473409542326298065643877545137006088212887701474762069727938533040741104382845811271000343936673939143062707339501812212873308519136652715365832114940814074060507109589308237016757815133389423892377705853667554934075587987160446057942415029630460798139488078236503075746137404703282672255130;
            6'd39: xpb[61] = 1024'd33894316704379156097089361784729132624417338515185589196939988054900763736021098225488723794960994862138529646479441342597531098475363919522250249893951921019112043214767950182418737151832703099598169547833375136387226041794076669045221130690167062523267060012563048704676090357820790203230200190585819455126;
            6'd40: xpb[61] = 1024'd88843756277058637119568108647974632349655559019100774309124129700016353081412802320251414421733852762719864763742436976711418698290135960726352105667582167606082646058293043641960603905874374903748721570664566226761107080141495176979832843903117516370938993808782357299970630553067137677441685504514561139453;
            6'd41: xpb[61] = 1024'd19726500165613376743247928106405699330195352397280275293176416280155047089495367504999033833849036353858050473547939176246242457263687667375293836424881373259362574332246919763872231468398840986589075985108517470770627268268016911949465987432838520951791024190884607865158642674384852134534480991817708339449;
            6'd42: xpb[61] = 1024'd74675939738292857765726674969651199055433572901195460405360557925270636434887071599761724460621894254439385590810934810360130057078459708579395692198511619846333177175772013223414098222440512790739628007939708561144508306615435419884077700645788974799462957987103916460453182869631199608745966305746450023776;
            6'd43: xpb[61] = 1024'd5558683626847597389406494428082266035973366279374961389412844505409330442969636784509343872737077845577571300616437009894953816052011415228337422955810825499613105449725889345325725784964978873579982422383659805154028494741957154853710844175509979380314988369206167025641194990948914065838761793049597223772;
            6'd44: xpb[61] = 1024'd60508123199527078411885241291327765761211586783290146501596986150524919788361340879272034499509935746158906417879432644008841415866783456432439278729441072086583708293250982804867592539006650677730534445214850895527909533089375662788322557388460433227986922165425475620935735186195261540050247106978338908099;
            6'd45: xpb[61] = 1024'd115457562772206559434363988154573265486449807287205331613781127795640509133753044974034725126282793646740241535142428278122729015681555497636541134503071318673554311136776076264409459293048322481881086468046041985901790571436794170722934270601410887075658855961644784216230275381441609014261732420907080592426;
            6'd46: xpb[61] = 1024'd46340306660761299058043807613004332466989600665384832597833414375779203141835610158782344538397977237878427244947930477657552774655107204285482865260370524326834239410729952386321086855572788564721440882489993229911310759563315905692567414131131891656510886343747034781418287502759323471354527908210227792422;
            6'd47: xpb[61] = 1024'd101289746233440780080522554476249832192227821169300017710017556020894792487227314253545035165170835138459762362210926111771440374469879245489584721034000770913804842254255045845862953609614460368871992905321184320285191797910734413627179127344082345504182820139966343376712827698005670945566013222138969476749;
            6'd48: xpb[61] = 1024'd32172490121995519704202373934680899172767614547479518694069842601033486495309879438292654577286018729597948072016428311306264133443430952138526451791299976567084770528208921967774581172138926451712347319765135564294711986037256148596812270873803350085034850522068593941900839819323385402658808709442116676745;
            6'd49: xpb[61] = 1024'd87121929694675000726681120797926398898005835051394703806253984246149075840701583533055345204058876630179283189279423945420151733258202993342628307564930223154055373371734015427316447926180598255862899342596326654668593024384674656531423984086753803932706784318287902537195380014569732876870294023370858361072;
            6'd50: xpb[61] = 1024'd18004673583229740350360940256357465878545628429574204790306270826287769848784148717802964616174060221317468899084926144954975492231754699991570038322229428807335301645687891549228075488705064338703253757040277898678113212511196391501057127616474808513558814700390153102383392135887447333963089510674005561068;
            6'd51: xpb[61] = 1024'd72954113155909221372839687119602965603783848933489389902490412471403359194175852812565655242946918121898804016347921779068863092046526741195671894095859675394305904489212985008769942242746736142853805779871468989051994250858614899435668840829425262361230748496609461697677932331133794808174574824602747245395;
            6'd52: xpb[61] = 1024'd3836857044463960996519506578034032584323642311668890886542699051542053202258417997313274655062101713036989726153423978603686851020078447844613624853158881047585832763166861130681569805271202225694160194315420233061514438985136634405301984359146266942082778878711712262865944452451509265267370311905894445391;
            6'd53: xpb[61] = 1024'd58786296617143442018998253441279532309561862815584075998726840696657642547650122092075965281834959613618324843416419612717574450834850489048715480626789127634556435606691954590223436559312874029844712217146611323435395477332555142339913697572096720789754712674931020858160484647697856739478855625834636129718;
            6'd54: xpb[61] = 1024'd113735736189822923041477000304525032034800083319499261110910982341773231893041826186838655908607817514199659960679415246831462050649622530252817336400419374221527038450217048049765303313354545833995264239977802413809276515679973650274525410785047174637426646471150329453455024842944204213690340939763377814045;
            6'd55: xpb[61] = 1024'd44618480078377662665156819762956099015339876697678762094963268921911925901124391371586275320723001105337845670484917446366285809623174236901759067157718579874806966724170924171676930875879011916835618654421753657818796703806495385244158554314768179218278676853252580018643036964261918670783136427066525014041;
            6'd56: xpb[61] = 1024'd99567919651057143687635566626201598740578097201593947207147410567027515246516095466348965947495859005919180787747913080480173409437946278105860922931348826461777569567696017631218797629920683720986170677252944748192677742153913893178770267527718633065950610649471888613937577159508266144994621740995266698368;
            6'd57: xpb[61] = 1024'd30450663539611883311315386084632665721117890579773448191199697147166209254598660651096585359611042597057366497553415280014997168411497984754802653688648032115057497841649893753130425192445149803826525091696895992202197930280435628148403411057439637646802641031574139179125589280825980602087417228298413898364;
            6'd58: xpb[61] = 1024'd85400103112291364333794132947878165446356111083688633303383838792281798599990364745859275986383900497638701614816410914128884768226270025958904509462278278702028100685174987212672291946486821607977077114528087082576078968627854136083015124270390091494474574827793447774420129476072328076298902542227155582691;
            6'd59: xpb[61] = 1024'd16282847000846103957473952406309232426895904461868134287436125372420492608072929930606895398499084088776887324621913113663708527199821732607846240219577484355308028959128863334583919509011287690817431528972038326585599156754375871052648267800111096075326605209895698339608141597390042533391698029530302782687;
            6'd60: xpb[61] = 1024'd71232286573525584979952699269554732152134124965783319399620267017536081953464634025369586025271941989358222441884908747777596127014593773811948095993207730942278631802653956794125786263052959494967983551803229416959480195101794378987259981013061549922998539006115006934902681792636390007603183343459044467014;
            6'd61: xpb[61] = 1024'd2115030462080324603632518727985799132673918343962820383672553597674775961547199210117205437387125580496408151690410947312419885988145480460889826750506936595558560076607832916037413825577425577808337966247180660969000383228316113956893124542782554503850569388217257500090693913954104464695978830762191667010;
            6'd62: xpb[61] = 1024'd57064470034759805626111265591231298857912138847878005495856695242790365306938903304879896064159983481077743268953406581426307485802917521664991682524137183182529162920132926375579280579619097381958889989078371751342881421575734621891504837755733008351522503184436566095385234109200451938907464144690933351337;
            6'd63: xpb[61] = 1024'd112013909607439286648590012454476798583150359351793190608040836887905954652330607399642586690932841381659078386216402215540195085617689562869093538297767429769499765763658019835121147333660769186109442011909562841716762459923153129826116550968683462199194436980655874690679774304446799413118949458619675035664;
        endcase
    end

    always_comb begin
        case(flag[20][16:12])
            5'd0: xpb[62] = 1024'd0;
            5'd1: xpb[62] = 1024'd42896653495994026272269831912907865563690152729972691592093123468044648660413172584390206103048024972797264096021904415075018844591241269518035269055066635422779694037611895957032774896185235268949796426353514085726282648049674864795749694498404466780046467362758125255867786425764513870211744945922822235660;
            5'd2: xpb[62] = 1024'd85793306991988052544539663825815731127380305459945383184186246936089297320826345168780412206096049945594528192043808830150037689182482539036070538110133270845559388075223791914065549792370470537899592852707028171452565296099349729591499388996808933560092934725516250511735572851529027740423489891845644471320;
            5'd3: xpb[62] = 1024'd4623264803857337418010568333909163946372031064182390648147515339157050643930378843155547094486400608948642880608219810645992692932503473998945682148868865334648407543264470533468085497038500085539191670673302410814487093928127821422270513811983951073319498674157317737496831203364908593516545011142872222649;
            5'd4: xpb[62] = 1024'd47519918299851363690280400246817029510062183794155082240240638807201699304343551427545753197534425581745906976630124225721011537523744743516980951203935500757428101580876366490500860393223735354488988097026816496540769741977802686218020208310388417853365966036915442993364617629129422463728289957065694458309;
            5'd5: xpb[62] = 1024'd90416571795845389962550232159724895073752336524127773832333762275246347964756724011935959300582450554543171072652028640796030382114986013035016220259002136180207795618488262447533635289408970623438784523380330582267052390027477551013769902808792884633412433399673568249232404054893936333940034902988516693969;
            5'd6: xpb[62] = 1024'd9246529607714674836021136667818327892744062128364781296295030678314101287860757686311094188972801217897285761216439621291985385865006947997891364297737730669296815086528941066936170994077000171078383341346604821628974187856255642844541027623967902146638997348314635474993662406729817187033090022285744445298;
            5'd7: xpb[62] = 1024'd52143183103708701108290968580726193456434214858337472888388154146358749948273930270701300292020826190694549857238344036367004230456248217515926633352804366092076509124140837023968945890262235440028179767700118907355256835905930507640290722122372368926685464711072760730861448832494331057244834968208566680958;
            5'd8: xpb[62] = 1024'd95039836599702727380560800493634059020124367588310164480481277614403398608687102855091506395068851163491813953260248451442023075047489487033961902407871001514856203161752732981001720786447470708977976194053632993081539483955605372436040416620776835706731932073830885986729235258258844927456579914131388916618;
            5'd9: xpb[62] = 1024'd13869794411572012254031705001727491839116093192547171944442546017471151931791136529466641283459201826845928641824659431937978078797510421996837046446606596003945222629793411600404256491115500256617575012019907232443461281784383464266811541435951853219958496022471953212490493610094725780549635033428616667947;
            5'd10: xpb[62] = 1024'd56766447907566038526301536914635357402806245922519863536535669485515800592204309113856847386507226799643192737846563847012996923388751691514872315501673231426724916667405307557437031387300735525567371438373421318169743929834058329062561235934356320000004963385230078468358280035859239650761379979351438903607;
            5'd11: xpb[62] = 1024'd99663101403560064798571368827543222966496398652492555128628792953560449252617481698247053489555251772440456833868468262088015767979992961032907584556739866849504610705017203514469806283485970794517167864726935403896026577883733193858310930432760786780051430747988203724226066461623753520973124925274261139267;
            5'd12: xpb[62] = 1024'd18493059215429349672042273335636655785488124256729562592590061356628202575721515372622188377945602435794571522432879242583970771730013895995782728595475461338593630173057882133872341988154000342156766682693209643257948375712511285689082055247935804293277994696629270949987324813459634374066180044571488890596;
            5'd13: xpb[62] = 1024'd61389712711423375944312105248544521349178276986702254184683184824672851236134687957012394480993627408591835618454783657658989616321255165513817997650542096761373324210669778090905116884339235611106563109046723728984231023762186150484831749746340271073324462059387396205855111239224148244277924990494311126256;
            5'd14: xpb[62] = 1024'd104286366207417402216581937161452386912868429716674945776776308292717499896547860541402600584041652381389099714476688072734008460912496435031853266705608732184153018248281674047937891780524470880056359535400237814710513671811861015280581444244744737853370929422145521461722897664988662114489669936417133361916;
            5'd15: xpb[62] = 1024'd23116324019286687090052841669545819731860155320911953240737576695785253219651894215777735472432003044743214403041099053229963464662517369994728410744344326673242037716322352667340427485192500427695958353366512054072435469640639107111352569059919755366597493370786588687484156016824542967582725055714361113245;
            5'd16: xpb[62] = 1024'd66012977515280713362322673582453685295550308050884644832830700163829901880065066800167941575480028017540478499063003468304982309253758639512763679799410962096021731753934248624373202381377735696645754779720026139798718117690313971907102263558324222146643960733544713943351942442589056837794470001637183348905;
            5'd17: xpb[62] = 1024'd108909631011274739634592505495361550859240460780857336424923823631874550540478239384558147678528052990337742595084907883380001153844999909030798948854477597518801425791546144581405977277562970965595551206073540225525000765739988836702851958056728688926690428096302839199219728868353570708006214947560005584565;
            5'd18: xpb[62] = 1024'd27739588823144024508063410003454983678232186385094343888885092034942303863582273058933282566918403653691857283649318863875956157595020843993674092893213192007890445259586823200808512982231000513235150024039814464886922563568766928533623082871903706439916992044943906424980987220189451561099270066857233335894;
            5'd19: xpb[62] = 1024'd70636242319138050780333241916362849241922339115067035480978215502986952523995445643323488669966428626489121379671223278950975002186262113511709361948279827430670139297198719157841287878416235782184946450393328550613205211618441793329372777370308173219963459407702031680848773645953965431311015012780055571554;
            5'd20: xpb[62] = 1024'd113532895815132077052603073829270714805612491845039727073071338971031601184408618227713694773014453599286385475693127694025993846777503383029744631003346462853449833334810615114874062774601471051134742876746842636339487859668116658125122471868712640000009926770460156936716560071718479301522759958702877807214;
            5'd21: xpb[62] = 1024'd32362853627001361926073978337364147624604217449276734537032607374099354507512651902088829661404804262640500164257538674521948850527524317992619775042082057342538852802851293734276598479269500598774341694713116875701409657496894749955893596683887657513236490719101224162477818423554360154615815078000105558543;
            5'd22: xpb[62] = 1024'd75259507122995388198343810250272013188294370179249426129125730842144003167925824486479035764452829235437764260279443089596967695118765587510655044097148692765318546840463189691309373375454735867724138121066630961427692305546569614751643291182292124293282958081859349418345604849318874024827560023922927794203;
            5'd23: xpb[62] = 1024'd118156160618989414470613642163179878751984522909222117721218854310188651828338997070869241867500854208235028356301347504671986539710006857028690313152215328188098240878075085648342148271639971136673934547420145047153974953596244479547392985680696591073329425444617474674213391275083387895039304969845750029863;
            5'd24: xpb[62] = 1024'd36986118430858699344084546671273311570976248513459125185180122713256405151443030745244376755891204871589143044865758485167941543460027791991565457190950922677187260346115764267744683976308000684313533365386419286515896751425022571378164110495871608586555989393258541899974649626919268748132360089142977781192;
            5'd25: xpb[62] = 1024'd79882771926852725616354378584181177134666401243431816777273246181301053811856203329634582858939229844386407140887662900242960388051269061509600726246017558099966954383727660224777458872493235953263329791739933372242179399474697436173913804994276075366602456756016667155842436052683782618344105035065800016852;
            5'd26: xpb[62] = 1024'd122779425422846751888624210497089042698356553973404508369366369649345702472269375914024788961987254817183671236909567315317979232642510331027635995301084193522746648421339556181810233768678471222213126218093447457968462047524372300969663499492680542146648924118774792411710222478448296488555849980988622252512;
            5'd27: xpb[62] = 1024'd41609383234716036762095115005182475517348279577641515833327638052413455795373409588399923850377605480537785925473978295813934236392531265990511139339819788011835667889380234801212769473346500769852725036059721697330383845353150392800434624307855559659875488067415859637471480830284177341648905100285850003841;
            5'd28: xpb[62] = 1024'd84506036730710063034364946918090341081038432307614207425420761520458104455786582172790129953425630453335050021495882710888953080983772535508546408394886423434615361926992130758245544369531736038802521462413235783056666493402825257596184318806260026439921955430173984893339267256048691211860650046208672239501;
            5'd29: xpb[62] = 1024'd3335994542579347907835851426183773900030157911851214889382029923525857778890615847165264841815981116689164710060293691384908084733793470471421552433622017923704381395032809377648080074199765586442120280379510022418588291231603349426955443621435043953148519378815052119100525607884572064953705165505899990830;
            5'd30: xpb[62] = 1024'd46232648038573374180105683339091639463720310641823906481475153391570506439303788431555470944864006089486428806082198106459926929325034739989456821488688653346484075432644705334680854970385000855391916706733024108144870939281278214222705138119839510733194986741573177374968312033649085935165450111428722226490;
            5'd31: xpb[62] = 1024'd89129301534567400452375515251999505027410463371796598073568276859615155099716961015945677047912031062283692902104102521534945773916276009507492090543755288769263769470256601291713629866570236124341713133086538193871153587330953079018454832618243977513241454104331302630836098459413599805377195057351544462150;
        endcase
    end

    always_comb begin
        case(flag[21][5:0])
            6'd0: xpb[63] = 1024'd0;
            6'd1: xpb[63] = 1024'd66012977515280713362322673582453685295550308050884644832830700163829901880065066800167941575480028017540478499063003468304982309253758639512763679799410962096021731753934248624373202381377735696645754779720026139798718117690313971907102263558324222146643960733544713943351942442589056837794470001637183348905;
            6'd2: xpb[63] = 1024'd7959259346436685325846419760092937846402188976033605537529545262682908422820994690320811936302381725637807590668513502030900777666296944470367234582490883258352788938297279911116165571238265671981311951052812433233075385159731170849225957433418995026468018052972369856597356811249480658470250176648772213479;
            6'd3: xpb[63] = 1024'd73972236861717398688169093342546623141952497026918250370360245426512810302886061490488753511782409743178286089731516970335883086920055583983130914381901845354374520692231528535489367952616001368627066730772838573031793502850045142756328220991743217173111978786517083799949299253838537496264720178285955562384;
            6'd4: xpb[63] = 1024'd15918518692873370651692839520185875692804377952067211075059090525365816845641989380641623872604763451275615181337027004061801555332593888940734469164981766516705577876594559822232331142476531343962623902105624866466150770319462341698451914866837990052936036105944739713194713622498961316940500353297544426958;
            6'd5: xpb[63] = 1024'd81931496208154084014015513102639560988354686002951855907889790689195718725707056180809565448084791468816093680400030472366783864586352528453498148964392728612727309630528808446605533523854267040608378681825651006264868888009776313605554178425162212199579996839489453656546656065088018154734970354934727775863;
            6'd6: xpb[63] = 1024'd23877778039310055977539259280278813539206566928100816612588635788048725268462984070962435808907145176913422772005540506092702332998890833411101703747472649775058366814891839733348496713714797015943935853158437299699226155479193512547677872300256985079404054158917109569792070433748441975410750529946316640437;
            6'd7: xpb[63] = 1024'd89890755554590769339861932862732498834756874978985461445419335951878627148528050871130377384387173194453901271068543974397684642252649472923865383546883611871080098568826088357721699095092532712589690632878463439497944273169507484454780135858581207226048014892461823513144012876337498813205220531583499989342;
            6'd8: xpb[63] = 1024'd31837037385746741303385679040371751385608755904134422150118181050731633691283978761283247745209526902551230362674054008123603110665187777881468938329963533033411155753189119644464662284953062687925247804211249732932301540638924683396903829733675980105872072211889479426389427244997922633881000706595088853916;
            6'd9: xpb[63] = 1024'd97850014901027454665708352622825436681159063955019066982948881214561535571349045561451189320689554920091708861737057476428585419918946417394232618129374495129432887507123368268837864666330798384571002583931275872731019658329238655304006093292000202252516032945434193369741369687586979471675470708232272202821;
            6'd10: xpb[63] = 1024'd39796296732183426629232098800464689232010944880168027687647726313414542114104973451604059681511908628189037953342567510154503888331484722351836172912454416291763944691486399555580827856191328359906559755264062166165376925798655854246129787167094975132340090264861849282986784056247403292351250883243861067395;
            6'd11: xpb[63] = 1024'd105809274247464139991554772382918374527561252931052672520478426477244443994170040251772001256991936645729516452405570978459486197585243361864599852711865378387785676445420648179954030237569064056552314534984088305964095043488969826153232050725419197278984050998406563226338726498836460130145720884881044416300;
            6'd12: xpb[63] = 1024'd47755556078620111955078518560557627078413133856201633225177271576097450536925968141924871617814290353826845544011081012185404665997781666822203407494945299550116733629783679466696993427429594031887871706316874599398452310958387025095355744600513970158808108317834219139584140867496883950821501059892633280874;
            6'd13: xpb[63] = 1024'd113768533593900825317401192143011312373963441907086278058007971739927352416991034942092813193294318371367324043074084480490386975251540306334967087294356261646138465383717928091070195808807329728533626486036900739197170428648700997002458008158838192305452069051378933082936083310085940788615971061529816629779;
            6'd14: xpb[63] = 1024'd55714815425056797280924938320650564924815322832235238762706816838780358959746962832245683554116672079464653134679594514216305443664078611292570642077436182808469522568080959377813158998667859703869183657369687032631527696118118195944581702033932965185276126370806588996181497678746364609291751236541405494353;
            6'd15: xpb[63] = 1024'd121727792940337510643247611903104250220365630883119883595537517002610260839812029632413625129596700097005131633742597982521287752917837250805334321876847144904491254322015208002186361380045595400514938437089713172430245813808432167851683965592257187331920087104351302939533440121335421447086221238178588843258;
            6'd16: xpb[63] = 1024'd63674074771493482606771358080743502771217511808268844300236362101463267382567957522566495490419053805102460725348108016247206221330375555762937876659927066066822311506378239288929324569906125375850495608422499465864603081277849366793807659467351960211744144423778958852778854489995845267762001413190177707832;
            6'd17: xpb[63] = 1024'd5620356602649454570295104258382755322069392733417805004935207200316273925323885412719365851241407513199789816953618049973124689742913860720541431443006987229153368690741270575672287759766655351186052779755285759298960348747266565735931353342446733091568201743206614766024268858656269088437781588201766572406;
            6'd18: xpb[63] = 1024'd71633334117930167932617777840836440617619700784302449837765907364146175805388952212887307426721435530740268316016621518278106998996672500233305111242417949325175100444675519200045490141144391047831807559475311899097678466437580537643033616900770955238212162476751328709376211301245325926232251589838949921311;
            6'd19: xpb[63] = 1024'd13579615949086139896141524018475693168471581709451410542464752462999182348144880103040177787543789238837597407622131552004025467409210805190908666025497870487506157629038550486788453331004921023167364730808098192532035733906997736585157310775865728118036219796178984622621625669905749746908031764850538785885;
            6'd20: xpb[63] = 1024'd79592593464366853258464197600929378464021889760336055375295452626829084228209946903208119363023817256378075906685135020309007776662969444703672345824908832583527889382972799111161655712382656719813119510528124332330753851597311708492259574334189950264680180529723698565973568112494806584702501766487722134790;
            6'd21: xpb[63] = 1024'd21538875295522825221987943778568631014873770685485016079994297725682090770965874793360989723846170964475404998290645054034926245075507749661275900607988753745858946567335830397904618902243186695148676681860910625765111119066728907434383268209284723144504237849151354479218982481155230405378281941499310999364;
            6'd22: xpb[63] = 1024'd87551852810803538584310617361022316310424078736369660912824997889511992651030941593528931299326198982015883497353648522339908554329266389174039580407399715841880678321270079022277821283620922391794431461580936765563829236757042879341485531767608945291148198582696068422570924923744287243172751943136494348269;
            6'd23: xpb[63] = 1024'd29498134641959510547834363538661568861275959661518621617523842988364999193786869483681801660148552690113212588959158556065827022741804694131643135190479637004211735505633110309020784473481452367129988632913723058998186504226460078283609225642703718170972255902123724335816339292404711063848532118148083212843;
            6'd24: xpb[63] = 1024'd95511112157240223910157037121115254156826267712403266450354543152194901073851936283849743235628580707653691088022162024370809331995563333644406814989890599100233467259567358933393986854859188063775743412633749198796904621916774050190711489201027940317616216635668438279168281734993767901643002119785266561748;
            6'd25: xpb[63] = 1024'd37457393988396195873680783298754506707678148637552227155053388251047907616607864174002613596450934415751020179627672058096727800408101638602010369772970520262564524443930390220136950044719718039111300583966535492231261889386191249132835183076122713197440273955096094192413696103654191722318782294796855426322;
            6'd26: xpb[63] = 1024'd103470371503676909236003456881208192003228456688436871987884088414877809496672930974170555171930962433291498678690675526401710109661860278114774049572381482358586256197864638844510152426097453735757055363686561632029980007076505221039937446634446935344084234688640808135765638546243248560113252296434038775227;
            6'd27: xpb[63] = 1024'd45416653334832881199527203058847444554080337613585832692582933513730816039428858864323425532753316141388827770296185560127628578074398583072377604355461403520917313382227670131253115615957983711092612535019347925464337274545922419982061140509541708223908292008068464049011052914903672380789032471445627639801;
            6'd28: xpb[63] = 1024'd111429630850113594561849876641301129849630645664470477525413633677560717919493925664491367108233344158929306269359189028432610887328157222585141284154872365616939045136161918755626317997335719407738367314739374065263055392236236391889163404067865930370552252741613177992362995357492729218583502473082810988706;
            6'd29: xpb[63] = 1024'd53375912681269566525373622818940382400482526589619438230112478776413724462249853554644237469055697867026635360964699062158529355740695527542744838937952286779270102320524950042369281187196249383073924486072160358697412659705653590831287097942960703250376310061040833905608409726153153039259282648094399853280;
            6'd30: xpb[63] = 1024'd119388890196550279887696296401394067696032834640504083062943178940243626342314920354812179044535725884567113860027702530463511664994454167055508518737363248875291834074459198666742483568573985079719679265792186498496130777395967562738389361501284925397020270794585547848960352168742209877053752649731583202185;
            6'd31: xpb[63] = 1024'd61335172027706251851220042579033320246884715565653043767642024039096632885070848244965049405358079592664442951633212564189430133406992472013112073520443170037622891258822229953485446758434515055055236437124972791930488044865384761680513055376379698276844328114013203762205766537402633697729532824743172066759;
            6'd32: xpb[63] = 1024'd3281453858862223814743788756672572797736596490802004472340869137949639427826776135117919766180433300761772043238722597915348601819530776970715628303523091199953948443185261240228409948295045030390793608457759085364845312334801960622636749251474471156668385433440859675451180906063057518405312999754760931333;
            6'd33: xpb[63] = 1024'd69294431374142937177066462339126258093286904541686649305171569301779541307891842935285861341660461318302250542301726066220330911073289416483479308102934053295975680197119509864601612329672780727036548388177785225163563430025115932529739012809798693303312346166985573618803123348652114356199783001391944280238;
            6'd34: xpb[63] = 1024'd11240713205298909140590208516765510644138785466835610009870414400632547850647770825438731702482815026399579633907236099946249379485827721441082862886013974458306737381482541151344575519533310702372105559510571518597920697494533131471862706684893466183136403486413229532048537717312538176875563176403533144812;
            6'd35: xpb[63] = 1024'd77253690720579622502912882099219195939689093517720254842701114564462449730712837625606673277962843043940058132970239568251231688739586360953846542685424936554328469135416789775717777900911046399017860339230597658396638815184847103378964970243217688329780364219957943475400480159901595014670033178040716493717;
            6'd36: xpb[63] = 1024'd19199972551735594466436628276858448490540974442869215547399959663315456273468765515759543638785196752037387224575749601977150157152124665911450097468504857716659526319779821062460741090771576374353417510563383951830996082654264302321088664118312461209604421539385599388645894528562018835345813353052305358291;
            6'd37: xpb[63] = 1024'd85212950067016307828759301859312133786091282493753860380230659827145358153533832315927485214265224769577865723638753070282132466405883305424213777267915819812681258073714069686833943472149312070999172290283410091629714200344578274228190927676636683356248382272930313331997836971151075673140283354689488707196;
            6'd38: xpb[63] = 1024'd27159231898172279792283048036951386336943163418902821084929504925998364696289760206080355575087578477675194815244263104008050934818421610381817332050995740975012315258077100973576906662009842046334729461616196385064071467813995473170314621551731456236072439592357969245243251339811499493816063529701077571770;
            6'd39: xpb[63] = 1024'd93172209413452993154605721619405071632493471469787465917760205089828266576354827006248297150567606495215673314307266572313033244072180249894581011850406703071034047012011349597950109043387577742980484241336222524862789585504309445077416885110055678382716400325902683188595193782400556331610533531338260920675;
            6'd40: xpb[63] = 1024'd35118491244608965118129467797044324183345352394936426622459050188681273119110754896401167511389960203313002405912776606038951712484718554852184566633486624233365104196374380884693072233248107718316041412669008818297146852973726644019540578985150451262540457645330339101840608151060980152286313706349849785249;
            6'd41: xpb[63] = 1024'd101131468759889678480452141379498009478895660445821071455289750352511174999175821696569109086869988220853480904975780074343934021738477194364948246432897586329386835950308629509066274614625843414961796192389034958095864970664040615926642842543474673409184418378875053045192550593650036990080783707987033134154;
            6'd42: xpb[63] = 1024'd43077750591045650443975887557137262029747541370970032159988595451364181541931749586721979447692341928950809996581290108069852490151015499322551801215977507491717893134671660795809237804486373390297353363721821251530222238133457814868766536418569446289008475698302708958437964962310460810756563882998621998728;
            6'd43: xpb[63] = 1024'd109090728106326363806298561139590947325297849421854676992819295615194083421996816386889921023172369946491288495644293576374834799404774138835315481015388469587739624888605909420182440185864109086943108143441847391328940355823771786775868799976893668435652436431847422901789907404899517648551033884635805347633;
            6'd44: xpb[63] = 1024'd51037009937482335769822307317230199876149730347003637697518140714047089964752744277042791383994723654588617587249803610100753267817312443792919035798468390750070682072968940706925403375724639062278665314774633684763297623293188985717992493851988441315476493751275078815035321773559941469226814059647394212207;
            6'd45: xpb[63] = 1024'd117049987452763049132144980899683885171700038397888282530348840877876991844817811077210732959474751672129096086312807078405735577071071083305682715597879352846092413826903189331298605757102374758924420094494659824562015740983502957625094757410312663462120454484819792758387264216148998307021284061284577561112;
            6'd46: xpb[63] = 1024'd58996269283919021095668727077323137722551919323037243235047685976729998387573738967363603320297105380226425177918317112131654045483609388263286270380959274008423471011266220618041568946962904734259977265827446117996373008452920156567218451285407436341944511804247448671632678584809422127697064236296166425686;
            6'd47: xpb[63] = 1024'd942551115074993059192473254962390273403800248186203939746531075583004930329666857516473681119459088323754269523827145857572513896147693220889825164039195170754528195629251904784532136823434709595534437160232411430730275922337355509342145160502209221768569123675104584878092953469845948372844411307755290260;
            6'd48: xpb[63] = 1024'd66955528630355706421515146837416075568954108299070848772577231239412906810394733657684415256599487105864232768586830614162554823149906332733653504963450157266776259949563500529157734518201170406241289216880258551229448393612651327416444408718826431368412529857219818528230035396058902786167314412944938639165;
            6'd49: xpb[63] = 1024'd8901810461511678385038893015055328119805989224219809477276076338265913353150661547837285617421840813961561860192340647888473291562444637691257059746530078429107317133926531815900697708061700381576846388213044844663805661082068526358568102593921204248236587176647474441475449764719326606843094587956527503739;
            6'd50: xpb[63] = 1024'd74914787976792391747361566597509013415356297275104454310106776502095815233215728348005227192901868831502040359255344116193455600816203277204020739545941040525129048887860780440273900089439436078222601167933070984462523778772382498265670366152245426394880547910192188384827392207308383444637564589593710852644;
            6'd51: xpb[63] = 1024'd16861069807948363710885312775148265966208178200253415014805621600948821775971656238158097553724222539599369450860854149919374069228741582161624294329020961687460106072223811727016863279299966053558158339265857277896881046241799697207794060027340199274704605229619844298072806575968807265313344764605299717218;
            6'd52: xpb[63] = 1024'd82874047323229077073207986357601951261758486251138059847636321764778723656036723038326039129204250557139847949923857618224356378482500221674387974128431923783481837826158060351390065660677701750203913118985883417695599163932113669114896323585664421421348565963164558241424749018557864103107814766242483066123;
            6'd53: xpb[63] = 1024'd24820329154385049036731732535241203812610367176287020552335166863631730198792650928478909490026604265237177041529367651950274846895038526631991528911511844945812895010521091638133028850538231725539470290318669711129956431401530868057020017460759194301172623282592214154670163387218287923783594941254071930697;
            6'd54: xpb[63] = 1024'd90833306669665762399054406117694889108160675227171665385165867027461632078857717728646851065506632282777655540592371120255257156148797166144755208710922807041834626764455340262506231231915967422185225070038695850928674549091844839964122281019083416447816584016136928098022105829807344761578064942891255279602;
            6'd55: xpb[63] = 1024'd32779588500821734362578152295334141659012556152320626089864712126314638621613645618799721426328985990874984632197881153981175624561335471102358763494002728204165683948818371549249194421776497397520782241371482144363031816561262038906245974894178189327640641335564584011267520198467768582253845117902844144176;
            6'd56: xpb[63] = 1024'd98792566016102447724900825877787826954562864203205270922695412290144540501678712418967663001809014008415463131260884622286157933815094110615122443293413690300187415702752620173622396803154233094166537021091508284161749934251576010813348238452502411474284602069109297954619462641056825420048315119540027493081;
            6'd57: xpb[63] = 1024'd40738847847258419688424572055427079505414745128354231627394257388997547044434640309120533362631367716512792222866394656012076402227632415572725998076493611462518472887115651460365359993014763069502094192424294577596107201720993209755471932327597184354108659388536953867864877009717249240724095294551616357655;
            6'd58: xpb[63] = 1024'd106751825362539133050747245637880764800965053179238876460224957552827448924499707109288474938111395734053270721929398124317058711481391055085489677875904573558540204641049900084738562374392498766147848972144320717394825319411307181662574195885921406500752620122081667811216819452306306078518565296188799706560;
            6'd59: xpb[63] = 1024'd48698107193695105014270991815520017351816934104387837164923802651680455467255634999441345298933749442150599813534908158042977179893929360043093232658984494720871261825412931371481525564253028741483406143477107010829182586880724380604697889761016179380576677441509323724462233820966729899194345471200388571134;
            6'd60: xpb[63] = 1024'd114711084708975818376593665397973702647367242155272481997754502815510357347320701799609286874413777459691078312597911626347959489147687999555856912458395456816892993579347179995854727945630764438129160923197133150627900704571038352511800153319340401527220638175054037667814176263555786736988815472837571920039;
            6'd61: xpb[63] = 1024'd56657366540131790340117411575612955198219123080421442702453347914363363890076629689762157235236131167788407404203421660073877957560226304513460467241475377979224050763710211282597691135491294413464718094529919444062257972040455551453923847194435174407044695494481693581059590632216210557664595647849160784613;
            6'd62: xpb[63] = 1024'd122670344055412503702440085158066640493769431131306087535284048078193265770141696489930098810716159185328885903266425128378860266813984944026224147040886340075245782517644459906970893516869030110110472874249945583860976089730769523361026110752759396553688656228026407524411533074805267395459065649486344133518;
            6'd63: xpb[63] = 1024'd64616625886568475665963831335705893044621312056455048239982893177046272312897624380082969171538512893426214994871935162104778735226523248983827701823966261237576839702007491193713856706729560085446030045582731877295333357200186722303149804627854169433512713547454063437656947443465691216134845824497932998092;
        endcase
    end

    always_comb begin
        case(flag[21][11:6])
            6'd0: xpb[64] = 1024'd0;
            6'd1: xpb[64] = 1024'd6562907717724447629487577513345145595473192981604008944681738275899278855653552270235839532360866601523544086477445195830697203639061553941431256607046182399907896886370522480456819896590090060781587216915518170729690624669603921245273498502948942313336770866881719350902361812126115036810625999509521862666;
            6'd2: xpb[64] = 1024'd13125815435448895258975155026690291190946385963208017889363476551798557711307104540471679064721733203047088172954890391661394407278123107882862513214092364799815793772741044960913639793180180121563174433831036341459381249339207842490546997005897884626673541733763438701804723624252230073621251999019043725332;
            6'd3: xpb[64] = 1024'd19688723153173342888462732540035436786419578944812026834045214827697836566960656810707518597082599804570632259432335587492091610917184661824293769821138547199723690659111567441370459689770270182344761650746554512189071874008811763735820495508846826940010312600645158052707085436378345110431877998528565587998;
            6'd4: xpb[64] = 1024'd26251630870897790517950310053380582381892771926416035778726953103597115422614209080943358129443466406094176345909780783322788814556246215765725026428184729599631587545482089921827279586360360243126348867662072682918762498678415684981093994011795769253347083467526877403609447248504460147242503998038087450664;
            6'd5: xpb[64] = 1024'd32814538588622238147437887566725727977365964908020044723408691379496394278267761351179197661804333007617720432387225979153486018195307769707156283035230911999539484431852612402284099482950450303907936084577590853648453123348019606226367492514744711566683854334408596754511809060630575184053129997547609313330;
            6'd6: xpb[64] = 1024'd39377446306346685776925465080070873572839157889624053668090429655395673133921313621415037194165199609141264518864671174984183221834369323648587539642277094399447381318223134882740919379540540364689523301493109024378143748017623527471640991017693653880020625201290316105414170872756690220863755997057131175996;
            6'd7: xpb[64] = 1024'd45940354024071133406413042593416019168312350871228062612772167931294951989574865891650876726526066210664808605342116370814880425473430877590018796249323276799355278204593657363197739276130630425471110518408627195107834372687227448716914489520642596193357396068172035456316532684882805257674381996566653038662;
            6'd8: xpb[64] = 1024'd52503261741795581035900620106761164763785543852832071557453906207194230845228418161886716258886932812188352691819561566645577629112492431531450052856369459199263175090964179843654559172720720486252697735324145365837524997356831369962187988023591538506694166935053754807218894497008920294485007996076174901328;
            6'd9: xpb[64] = 1024'd59066169459520028665388197620106310359258736834436080502135644483093509700881970432122555791247799413711896778297006762476274832751553985472881309463415641599171071977334702324111379069310810547034284952239663536567215622026435291207461486526540480820030937801935474158121256309135035331295633995585696763994;
            6'd10: xpb[64] = 1024'd65629077177244476294875775133451455954731929816040089446817382758992788556535522702358395323608666015235440864774451958306972036390615539414312566070461823999078968863705224804568198965900900607815872169155181707296906246696039212452734985029489423133367708668817193509023618121261150368106259995095218626660;
            6'd11: xpb[64] = 1024'd72191984894968923924363352646796601550205122797644098391499121034892067412189074972594234855969532616758984951251897154137669240029677093355743822677508006398986865750075747285025018862490990668597459386070699878026596871365643133698008483532438365446704479535698912859925979933387265404916885994604740489326;
            6'd12: xpb[64] = 1024'd78754892612693371553850930160141747145678315779248107336180859310791346267842627242830074388330399218282529037729342349968366443668738647297175079284554188798894762636446269765481838759081080729379046602986218048756287496035247054943281982035387307760041250402580632210828341745513380441727511994114262351992;
            6'd13: xpb[64] = 1024'd85317800330417819183338507673486892741151508760852116280862597586690625123496179513065913920691265819806073124206787545799063647307800201238606335891600371198802659522816792245938658655671170790160633819901736219485978120704850976188555480538336250073378021269462351561730703557639495478538137993623784214658;
            6'd14: xpb[64] = 1024'd91880708048142266812826085186832038336624701742456125225544335862589903979149731783301753453052132421329617210684232741629760850946861755180037592498646553598710556409187314726395478552261260850942221036817254390215668745374454897433828979041285192386714792136344070912633065369765610515348763993133306077324;
            6'd15: xpb[64] = 1024'd98443615765866714442313662700177183932097894724060134170226074138489182834803284053537592985412999022853161297161677937460458054585923309121468849105692735998618453295557837206852298448851350911723808253732772560945359370044058818679102477544234134700051563003225790263535427181891725552159389992642827939990;
            6'd16: xpb[64] = 1024'd105006523483591162071801240213522329527571087705664143114907812414388461690456836323773432517773865624376705383639123133291155258224984863062900105712738918398526350181928359687309118345441440972505395470648290731675049994713662739924375976047183077013388333870107509614437788994017840588970015992152349802656;
            6'd17: xpb[64] = 1024'd111569431201315609701288817726867475123044280687268152059589550690287740546110388594009272050134732225900249470116568329121852461864046417004331362319785100798434247068298882167765938242031531033286982687563808902404740619383266661169649474550132019326725104736989228965340150806143955625780641991661871665322;
            6'd18: xpb[64] = 1024'd118132338919040057330776395240212620718517473668872161004271288966187019401763940864245111582495598827423793556594013524952549665503107970945762618926831283198342143954669404648222758138621621094068569904479327073134431244052870582414922973053080961640061875603870948316242512618270070662591267991171393527988;
            6'd19: xpb[64] = 1024'd628550952639763561465045348743333569292239524740485820821172177109402920108354224465879900198791119504188235613965286204183028300949190332033750517546424664559366271468709791049338843694505433539959513007605397499761018501577730695217901872800454686578743056635609637038346356467552682283204164055320906323;
            6'd20: xpb[64] = 1024'd7191458670364211190952622862088479164765432506344494765502910453008681775761906494701719432559657721027732322091410482034880231940010744273465007124592607064467263157839232271506158740284595494321546729923123568229451643171181651940491400375749396999915513923517328987940708168593667719093830163564842768989;
            6'd21: xpb[64] = 1024'd13754366388088658820440200375433624760238625487948503710184648728907960631415458764937558964920524322551276408568855677865577435579072298214896263731638789464375160044209754751962978636874685555103133946838641738959142267840785573185764898878698339313252284790399048338843069980719782755904456163074364631655;
            6'd22: xpb[64] = 1024'd20317274105813106449927777888778770355711818469552512654866387004807239487069011035173398497281390924074820495046300873696274639218133852156327520338684971864283056930580277232419798533464775615884721163754159909688832892510389494431038397381647281626589055657280767689745431792845897792715082162583886494321;
            6'd23: xpb[64] = 1024'd26880181823537554079415355402123915951185011451156521599548125280706518342722563305409238029642257525598364581523746069526971842857195406097758776945731154264190953816950799712876618430054865676666308380669678080418523517179993415676311895884596223939925826524162487040647793604972012829525708162093408356987;
            6'd24: xpb[64] = 1024'd33443089541262001708902932915469061546658204432760530544229863556605797198376115575645077562003124127121908668001191265357669046496256960039190033552777336664098850703321322193333438326644955737447895597585196251148214141849597336921585394387545166253262597391044206391550155417098127866336334161602930219653;
            6'd25: xpb[64] = 1024'd40005997258986449338390510428814207142131397414364539488911601832505076054029667845880917094363990728645452754478636461188366250135318513980621290159823519064006747589691844673790258223235045798229482814500714421877904766519201258166858892890494108566599368257925925742452517229224242903146960161112452082319;
            6'd26: xpb[64] = 1024'd46568904976710896967878087942159352737604590395968548433593340108404354909683220116116756626724857330168996840956081657019063453774380067922052546766869701463914644476062367154247078119825135859011070031416232592607595391188805179412132391393443050879936139124807645093354879041350357939957586160621973944985;
            6'd27: xpb[64] = 1024'd53131812694435344597365665455504498333077783377572557378275078384303633765336772386352596159085723931692540927433526852849760657413441621863483803373915883863822541362432889634703898016415225919792657248331750763337286015858409100657405889896391993193272909991689364444257240853476472976768212160131495807651;
            6'd28: xpb[64] = 1024'd59694720412159792226853242968849643928550976359176566322956816660202912620990324656588435691446590533216085013910972048680457861052503175804915059980962066263730438248803412115160717913005315980574244465247268934066976640528013021902679388399340935506609680858571083795159602665602588013578838159641017670317;
            6'd29: xpb[64] = 1024'd66257628129884239856340820482194789524024169340780575267638554936102191476643876926824275223807457134739629100388417244511155064691564729746346316588008248663638335135173934595617537809595406041355831682162787104796667265197616943147952886902289877819946451725452803146061964477728703050389464159150539532983;
            6'd30: xpb[64] = 1024'd72820535847608687485828397995539935119497362322384584212320293212001470332297429197060114756168323736263173186865862440341852268330626283687777573195054431063546232021544457076074357706185496102137418899078305275526357889867220864393226385405238820133283222592334522496964326289854818087200090158660061395649;
            6'd31: xpb[64] = 1024'd79383443565333135115315975508885080714970555303988593157002031487900749187950981467295954288529190337786717273343307636172549471969687837629208829802100613463454128907914979556531177602775586162919006115993823446256048514536824785638499883908187762446619993459216241847866688101980933124010716158169583258315;
            6'd32: xpb[64] = 1024'd85946351283057582744803553022230226310443748285592602101683769763800028043604533737531793820890056939310261359820752832003246675608749391570640086409146795863362025794285502036987997499365676223700593332909341616985739139206428706883773382411136704759956764326097961198769049914107048160821342157679105120981;
            6'd33: xpb[64] = 1024'd92509259000782030374291130535575371905916941267196611046365508039699306899258086007767633353250923540833805446298198027833943879247810945512071343016192978263269922680656024517444817395955766284482180549824859787715429763876032628129046880914085647073293535192979680549671411726233163197631968157188626983647;
            6'd34: xpb[64] = 1024'd99072166718506478003778708048920517501390134248800619991047246315598585754911638278003472885611790142357349532775643223664641082886872499453502599623239160663177819567026546997901637292545856345263767766740377958445120388545636549374320379417034589386630306059861399900573773538359278234442594156698148846313;
            6'd35: xpb[64] = 1024'd105635074436230925633266285562265663096863327230404628935728984591497864610565190548239312417972656743880893619253088419495338286525934053394933856230285343063085716453397069478358457189135946406045354983655896129174811013215240470619593877919983531699967076926743119251476135350485393271253220156207670708979;
            6'd36: xpb[64] = 1024'd112197982153955373262753863075610808692336520212008637880410722867397143466218742818475151950333523345404437705730533615326035490164995607336365112837331525462993613339767591958815277085726036466826942200571414299904501637884844391864867376422932474013303847793624838602378497162611508308063846155717192571645;
            6'd37: xpb[64] = 1024'd118760889871679820892241440588955954287809713193612646825092461143296422321872295088710991482694389946927981792207978811156732693804057161277796369444377707862901510226138114439272096982316126527608529417486932470634192262554448313110140874925881416326640618660506557953280858974737623344874472155226714434311;
            6'd38: xpb[64] = 1024'd1257101905279527122930090697486667138584479049480971641642344354218805840216708448931759800397582239008376471227930572408366056601898380664067501035092849329118732542937419582098677687389010867079919026015210794999522037003155461390435803745600909373157486113271219274076692712935105364566408328110641812646;
            6'd39: xpb[64] = 1024'd7820009623003974752417668210831812734057672031084980586324082630118084695870260719167599332758448840531920557705375768239063260240959934605498757642139031729026629429307942062555497583979100927861506242930728965729212661672759382635709302248549851686494256980152938624979054525061220401377034327620163675312;
            6'd40: xpb[64] = 1024'd14382917340728422381905245724176958329530865012688989531005820906017363551523812989403438865119315442055464644182820964069760463880021488546930014249185214128934526315678464543012317480569190988643093459846247136458903286342363303880982800751498793999831027847034657975881416337187335438187660327129685537978;
            6'd41: xpb[64] = 1024'd20945825058452870011392823237522103925004057994292998475687559181916642407177365259639278397480182043579008730660266159900457667519083042488361270856231396528842423202048987023469137377159281049424680676761765307188593911011967225126256299254447736313167798713916377326783778149313450474998286326639207400644;
            6'd42: xpb[64] = 1024'd27508732776177317640880400750867249520477250975897007420369297457815921262830917529875117929841048645102552817137711355731154871158144596429792527463277578928750320088419509503925957273749371110206267893677283477918284535681571146371529797757396678626504569580798096677686139961439565511808912326148729263310;
            6'd43: xpb[64] = 1024'd34071640493901765270367978264212395115950443957501016365051035733715200118484469800110957462201915246626096903615156551561852074797206150371223784070323761328658216974790031984382777170339461170987855110592801648647975160351175067616803296260345620939841340447679816028588501773565680548619538325658251125976;
            6'd44: xpb[64] = 1024'd40634548211626212899855555777557540711423636939105025309732774009614478974138022070346796994562781848149640990092601747392549278436267704312655040677369943728566113861160554464839597066929551231769442327508319819377665785020778988862076794763294563253178111314561535379490863585691795585430164325167772988642;
            6'd45: xpb[64] = 1024'd47197455929350660529343133290902686306896829920709034254414512285513757829791574340582636526923648449673185076570046943223246482075329258254086297284416126128474010747531076945296416963519641292551029544423837990107356409690382910107350293266243505566514882181443254730393225397817910622240790324677294851308;
            6'd46: xpb[64] = 1024'd53760363647075108158830710804247831902370022902313043199096250561413036685445126610818476059284515051196729163047492139053943685714390812195517553891462308528381907633901599425753236860109731353332616761339356160837047034359986831352623791769192447879851653048324974081295587209944025659051416324186816713974;
            6'd47: xpb[64] = 1024'd60323271364799555788318288317592977497843215883917052143777988837312315541098678881054315591645381652720273249524937334884640889353452366136948810498508490928289804520272121906210056756699821414114203978254874331566737659029590752597897290272141390193188423915206693432197949022070140695862042323696338576640;
            6'd48: xpb[64] = 1024'd66886179082524003417805865830938123093316408865521061088459727113211594396752231151290155124006248254243817336002382530715338092992513920078380067105554673328197701406642644386666876653289911474895791195170392502296428283699194673843170788775090332506525194782088412783100310834196255732672668323205860439306;
            6'd49: xpb[64] = 1024'd73449086800248451047293443344283268688789601847125070033141465389110873252405783421525994656367114855767361422479827726546035296631575474019811323712600855728105598293013166867123696549880001535677378412085910673026118908368798595088444287278039274819861965648970132134002672646322370769483294322715382301972;
            6'd50: xpb[64] = 1024'd80011994517972898676781020857628414284262794828729078977823203665010152108059335691761834188727981457290905508957272922376732500270637027961242580319647038128013495179383689347580516446470091596458965629001428843755809533038402516333717785780988217133198736515851851484905034458448485806293920322224904164638;
            6'd51: xpb[64] = 1024'd86574902235697346306268598370973559879735987810333087922504941940909430963712887961997673721088848058814449595434718118207429703909698581902673836926693220527921392065754211828037336343060181657240552845916947014485500157708006437578991284283937159446535507382733570835807396270574600843104546321734426027304;
            6'd52: xpb[64] = 1024'd93137809953421793935756175884318705475209180791937096867186680216808709819366440232233513253449714660337993681912163314038126907548760135844105093533739402927829288952124734308494156239650271718022140062832465185215190782377610358824264782786886101759872278249615290186709758082700715879915172321243947889970;
            6'd53: xpb[64] = 1024'd99700717671146241565243753397663851070682373773541105811868418492707988675019992502469352785810581261861537768389608509868824111187821689785536350140785585327737185838495256788950976136240361778803727279747983355944881407047214280069538281289835044073209049116497009537612119894826830916725798320753469752636;
            6'd54: xpb[64] = 1024'd106263625388870689194731330911008996666155566755145114756550156768607267530673544772705192318171447863385081854867053705699521314826883243726967606747831767727645082724865779269407796032830451839585314496663501526674572031716818201314811779792783986386545819983378728888514481706952945953536424320262991615302;
            6'd55: xpb[64] = 1024'd112826533106595136824218908424354142261628759736749123701231895044506546386327097042941031850532314464908625941344498901530218518465944797668398863354877950127552979611236301749864615929420541900366901713579019697404262656386422122560085278295732928699882590850260448239416843519079060990347050319772513477968;
            6'd56: xpb[64] = 1024'd119389440824319584453706485937699287857101952718353132645913633320405825241980649313176871382893181066432170027821944097360915722105006351609830119961924132527460876497606824230321435826010631961148488930494537868133953281056026043805358776798681871013219361717142167590319205331205176027157676319282035340634;
            6'd57: xpb[64] = 1024'd1885652857919290684395136046230000707876718574221457462463516531328208760325062673397639700596373358512564706841895858612549084902847570996101251552639273993678098814406129373148016531083516300619878539022816192499283055504733192085653705618401364059736229169906828911115039069402658046849612492165962718969;
            6'd58: xpb[64] = 1024'd8448560575643738313882713559575146303349911555825466407145254807227487615978614943633479232957239960036108793319341054443246288541909124937532508159685456393585995700776651853604836427673606361401465755938334363228973680174337113330927204121350306373073000036788548262017400881528773083660238491675484581635;
            6'd59: xpb[64] = 1024'd15011468293368185943370291072920291898823104537429475351826993083126766471632167213869318765318106561559652879796786250273943492180970678878963764766731638793493892587147174334061656324263696422183052972853852533958664304843941034576200702624299248686409770903670267612919762693654888120470864491185006444301;
            6'd60: xpb[64] = 1024'd21574376011092633572857868586265437494296297519033484296508731359026045327285719484105158297678973163083196966274231446104640695820032232820395021373777821193401789473517696814518476220853786482964640189769370704688354929513544955821474201127248190999746541770551986963822124505781003157281490490694528306967;
            6'd61: xpb[64] = 1024'd28137283728817081202345446099610583089769490500637493241190469634925324182939271754340997830039839764606741052751676641935337899459093786761826277980824003593309686359888219294975296117443876543746227406684888875418045554183148877066747699630197133313083312637433706314724486317907118194092116490204050169633;
            6'd62: xpb[64] = 1024'd34700191446541528831833023612955728685242683482241502185872207910824603038592824024576837362400706366130285139229121837766035103098155340703257534587870185993217583246258741775432116014033966604527814623600407046147736178852752798312021198133146075626420083504315425665626848130033233230902742489713572032299;
            6'd63: xpb[64] = 1024'd41263099164265976461320601126300874280715876463845511130553946186723881894246376294812676894761572967653829225706567033596732306737216894644688791194916368393125480132629264255888935910624056665309401840515925216877426803522356719557294696636095017939756854371197145016529209942159348267713368489223093894965;
        endcase
    end

    always_comb begin
        case(flag[21][16:12])
            5'd0: xpb[65] = 1024'd0;
            5'd1: xpb[65] = 1024'd47826006881990424090808178639646019876189069445449520075235684462623160749899928565048516427122439569177373312184012229427429510376278448586120047801962550793033377018999786736345755807214146726090989057431443387607117428191960640802568195139043960253093625238078864367431571754285463304523994488732615757631;
            5'd2: xpb[65] = 1024'd95652013763980848181616357279292039752378138890899040150471368925246321499799857130097032854244879138354746624368024458854859020752556897172240095603925101586066754037999573472691511614428293452181978114862886775214234856383921281605136390278087920506187250476157728734863143508570926609047988977465231515262;
            5'd3: xpb[65] = 1024'd19411324961846530873625608514123626883868781210612876097575198322892586912390646785130478066709644398088970529094543253703224690287615011203200018389556611445409456487428142871407028230125234456962769563907090316456991434354985149442726015733902431492460972300119535072188187188927756896453293639572252788562;
            5'd4: xpb[65] = 1024'd67237331843836954964433787153769646760057850656062396172810882785515747662290575350178994493832083967266343841278555483130654200663893459789320066191519162238442833506427929607752784037339381183053758621338533704064108862546945790245294210872946391745554597538198399439619758943213220200977288128304868546193;
            5'd5: xpb[65] = 1024'd115063338725827379055241965793415666636246920101511916248046567248138908412190503915227510920954523536443717153462567712558083711040171908375440113993481713031476210525427716344098539844553527909144747678769977091671226290738906431047862406011990351998648222776277263807051330697498683505501282617037484303824;
            5'd6: xpb[65] = 1024'd38822649923693061747251217028247253767737562421225752195150396645785173824781293570260956133419288796177941058189086507406449380575230022406400036779113222890818912974856285742814056460250468913925539127814180632913982868709970298885452031467804862984921944600239070144376374377855513792906587279144505577124;
            5'd7: xpb[65] = 1024'd86648656805683485838059395667893273643926631866675272270386081108408334574681222135309472560541728365355314370373098736833878890951508470992520084581075773683852289993856072479159812267464615640016528185245624020521100296901930939688020226606848823238015569838317934511807946132140977097430581767877121334755;
            5'd8: xpb[65] = 1024'd10407968003549168530068646902724860775417274186389108217489910506054599987272011790342917773006493625089538275099617531682244560486566585023480007366707283543194992443284641877875328883161556644797319634289827561763856874872994807525609852062663334224289291662279740849132989812497807384835886429984142608055;
            5'd9: xpb[65] = 1024'd58233974885539592620876825542370880651606343631838628292725594968677760737171940355391434200128933194266911587283629761109674070862845033609600055168669834336228369462284428614221084690375703370888308691721270949370974303064955448328178047201707294477382916900358605216564561566783270689359880918716758365686;
            5'd10: xpb[65] = 1024'd106059981767530016711685004182016900527795413077288148367961279431300921487071868920439950627251372763444284899467641990537103581239123482195720102970632385129261746481284215350566840497589850096979297749152714336978091731256916089130746242340751254730476542138437469583996133321068733993883875407449374123317;
            5'd11: xpb[65] = 1024'd29819292965395699403694255416848487659286055397001984315065108828947186899662658575473395839716138023178508804194160785385469250774181596226680025756263894988604448930712784749282357113286791101760089198196917878220848309227979956968335867796565765716750263962399275921321177001425564281289180069556395396617;
            5'd12: xpb[65] = 1024'd77645299847386123494502434056494507535475124842451504390300793291570347649562587140521912266838577592355882116378173014812898761150460044812800073558226445781637825949712571485628112920500937827851078255628361265827965737419940597770904062935609725969843889200478140288752748755711027585813174558289011154248;
            5'd13: xpb[65] = 1024'd1404611045251806186511685291326094666965767162165340337404622689216613062153376795555357479303342852090106021104691809661264430685518158843759996343857955640980528399141140884343629536197878832631869704672564807070722315391004465608493688391424236956117611024439946626077792436067857873218479220396032427548;
            5'd14: xpb[65] = 1024'd49230617927242230277319863930972114543154836607614860412640307151839773812053305360603873906425782421267479333288704039088693941061796607429880044145820506434013905418140927620689385343412025558722858762104008194677839743582965106411061883530468197209211236262518810993509364190353321177742473709128648185179;
            5'd15: xpb[65] = 1024'd97056624809232654368128042570618134419343906053064380487875991614462934561953233925652390333548221990444852645472716268516123451438075056016000091947783057227047282437140714357035141150626172284813847819535451582284957171774925747213630078669512157462304861500597675360940935944638784482266468197861263942810;
            5'd16: xpb[65] = 1024'd20815936007098337060137293805449721550834548372778216434979821012109199974544023580685835546012987250179076550199235063364489120973133170046960014733414567086389984886569283755750657766323113289594639268579655123527713749745989615051219704125326668448578583324559481698265979624995614769671772859968285216110;
            5'd17: xpb[65] = 1024'd68641942889088761150945472445095741427023617818227736510215505474732360724443952145734351973135426819356449862383247292791918631349411618633080062535377117879423361905569070492096413573537260015685628326011098511134831177937950255853787899264370628701672208562638346065697551379281078074195767348700900973741;
            5'd18: xpb[65] = 1024'd116467949771079185241753651084741761303212687263677256585451189937355521474343880710782868400257866388533823174567259522219348141725690067219200110337339668672456738924568857228442169380751406741776617383442541898741948606129910896656356094403414588954765833800717210433129123133566541378719761837433516731372;
            5'd19: xpb[65] = 1024'd40227260968944867933762902319573348434703329583391092532555019335001786886934670365816313612722631648268047079293778317067713811260748181250160033122971178531799441373997426627157685996448347746557408832486745439984705184100974764493945719859229099941039555624679016770454166813923371666125066499540538004672;
            5'd20: xpb[65] = 1024'd88053267850935292024571080959219368310892399028840612607790703797624947636834598930864830039845071217445420391477790546495143321637026629836280080924933729324832818392997213363503441803662494472648397889918188827591822612292935405296513914998273060194133180862757881137885738568208834970649060988273153762303;
            5'd21: xpb[65] = 1024'd11812579048800974716580332194050955442383041348554448554894533195271213049425388585898275252309836477179644296204309341343508991172084743867240003710565239184175520842425782762218958419359435477429189338962392368834579190263999273134103540454087571180406902686719687475210782248565665258054365650380175035603;
            5'd22: xpb[65] = 1024'd59638585930791398807388510833696975318572110794003968630130217657894373799325317150946791679432276046357017608388321570770938501548363192453360051512527789977208897861425569498564714226573582203520178396393835756441696618455959913936671735593131531433500527924798551842642354002851128562578360139112790793234;
            5'd23: xpb[65] = 1024'd107464592812781822898196689473342995194761180239453488705365902120517534549225245715995308106554715615534390920572333800198368011924641641039480099314490340770242274880425356234910470033787728929611167453825279144048814046647920554739239930732175491686594153162877416210073925757136591867102354627845406550865;
            5'd24: xpb[65] = 1024'd31223904010647505590205940708174582326251822559167324652469731518163799961816035371028753319019480875268614825298852595046733681459699755070440022100121850629584977329853925633625986649484669934391958902869482685291570624618984422576829556187990002672867874986839222547398969437493422154507659289952427824165;
            5'd25: xpb[65] = 1024'd79049910892637929681014119347820602202440892004616844727705415980786960711715963936077269746141920444445988137482864824474163191835978203656560069902084401422618354348853712369971742456698816660482947960300926072898688052810945063379397751327033962925961500224918086914830541191778885459031653778685043581796;
            5'd26: xpb[65] = 1024'd2809222090503612373023370582652189333931534324330680674809245378433226124306753591110714958606685704180212042209383619322528861371036317687519992687715911281961056798282281768687259072395757665263739409345129614141444630782008931216987376782848473912235222048879893252155584872135715746436958440792064855096;
            5'd27: xpb[65] = 1024'd50635228972494036463831549222298209210120603769780200750044929841056386874206682156159231385729125273357585354393395848749958371747314766273640040489678462074994433817282068505033014879609904391354728466776573001748562058973969572019555571921892434165328847286958757619587156626421179050960952929524680612727;
            5'd28: xpb[65] = 1024'd98461235854484460554639727861944229086309673215229720825280614303679547624106610721207747812851564842534958666577408078177387882123593214859760088291641012868027810836281855241378770686824051117445717524208016389355679487165930212822123767060936394418422472525037621987018728380706642355484947418257296370358;
            5'd29: xpb[65] = 1024'd22220547052350143246648979096775816217800315534943556772384443701325813036697400376241193025316330102269182571303926873025753551658651328890720011077272522727370513285710424640094287302520992122226508973252219930598436065136994080659713392516750905404696194348999428324343772061063472642890252080364317643658;
            5'd30: xpb[65] = 1024'd70046553934340567337457157736421836093989384980393076847620128163948973786597328941289709452438769671446555883487939102453183062034929777476840058879235073520403890304710211376440043109735138848317498030683663318205553493328954721462281587655794865657789819587078292691775343815348935947414246569096933401289;
            5'd31: xpb[65] = 1024'd117872560816330991428265336376067855970178454425842596922855812626572134536497257506338225879561209240623929195671951331880612572411208226062960106681197624313437267323709998112785798916949285574408487088115106705812670921520915362264849782794838825910883444825157157059206915569634399251938241057829549158920;
        endcase
    end

    always_comb begin
        case(flag[22][5:0])
            6'd0: xpb[66] = 1024'd0;
            6'd1: xpb[66] = 1024'd20815936007098337060137293805449721550834548372778216434979821012109199974544023580685835546012987250179076550199235063364489120973133170046960014733414567086389984886569283755750657766323113289594639268579655123527713749745989615051219704125326668448578583324559481698265979624995614769671772859968285216110;
            6'd2: xpb[66] = 1024'd41631872014196674120274587610899443101669096745556432869959642024218399949088047161371671092025974500358153100398470126728978241946266340093920029466829134172779969773138567511501315532646226579189278537159310247055427499491979230102439408250653336897157166649118963396531959249991229539343545719936570432220;
            6'd3: xpb[66] = 1024'd62447808021295011180411881416349164652503645118334649304939463036327599923632070742057506638038961750537229650597705190093467362919399510140880044200243701259169954659707851267251973298969339868783917805738965370583141249237968845153659112375980005345735749973678445094797938874986844309015318579904855648330;
            6'd4: xpb[66] = 1024'd83263744028393348240549175221798886203338193491112865739919284048436799898176094322743342184051949000716306200796940253457956483892532680187840058933658268345559939546277135023002631065292453158378557074318620494110854998983958460204878816501306673794314333298237926793063918499982459078687091439873140864440;
            6'd5: xpb[66] = 1024'd104079680035491685300686469027248607754172741863891082174899105060545999872720117903429177730064936250895382750996175316822445604865665850234800073667072835431949924432846418778753288831615566447973196342898275617638568748729948075256098520626633342242892916622797408491329898124978073848358864299841426080550;
            6'd6: xpb[66] = 1024'd828920358465280962024835427883896560308863110933614481747071007678304509955002574099942061420249191631309893737916945607870884997578685726599963384156361584649234749844485196873707406421474016257638003090690894801921648255040917342339655068730561424651596533239832159489349676045055600911947333184116812329;
            6'd7: xpb[66] = 1024'd21644856365563618022162129233333618111143411483711830916726892019787504484499026154785777607433236441810386443937152008972360005970711855773559978117570928671039219636413768952624365172744587305852277271670346018329635398001030532393559359194057229873230179857799313857755329301040670370583720193152402028439;
            6'd8: xpb[66] = 1024'd42460792372661955082299423038783339661977959856490047351706713031896704459043049735471613153446223691989462994136387072336849126943845025820519992850985495757429204522983052708375022939067700595446916540250001141857349147747020147444779063319383898321808763182358795556021308926036285140255493053120687244549;
            6'd9: xpb[66] = 1024'd63276728379760292142436716844233061212812508229268263786686534044005904433587073316157448699459210942168539544335622135701338247916978195867480007584400062843819189409552336464125680705390813885041555808829656265385062897493009762495998767444710566770387346506918277254287288551031899909927265913088972460659;
            6'd10: xpb[66] = 1024'd84092664386858629202574010649682782763647056602046480221666355056115104408131096896843284245472198192347616094534857199065827368890111365914440022317814629930209174296121620219876338471713927174636195077409311388912776647238999377547218471570037235218965929831477758952553268176027514679599038773057257676769;
            6'd11: xpb[66] = 1024'd104908600393956966262711304455132504314481604974824696656646176068224304382675120477529119791485185442526692644734092262430316489863244535961400037051229197016599159182690903975626996238037040464230834345988966512440490396984988992598438175695363903667544513156037240650819247801023129449270811633025542892879;
            6'd12: xpb[66] = 1024'd1657840716930561924049670855767793120617726221867228963494142015356609019910005148199884122840498383262619787475833891215741769995157371453199926768312723169298469499688970393747414812842948032515276006181381789603843296510081834684679310137461122849303193066479664318978699352090111201823894666368233624658;
            6'd13: xpb[66] = 1024'd22473776724028898984186964661217514671452274594645445398473963027465808994454028728885719668853485633441696337675068954580230890968290541500159941501727290255688454386258254149498072579166061322109915274761036913131557046256071449735899014262787791297881776391039146017244678977085725971495667526336518840768;
            6'd14: xpb[66] = 1024'd43289712731127236044324258466667236222286822967423661833453784039575008968998052309571555214866472883620772887874304017944720011941423711547119956235141857342078439272827537905248730345489174611704554543340692036659270796002061064787118718388114459746460359715598627715510658602081340741167440386304804056878;
            6'd15: xpb[66] = 1024'd64105648738225573104461552272116957773121371340201878268433605051684208943542075890257390760879460133799849438073539081309209132914556881594079970968556424428468424159396821660999388111812287901299193811920347160186984545748050679838338422513441128195038943040158109413776638227076955510839213246273089272988;
            6'd16: xpb[66] = 1024'd84921584745323910164598846077566679323955919712980094703413426063793408918086099470943226306892447383978925988272774144673698253887690051641039985701970991514858409045966105416750045878135401190893833080500002283714698295494040294889558126638767796643617526364717591112042617852072570280510986106241374489098;
            6'd17: xpb[66] = 1024'd105737520752422247224736139883016400874790468085758311138393247075902608892630123051629061852905434634158002538472009208038187374860823221688000000435385558601248393932535389172500703644458514480488472349079657407242412045240029909940777830764094465092196109689277072810308597477068185050182758966209659705208;
            6'd18: xpb[66] = 1024'd2486761075395842886074506283651689680926589332800843445241213023034913529865007722299826184260747574893929681213750836823612654992736057179799890152469084753947704249533455590621122219264422048772914009272072684405764944765122752027018965206191684273954789599719496478468049028135166802735841999552350436987;
            6'd19: xpb[66] = 1024'd23302697082494179946211800089101411231761137705579059880221034035144113504409031302985661730273734825073006231412985900188101775965869227226759904885883651840337689136102739346371779985587535338367553277851727807933478694511112367078238669331518352722533372924278978176734028653130781572407614859520635653097;
            6'd20: xpb[66] = 1024'd44118633089592517006349093894551132782595686078357276315200855047253313478953054883671497276286722075252082781612220963552590896939002397273719919619298218926727674022672023102122437751910648627962192546431382931461192444257101982129458373456845021171111956248838459875000008278126396342079387719488920869207;
            6'd21: xpb[66] = 1024'd64934569096690854066486387700000854333430234451135492750180676059362513453497078464357332822299709325431159331811456026917080017912135567320679934352712786013117658909241306857873095518233761917556831815011038054988906194003091597180678077582171689619690539573397941573265987903122011111751160579457206085317;
            6'd22: xpb[66] = 1024'd85750505103789191126623681505450575884264782823913709185160497071471713428041102045043168368312696575610235882010691090281569138885268737367639949086127353099507643795810590613623753284556875207151471083590693178516619943749081212231897781707498358068269122897957423271531967528117625881422933439425491301427;
            6'd23: xpb[66] = 1024'd106566441110887528186760975310900297435099331196691925620140318083580913402585125625729003914325683825789312432209926153646058259858401907414599963819541920185897628682379874369374411050879988496746110352170348302044333693495070827283117485832825026516847706222516904969797947153113240651094706299393776517537;
            6'd24: xpb[66] = 1024'd3315681433861123848099341711535586241235452443734457926988284030713218039820010296399768245680996766525239574951667782431483539990314742906399853536625446338596938999377940787494829625685896065030552012362763579207686593020163669369358620274922245698606386132959328637957398704180222403647789332736467249316;
            6'd25: xpb[66] = 1024'd24131617440959460908236635516985307792070000816512674361968105042822418014364033877085603791693984016704316125150902845795972660963447912953359868270040013424986923885947224543245487392009009354625191280942418702735400342766153284420578324400248914147184969457518810336223378329175837173319562192704752465426;
            6'd26: xpb[66] = 1024'd44947553448057797968373929322435029342904549189290890796947926054931617988908057457771439337706971266883392675350137909160461781936581083000319883003454580511376908772516508298996145158332122644219830549522073826263114092512142899471798028525575582595763552782078292034489357954171451942991335052673037681536;
            6'd27: xpb[66] = 1024'd65763489455156135028511223127884750893739097562069107231927747067040817963452081038457274883719958517062469225549372972524950902909714253047279897736869147597766893659085792054746802924655235933814469818101728949790827842258132514523017732650902251044342136106637773732755337579167066712663107912641322897646;
            6'd28: xpb[66] = 1024'd86579425462254472088648516933334472444573645934847323666907568079150017937996104619143110429732945767241545775748608035889440023882847423094239912470283714684156878545655075810497460690978349223409109086681384073318541592004122129574237436776228919492920719431197255431021317204162681482334880772609608113756;
            6'd29: xpb[66] = 1024'd107395361469352809148785810738784193995408194307625540101887389091259217912540128199828945975745933017420622325947843099253929144855980593141199927203698281770546863432224359566248118457301462513003748355261039196846255341750111744625457140901555587941499302755756737129287296829158296252006653632577893329866;
            6'd30: xpb[66] = 1024'd4144601792326404810124177139419482801544315554668072408735355038391522549775012870499710307101245958156549468689584728039354424987893428632999816920781807923246173749222425984368537032107370081288190015453454474009608241275204586711698275343652807123257982666199160797446748380225278004559736665920584061645;
            6'd31: xpb[66] = 1024'd24960537799424741870261470944869204352378863927446288843715176050500722524319036451185545853114233208335626018888819791403843545961026598679959831654196375009636158635791709740119194798430483370882829284033109597537321991021194201762917979468979475571836565990758642495712728005220892774231509525888869277755;
            6'd32: xpb[66] = 1024'd45776473806523078930398764750318925903213412300224505278694997062609922498863060031871381399127220458514702569088054854768332666934159768726919846387610942096026143522360993495869852564753596660477468552612764721065035740767183816814137683594306144020415149315318124193978707630216507543903282385857154493865;
            6'd33: xpb[66] = 1024'd66592409813621415990536058555768647454047960673002721713674818074719122473407083612557216945140207708693779119287289918132821787907292938773879861121025509182416128408930277251620510331076709950072107821192419844592749490513173431865357387719632812468993732639877605892244687255212122313575055245825439709975;
            6'd34: xpb[66] = 1024'd87408345820719753050673352361218369004882509045780938148654639086828322447951107193243052491153194958872855669486524981497310908880426108820839875854440076268806113295499561007371168097399823239666747089772074968120463240259163046916577091844959480917572315964437087590510666880207737083246828105793724926085;
            6'd35: xpb[66] = 1024'd108224281827818090110810646166668090555717057418559154583634460098937522422495130773928888037166182209051932219685760044861800029853559278867799890587854643355196098182068844763121825863722936529261386358351730091648176990005152661967796795970286149366150899288996569288776646505203351852918600965762010142195;
            6'd36: xpb[66] = 1024'd4973522150791685772149012567303379361853178665601686890482426046069827059730015444599652368521495149787859362427501673647225309985472114359599780304938169507895408499066911181242244438528844097545828018544145368811529889530245504054037930412383368547909579199438992956936098056270333605471683999104700873974;
            6'd37: xpb[66] = 1024'd25789458157890022832286306372753100912687727038379903325462247058179027034274039025285487914534482399966935912626736737011714430958605284406559795038352736594285393385636194936992902204851957387140467287123800492339243639276235119105257634537710036996488162523998474655202077681265948375143456859072986090084;
            6'd38: xpb[66] = 1024'd46605394164988359892423600178202822463522275411158119760442068070288227008818062605971323460547469650146012462825971800376203551931738454453519809771767303680675378272205478692743559971175070676735106555703455615866957389022224734156477338663036705445066745848557956353468057306261563144815229719041271306194;
            6'd39: xpb[66] = 1024'd67421330172086696952560893983652544014356823783936336195421889082397426983362086186657159006560456900325089013025206863740692672904871624500479824505181870767065363158774762448494217737498183966329745824283110739394671138768214349207697042788363373893645329173117438051734036931257177914487002579009556522304;
            6'd40: xpb[66] = 1024'd88237266179185034012698187789102265565191372156714552630401710094506626957906109767342994552573444150504165563224441927105181793878004794547439839238596437853455348045344046204244875503821297255924385092862765862922384888514203964258916746913690042342223912497676919750000016556252792684158775438977841738414;
            6'd41: xpb[66] = 1024'd109053202186283371072835481594551987116025920529492769065381531106615826932450133348028830098586431400683242113423676990469670914851137964594399853972011004939845332931913329959995533270144410545519024361442420986450098638260193579310136451039016710790802495822236401448265996181248407453830548298946126954524;
            6'd42: xpb[66] = 1024'd5802442509256966734173847995187275922162041776535301372229497053748131569685018018699594429941744341419169256165418619255096194983050800086199743689094531092544643248911396378115951844950318113803466021634836263613451537785286421396377585481113929972561175732678825116425447732315389206383631332288817686303;
            6'd43: xpb[66] = 1024'd26618378516355303794311141800636997472996590149313517807209318065857331544229041599385429975954731591598245806364653682619585315956183970133159758422509098178934628135480680133866609611273431403398105290214491387141165287531276036447597289606440598421139759057238306814691427357311003976055404192257102902413;
            6'd44: xpb[66] = 1024'd47434314523453640854448435606086719023831138522091734242189139077966531518773065180071265521967718841777322356563888745984074436929317140180119773155923665265324613022049963889617267377596544692992744558794146510668879037277265651498816993731767266869718342381797788512957406982306618745727177052225388118523;
            6'd45: xpb[66] = 1024'd68250250530551977914585729411536440574665686894869950677168960090075731493317088760757101067980706091956398906763123809348563557902450310227079787889338232351714597908619247645367925143919657982587383827373801634196592787023255266550036697857093935318296925706357270211223386607302233515398949912193673334633;
            6'd46: xpb[66] = 1024'd89066186537650314974723023216986162125500235267648167112148781102184931467861112341442936613993693342135475456962358872713052678875583480274039802622752799438104582795188531401118582910242771272182023095953456757724306536769244881601256401982420603766875509030916751909489366232297848285070722772161958550743;
            6'd47: xpb[66] = 1024'd109882122544748652034860317022435883676334783640426383547128602114294131442405135922128772160006680592314552007161593936077541799848716650320999817356167366524494567681757815156869240676565884561776662364533111881252020286515234496652476106107747272215454092355476233607755345857293463054742495632130243766853;
            6'd48: xpb[66] = 1024'd6631362867722247696198683423071172482470904887468915853976568061426436079640020592799536491361993533050479149903335564862967079980629485812799707073250892677193877998755881574989659251371792130061104024725527158415373186040327338738717240549844491397212772265918657275914797408360444807295578665472934498632;
            6'd49: xpb[66] = 1024'd27447298874820584756335977228520894033305453260247132288956389073535636054184044173485372037374980783229555700102570628227456200953762655859759721806665459763583862885325165330740317017694905419655743293305182281943086935786316953789936944675171159845791355590478138974180777033356059576967351525441219714742;
            6'd50: xpb[66] = 1024'd48263234881918921816473271033970615584140001633025348723936210085644836028728067754171207583387968033408632250301805691591945321926895825906719736540080026849973847771894449086490974784018018709250382561884837405470800685532306568841156648800497828294369938915037620672446756658351674346639124385409504930852;
            6'd51: xpb[66] = 1024'd69079170889017258876610564839420337134974550005803565158916031097754036003272091334857043129400955283587708800501040754956434442900028995953679751273494593936363832658463732842241632550341131998845021830464492528998514435278296183892376352925824496742948522239597102370712736283347289116310897245377790146962;
            6'd52: xpb[66] = 1024'd89895106896115595936747858644870058685809098378581781593895852109863235977816114915542878675413942533766785350700275818320923563873162166000639766006909161022753817545033016597992290316664245288439661099044147652526228185024285798943596057051151165191527105564156584068978715908342903885982670105346075363072;
            6'd53: xpb[66] = 1024'd110711042903213932996885152450319780236643646751359998028875673121972435952360138496228714221426929783945861900899510881685412684846295336047599780740323728109143802431602300353742948082987358578034300367623802776053941934770275413994815761176477833640105688888716065767244695533338518655654442965314360579182;
            6'd54: xpb[66] = 1024'd7460283226187528658223518850955069042779767998402530335723639069104740589595023166899478552782242724681789043641252510470837964978208171539399670457407254261843112748600366771863366657793266146318742027816218053217294834295368256081056895618575052821864368799158489435404147084405500408207525998657051310961;
            6'd55: xpb[66] = 1024'd28276219233285865718360812656404790593614316371180746770703460081213940564139046747585314098795229974860865593840487573835327085951341341586359685190821821348233097635169650527614024424116379435913381296395873176745008584041357871132276599743901721270442952123717971133670126709401115177879298858625336527071;
            6'd56: xpb[66] = 1024'd49092155240384202778498106461854512144448864743958963205683281093323140538683070328271149644808217225039942144039722637199816206924474511633319699924236388434623082521738934283364682190439492725508020564975528300272722333787347486183496303869228389719021535448277452831936106334396729947551071718593621743181;
            6'd57: xpb[66] = 1024'd69908091247482539838635400267304233695283413116737179640663102105432340513227093908956985190821204475219018694238957700564305327897607681680279714657650955521013067408308218039115339956762606015102659833555183423800436083533337101234716007994555058167600118772836934530202085959392344717222844578561906959291;
            6'd58: xpb[66] = 1024'd90724027254580876898772694072753955246117961489515396075642923117541540487771117489642820736834191725398095244438192763928794448870740851727239729391065522607403052294877501794865997723085719304697299102134838547328149833279326716285935712119881726616178702097396416228468065584387959486894617438530192175401;
            6'd59: xpb[66] = 1024'd111539963261679213958909987878203676796952509862293612510622744129650740462315141070328656282847178975577171794637427827293283569843874021774199744124480089693793037181446785550616655489408832594291938370714493670855863583025316331337155416245208395064757285421955897926734045209383574256566390298498477391511;
            6'd60: xpb[66] = 1024'd8289203584652809620248354278838965603088631109336144817470710076783045099550025740999420614202491916313098937379169456078708849975786857265999633841563615846492347498444851968737074064214740162576380030906908948019216482550409173423396550687305614246515965332398321594893496760450556009119473331841168123290;
            6'd61: xpb[66] = 1024'd29105139591751146680385648084288687153923179482114361252450531088892245074094049321685256160215479166492175487578404519443197970948920027312959648574978182932882332385014135724487731830537853452171019299486564071546930232296398788474616254812632282695094548656957803293159476385446170778791246191809453339400;
            6'd62: xpb[66] = 1024'd49921075598849483740522941889738408704757727854892577687430352101001445048638072902371091706228466416671252037777639582807687091922053197359919663308392750019272317271583419480238389596860966741765658568066219195074643982042388403525835958937958951143673131981517284991425456010441785548463019051777738555510;
            6'd63: xpb[66] = 1024'd70737011605947820800660235695188130255592276227670794122410173113110645023182096483056927252241453666850328587976874646172176212895186367406879678041807317105662302158152703235989047363184080031360297836645874318602357731788378018577055663063285619592251715306076766689691435635437400318134791911746023771620;
        endcase
    end

    always_comb begin
        case(flag[22][11:6])
            6'd0: xpb[67] = 1024'd0;
            6'd1: xpb[67] = 1024'd91552947613046157860797529500637851806426824600449010557389994125219844997726120063742762798254440917029405138176109709536665333868319537453839692775221884192052287044721986991739705129507193320954937105225529442130071481534367633628275367188612288040830298630636248387957415260433015087806564771714308987730;
            6'd2: xpb[67] = 1024'd59039199541967574322796131596461270868155222075162336986648133185462794658143101217470454381851207524615660868894725984494266826895418740352519260534112727450413899519872756645849171067497180920599676602063819037895782112847838494291572164693995126814840693847155438745808302446937397158494439716803023491129;
            6'd3: xpb[67] = 1024'd26525451470888990784794733692284689929883619549875663415906272245705744318560082371198145965447974132201916599613342259451868319922517943251198828293003570708775511995023526299958637005487168520244416098902108633661492744161309354954868962199377965588851089063674629103659189633441779229182314661891737994528;
            6'd4: xpb[67] = 1024'd118078399083935148645592263192922541736310444150324673973296266370925589316286202434940908763702415049231321737789451968988533653790837480705038521068225454900827799039745513291698342134994361841199353204127638075791564225695676988583144329387990253629681387694310877491616604893874794316988879433606046982258;
            6'd5: xpb[67] = 1024'd85564651012856565107590865288745960798038841625038000402554405431168538976703183588668600347299181656817577468508068243946135146817936683603718088827116298159189411514896282945807808072984349440844092700965927671557274857009147849246441126893373092403691782910830067849467492080379176387676754378694761485657;
            6'd6: xpb[67] = 1024'd53050902941777981569589467384569379859767239099751326831812544491411488637120164742396291930895948264403833199226684518903736639845035886502397656586007141417551023990047052599917274010974337040488832197804217267322985488322618709909737924398755931177702178127349258207318379266883558458364629323783475989056;
            6'd7: xpb[67] = 1024'd20537154870699398031588069480392798921495636574464653261070683551654438297537145896123983514492714871990088929945300793861338132872135089401077224344897984675912636465197822254026739948964324640133571694642506863088696119636089570573034721904138769951712573343868448565169266453387940529052504268872190492455;
            6'd8: xpb[67] = 1024'd112090102483745555892385598981030650727922461174913663818460677676874283295263265959866746312747155789019494068121410503398003466740454626854916917120119868867964923509919809245766445078471517961088508799868036305218767601170457204201310089092751057992542871974504696953126681713820955616859069040586499480185;
            6'd9: xpb[67] = 1024'd79576354412666972354384201076854069789650858649626990247718816737117232955680247113594437896343922396605749798840026778355604959767553829753596484879010712126326535985070578899875911016461505560733248296706325900984478232483928064864606886598133896766553267191023887310977568900325337687546943985675213983584;
            6'd10: xpb[67] = 1024'd47062606341588388816382803172677488851379256124340316676976955797360182616097228267322129479940689004192005529558643053313206452794653032652276052637901555384688148460221348553985376954451493160377987793544615496750188863797398925527903684103516735540563662407543077668828456086829719758234818930763928486983;
            6'd11: xpb[67] = 1024'd14548858270509805278381405268500907913107653599053643106235094857603132276514209421049821063537455611778261260277259328270807945821752235550955620396792398643049760935372118208094842892441480760022727290382905092515899495110869786191200481608899574314574057624062268026679343273334101828922693875852642990382;
            6'd12: xpb[67] = 1024'd106101805883555963139178934769138759719534478199502653663625088982822977274240329484792583861791896528807666398453369037807473279690071773004795313172014282835102047980094105199834548021948674080977664395608434534645970976645237419819475848797511862355404356254698516414636758533767116916729258647566951978112;
            6'd13: xpb[67] = 1024'd73588057812477379601177536864962178781262875674215980092883228043065926934657310638520275445388663136393922129171985312765074772717170975903474880930905126093463660455244874853944013959938661680622403892446724130411681607958708280482772646302894701129414751471217706772487645720271498987417133592655666481511;
            6'd14: xpb[67] = 1024'd41074309741398796063176138960785597842991273148929306522141367103308876595074291792247967028985429743980177859890601587722676265744270178802154448689795969351825272930395644508053479897928649280267143389285013726177392239272179141146069443808277539903425146687736897130338532906775881058105008537744380984910;
            6'd15: xpb[67] = 1024'd8560561670320212525174741056609016904719670623642632951399506163551826255491272945975658612582196351566433590609217862680277758771369381700834016448686812610186885405546414162162945835918636879911882886123303321943102870585650001809366241313660378677435541904256087488189420093280263128792883482833095488309;
            6'd16: xpb[67] = 1024'd100113509283366370385972270557246868711146495224091643508789500288771671253217393009718421410836637268595838728785327572216943092639688919154673709223908696802239172450268401153902650965425830200866819991348832764073174352120017635437641608502272666718265840534892335876146835353713278216599448254547404476039;
            6'd17: xpb[67] = 1024'd67599761212287786847970872653070287772874892698804969938047639349014620913634374163446112994433403876182094459503943847174544585666788122053353276982799540060600784925419170808012116903415817800511559488187122359838884983433488496100938406007655505492276235751411526233997722540217660287287323199636118979438;
            6'd18: xpb[67] = 1024'd35086013141209203309969474748893706834603290173518296367305778409257570574051355317173804578030170483768350190222560122132146078693887324952032844741690383318962397400569940462121582841405805400156298985025411955604595614746959356764235203513038344266286630967930716591848609726722042357975198144724833482837;
            6'd19: xpb[67] = 1024'd2572265070130619771968076844717125896331687648231622796563917469500520234468336470901496161626937091354605920941176397089747571720986527850712412500581226577324009875720710116231048779395792999801038481863701551370306246060430217427532001018421183040297026184449906949699496913226424428663073089813547986236;
            6'd20: xpb[67] = 1024'd94125212683176777632765606345354977702758512248680633353953911594720365232194456534644258959881378008384011059117286106626412905589306065304552105275803110769376296920442697107970753908902986320755975587089230993500377727594797851055807368207033471081127324815086155337656912173659439516469637861527856973966;
            6'd21: xpb[67] = 1024'd61611464612098194094764208441178396764486909723393959783212050654963314892611437688371950543478144615970266789835902381584014398616405268203231673034693954027737909395593466762080219846892973920400715083927520589266088358908268711719104165712416309855137720031605345695507799360163821587157512806616571477365;
            6'd22: xpb[67] = 1024'd29097716541019610556762810537001815826215307198107286212470189715206264553028418842099642127074911223556522520554518656541615891643504471101911240793584797286099521870744236416189685784882961520045454580765810185031798990221739572382400963217799148629148115248124536053358686546668203657845387751705285980764;
            6'd23: xpb[67] = 1024'd120650664154065768417560340037639667632642131798556296769860183840426109550754538905842404925329352140585927658730628366078281225511824008555750933568806681478151808915466223407929390914390154841000391685991339627161870471756107206010676330406411436669978413878760784441316101807101218745651952523419594968494;
            6'd24: xpb[67] = 1024'd88136916082987184879558942133463086694370529273269623199118322900669059211171520059570096508926118748172183389449244641035882718538923211454430501327697524736513421390616993062038856852380142440645131182829629222927581103069578066673973127911794275443988809095279974799166988993605600816339827468508309471893;
            6'd25: xpb[67] = 1024'd55623168011908601341557544229286505756098926747982949628376461960912008871588501213297788092522885355758439120167860915993484211566022414353110069086588367994875033865767762716148322790370130040289870679667918818693291734383048927337269925417177114217999204311799165157017876180109982887027702413597023975292;
            6'd26: xpb[67] = 1024'd23109419940830017803556146325109924817827324222696276057634601021154958532005482367025479676119651963344694850886477190951085704593121617251789636845479211253236646340918532370257788728360117639934610176506208414459002365696519788000566722922559952992009599528318355514868763366614364957715577358685738478691;
            6'd27: xpb[67] = 1024'd114662367553876175664353675825747776624254148823145286615024595146374803529731602430768242474374092880374099989062586900487751038461441154705629329620701095445288933385640519361997493857867310960889547281731737856589073847230887421628842090111172241032839898158954603902826178627047380045522142130400047466421;
            6'd28: xpb[67] = 1024'd82148619482797592126352277921571195685982546297858613044282734206617753190148583584495934057970859487960355719781203175445352531488540357604308897379591938703650545860791289016106959795857298560534286778570027452354784478544358282292138887616555079806850293375473794260677065813551762116210017075488761969820;
            6'd29: xpb[67] = 1024'd49634871411719008588350880017394614747710943772571939473540873266860702850565564738223625641567626095546611450499819450402954024515639560502988465138482781962012158335942058670216425733847286160179026275408317048120495109857829142955435685121937918580860688591992984618527953000056144186897892020577476473219;
            6'd30: xpb[67] = 1024'd17121123340640425050349482113218033809439341247285265902799012327103652510982545891951317225164392703132867181218435725360555517542738763401668032897373625220373770811092828324325891671837273759823765772246606643886205741171300003618732482627320757354871083808512174976378840186560526257585766965666190976618;
            6'd31: xpb[67] = 1024'd108674070953686582911147011613855885615866165847734276460189006452323497508708665955694080023418833620162272319394545434897220851411058300855507725672595509412426057855814815316065596801344467080778702877472136086016277222705667637247007849815933045395701382439148423364336255446993541345392331737380499964348;
            6'd32: xpb[67] = 1024'd76160322882607999373145613709679304677594563322447602889447145512566447169125647109421771607015600227748528050113161709854822344438157503754187293431486352670787670330965584970175062739334454680423442374310425681781987854019138497910304647321315884169711777655667613722187142633497923416080206682469214467747;
            6'd33: xpb[67] = 1024'd43646574811529415835144215805502723739322960797160929318705284572809396829542628263149463190612366835334783780831777984812423837465256706652866861190377195929149282806116354624284528677324442280068181871148715277547698485332609358573601444826698722943722172872186804080038029820002305486768081627557928971146;
            6'd34: xpb[67] = 1024'd11132826740450832297142817901326142801051358271874255747963423633052346489959609416877154774209133442921039511550394259770025330492355909551546428949268039187510895281267124278393994615314429879712921367987004873313409116646080219236898242332081561717732568088705994437888917006506687557455956572646643474545;
            6'd35: xpb[67] = 1024'd102685774353496990157940347401963994607478182872323266305353417758272191487685729480619917572463574359950444649726503969306690664360675447005386121724489923379563182325989111270133699744821623200667858473212534315443480598180447852865173609520693849758562866719342242825846332266939702645262521344360952462275;
            6'd36: xpb[67] = 1024'd70172026282418406619938949497787413669206580347036592734611556818515141148102710634347609156060340967536700380445120244264292157387774649904065689483380766637924794801139880924243165682811610800312597970050823911209191229493918713528470407026076688532573261935861433183697219453444084715950396289449666965674;
            6'd37: xpb[67] = 1024'd37658278211339823081937551593610832730934977821749919163869695878758090808519691788075300739657107575122956111163736519221893650414873852802745257242271609896286407276290650578352631620801598399957337466889113506974901860807389574191767204531459527306583657152380623541548106639948466786638271234538381469073;
            6'd38: xpb[67] = 1024'd5144530140261239543936153689434251792663375296463245593127834939001040468936672941802992323253874182709211841882352794179495143441973055701424825001162453154648019751441420232462097558791585999602076963727403102740612492120860434855064002036842366080594052368899813899398993826452848857326146179627095972472;
            6'd39: xpb[67] = 1024'd96697477753307397404733683190072103599090199896912256150517829064220885466662793005545755121508315099738616980058462503716160477310292593155264517776384337346700306796163407224201802688298779320557014068952932544870683973655228068483339369225454654121424350999536062287356409086885863945132710951341404960202;
            6'd40: xpb[67] = 1024'd64183729682228813866732285285895522660818597371625582579775968124463835127079774159273446705105081707324872710777078778673761970337391796053944085535275180605061919271314176878311268626288766920201753565791222140636394604968698929146636166730837492895434746216055252645207296273390246015820585896430119463601;
            6'd41: xpb[67] = 1024'd31669981611150230328730887381718941722546994846338909009034107184706784787496755313001138288701848314911128441495695053631363463364490998952623653294166023863423531746464946532420734564278754519846493062629511736402105236282169789809932964236220331669445141432574443003058183459894628086508460841518833967000;
            6'd42: xpb[67] = 1024'd123222929224196388189528416882356793528973819446787919566424101309926629785222875376743901086956289231940533579671804763168028797232810536406463346069387908055475818791186933524160439693785947840801430167855041178532176717816537423438208331424832619710275440063210691391015598720327643174315025613233142954730;
            6'd43: xpb[67] = 1024'd90709181153117804651527018978180212590702216921501245995682240370169579445639856530471592670553055839526789310390421038125630290259909739305142913828278751313837431266337703178269905631775935440446169664693330774297887349130008284101505128930215458484285835279729881748866485906832025245002900558321857458129;
            6'd44: xpb[67] = 1024'd58195433082039221113525621074003631652430614396214572424940379430412529106056837684199284254149822447113045041109037313083231783287008942203822481587169594572199043741488472832379371569765923040090909161531620370063597980443479144764801926435598297258296230496249072106717373093336407315690775503410571961528;
            6'd45: xpb[67] = 1024'd25681685010960637575524223169827050714159011870927898854198518490655478766473818837926975837746589054699300771827653588040833276314108145102502049346060437830560656216639242486488837507755910639735648658369909965829308611756950005428098723940981136032306625712768262464568260279840789386378650448499286464927;
            6'd46: xpb[67] = 1024'd117234632624006795436321752670464902520585836471376909411588512615875323764199938901669738636001029971728705910003763297577498610182427682556341742121282322022612943261361229478228542637263103960690585763595439407959380093291317639056374091129593424073136924343404510852525675540273804474185215220213595452657;
            6'd47: xpb[67] = 1024'd84720884552928211898320354766288321582314233946090235840846651676118273424616920055397430219597796579314961640722379572535100103209526885455021309880173165280974555736511999132338008575253091560335325260433729003725090724604788499719670888634976262847147319559923701210376562726778186544873090165302309956056;
            6'd48: xpb[67] = 1024'd52207136481849628360318956862111740644042631420803562270104790736361223085033901209125121803194563186901217371440995847492701596236626088353700877639064008539336168211662768786447474513243079159980064757272018599490801355918259360382967686140359101621157714776442891568227449913282568615560965110391024459455;
            6'd49: xpb[67] = 1024'd19693388410771044822317558957935159705771028895516888699362929796604172745450882362852813386791329794487473102159612122450303089263725291252380445397954851797697780686813538440556940451233066759624804254110308195256511987231730221046264483645741940395168109992962081926078337099786950686248840055479738962854;
            6'd50: xpb[67] = 1024'd111246336023817202683115088458573011512197853495965899256752923921824017743177002426595576185045770711516878240335721831986968423132044828706220138173176735989750067731535525432296645580740260080579741359335837637386583468766097854674539850834354228435998408623598330314035752360219965774055404827194047950584;
            6'd51: xpb[67] = 1024'd78732587952738619145113690554396430573926250970679225686011062982066967403593983580323267768642537319103133971054338106944569916159144031604899705932067579248111680206686295086406111518730247680224480856174127233152294100079568715337836648339737067210008803840117520671886639546724347844743279772282762453983;
            6'd52: xpb[67] = 1024'd46218839881660035607112292650219849635654648445392552115269202042309917064010964734050959352239303926689389701772954381902171409186243234503579273690958422506473292681837064740515577456720235279869220353012416828918004731393039576001133445845119905984019199056636711029737526733228729915431154717371476957382;
            6'd53: xpb[67] = 1024'd13705091810581452069110894746043268697383045920105878544527341102552866724427945887778650935836070534275645432491570656859772902213342437402258841449849265764834905156987834394625043394710222879513959849850706424683715362706510436664430243350502744758029594273155901387588413919733111986119029662460191460781;
            6'd54: xpb[67] = 1024'd105258039423627609929908424246681120503809870520554889101917335227772711722154065951521413734090511451305050570667680366396438236081661974856098534225071149956887192201709821386364748524217416200468896955076235866813786844240878070292705610539115032798859892903792149775545829180166127073925594434174500448511;
            6'd55: xpb[67] = 1024'd72744291352549026391907026342504539565538267995268215531175474288015661382571047105249105317687278058891306301386296641354039729108761177754778101983961993215248804676860591040474214462207403800113636451914525462579497475554348930956002408044497871572870288120311340133396716366670509144613469379263214951910;
            6'd56: xpb[67] = 1024'd40230543281470442853905628438327958627266665469981541960433613348258611042988028258976796901284044666477562032104912916311641222135860380653457669742852836473610417152011360694583680400197391399758375948752815058345208106867819791619299205549880710346880683336830530491247603553174891215301344324351929455309;
            6'd57: xpb[67] = 1024'd7716795210391859315904230534151377688995062944694868389691752408501560703405009412704488484880811274063817762823529191269242715162959583552137237501743679731972029627162130348693146338187378999403115445591104654110918738181290652282596003055263549120891078553349720849098490739679273285989219269440643958708;
            6'd58: xpb[67] = 1024'd99269742823438017176701760034789229495421887545143878947081746533721405701131129476447251283135252191093222900999638900805908049031279121005976930276965563924024316671884117340432851467694572320358052550816634096240990219715658285910871370243875837161721377183985969237055906000112288373795784041154952946438;
            6'd59: xpb[67] = 1024'd66755994752359433638700362130612648557150285019857205376339885593964355361548110630174942866732018798679478631718255175763509542058378323904656498035856407182385929147034886994542317405684559920002792047654923692006700851029129146574168167749258675935731772400505159594906793186616670444483658986243667449837;
            6'd60: xpb[67] = 1024'd34242246681280850100698964226436067618878682494570531805598024654207305021965091783902634450328785406265734362436871450721111035085477526803336065794747250440747541622185656648651783343674547519647531544493213287772411482342600007237464965254641514709742167617024349952757680373121052515171533931332381953236;
            6'd61: xpb[67] = 1024'd1728498610202266562697566322259486680607079969283858234856163714450254682382072937630326033925552013851990093155487725678712528112576729702015633553638093699109154097336426302761249281664535119292271041331502883538122113656070867900761762760024353483752562833543540310608567559625434585859408876421096456635;
            6'd62: xpb[67] = 1024'd93281446223248424423495095822897338487033904569732868792246157839670099680108193001373088832179992930881395231331597435215377861980896267155855326328859977891161441142058413294500954411171728440247208146557032325668193595190438501529037129948636641524582861464179788698565982820058449673665973648135405444365;
            6'd63: xpb[67] = 1024'd60767698152169840885493697918720757548762302044446195221504296899913049340525174155100780415776759538467650962050213710172979355007995470054534894087750821149523053617209182948610420349161716039891947643395321921433904226503909362192333927454019480298593256680698979056416870006562831744353848593224119947764;
        endcase
    end

    always_comb begin
        case(flag[22][16:12])
            5'd0: xpb[68] = 1024'd0;
            5'd1: xpb[68] = 1024'd28253950081091257347492300014544176610490699519159521650762435960155999000942155308828471999373526146053906692768829985130580848035094672953214461846641664407884666092359952602719886287151703639536687140233611517199614857817380222855630724959402319072603651897218169414267757193067213815041723538312834451163;
            5'd2: xpb[68] = 1024'd56507900162182514694984600029088353220981399038319043301524871920311998001884310617656943998747052292107813385537659970261161696070189345906428923693283328815769332184719905205439772574303407279073374280467223034399229715634760445711261449918804638145207303794436338828535514386134427630083447076625668902326;
            5'd3: xpb[68] = 1024'd84761850243273772042476900043632529831472098557478564952287307880467997002826465926485415998120578438161720078306489955391742544105284018859643385539924993223653998277079857808159658861455110918610061420700834551598844573452140668566892174878206957217810955691654508242803271579201641445125170614938503353489;
            5'd4: xpb[68] = 1024'd113015800324365029389969200058176706441962798076638086603049743840623996003768621235313887997494104584215626771075319940522323392140378691812857847386566657631538664369439810410879545148606814558146748560934446068798459431269520891422522899837609276290414607588872677657071028772268855260166894153251337804652;
            5'd5: xpb[68] = 1024'd17203054721331545338662572667906450307755070470061924125680324735803099667401637634127288782209956420826384056386656491073840399334253030210912184216877281105732655892228545675969192244241312476373238092780817739633713438866004341313175055113782146096198356071973789041232257891407436058089927864938577771484;
            5'd6: xpb[68] = 1024'd45457004802422802686154872682450626918245769989221445776442760695959098668343792942955760781583482566880290749155486476204421247369347703164126646063518945513617321984588498278689078531393016115909925233014429256833328296683384564168805780073184465168802007969191958455500015084474649873131651403251412222647;
            5'd7: xpb[68] = 1024'd73710954883514060033647172696994803528736469508380967427205196656115097669285948251784232780957008712934197441924316461335002095404442376117341107910160609921501988076948450881408964818544719755446612373248040774032943154500764787024436505032586784241405659866410127869767772277541863688173374941564246673810;
            5'd8: xpb[68] = 1024'd101964904964605317381139472711538980139227169027540489077967632616271096670228103560612704780330534858988104134693146446465582943439537049070555569756802274329386654169308403484128851105696423394983299513481652291232558012318145009880067229991989103314009311763628297284035529470609077503215098479877081124973;
            5'd9: xpb[68] = 1024'd6152159361571833329832845321268724005019441420964326600598213511450200333861119959426105565046386695598861420004482997017099950633411387468609906587112897803580645692097138749218498201330921313209789045328023962067812019914628459770719385268161973119793060246729408668196758589747658301138132191564321091805;
            5'd10: xpb[68] = 1024'd34406109442663090677325145335812900615510140940123848251360649471606199334803275268254577564419912841652768112773312982147680798668506060421824368433754562211465311784457091351938384488482624952746476185561635479267426877732008682626350110227564292192396712143947578082464515782814872116179855729877155542968;
            5'd11: xpb[68] = 1024'd62660059523754348024817445350357077226000840459283369902123085431762198335745430577083049563793438987706674805542142967278261646703600733375038830280396226619349977876817043954658270775634328592283163325795246996467041735549388905481980835186966611265000364041165747496732272975882085931221579268189989994131;
            5'd12: xpb[68] = 1024'd90914009604845605372309745364901253836491539978442891552885521391918197336687585885911521563166965133760581498310972952408842494738695406328253292127037891027234643969176996557378157062786032231819850466028858513666656593366769128337611560146368930337604015938383916911000030168949299746263302806502824445294;
            5'd13: xpb[68] = 1024'd119167959685936862719802045379445430446982239497602413203647957352074196337629741194739993562540491279814488191079802937539423342773790079281467753973679555435119310061536949160098043349937735871356537606262470030866271451184149351193242285105771249410207667835602086325267787362016513561305026344815658896457;
            5'd14: xpb[68] = 1024'd23355214082903378668495417989175174312774511891026250726278538247253300001262757593553394347256343116425245476391139488090940349967664417679522090803990178909313301584325684425187690445572233789583027138108841701701525458780632801083894440381944119215991416318703197709429016481155094359228060056502898863289;
            5'd15: xpb[68] = 1024'd51609164163994636015987718003719350923265211410185772377040974207409299002204912902381866346629869262479152169159969473221521198002759090632736552650631843317197967676685637027907576732723937429119714278342453218901140316598013023939525165341346438288595068215921367123696773674222308174269783594815733314452;
            5'd16: xpb[68] = 1024'd79863114245085893363480018018263527533755910929345294027803410167565298003147068211210338346003395408533058861928799458352102046037853763585951014497273507725082633769045589630627463019875641068656401418576064736100755174415393246795155890300748757361198720113139536537964530867289521989311507133128567765615;
            5'd17: xpb[68] = 1024'd108117064326177150710972318032807704144246610448504815678565846127721297004089223520038810345376921554586965554697629443482682894072948436539165476343915172132967299861405542233347349307027344708193088558809676253300370032232773469650786615260151076433802372010357705952232288060356735804353230671441402216778;
            5'd18: xpb[68] = 1024'd12304318723143666659665690642537448010038882841928653201196427022900400667722239918852211130092773391197722840008965994034199901266822774937219813174225795607161291384194277498436996402661842626419578090656047924135624039829256919541438770536323946239586120493458817336393517179495316602276264383128642183610;
            5'd19: xpb[68] = 1024'd40558268804234924007157990657081624620529582361088174851958862983056399668664395227680683129466299537251629532777795979164780749301917447890434275020867460015045957476554230101156882689813546265956265230889659441335238897646637142397069495495726265312189772390676986750661274372562530417317987921441476634773;
            5'd20: xpb[68] = 1024'd68812218885326181354650290671625801231020281880247696502721298943212398669606550536509155128839825683305536225546625964295361597337012120843648736867509124422930623568914182703876768976965249905492952371123270958534853755464017365252700220455128584384793424287895156164929031565629744232359711459754311085936;
            5'd21: xpb[68] = 1024'd97066168966417438702142590686169977841510981399407218153483734903368397670548705845337627128213351829359442918315455949425942445372106793796863198714150788830815289661274135306596655264116953545029639511356882475734468613281397588108330945414530903457397076185113325579196788758696958047401434998067145537099;
            5'd22: xpb[68] = 1024'd1253423363383954650835963295899721707303253792831055676114315798547501334181722244151027912929203665970200203626792499977459452565981132194917535544461412305009281184062870571686302359751451463256129043203254146569722620877881037998983100690703773263180824668214436963358017877835538845324468709754385503931;
            5'd23: xpb[68] = 1024'd29507373444475211998328263310443898317793953311990577326876751758703500335123877552979499912302729812024106896395622485108040300601075805148131997391103076712893947276422823174406188646903155102792816183436865663769337478695261260854613825650106092335784476565432606377625775070902752660366192248067219955094;
            5'd24: xpb[68] = 1024'd57761323525566469345820563324988074928284652831150098977639187718859499336066032861807971911676255958078013589164452470238621148636170478101346459237744741120778613368782775777126074934054858742329503323670477180968952336512641483710244550609508411408388128462650775791893532263969966475407915786380054406257;
            5'd25: xpb[68] = 1024'd86015273606657726693312863339532251538775352350309620628401623679015498337008188170636443911049782104131920281933282455369201996671265151054560921084386405528663279461142728379845961221206562381866190463904088698168567194330021706565875275568910730480991780359868945206161289457037180290449639324692888857420;
            5'd26: xpb[68] = 1024'd114269223687748984040805163354076428149266051869469142279164059639171497337950343479464915910423308250185826974702112440499782844706359824007775382931028069936547945553502680982565847508358266021402877604137700215368182052147401929421506000528313049553595432257087114620429046650104394105491362863005723308583;
            5'd27: xpb[68] = 1024'd18456478084715499989498535963806172015058324262892979801794640534350601001583359878278316695139160086796584260013448991051299851900234162405829719761338693410741937076291416247655494603992763939629367135984071886203436059743885379312158155804485919359379180740188226004590275769242974903414396574692963275415;
            5'd28: xpb[68] = 1024'd46710428165806757336990835978350348625549023782052501452557076494506600002525515187106788694512686232850490952782278976181880699935328835359044181607980357818626603168651368850375380891144467579166054276217683403403050917561265602167788880763888238431982832637406395418858032962310188718456120113005797726578;
            5'd29: xpb[68] = 1024'd74964378246898014684483135992894525236039723301212023103319512454662599003467670495935260693886212378904397645551108961312461547970423508312258643454622022226511269261011321453095267178296171218702741416451294920602665775378645825023419605723290557504586484534624564833125790155377402533497843651318632177741;
            5'd30: xpb[68] = 1024'd103218328327989272031975436007438701846530422820371544754081948414818598004409825804763732693259738524958304338319938946443042396005518181265473105301263686634395935353371274055815153465447874858239428556684906437802280633196026047879050330682692876577190136431842734247393547348444616348539567189631466628904;
            5'd31: xpb[68] = 1024'd7405582724955787980668808617168445712322695213795382276712529309997701668042842203577133477975590361569061623631275496994559403199392519663527442131574310108589926876160009320904800561082372776465918088531278108637534640792509497769702485958865746382973884914943845631554776467583197146462600901318706595736;
        endcase
    end

    always_comb begin
        case(flag[23][5:0])
            6'd0: xpb[69] = 1024'd0;
            6'd1: xpb[69] = 1024'd79863114245085893363480018018263527533755910929345294027803410167565298003147068211210338346003395408533058861928799458352102046037853763585951014497273507725082633769045589630627463019875641068656401418576064736100755174415393246795155890300748757361198720113139536537964530867289521989311507133128567765615;
            6'd2: xpb[69] = 1024'd35659532806047045328161108631712622322813394732954903927474965270153700668984997512405605477349116507622968316400105482125140251234487192616741903978215974516474592968519961923624686848234076416002605228764889625837149498609889720625333210918268065455577536812162015045822533660650410961504324439631541046899;
            6'd3: xpb[69] = 1024'd115522647051132938691641126649976149856569305662300197955278375437718998672132065723615943823352511916156027178328904940477242297272340956202692918475489482241557226737565551554252149868109717484659006647340954361937904673025282967420489101219016822816776256925301551583787064527939932950815831572760108812514;
            6'd4: xpb[69] = 1024'd71319065612094090656322217263425244645626789465909807854949930540307401337969995024811210954698233015245936632800210964250280502468974385233483807956431949032949185937039923847249373696468152832005210457529779251674298997219779441250666421836536130911155073624324030091645067321300821923008648879263082093798;
            6'd5: xpb[69] = 1024'd27115484173055242621003307876874339434684273269519417754621485642895804003807924326006478086043954114335846087271516988023318707665607814264274697437374415824341145136514296140246597524826588179351414267718604141410693321414275915080843742454055439005533890323346508599503070114661710895201466185766055375082;
            6'd6: xpb[69] = 1024'd106978598418141135984483325895137866968440184198864711782424895810461102006954992537216816432047349522868904949200316446375420753703461577850225711934647923549423778905559885770874060544702229248007815686294668877511448495829669161875999632754804196366732610436486045137467600981951232884512973318894623140697;
            6'd7: xpb[69] = 1024'd62775016979102287949164416508586961757497668002474321682096450913049504672792921838412083563393070621958814403671622470148458958900095006881016601415590390340815738105034258063871284373060664595354019496483493767247842820024165635706176953372323504461111427135508523645325603775312121856705790625397596421981;
            6'd8: xpb[69] = 1024'd18571435540063439913845507122036056546555151806083931581768006015637907338630851139607350694738791721048723858142928493921497164096728435911807490896532857132207697304508630356868508201419099942700223306672318656984237144218662109536354273989842812555490243834531002153183606568673010828898607931900569703265;
            6'd9: xpb[69] = 1024'd98434549785149333277325525140299584080311062735429225609571416183203205341777919350817689040742187129581782720071727952273599210134582199497758505393806364857290331073554219987495971221294741011356624725248383393084992318634055356331510164290591569916688963947670538691148137435962532818210115065029137468880;
            6'd10: xpb[69] = 1024'd54230968346110485242006615753748678869368546539038835509242971285791608007615848652012956172087908228671692174543033976046637415331215628528549394874748831648682290273028592280493195049653176358702828535437208282821386642828551830161687484908110878011067780646693017199006140229323421790402932371532110750164;
            6'd11: xpb[69] = 1024'd10027386907071637206687706367197773658426030342648445408914526388380010673453777953208223303433629327761601629014339999819675620527849057559340284355691298440074249472502964573490418878011611706049032345626033172557780967023048303991864805525630186105446597345715495706864143022684310762595749678035084031448;
            6'd12: xpb[69] = 1024'd89890501152157530570167724385461301192181941271993739436717936555945308676600846164418561649437024736294660490943139458171777666565702821145291298852964806165156883241548554204117881897887252774705433764202097908658536141438441550787020695826378943466645317458855032244828673889973832751907256811163651797063;
            6'd13: xpb[69] = 1024'd45686919713118682534848814998910395981239425075603349336389491658533711342438775465613828780782745835384569945414445481944815871762336250176082188333907272956548842441022926497115105726245688122051637574390922798394930465632938024617198016443898251561024134157877510752686676683334721724100074117666625078347;
            6'd14: xpb[69] = 1024'd1483338274079834499529905612359490770296908879212959236061046761122114008276704766809095912128466934474479399885751505717854076958969679206873077814849739747940801640497298790112329554604123469397841384579747688131324789827434498447375337061417559655402950856899989260544679476695610696292891424169598359631;
            6'd15: xpb[69] = 1024'd81346452519165727863009923630623018304052819808558253263864456928687412011423772978019434258131862343007538261814550964069956122996823442792824092312123247473023435409542888420739792574479764538054242803155812424232079964242827745242531227362166317016601670970039525798509210343985132685604398557298166125246;
            6'd16: xpb[69] = 1024'd37142871080126879827691014244072113093110303612167863163536012031275814677261702279214701389477583442097447716285856987842994328193456871823614981793065714264415394609017260713737016402838199885400446613344637313968474288437324219072708547979685625110980487669062004306367213137346021657797215863801139406530;
            6'd17: xpb[69] = 1024'd117005985325212773191171032262335640626866214541513157191339422198841112680408770490425039735480978850630506578214656446195096374231310635409565996290339221989498028378062850344364479422713840954056848031920702050069229462852717465867864438280434382472179207782201540844331744004635543647108722996929707172145;
            6'd18: xpb[69] = 1024'd72802403886173925155852122875784735415923698345122767091010977301429515346246699791620306866826699949720416032685962469968134579427944064440356885771281688780889987577537222637361703251072276301403051842109526939805623787047213939698041758897953690566558024481224019352189746797996432619301540303432680453429;
            6'd19: xpb[69] = 1024'd28598822447135077120533213489233830204981182148732376990682532404017918012084629092815573998172421048810325487157268493741172784624577493471147775252224155572281946777011594930358927079430711648749255652298351829542018111241710413528219079515472998660936841180246497860047749591357321591494357609935653734713;
            6'd20: xpb[69] = 1024'd108461936692220970484013231507497357738737093078077671018485942571583216015231697304025912344175816457343384349086067952093274830662431257057098789749497663297364580546057184560986390099306352717405657070874416565642773285657103660323374969816221756022135561293386034398012280458646843580805864743064221500328;
            6'd21: xpb[69] = 1024'd64258355253182122448694322120946452527794576881687280918157497674171618681069626605221179475521537556433293803557373975866313035859064686087889679230440130088756539745531556853983613927664788064751860881063241455379167609851600134153552290433741064116514377992408512905870283252007732552998682049567194781612;
            6'd22: xpb[69] = 1024'd20054773814143274413375412734395547316852060685296890817829052776760021346907555906416446606867258655523203258028679999639351241055698115118680568711382596880148498945005929146980837756023223412098064691252066345115561934046096607983729611051260372210893194691430991413728286045368621525191499356070168062896;
            6'd23: xpb[69] = 1024'd99917888059229167776855430752659074850607971614642184845632462944325319350054624117626784952870654064056262119957479457991453287093551878704631583208656104605231132714051518777608300775898864480754466109828131081216317108461489854778885501352009129572091914804570527951692816912658143514503006489198735828511;
            6'd24: xpb[69] = 1024'd55714306620190319741536521366108169639665455418251794745304018046913722015892553418822052084216375163146171574428785481764491492290185307735422472689598571396623091913525891070605524604257299828100669920016955970952711432655986328609062821969528437666470731503593006459550819706019032486695823795701709109795;
            6'd25: xpb[69] = 1024'd11510725181151471706217611979557264428722939221861404644975573149502124681730482720017319215562096262236081028900091505537529697486818736766213362170541038188015051113000263363602748432615735175446873730205780860689105756850482802439240142587047745760849548202615484967408822499379921458888641102204682391079;
            6'd26: xpb[69] = 1024'd91373839426237365069697629997820791962478850151206698672778983317067422684877550931227657561565491670769139890828890963889631743524672500352164376667814545913097684882045852994230211452491376244103275148781845596789860931265876049234396032887796503122048268315755021505373353366669443448200148235333250156694;
            6'd27: xpb[69] = 1024'd47170257987198517034378720611269886751536333954816308572450538419655825350715480232422924692911212769859049345300196987662669948721305929382955266148757012704489644081520225287227435280849811591449478958970670486526255255460372523064573353505315811216427085014777500013231356160030332420392965541836223437978;
            6'd28: xpb[69] = 1024'd2966676548159668999059811224718981540593817758425918472122093522244228016553409533618191824256933868948958799771503011435708153917939358413746155629699479495881603280994597580224659109208246938795682769159495376262649579654868996894750674122835119310805901713799978521089358953391221392585782848339196719262;
            6'd29: xpb[69] = 1024'd82829790793245562362539829242982509074349728687771212499925503689809526019700477744828530170260329277482017661700302469787810199955793121999697170126972987220964237050040187210852122129083888007452084187735560112363404754070262243689906564423583876672004621826939515059053889820680743381897289981467764484877;
            6'd30: xpb[69] = 1024'd38626209354206714327220919856431603863407212491380822399597058792397928685538407046023797301606050376571927116171608493560848405152426551030488059607915454012356196249514559503849345957442323354798287997924385002099799078264758717520083885041103184766383438525961993566911892614041632354090107287970737766161;
            6'd31: xpb[69] = 1024'd118489323599292607690700937874695131397163123420726116427400468959963226688685475257234135647609445785104985978100407951912950451190280314616439074105188961737438830018560149134476808977317964423454689416500449738200554252680151964315239775341851942127582158639101530104876423481331154343401614421099305531776;
            6'd32: xpb[69] = 1024'd74285742160253759655382028488144226186220607224335726327072024062551629354523404558429402778955166884194895432571713975685988656386913743647229963586131428528830789218034521427474032805676399770800893226689274627936948576874648438145417095959371250221960975338124008612734426274692043315594431727602278813060;
            6'd33: xpb[69] = 1024'd30082160721214911620063119101593320975278091027945336226743579165140032020361333859624669910300887983284804887043019999459026861583547172678020853067073895320222748417508893720471256634034835118147097036878099517673342901069144911975594416576890558316339792037146487120592429068052932287787249034105252094344;
            6'd34: xpb[69] = 1024'd109945274966300804983543137119856848509034001957290630254546989332705330023508402070835008256304283391817863748971819457811128907621400936263971867564347403045305382186554483351098719653910476186803498455454164253774098075484538158770750306877639315677538512150286023658556959935342454277098756167233819859959;
            6'd35: xpb[69] = 1024'd65741693527261956948224227733305943298091485760900240154218544435293732689346331372030275387650004490907773203443125481584167112818034365294762757045289869836697341386028855644095943482268911534149702265642989143510492399679034632600927627495158623771917328849308502166414962728703343249291573473736793141243;
            6'd36: xpb[69] = 1024'd21538112088223108912905318346755038087148969564509850053890099537882135355184260673225542518995725589997682657914431505357205318014667794325553646526232336628089300585503227937093167310627346881495906075831814033246886723873531106431104948112677931866296145548330980674272965522064232221484390780239766422527;
            6'd37: xpb[69] = 1024'd101401226333309002276385336365018565620904880493855144081693509705447433358331328884435880864999120998530741519843230963709307364052521557911504661023505844353171934354548817567720630330502987950152307494407878769347641898288924353226260838413426689227494865661470517212237496389353754210795897913368334188142;
            6'd38: xpb[69] = 1024'd57197644894270154241066426978467660409962364297464753981365064808035836024169258185631147996344842097620650974314536987482345569249154986942295550504448311144563893554023189860717854158861423297498511304596703659084036222483420827056438159030945997321873682360492995720095499182714643182988715219871307469426;
            6'd39: xpb[69] = 1024'd12994063455231306205747517591916755199019848101074363881036619910624238690007187486826415127690563196710560428785843011255383774445788415973086439985390777935955852753497562153715077987219858644844715114785528548820430546677917300886615479648465305416252499059515474227953501976075532155181532526374280750710;
            6'd40: xpb[69] = 1024'd92857177700317199569227535610180282732775759030419657908840030078189536693154255698036753473693958605243619290714642469607485820483642179559037454482664285661038486522543151784342541007095499713501116533361593284921185721093310547681771369949214062777451219172655010765918032843365054144493039659502848516325;
            6'd41: xpb[69] = 1024'd48653596261278351533908626223629377521833242834029267808511585180777939358992184999232020605039679704333528745185948493380524025680275608589828343963606752452430445722017524077339764835453935060847320343550418174657580045287807021511948690566733370871830035871677489273776035636725943116685856966005821797609;
            6'd42: xpb[69] = 1024'd4450014822239503498589716837078472310890726637638877708183140283366342024830114300427287736385400803423438199657254517153562230876909037620619233444549219243822404921491896370336988663812370408193524153739243064393974369482303495342126011184252678966208852570699967781634038430086832088878674272508795078893;
            6'd43: xpb[69] = 1024'd84313129067325396862069734855341999844646637566984171735986550450931640027977182511637626082388796211956497061586053975505664276914762801206570247941822726968905038690537486000964451683688011476849925572315307800494729543897696742137281901485001436327407572683839504319598569297376354078190181405637362844508;
            6'd44: xpb[69] = 1024'd40109547628286548826750825468791094633704121370593781635658105553520042693815111812832893213734517311046406516057359999278702482111396230237361137422765193760296997890011858293961675512046446824196129382504132690231123868092193215967459222102520744421786389382861982827456572090737243050382998712140336125792;
            6'd45: xpb[69] = 1024'd119972661873372442190230843487054622167460032299939075663461515721085340696962180024043231559737912719579465377986159457630804528149249993823312151920038701485379631659057447924589138531922087892852530801080197426331879042507586462762615112403269501782985109496001519365421102958026765039694505845268903891407;
            6'd46: xpb[69] = 1024'd75769080434333594154911934100503716956517516103548685563133070823673743362800109325238498691083633818669374832457465481403842733345883422854103041400981168276771590858531820217586362360280523240198734611269022316068273366702082936592792433020788809877363926195023997873279105751387654011887323151771877172691;
            6'd47: xpb[69] = 1024'd31565498995294746119593024713952811745574999907158295462804625926262146028638038626433765822429354917759284286928771505176880938542516851884893930881923635068163550058006192510583586188638958587544938421457847205804667690896579410422969753638308117971742742894046476381137108544748542984080140458274850453975;
            6'd48: xpb[69] = 1024'd111428613240380639483073042732216339279330910836503589490608036093827444031785106837644104168432750326292343148857570963528982984580370615470844945379197142793246183827051782141211049208514599656201339840033911941905422865311972657218125643939056875332941463007186012919101639412038064973391647591403418219590;
            6'd49: xpb[69] = 1024'd67225031801341791447754133345665434068388394640113199390279591196415846697623036138839371299778471425382252603328876987302021189777004044501635834860139609584638143026526154434208273036873035003547543650222736831641817189506469131048302964556576183427320279706208491426959642205398953945584464897906391500874;
            6'd50: xpb[69] = 1024'd23021450362302943412435223959114528857445878443722809289951146299004249363460965440034638431124192524472162057800183011075059394973637473532426724341082076376030102226000526727205496865231470350893747460411561721378211513700965604878480285174095491521699096405230969934817644998759842917777282204409364782158;
            6'd51: xpb[69] = 1024'd102884564607388836775915241977378056391201789373068103317754556466569547366608033651244976777127587933005220919728982469427161441011491237118377738838355584101112735995046116357832959885107111419550148878987626457478966688116358851673636175474844248882897816518370506472782175866049364907088789337537932547773;
            6'd52: xpb[69] = 1024'd58680983168349988740596332590827151180259273176677713217426111569157950032445962952440243908473309032095130374200288493200199646208124666149168628319298050892504695194520488650830183713465546766896352689176451347215361012310855325503813496092363556977276633217392984980640178659410253879281606644040905829057;
            6'd53: xpb[69] = 1024'd14477401729311140705277423204276245969316756980287323117097666671746352698283892253635511039819030131185039828671594516973237851404758095179959517800240517683896654393994860943827407541823982114242556499365276236951755336505351799333990816709882865071655449916415463488498181452771142851474423950543879110341;
            6'd54: xpb[69] = 1024'd94340515974397034068757441222539773503072667909632617144901076839311650701430960464845849385822425539718098690600393975325339897442611858765910532297514025408979288163040450574454870561699623182898957917941340973052510510920745046129146707010631622432854170029555000026462712320060664840785931083672446875956;
            6'd55: xpb[69] = 1024'd50136934535358186033438531835988868292130151713242227044572631941900053367268889766041116517168146638808008145071699999098378102639245287796701421778456492200371247362514822867452094390058058530245161728130165862788904835115241519959324027628150930527232986728577478534320715113421553812978748390175420157240;
            6'd56: xpb[69] = 1024'd5933353096319337998119622449437963081187635516851836944244187044488456033106819067236383648513867737897917599543006022871416307835878716827492311259398958991763206561989195160449318218416493877591365538318990752525299159309737993789501348245670238621611803427599957042178717906782442785171565696678393438524;
            6'd57: xpb[69] = 1024'd85796467341405231361599640467701490614943546446197130972047597212053754036253887278446721994517263146430976461471805481223518353873732480413443325756672466716845840331034784791076781238292134946247766956895055488626054333725131240584657238546418995982810523540739493580143248774071964774483072829806961204139;
            6'd58: xpb[69] = 1024'd41592885902366383326280731081150585404001030249806740871719152314642156702091816579641989125862984245520885915943111504996556559070365909444234215237614933508237799530509157084074005066650570293593970767083880378362448657919627714414834559163938304077189340239761972088001251567432853746675890136309934485423;
            6'd59: xpb[69] = 1024'd121456000147452276689760749099414112937756941179152034899522562482207454705238884790852327471866379654053944777871910963348658605108219673030185229734888441233320433299554746714701468086526211362250372185659945114463203832335020961209990449464687061438388060352901508625965782434722375735987397269438502251038;
            6'd60: xpb[69] = 1024'd77252418708413428654441839712863207726814424982761644799194117584795857371076814092047594603212100753143854232343216987121696810304853102060976119215830908024712392499029119007698691914884646709596575995848770004199598156529517435040167770082206369532766877051923987133823785228083264708180214575941475532322;
            6'd61: xpb[69] = 1024'd33048837269374580619122930326312302515871908786371254698865672687384260036914743393242861734557821852233763686814523010894735015501486531091767008696773374816104351698503491300695915743243082056942779806037594893935992480724013908870345090699725677627145693750946465641681788021444153680373031882444448813606;
            6'd62: xpb[69] = 1024'd112911951514460473982602948344575830049627819715716548726669082854949558040061811604453200080561217260766822548743322469246837061539340294677718023194046882541186985467549080931323378763118723125599181224613659630036747655139407155665500981000474434988344413864086002179646318888733675669684539015573016579221;
            6'd63: xpb[69] = 1024'd68708370075421625947284038958024924838685303519326158626340637957537960705899740905648467211906938359856732003214628493019875266735973723708508912674989349332578944667023453224320602591477158472945385034802484519773141979333903629495678301617993743082723230563108480687504321682094564641877356322075989860505;
        endcase
    end

    always_comb begin
        case(flag[23][11:6])
            6'd0: xpb[70] = 1024'd0;
            6'd1: xpb[70] = 1024'd24504788636382777911965129571474019627742787322935768526012193060126363371737670206843734343252659458946641457685934516792913471932607152739299802155931816123970903866497825517317826419835593820291588844991309409509536303528400103325855622235513051177102047262130959195362324475455453614070173628578963141789;
            6'd2: xpb[70] = 1024'd49009577272765555823930259142948039255485574645871537052024386120252726743475340413687468686505318917893282915371869033585826943865214305478599604311863632247941807732995651034635652839671187640583177689982618819019072607056800206651711244471026102354204094524261918390724648950910907228140347257157926283578;
            6'd3: xpb[70] = 1024'd73514365909148333735895388714422058883228361968807305578036579180379090115213010620531203029757978376839924373057803550378740415797821458217899406467795448371912711599493476551953479259506781460874766534973928228528608910585200309977566866706539153531306141786392877586086973426366360842210520885736889425367;
            6'd4: xpb[70] = 1024'd98019154545531111647860518285896078510971149291743074104048772240505453486950680827374937373010637835786565830743738067171653887730428610957199208623727264495883615465991302069271305679342375281166355379965237638038145214113600413303422488942052204708408189048523836781449297901821814456280694514315852567156;
            6'd5: xpb[70] = 1024'd122523943181913889559825647857370098138713936614678842630060965300631816858688351034218671716263297294733207288429672583964567359663035763696499010779659080619854519332489127586589132099177969101457944224956547047547681517642000516629278111177565255885510236310654795976811622377277268070350868142894815708945;
            6'd6: xpb[70] = 1024'd22962036134171926072991850024029685021758296811878927027941303295781284893116882331047334844858282444236699338658113666178416990754422581880638687919259855810134748629415735766276719327496357200439335461560616610692856970949503846990155163729848857795792380158668697142067418778804088667302351944848184366403;
            6'd7: xpb[70] = 1024'd47466824770554703984956979595503704649501084134814695553953496355907648264854552537891069188110941903183340796344048182971330462687029734619938490075191671934105652495913561283594545747331951020730924306551926020202393274477903950316010785965361908972894427420799656337429743254259542281372525573427147508192;
            6'd8: xpb[70] = 1024'd71971613406937481896922109166977724277243871457750464079965689416034011636592222744734803531363601362129982254029982699764243934619636887359238292231123488058076556362411386800912372167167544841022513151543235429711929578006304053641866408200874960149996474682930615532792067729714995895442699202006110649981;
            6'd9: xpb[70] = 1024'd96476402043320259808887238738451743904986658780686232605977882476160375008329892951578537874616260821076623711715917216557157406552244040098538094387055304182047460228909212318230198587003138661314101996534544839221465881534704156967722030436388011327098521945061574728154392205170449509512872830585073791770;
            6'd10: xpb[70] = 1024'd120981190679703037720852368309925763532729446103622001131990075536286738380067563158422272217868920280023265169401851733350070878484851192837837896542987120306018364095407037835548025006838732481605690841525854248731002185063104260293577652671901062504200569207192533923516716680625903123583046459164036933559;
            6'd11: xpb[70] = 1024'd21419283631961074234018570476585350415773806300822085529870413531436206414496094455250935346463905429526757219630292815563920509576238011021977573682587895496298593392333646015235612235157120580587082078129923811876177638370607590654454705224184664414482713055206435088772513082152723720534530261117405591017;
            6'd12: xpb[70] = 1024'd45924072268343852145983700048059370043516593623757854055882606591562569786233764662094669689716564888473398677316227332356833981508845163761277375838519711620269497258831471532553438654992714400878670923121233221385713941899007693980310327459697715591584760317337394284134837557608177334604703889696368732806;
            6'd13: xpb[70] = 1024'd70428860904726630057948829619533389671259380946693622581894799651688933157971434868938404032969224347420040135002161849149747453441452316500577177994451527744240401125329297049871265074828308221170259768112542630895250245427407797306165949695210766768686807579468353479497162033063630948674877518275331874595;
            6'd14: xpb[70] = 1024'd94933649541109407969913959191007409299002168269629391107906992711815296529709105075782138376221883806366681592688096365942660925374059469239876980150383343868211304991827122567189091494663902041461848613103852040404786548955807900632021571930723817945788854841599312674859486508519084562745051146854295016384;
            6'd15: xpb[70] = 1024'd119438438177492185881879088762481428926744955592565159633919185771941659901446775282625872719474543265313323050374030882735574397306666621979176782306315159992182208858324948084506917914499495861753437458095161449914322852484208003957877194166236869122890902103730271870221810983974538176815224775433258158173;
            6'd16: xpb[70] = 1024'd19876531129750222395045290929141015809789315789765244031799523767091127935875306579454535848069528414816815100602471964949424028398053440163316459445915935182462438155251556264194505142817883960734828694699231013059498305791711334318754246718520471033173045951744173035477607385501358773766708577386626815631;
            6'd17: xpb[70] = 1024'd44381319766133000307010420500615035437532103112701012557811716827217491307612976786298270191322187873763456558288406481742337500330660592902616261601847751306433342021749381781512331562653477781026417539690540422569034609320111437644609868954033522210275093213875132230839931860956812387836882205965589957420;
            6'd18: xpb[70] = 1024'd68886108402515778218975550072089055065274890435636781083823909887343854679350646993142004534574847332710098015974340998535250972263267745641916063757779567430404245888247207298830157982489071601318006384681849832078570912848511540970465491189546573387377140476006091426202256336412266001907055834544553099209;
            6'd19: xpb[70] = 1024'd93390897038898556130940679643563074693017677758572549609836102947470218051088317199985738877827506791656739473660275515328164444195874898381215865913711383554375149754745032816147984402324665421609595229673159241588107216376911644296321113425059624564479187738137050621564580811867719615977229463123516240998;
            6'd20: xpb[70] = 1024'd117895685675281334042905809215037094320760465081508318135848296007596581422825987406829473221080166250603380931346210032121077916128482051120515668069643199678346053621242858333465810822160259241901184074664468651097643519905311747622176735660572675741581235000268009816926905287323173230047403091702479382787;
            6'd21: xpb[70] = 1024'd18333778627539370556072011381696681203804825278708402533728634002746049457254518703658136349675151400106872981574651114334927547219868869304655345209243974868626282918169466513153398050478647340882575311268538214242818973212815077983053788212856277651863378848281910982182701688849993826998886893655848040245;
            6'd22: xpb[70] = 1024'd42838567263922148468037140953170700831547612601644171059740827062872412828992188910501870692927810859053514439260585631127841019152476022043955147365175790992597186784667292030471224470314241161174164156259847623752355276741215181308909410448369328828965426110412870177545026164305447441069060522234811182034;
            6'd23: xpb[70] = 1024'd67343355900304926380002270524644720459290399924579939585753020122998776200729859117345605036180470318000155896946520147920754491085083174783254949521107607116568090651165117547789050890149834981465753001251157033261891580269615284634765032683882380006067473372543829372907350639760901055139234150813774323823;
            6'd24: xpb[70] = 1024'd91848144536687704291967400096118740087033187247515708111765213183125139572467529324189339379433129776946797354632454664713667963017690327522554751677039423240538994517662943065106877309985428801757341846242466442771427883798015387960620654919395431183169520634674788568269675115216354669209407779392737465612;
            6'd25: xpb[70] = 1024'd116352933173070482203932529667592759714775974570451476637777406243251502944205199531033073722685789235893438812318389181506581434950297480261854553832971239364509898384160768582424703729821022622048930691233775852280964187326415491286476277154908482360271567896805747763631999590671808283279581407971700607401;
            6'd26: xpb[70] = 1024'd16791026125328518717098731834252346597820334767651561035657744238400970978633730827861736851280774385396930862546830263720431066041684298445994230972572014554790127681087376762112290958139410721030321927837845415426139640633918821647353329707192084270553711744819648928887795992198628880231065209925069264859;
            6'd27: xpb[70] = 1024'd41295814761711296629063861405726366225563122090587329561669937298527334350371401034705471194533433844343572320232764780513344537974291451185294033128503830678761031547585202279430117377975004541321910772829154824935675944162318924973208951942705135447655759006950608124250120467654082494301238838504032406648;
            6'd28: xpb[70] = 1024'd65800603398094074541028990977200385853305909413523098087682130358653697722109071241549205537786093303290213777918699297306258009906898603924593835284435646802731935414083027796747943797810598361613499617820464234445212247690719028299064574178218186624757806269081567319612444943109536108371412467082995548437;
            6'd29: xpb[70] = 1024'd90305392034476852452994120548674405481048696736458866613694323418780061093846741448392939881038752762236855235604633814099171481839505756663893637440367462926702839280580853314065770217646192181905088462811773643954748551219119131624920196413731237801859853531212526514974769418564989722441586095661958690226;
            6'd30: xpb[70] = 1024'd114810180670859630364959250120148425108791484059394635139706516478906424465584411655236674224291412221183496693290568330892084953772112909403193439596299279050673743147078678831383596637481786002196677307803083053464284854747519234950775818649244288978961900793343485710337093894020443336511759724240921832015;
            6'd31: xpb[70] = 1024'd15248273623117666878125452286808011991835844256594719537586854474055892500012942952065337352886397370686988743519009413105934584863499727587333116735900054240953972444005287011071183865800174101178068544407152616609460308055022565311652871201527890889244044641357386875592890295547263933463243526194290489473;
            6'd32: xpb[70] = 1024'd39753062259500444790090581858282031619578631579530488063599047534182255871750613158909071696139056829633630201204943929898848056796106880326632918891831870364924876310503112528389010285635767921469657389398462026118996611583422668637508493437040942066346091903488346070955214771002717547533417154773253631262;
            6'd33: xpb[70] = 1024'd64257850895883222702055711429756051247321418902466256589611240594308619243488283365752806039391716288580271658890878446691761528728714033065932721047763686488895780177000938045706836705471361741761246234389771435628532915111822771963364115672553993243448139165619305266317539246458171161603590783352216773051;
            6'd34: xpb[70] = 1024'd88762639532266000614020841001230070875064206225402025115623433654434982615225953572596540382644375747526913116576812963484675000661321185805232523203695502612866684043498763563024663125306955562052835079381080845138069218640222875289219737908067044420550186427750264461679863721913624775673764411931179914840;
            6'd35: xpb[70] = 1024'd113267428168648778525985970572704090502806993548337793641635626714561345986963623779440274725897035206473554574262747480277588472593928338544532325359627318736837587909996589080342489545142549382344423924372390254647605522168622978615075360143580095597652233689881223657042188197369078389743938040510143056629;
            6'd36: xpb[70] = 1024'd13705521120906815039152172739363677385851353745537878039515964709710814021392155076268937854492020355977046624491188562491438103685315156728672002499228093927117817206923197260030076773460937481325815160976459817792780975476126308975952412695863697507934377537895124822297984598895898986695421842463511714087;
            6'd37: xpb[70] = 1024'd38210309757289592951117302310837697013594141068473646565528157769837177393129825283112672197744679814923688082177123079284351575617922309467971804655159910051088721073421022777347903193296531301617404005967769227302317279004526412301808034931376748685036424800026084017660309074351352600765595471042474855876;
            6'd38: xpb[70] = 1024'd62715098393672370863082431882311716641336928391409415091540350829963540764867495489956406540997339273870329539863057596077265047550529462207271606811091726175059624939918848294665729613132125121908992850959078636811853582532926515627663657166889799862138472062157043213022633549806806214835769099621437997665;
            6'd39: xpb[70] = 1024'd87219887030055148775047561453785736269079715714345183617552543890089904136605165696800140884249998732816970997548992112870178519483136614946571408967023542299030528806416673811983556032967718942200581695950388046321389886061326618953519279402402851039240519324288002408384958025262259828905942728200401139454;
            6'd40: xpb[70] = 1024'd111724675666437926687012691025259755896822503037280952143564736950216267508342835903643875227502658191763612455234926629663091991415743767685871211122955358423001432672914499329301382452803312762492170540941697455830926189589726722279374901637915902216342566586418961603747282500717713442976116356779364281243;
            6'd41: xpb[70] = 1024'd12162768618695963200178893191919342779866863234481036541445074945365735542771367200472538356097643341267104505463367711876941622507130585870010888262556133613281661969841107508988969681121700861473561777545767018976101642897230052640251954190199504126624710434432862769003078902244534039927600158732732938701;
            6'd42: xpb[70] = 1024'd36667557255078741112144022763393362407609650557416805067457268005492098914509037407316272699350302800213745963149302228669855094439737738609310690418487949737252565836338933026306796100957294681765150622537076428485637946425630155966107576425712555303726757696563821964365403377699987653997773787311696080490;
            6'd43: xpb[70] = 1024'd61172345891461519024109152334867382035352437880352573593469461065618462286246707614160007042602962259160387420835236745462768566372344891348610492574419765861223469702836758543624622520792888502056739467528385837995174249954030259291963198661225606480828804958694781159727727853155441268067947415890659222279;
            6'd44: xpb[70] = 1024'd85677134527844296936074281906341401663095225203288342119481654125744825657984377821003741385855621718107028878521171262255682038304952044087910294730351581985194373569334584060942448940628482322348328312519695247504710553482430362617818820896738657657930852220825740355090052328610894882138121044469622364068;
            6'd45: xpb[70] = 1024'd110181923164227074848039411477815421290838012526224110645493847185871189029722048027847475729108281177053670336207105779048595510237559196827210096886283398109165277435832409578260275360464076142639917157511004657014246857010830465943674443132251708835032899482956699550452376804066348496208294673048585505857;
            6'd46: xpb[70] = 1024'd10620016116485111361205613644475008173882372723424195043374185181020657064150579324676138857703266326557162386435546861262445141328946015011349774025884173299445506732759017757947862588782464241621308394115074220159422310318333796304551495684535310745315043330970600715708173205593169093159778475001954163315;
            6'd47: xpb[70] = 1024'd35124804752867889273170743215949027801625160046359963569386378241147020435888249531519873200955925785503803844121481378055358613261553167750649576181815989423416410599256843275265689008618058061912897239106383629668958613846733899630407117920048361922417090593101559911070497681048622707229952103580917305104;
            6'd48: xpb[70] = 1024'd59629593389250667185135872787423047429367947369295732095398571301273383807625919738363607544208585244450445301807415894848272085194160320489949378337747805547387314465754668792583515428453651882204486084097693039178494917375134002956262740155561413099519137855232519106432822156504076321300125732159880446893;
            6'd49: xpb[70] = 1024'd84134382025633445097101002358897067057110734692231500621410764361399747179363589945207341887461244703397086759493350411641185557126767473229249180493679621671358218332252494309901341848289245702496074929089002448688031220903534106282118362391074464276621185117363478301795146631959529935370299360738843588682;
            6'd50: xpb[70] = 1024'd108639170662016223009066131930371086684853522015167269147422957421526110551101260152051076230713904162343728217179284928434099029059374625968548982649611437795329122198750319827219168268124839522787663774080311858197567524431934209607973984626587515453723232379494437497157471107414983549440472989317806730471;
            6'd51: xpb[70] = 1024'd9077263614274259522232334097030673567897882212367353545303295416675578585529791448879739359308889311847220267407726010647948660150761444152688659789212212985609351495676928006906755496443227621769055010684381421342742977739437539968851037178871117364005376227508338662413267508941804146391956791271175387929;
            6'd52: xpb[70] = 1024'd33582052250657037434197463668504693195640669535303122071315488476801941957267461655723473702561548770793861725093660527440862132083368596891988461945144029109580255362174753524224581916278821442060643855675690830852279281267837643294706659414384168541107423489639297857775591984397257760462130419850138529718;
            6'd53: xpb[70] = 1024'd58086840887039815346162593239978712823383456858238890597327681536928305329005131862567208045814208229740503182779595044233775604015975749631288264101075845233551159228672579041542408336114415262352232700667000240361815584796237746620562281649897219718209470751770257053137916459852711374532304048429101671507;
            6'd54: xpb[70] = 1024'd82591629523422593258127722811452732451126244181174659123339874597054668700742802069410942389066867688687144640465529561026689075948582902370588066257007661357522063095170404558860234755950009082643821545658309649871351888324637849946417903885410270895311518013901216248500240935308164988602477677008064813296;
            6'd55: xpb[70] = 1024'd107096418159805371170092852382926752078869031504110427649352067657181032072480472276254676732319527147633786098151464077819602547881190055109887868412939477481492966961668230076178061175785602902935410390649619059380888191853037953272273526120923322072413565276032175443862565410763618602672651305587027955085;
            6'd56: xpb[70] = 1024'd7534511112063407683259054549586338961913391701310512047232405652330500106909003573083339860914512297137278148379905160033452178972576873294027545552540252671773196258594838255865648404103991001916801627253688622526063645160541283633150578673206923982695709124046076609118361812290439199624135107540396612543;
            6'd57: xpb[70] = 1024'd32039299748446185595224184121060358589656179024246280573244598712456863478646673779927074204167171756083919606065839676826365650905184026033327347708472068795744100125092663773183474823939584822208390472244998032035599948688941386959006200908719975159797756386177035804480686287745892813694308736119359754332;
            6'd58: xpb[70] = 1024'd56544088384828963507189313692534378217398966347182049099256791772583226850384343986770808547419831215030561063751774193619279122837791178772627149864403884919715003991590489290501301243775178642499979317236307441545136252217341490284861823144233026336899803648307994999843010763201346427764482364698322896121;
            6'd59: xpb[70] = 1024'd81048877021211741419154443264008397845141753670117817625268984832709590222122014193614542890672490673977202521437708710412192594770398331511926952020335701043685907858088314807819127663610772462791568162227616851054672555745741593610717445379746077514001850910438954195205335238656800041834655993277286037910;
            6'd60: xpb[70] = 1024'd105553665657594519331119572835482417472884540993053586151281177892835953593859684400458277233925150132923843979123643227205106066703005484251226754176267517167656811724586140325136954083446366283083157007218926260564208859274141696936573067615259128691103898172569913390567659714112253655904829621856249179699;
            6'd61: xpb[70] = 1024'd5991758609852555844285775002142004355928901190253670549161515887985421628288215697286940362520135282427336029352084309418955697794392302435366431315868292357937041021512748504824541311764754382064548243822995823709384312581645027297450120167542730601386042020583814555823456115639074252856313423809617837157;
            6'd62: xpb[70] = 1024'd30496547246235333756250904573616023983671688513189439075173708948111785000025885904130674705772794741373977487038018826211869169726999455174666233471800108481907944888010574022142367731600348202356137088814305233218920616110045130623305742403055781778488089282714773751185780591094527866926487052388580978946;
            6'd63: xpb[70] = 1024'd55001335882618111668216034145090043611414475836125207601185902008238148371763556110974409049025454200320618944723953343004782641659606607913966035627731924605878848754508399539460194151435942022647725933805614642728456919638445233949161364638568832955590136544845732946548105066549981480996660680967544120735;
        endcase
    end

    always_comb begin
        case(flag[23][16:12])
            5'd0: xpb[71] = 1024'd0;
            5'd1: xpb[71] = 1024'd79506124519000889580181163716564063239157263159060976127198095068364511743501226317818143392278113659267260402409887859797696113592213760653265837783663740729849752621006225056778020571271535842939314778796924052237993223166845337275016986874081884132692183806976692141910429542005435095066834309546507262524;
            5'd2: xpb[71] = 1024'd34945553353877037761563400028313693733616099192386268126264335071752128149693313725621215569898553009091371397362282285016328386343207186751371550550996440526008830672441232775925801951025865964568431949206608258111625596112793901585055404064934318998564464199836326253714331010082237173014978792467420040717;
            5'd3: xpb[71] = 1024'd114451677872877927341744563744877756972773362351447244253462430140116639893194540043439358962176666668358631799772170144814024499935420947404637388334660181255858583293447457832703822522297401807507746728003532310349618819279639238860072390939016203131256648006813018395624760552087672268081813102013927303241;
            5'd4: xpb[71] = 1024'd69891106707754075523126800056627387467232198384772536252528670143504256299386627451242431139797106018182742794724564570032656772686414373502743101101992881052017661344882465551851603902051731929136863898413216516223251192225587803170110808129868637997128928399672652507428662020164474346029957584934840081434;
            5'd5: xpb[71] = 1024'd25330535542630223704509036368377017961691034418097828251594910146891872705578714859045503317417545368006853789676958995251289045437407799600848813869325580848176739396317473270999385281806062050765981068822900722096883565171536367480149225320721072863001208792532286619232563488241276423978102067855752859627;
            5'd6: xpb[71] = 1024'd104836660061631113284690200084941081200848297577158804378793005215256384449079941176863646709695659027274114192086846855048985159029621560254114651652989321578026492017323698327777405853077597893705295847619824774334876788338381704755166212194802956995693392599508978761142993030246711519044936377402260122151;
            5'd7: xpb[71] = 1024'd60276088896507261466072436396690711695307133610484096377859245218644000855272028584666718887316098377098225187039241280267617431780614986352220364420322021374185570068758706046925187232831928015334413018029508980208509161284330269065204629385655391861565672992368612872946894498323513596993080860323172900344;
            5'd8: xpb[71] = 1024'd15715517731383409647454672708440342189765969643809388376925485222031617261464115992469791064936537726922336181991635705486249704531608412450326077187654721170344648120193713766072968612586258136963530188439193186082141534230278833375243046576507826727437953385228246984750795966400315674941225343244085678537;
            5'd9: xpb[71] = 1024'd95221642250384299227635836425004405428923232802870364504123580290396129004965342310287934457214651386189596584401523565283945818123822173103591914971318461900194400741199938822850989183857793979902844967236117238320134757397124170650260033450589710860130137192204939126661225508405750770008059652790592941061;
            5'd10: xpb[71] = 1024'd50661071085260447409018072736754035923382068836195656503189820293783745411157429718091006634835090736013707579353917990502578090874815599201697627738651161696353478792634946541998770563612124101531962137645801444193767130343072734960298450641442145726002417585064573238465126976482552847956204135711505719254;
            5'd11: xpb[71] = 1024'd6100499920136595590400309048503666417840904869520948502256060297171361817349517125894078812455530085837818574306312415721210363625809025299803340505983861492512556844069954261146551943366454223161079308055485650067399503289021299270336867832294580591874697977924207350269028444559354925904348618632418497447;
            5'd12: xpb[71] = 1024'd85606624439137485170581472765067729656998168028581924629454155365535873560850743443712222204733643745105078976716200275518906477218022785953069178289647602222362309465076179317924572514637990066100394086852409702305392726455866636545353854706376464724566881784900899492179457986564790020971182928178925759971;
            5'd13: xpb[71] = 1024'd41046053274013633351963709076817360151457004061907216628520395368923489967042830851515294382354083094929189971668594700737538749969016212051174891056980302018521387516511187037072353894392320187729511257262093908179025099401815200855392271897228899590439162177760533603983359454641592098919327411099838538164;
            5'd14: xpb[71] = 1024'd120552177793014522932144872793381423390614267220968192755718490437288001710544057169333437774632196754196450374078482560535234863561229972704440728840644042748371140137517412093850374465663856030668826036059017960417018322568660538130409258771310783723131345984737225745893788996647027193986161720646345800688;
            5'd15: xpb[71] = 1024'd75991606627890671113527109105131053885073103254293484754784730440675618116736144577136509952252636104020561369030876985753867136312223398802546441607976742544530218188952419812998155845418186152297943206468702166290650695514609102440447675962163218589003626377596859857697690464723829271934306203567258578881;
            5'd16: xpb[71] = 1024'd31431035462766819294909345416880684379531939287618776753850970444063234522928231984939582129873075453844672363983271410972499409063216824900652154375309442340689296240387427532145937225172516273927060376878386372164283068460557666750486093153015653454875906770456493969501591932800631349882450686488171357074;
            5'd17: xpb[71] = 1024'd110937159981767708875090509133444747618689202446679752881049065512427746266429458302757725522151189113111932766393159270770195522655430585553917992158973183070539048861393652588923957796444052116866375155675310424402276291627403004025503080027097537587568090577433186111412021474806066444949284996034678619598;
            5'd18: xpb[71] = 1024'd66376588816643857056472745445194378113148038480005044880115305515815362672621545710560797699771628462936043761345553695988827795406424011652023704926305882866698126912828660308071739176198382238495492326084994630275908664573351568335541497217949972453440370970292820223215922942882868522897429478955591397791;
            5'd19: xpb[71] = 1024'd21816017651520005237854981756944008607606874513330336879181545519202979078813633118363869877392067812760154756297948121207460068157417437750129417693638582662857204964263668027219520555952712360124609496494678836149541037519300132645579914408802407319312651363152454335019824410959670600845573961876504175984;
            5'd20: xpb[71] = 1024'd101322142170520894818036145473508071846764137672391313006379640587567490822314859436182013269670181472027415158707835981005156181749631198403395255477302323392706957585269893083997541127224248203063924275291602888387534260686145469920596901282884291452004835170129146476930253952965105695912408271423011438508;
            5'd21: xpb[71] = 1024'd56761571005397042999418381785257702341222973705716605005445880590955107228506946843985085447290620821851526153660230406223788454500624624501500968244635023188866035636704900803145322506978578324693041445701287094261166633632094034230635318473736726317877115562988780588734155421041907773860552754343924216701;
            5'd22: xpb[71] = 1024'd12200999840273191180800618097007332835681809739041897004512120594342723634699034251788157624911060171675637148612624831442420727251618050599606681011967722985025113688139908522293103886732908446322158616110971300134799006578042598540673735664589161183749395955848414700538056889118709851808697237264836994894;
            5'd23: xpb[71] = 1024'd91707124359274080760981781813571396074839072898102873131710215662707235378200260569606301017189173830942897551022512691240116840843831811252872518795631463714874866309146133579071124458004444289261473394907895352372792229744887935815690722538671045316441579762825106842448486431124144946875531546811344257418;
            5'd24: xpb[71] = 1024'd47146553194150228942364018125321026569297908931428165130776455666094851784392347977409373194809613180767008545974907116458749113594825237350978231562964163511033944360581141298218905837758774410890590565317579558246424602690836500125729139729523480182313860155684740954252387899200947024823676029732257035611;
            5'd25: xpb[71] = 1024'd2585982029026377123746254437070657063756744964753457129842695669482468190584435385212445372430052530591119540927301541677381386345818663449083944330296863307193022412016149017366687217513104532519707735727263764120056975636785064435767556920375915048186140548544375066056289367277749102771820512653169813804;
            5'd26: xpb[71] = 1024'd82092106548027266703927418153634720302914008123814433257040790737846979934085661703030588764708166189858379943337189401475077499938032424102349782113960604037042775033022374074144707788784640375459022514524187816358050198803630401710784543794457799180878324355521067207966718909283184197838654822199677076328;
            5'd27: xpb[71] = 1024'd37531535382903414885309654465384350797372844157139725256107030741234596340277749110833660942328605539682490938289583826693709772689025850200455494881293303833201853084457381793292489168538970497088139684933872022231682571749578966020822960985310234046750604748380701319770620377359986275786799305120589854521;
            5'd28: xpb[71] = 1024'd117037659901904304465490818181948414036530107316200701383305125809599108083778975428651804334606719198949751340699471686491405886281239610853721332664957044563051605705463606850070509739810506340027454463730796074469675794916424303295839947859392118179442788555357393461681049919365421370853633614667097117045;
            5'd29: xpb[71] = 1024'd72477088736780452646873054493698044530988943349525993382371365812986724489971062836454876512227158548773862335651866111710038159032233036951827045432289744359210683756898614569218291119564836461656571634140480280343308167862372867605878365050244553045315068948217027573484951387442223448801778097588009895238;
            5'd30: xpb[71] = 1024'd27916517571656600828255290805447675025447779382851285381437605816374340896163150244257948689847597898597973330604260536928670431783226463049932758199622444155369761808333622288366072499319166583285688804550164486216940540808321431915916782241096987911187349341076661685288852855519025526749922580508922673431;
            5'd31: xpb[71] = 1024'd107422642090657490408436454522011738264605042541912261508635700884738852639664376562076092082125711557865233733014148396726366545375440223703198595983286184885219514429339847345144093070590702426225003583347088538454933763975166769190933769115178872043879533148053353827199282397524460621816756890055429935955;
        endcase
    end

    always_comb begin
        case(flag[24][5:0])
            6'd0: xpb[72] = 1024'd0;
            6'd1: xpb[72] = 1024'd31431035462766819294909345416880684379531939287618776753850970444063234522928231984939582129873075453844672363983271410972499409063216824900652154375309442340689296240387427532145937225172516273927060376878386372164283068460557666750486093153015653454875906770456493969501591932800631349882450686488171357074;
            6'd2: xpb[72] = 1024'd62862070925533638589818690833761368759063878575237553507701940888126469045856463969879164259746150907689344727966542821944998818126433649801304308750618884681378592480774855064291874450345032547854120753756772744328566136921115333500972186306031306909751813540912987939003183865601262699764901372976342714148;
            6'd3: xpb[72] = 1024'd94293106388300457884728036250642053138595817862856330261552911332189703568784695954818746389619226361534017091949814232917498227189650474701956463125928327022067888721162282596437811675517548821781181130635159116492849205381673000251458279459046960364627720311369481908504775798401894049647352059464514071222;
            6'd4: xpb[72] = 1024'd1657446166942535780838454262708304773429330024739422887272026711276042754403789029743257304834627505935540048475592209310933795411646965047448492484906728429066510391978492790953509709172859374398043899126305642292771423621333894036965802928833164552683723667708917847899839657273892382411112919327090943965;
            6'd5: xpb[72] = 1024'd33088481629709355075747799679588989152961269312358199641122997155339277277332021014682839434707702959780212412458863620283433204474863789948100646860216170769755806632365920323099446934345375648325104276004692014457054492081891560787451896081848818007559630438165411817401431590074523732293563605815262301039;
            6'd6: xpb[72] = 1024'd64519517092476174370657145096469673532493208599976976394973967599402511800260252999622421564580778413624884776442135031255932613538080614848752801235525613110445102872753347855245384159517891922252164652883078386621337560542449227537937989234864471462435537208621905786903023522875155082176014292303433658113;
            6'd7: xpb[72] = 1024'd95950552555242993665566490513350357912025147887595753148824938043465746323188484984562003694453853867469557140425406442228432022601297439749404955610835055451134399113140775387391321384690408196179225029761464758785620629003006894288424082387880124917311443979078399756404615455675786432058464978791605015187;
            6'd8: xpb[72] = 1024'd3314892333885071561676908525416609546858660049478845774544053422552085508807578059486514609669255011871080096951184418621867590823293930094896984969813456858133020783956985581907019418345718748796087798252611284585542847242667788073931605857666329105367447335417835695799679314547784764822225838654181887930;
            6'd9: xpb[72] = 1024'd34745927796651890856586253942297293926390599337097622528395023866615320031735810044426096739542330465715752460934455829594366999886510754995549139345122899198822317024344413114052956643518235022723148175130997656749825915703225454824417699010681982560243354105874329665301271247348416114704676525142353245004;
            6'd10: xpb[72] = 1024'd66176963259418710151495599359177978305922538624716399282245994310678554554664042029365678869415405919560424824917727240566866408949727579896201293720432341539511613264731840646198893868690751296650208552009384028914108984163783121574903792163697636015119260876330823634802863180149047464587127211630524602078;
            6'd11: xpb[72] = 1024'd97607998722185529446404944776058662685454477912335176036096964754741789077592274014305260999288481373405097188900998651539365818012944404796853448095741783880200909505119268178344831093863267570577268928887770401078392052624340788325389885316713289469995167646787317604304455112949678814469577898118695959152;
            6'd12: xpb[72] = 1024'd4972338500827607342515362788124914320287990074218268661816080133828128263211367089229771914503882517806620145426776627932801386234940895142345477454720185287199531175935478372860529127518578123194131697378916926878314270864001682110897408786499493658051171003126753543699518971821677147233338757981272831895;
            6'd13: xpb[72] = 1024'd36403373963594426637424708205005598699819929361837045415667050577891362786139599074169354044376957971651292509410048038905300795298157720042997631830029627627888827416322905905006466352691094397121192074257303299042597339324559348861383501939515147112927077773583247513201110904622308497115789444469444188969;
            6'd14: xpb[72] = 1024'd67834409426361245932334053621886283079351868649455822169518021021954597309067831059108936174250033425495964873393319449877800204361374544943649786205339069968578123656710333437152403577863610671048252451135689671206880407785117015611869595092530800567802984544039741482702702837422939846998240130957615546043;
            6'd15: xpb[72] = 1024'd99265444889128065227243399038766967458883807937074598923368991466017831831996063044048518304123108879340637237376590860850299613424591369844301940580648512309267419897097760969298340803036126944975312828014076043371163476245674682362355688245546454022678891314496235452204294770223571196880690817445786903117;
            6'd16: xpb[72] = 1024'd6629784667770143123353817050833219093717320098957691549088106845104171017615156118973029219338510023742160193902368837243735181646587860189793969939626913716266041567913971163814038836691437497592175596505222569171085694485335576147863211715332658210734894670835671391599358629095569529644451677308363775860;
            6'd17: xpb[72] = 1024'd38060820130536962418263162467713903473249259386576468302939077289167405540543388103912611349211585477586832557885640248216234590709804685090446124314936356056955337808301398695959976061863953771519235973383608941335368762945893242898349304868348311665610801441292165361100950561896200879526902363796535132934;
            6'd18: xpb[72] = 1024'd69491855593303781713172507884594587852781198674195245056790047733230640063471620088852193479084660931431504921868911659188733999773021509991098278690245798397644634048688826228105913287036470045446296350261995313499651831406450909648835398021363965120486708211748659330602542494696832229409353050284706490008;
            6'd19: xpb[72] = 1024'd100922891056070601008081853301475272232313137961814021810641018177293874586399852073791775608957736385276177285852183070161233408836238334891750433065555240738333930289076253760251850512208986319373356727140381685663934899867008576399321491174379618575362614982205153300104134427497463579291803736772877847082;
            6'd20: xpb[72] = 1024'd8287230834712678904192271313541523867146650123697114436360133556380213772018945148716286524173137529677700242377961046554668977058234825237242462424533642145332551959892463954767548545864296871990219495631528211463857118106669470184829014644165822763418618338544589239499198286369461912055564596635454719825;
            6'd21: xpb[72] = 1024'd39718266297479498199101616730422208246678589411315891190211104000443448294947177133655868654046212983522372606361232457527168386121451650137894616799843084486021848200279891486913485771036813145917279872509914583628140186567227136935315107797181476218294525109001083209000790219170093261938015283123626076899;
            6'd22: xpb[72] = 1024'd71149301760246317494010962147302892626210528698934667944062074444506682817875409118595450783919288437367044970344503868499667795184668475038546771175152526826711144440667319019059422996209329419844340249388300955792423255027784803685801200950197129673170431879457577178502382151970724611820465969611797433973;
            6'd23: xpb[72] = 1024'd102580337223013136788920307564183577005742467986553444697913044888569917340803641103535032913792363891211717334327775279472167204247885299939198925550461969167400440681054746551205360221381845693771400626266687327956706323488342470436287294103212783128046338649914071148003974084771355961702916656099968791047;
            6'd24: xpb[72] = 1024'd9944677001655214685030725576249828640575980148436537323632160267656256526422734178459543829007765035613240290853553255865602772469881790284690954909440370574399062351870956745721058255037156246388263394757833853756628541728003364221794817572998987316102342006253507087399037943643354294466677515962545663790;
            6'd25: xpb[72] = 1024'd41375712464422033979940070993130513020107919436055314077483130711719491049350966163399125958880840489457912654836824666838102181533098615185343109284749812915088358592258384277866995480209672520315323771636220225920911610188561030972280910726014640770978248776710001056900629876443985644349128202450717020864;
            6'd26: xpb[72] = 1024'd72806747927188853274849416410011197399639858723674090831334101155782725572279198148338708088753915943302585018820096077810601590596315440085995263660059255255777654832645811810012932705382188794242384148514606598085194678649118697722767003879030294225854155547166495026402221809244616994231578888938888377938;
            6'd27: xpb[72] = 1024'd104237783389955672569758761826891881779171798011292867585185071599845960095207430133278290218626991397147257382803367488783100999659532264986647418035368697596466951073033239342158869930554705068169444525392992970249477747109676364473253097032045947680730062317622988995903813742045248344114029575427059735012;
            6'd28: xpb[72] = 1024'd11602123168597750465869179838958133414005310173175960210904186978932299280826523208202801133842392541548780339329145465176536567881528755332139447394347099003465572743849449536674567964210015620786307293884139496049399965349337258258760620501832151868786065673962424935298877600917246676877790435289636607755;
            6'd29: xpb[72] = 1024'd43033158631364569760778525255838817793537249460794736964755157422995533803754755193142383263715467995393452703312416876149035976944745580232791601769656541344154868984236877068820505189382531894713367670762525868213683033809894925009246713654847805323661972444418918904800469533717878026760241121777807964829;
            6'd30: xpb[72] = 1024'd74464194094131389055687870672719502173069188748413513718606127867058768326682987178081965393588543449238125067295688287121535386007962405133443756144965983684844165224624304600966442414555048168640428047640912240377966102270452591759732806807863458778537879214875412874302061466518509376642691808265979321903;
            6'd31: xpb[72] = 1024'd105895229556898208350597216089600186552601128036032290472457098311122002849611219163021547523461618903082797431278959698094034795071179230034095910520275426025533461465011732133112379639727564442567488424519298612542249170731010258510218899960879112233413785985331906843803653399319140726525142494754150678977;
            6'd32: xpb[72] = 1024'd13259569335540286246707634101666438187434640197915383098176213690208342035230312237946058438677020047484320387804737674487470363293175720379587939879253827432532083135827942327628077673382874995184351193010445138342171388970671152295726423430665316421469789341671342783198717258191139059288903354616727551720;
            6'd33: xpb[72] = 1024'd44690604798307105541616979518547122566966579485534159852027184134271576558158544222885640568550095501328992751788009085459969772356392545280240094254563269773221379376215369859774014898555391269111411569888831510506454457431228819046212516583680969876345696112127836752700309190991770409171354041104898908794;
            6'd34: xpb[72] = 1024'd76121640261073924836526324935427806946498518773152936605878154578334811081086776207825222698423170955173665115771280496432469181419609370180892248629872712113910675616602797391919952123727907543038471946767217882670737525891786485796698609736696623331221602882584330722201901123792401759053804727593070265868;
            6'd35: xpb[72] = 1024'd107552675723840744131435670352308491326030458060771713359729125022398045604015008192764804828296246409018337479754551907404968590482826195081544403005182154454599971856990224924065889348900423816965532323645604254835020594352344152547184702889712276786097509653040824691703493056593033108936255414081241622942;
            6'd36: xpb[72] = 1024'd14917015502482822027546088364374742960863970222654805985448240401484384789634101267689315743511647553419860436280329883798404158704822685427036432364160555861598593527806435118581587382555734369582395092136750780634942812592005046332692226359498480974153513009380260631098556915465031441700016273943818495685;
            6'd37: xpb[72] = 1024'd46348050965249641322455433781255427340395909510273582739299210845547619312562333252628897873384723007264532800263601294770903567768039510327688586739469998202287889768193862650727524607728250643509455469015137152799225881052562713083178319512514134429029419779836754600600148848265662791582466960431989852759;
            6'd38: xpb[72] = 1024'd77779086428016460617364779198136111719927848797892359493150181289610853835490565237568480003257798461109205164246872705743402976831256335228340741114779440542977186008581290182873461832900766917436515845893523524963508949513120379833664412665529787883905326550293248570101740781066294141464917646920161209833;
            6'd39: xpb[72] = 1024'd109210121890783279912274124615016796099459788085511136247001151733674088358418797222508062133130873914953877528230144116715902385894473160128992895490088882883666482248968717715019399058073283191363576222771909897127792017973678046584150505818545441338781233320749742539603332713866925491347368333408332566907;
            6'd40: xpb[72] = 1024'd16574461669425357808384542627083047734293300247394228872720267112760427544037890297432573048346275059355400484755922093109337954116469650474484924849067284290665103919784927909535097091728593743980438991263056422927714236213338940369658029288331645526837236677089178478998396572738923824111129193270909439650;
            6'd41: xpb[72] = 1024'd48005497132192177103293888043963732113825239535013005626571237556823662066966122282372155178219350513200072848739193504081837363179686475375137079224376726631354400160172355441681034316901110017907499368141442795091997304673896607120144122441347298981713143447545672448499988505539555173993579879759080796724;
            6'd42: xpb[72] = 1024'd79436532594958996398203233460844416493357178822631782380422208000886896589894354267311737308092425967044745212722464915054336772242903300275789233599686168972043696400559782973826971542073626291834559745019829167256280373134454273870630215594362952436589050218002166418001580438340186523876030566247252153798;
            6'd43: xpb[72] = 1024'd110867568057725815693112578877725100872889118110250559134273178444950131112822586252251319437965501420889417576705736326026836181306120125176441387974995611312732992640947210505972908767246142565761620121898215539420563441595011940621116308747378605891464956988458660387503172371140817873758481252735423510872;
            6'd44: xpb[72] = 1024'd18231907836367893589222996889791352507722630272133651759992293824036470298441679327175830353180902565290940533231514302420271749528116615521933417333974012719731614311763420700488606800901453118378482890389362065220485659834672834406623832217164810079520960344798096326898236230012816206522242112598000383615;
            6'd45: xpb[72] = 1024'd49662943299134712884132342306672036887254569559752428513843264268099704821369911312115412483053978019135612897214785713392771158591333440422585571709283455060420910552150848232634544026073969392305543267267748437384768728295230501157109925370180463534396867115254590296399828162813447556404692799086171740689;
            6'd46: xpb[72] = 1024'd81093978761901532179041687723552721266786508847371205267694234712162939344298143297054994612927053472980285261198057124365270567654550265323237726084592897401110206792538275764780481251246485666232603644146134809549051796755788167907596018523196116989272773885711084265901420095614078906287143485574343097763;
            6'd47: xpb[72] = 1024'd112525014224668351473951033140433405646318448134989982021545205156226173867226375281994576742800128926824957625181328535337769976717767090223889880459902339741799503032925703296926418476419001940159664021024521181713334865216345834658082111676211770444148680656167578235403012028414710256169594172062514454837;
            6'd48: xpb[72] = 1024'd19889354003310429370061451152499657281151960296873074647264320535312513052845468356919087658015530071226480581707106511731205544939763580569381909818880741148798124703741913491442116510074312492776526789515667707513257083456006728443589635145997974632204684012507014174798075887286708588933355031925091327580;
            6'd49: xpb[72] = 1024'd51320389466077248664970796569380341660683899584491851401115290979375747575773700341858669787888605525071152945690377922703704954002980405470034064194190183489487420944129341023588053735246828766703587166394054079677540151916564395194075728299013628087080590782963508144299667820087339938815805718413262684654;
            6'd50: xpb[72] = 1024'd82751424928844067959880141986261026040215838872110628154966261423438982098701932326798251917761680978915825309673649333676204363066197230370686218569499625830176717184516768555733990960419345040630647543272440451841823220377122061944561821452029281541956497553420002113801259752887971288698256404901434041728;
            6'd51: xpb[72] = 1024'd114182460391610887254789487403141710419747778159729404908817231867502216621630164311737834047634756432760497673656920744648703772129414055271338372944809068170866013424904196087879928185591861314557707920150826824006106288837679728695047914605044934996832404323876496083302851685688602638580707091389605398802;
            6'd52: xpb[72] = 1024'd21546800170252965150899905415207962054581290321612497534536347246588555807249257386662344962850157577162020630182698721042139340351410545616830402303787469577864635095720406282395626219247171867174570688641973349806028507077340622480555438074831139184888407680215932022697915544560600971344467951252182271545;
            6'd53: xpb[72] = 1024'd52977835633019784445809250832088646434113229609231274288387317690651790330177489371601927092723233031006692994165970132014638749414627370517482556679096911918553931336107833814541563444419688141101631065520359721970311575537898289231041531227846792639764314450672425992199507477361232321226918637740353628619;
            6'd54: xpb[72] = 1024'd84408871095786603740718596248969330813645168896850051042238288134715024853105721356541509222596308484851365358149241542987138158477844195418134711054406354259243227576495261346687500669592204415028691442398746094134594643998455955981527624380862446094640221221128919961701099410161863671109369324228524985693;
            6'd55: xpb[72] = 1024'd115839906558553423035627941665850015193177108184468827796089258578778259376033953341481091352469383938696037722132512953959637567541061020318786865429715796599932523816882688878833437894764720688955751819277132466298877712459013622732013717533878099549516127991585413931202691342962495020991820010716696342767;
            6'd56: xpb[72] = 1024'd23204246337195500931738359677916266828010620346351920421808373957864598561653046416405602267684785083097560678658290930353073135763057510664278894788694198006931145487698899073349135928420031241572614587768278992098799930698674516517521241003664303737572131347924849870597755201834493353755580870579273215510;
            6'd57: xpb[72] = 1024'd54635281799962320226647705094796951207542559633970697175659344401927833084581278401345184397557860536942233042641562341325572544826274335564931049164003640347620441728086326605495073153592547515499674964646665364263082999159232183268007334156679957192448038118381343840099347134635124703638031557067444572584;
            6'd58: xpb[72] = 1024'd86066317262729139521557050511677635587074498921589473929510314845991067607509510386284766527430935990786905406624833752298071953889491160465583203539313082688309737968473754137641010378765063789426735341525051736427366067619789850018493427309695610647323944888837837809600939067435756053520482243555615929658;
            6'd59: xpb[72] = 1024'd117497352725495958816466395928558319966606438209208250683361285290054302130437742371224348657304011444631577770608105163270571362952707985366235357914622525028999034208861181669786947603937580063353795718403438108591649136080347516768979520462711264102199851659294331779102531000236387403402932930043787286732;
            6'd60: xpb[72] = 1024'd24861692504138036712576813940624571601439950371091343309080400669140641316056835446148859572519412589033100727133883139664006931174704475711727387273600926435997655879677391864302645637592890615970658486894584634391571354320008410554487043932497468290255855015633767718497594859108385736166693789906364159475;
            6'd61: xpb[72] = 1024'd56292727966904856007486159357505255980971889658710120062931371113203875838985067431088441702392488042877773091117154550636506340237921300612379541648910368776686952120064819396448582862765406889897718863772971006555854422780566077304973137085513121745131761786090261687999186791909017086049144476394535516549;
            6'd62: xpb[72] = 1024'd87723763429671675302395504774385940360503828946328896816782341557267110361913299416028023832265563496722445455100425961609005749301138125513031696024219811117376248360452246928594520087937923163824779240651357378720137491241123744055459230238528775200007668556546755657500778724709648435931595162882706873623;
            6'd63: xpb[72] = 1024'd119154798892438494597304850191266624740035768233947673570633312001330344884841531400967605962138638950567117819083697372581505158364354950413683850399529253458065544600839674460740457313110439437751839617529743750884420559701681410805945323391544428654883575327003249627002370657510279785814045849370878230697;
        endcase
    end

    always_comb begin
        case(flag[24][11:6])
            6'd0: xpb[73] = 1024'd0;
            6'd1: xpb[73] = 1024'd26519138671080572493415268203332876374869280395830766196352427380416684070460624475892116877354040094968640775609475348974940726586351440759175879758507654865064166271655884655256155346765749990368702386020890276684342777941342304591452846861330632842939578683342685566397434516382278118577806709233455103440;
            6'd2: xpb[73] = 1024'd53038277342161144986830536406665752749738560791661532392704854760833368140921248951784233754708080189937281551218950697949881453172702881518351759517015309730128332543311769310512310693531499980737404772041780553368685555882684609182905693722661265685879157366685371132794869032764556237155613418466910206880;
            6'd3: xpb[73] = 1024'd79557416013241717480245804609998629124607841187492298589057282141250052211381873427676350632062120284905922326828426046924822179759054322277527639275522964595192498814967653965768466040297249971106107158062670830053028333824026913774358540583991898528818736050028056699192303549146834355733420127700365310320;
            6'd4: xpb[73] = 1024'd106076554684322289973661072813331505499477121583323064785409709521666736281842497903568467509416160379874563102437901395899762906345405763036703519034030619460256665086623538621024621387062999961474809544083561106737371111765369218365811387445322531371758314733370742265589738065529112474311226836933820413760;
            6'd5: xpb[73] = 1024'd8528997671278121068277413611849949129647974853418146853630281837106525014993983469445513172112526165400054470589883310295639792090536869240719273776207233391630156788708205938650537542311544230533314321717211537057353039485814749992285664623423714947877990002596369801880644507982757575770343719541681032869;
            6'd6: xpb[73] = 1024'd35048136342358693561692681815182825504517255249248913049982709217523209085454607945337630049466566260368695246199358659270580518676888309999895153534714888256694323060364090593906692889077294220902016707738101813741695817427157054583738511484754347790817568685939055368278079024365035694348150428775136136309;
            6'd7: xpb[73] = 1024'd61567275013439266055107950018515701879386535645079679246335136597939893155915232421229746926820606355337336021808834008245521245263239750759071033293222543121758489332019975249162848235843044211270719093758992090426038595368499359175191358346084980633757147369281740934675513540747313812925957138008591239749;
            6'd8: xpb[73] = 1024'd88086413684519838548523218221848578254255816040910445442687563978356577226375856897121863804174646450305976797418309357220461971849591191518246913051730197986822655603675859904419003582608794201639421479779882367110381373309841663766644205207415613476696726052624426501072948057129591931503763847242046343189;
            6'd9: xpb[73] = 1024'd114605552355600411041938486425181454629125096436741211639039991358773261296836481373013980681528686545274617573027784706195402698435942632277422792810237852851886821875331744559675158929374544192008123865800772643794724151251183968358097052068746246319636304735967112067470382573511870050081570556475501446629;
            6'd10: xpb[73] = 1024'd17057995342556242136554827223699898259295949706836293707260563674213050029987966938891026344225052330800108941179766620591279584181073738481438547552414466783260313577416411877301075084623088461066628643434423074114706078971629499984571329246847429895755980005192739603761289015965515151540687439083362065738;
            6'd11: xpb[73] = 1024'd43577134013636814629970095427032774634165230102667059903612991054629734100448591414783143221579092425768749716789241969566220310767425179240614427310922121648324479849072296532557230431388838451435331029455313350799048856912971804576024176108178062738695558688535425170158723532347793270118494148316817169178;
            6'd12: xpb[73] = 1024'd70096272684717387123385363630365651009034510498497826099965418435046418170909215890675260098933132520737390492398717318541161037353776619999790307069429776513388646120728181187813385778154588441804033415476203627483391634854314109167477022969508695581635137371878110736556158048730071388696300857550272272618;
            6'd13: xpb[73] = 1024'd96615411355797959616800631833698527383903790894328592296317845815463102241369840366567376976287172615706031268008192667516101763940128060758966186827937431378452812392384065843069541124920338432172735801497093904167734412795656413758929869830839328424574716055220796302953592565112349507274107566783727376058;
            6'd14: xpb[73] = 1024'd123134550026878532110215900037031403758773071290159358492670273195879786311830464842459493853641212710674672043617668016491042490526479501518142066586445086243516978664039950498325696471686088422541438187517984180852077190736998718350382716692169961267514294738563481869351027081494627625851914276017182479498;
            6'd15: xpb[73] = 1024'd25586993013834363204832240835549847388943924560254440560890845511319575044981950408336539516337578496200163411769649930886919376271610607722157821328621700174890470366124617815951612626934632691599942965151634611172059118457444249976856993870271144843633970007789109405641933523948272727311031158625043098607;
            6'd16: xpb[73] = 1024'd52106131684914935698247509038882723763813204956085206757243272891736259115442574884228656393691618591168804187379125279861860102857962048481333701087129355039954636637780502471207767973700382681968645351172524887856401896398786554568309840731601777686573548691131794972039368040330550845888837867858498202047;
            6'd17: xpb[73] = 1024'd78625270355995508191662777242215600138682485351915972953595700272152943185903199360120773271045658686137444962988600628836800829444313489240509580845637009905018802909436387126463923320466132672337347737193415164540744674340128859159762687592932410529513127374474480538436802556712828964466644577091953305487;
            6'd18: xpb[73] = 1024'd105144409027076080685078045445548476513551765747746739149948127652569627256363823836012890148399698781106085738598075977811741556030664929999685460604144664770082969181092271781720078667231882662706050123214305441225087452281471163751215534454263043372452706057817166104834237073095107083044451286325408408927;
            6'd19: xpb[73] = 1024'd7596852014031911779694386244066920143722619017841821218168699968009415989515309401889935811096064566631577106750057892207618441775796036203701215346321278701456460883176939099345994822480426931764554900847955871545069380001916695377689811632364226948572381327042793641125143515548752184503568168933269028036;
            6'd20: xpb[73] = 1024'd34115990685112484273109654447399796518591899413672587414521127348426100059975933877782052688450104661600217882359533241182559168362147476962877095104828933566520627154832823754602150169246176922133257286868846148229412157943258999969142658493694859791511960010385479207522578031931030303081374878166724131476;
            6'd21: xpb[73] = 1024'd60635129356193056766524922650732672893461179809503353610873554728842784130436558353674169565804144756568858657969008590157499894948498917722052974863336588431584793426488708409858305516011926912501959672889736424913754935884601304560595505355025492634451538693728164773920012548313308421659181587400179234916;
            6'd22: xpb[73] = 1024'd87154268027273629259940190854065549268330460205334119807225982109259468200897182829566286443158184851537499433578483939132440621534850358481228854621844243296648959698144593065114460862777676902870662058910626701598097713825943609152048352216356125477391117377070850340317447064695586540236988296633634338356;
            6'd23: xpb[73] = 1024'd113673406698354201753355459057398425643199740601164886003578409489676152271357807305458403320512224946506140209187959288107381348121201799240404734380351898161713125969800477720370616209543426893239364444931516978282440491767285913743501199077686758320330696060413535906714881581077864658814795005867089441796;
            6'd24: xpb[73] = 1024'd16125849685310032847971799855916869273370593871259968071798981805115941004509292871335448983208590732031631577339941202503258233866332905444420489122528512093086617671885145037996532364791971162297869222565167408602422419487731445369975476255787941896450371329639163443005788023531509760273911888474950060905;
            6'd25: xpb[73] = 1024'd42644988356390605341387068059249745648239874267090734268151409185532625074969917347227565860562630827000272352949416551478198960452684346203596368881036166958150783943541029693252687711557721152666571608586057685286765197429073749961428323117118574739389950012981849009403222539913787878851718597708405164345;
            6'd26: xpb[73] = 1024'd69164127027471177834802336262582622023109154662921500464503836565949309145430541823119682737916670921968913128558891900453139687039035786962772248639543821823214950215196914348508843058323471143035273994606947961971107975370416054552881169978449207582329528696324534575800657056296065997429525306941860267785;
            6'd27: xpb[73] = 1024'd95683265698551750328217604465915498397978435058752266660856263946365993215891166299011799615270711016937553904168367249428080413625387227721948128398051476688279116486852799003764998405089221133403976380627838238655450753311758359144334016839779840425269107379667220142198091572678344116007332016175315371225;
            6'd28: xpb[73] = 1024'd122202404369632322821632872669248374772847715454583032857208691326782677286351790774903916492624751111906194679777842598403021140211738668481124008156559131553343282758508683659021153751854971123772678766648728515339793531253100663735786863701110473268208686063009905708595526089060622234585138725408770474665;
            6'd29: xpb[73] = 1024'd24654847356588153916249213467766818403018568724678114925429263642222466019503276340780962155321116897431686047929824512798898025956869774685139762898735745484716774460593350976647069907103515392831183544282378945659775458973546195362261140879211656844328361332235533244886432531514267336044255608016631093774;
            6'd30: xpb[73] = 1024'd51173986027668726409664481671099694777887849120508881121781691022639150089963900816673079032675156992400326823539299861773838752543221215444315642657243400349780940732249235631903225253869265383199885930303269222344118236914888499953713987740542289687267940015578218811283867047896545454622062317250086197214;
            6'd31: xpb[73] = 1024'd77693124698749298903079749874432571152757129516339647318134118403055834160424525292565195910029197087368967599148775210748779479129572656203491522415751055214845107003905120287159380600635015373568588316324159499028461014856230804545166834601872922530207518698920904377681301564278823573199869026483541300654;
            6'd32: xpb[73] = 1024'd104212263369829871396495018077765447527626409912170413514486545783472518230885149768457312787383237182337608374758250559723720205715924096962667402174258710079909273275561004942415535947400765363937290702345049775712803792797573109136619681463203555373147097382263589944078736080661101691777675735716996404094;
            6'd33: xpb[73] = 1024'd6664706356785702491111358876283891157797263182265495582707118098912306964036635334334358450079602967863099742910232474119597091461055203166683156916435324011282764977645672260041452102649309632995795479978700206032785720518018640763093958641304738949266772651489217480369642523114746793236792618324857023203;
            6'd34: xpb[73] = 1024'd33183845027866274984526627079616767532666543578096261779059545479328991034497259810226475327433643062831740518519707823094537818047406643925859036674942978876346931249301556915297607449415059623364497865999590482717128498459360945354546805502635371792206351334831903046767077039497024911814599327558312126643;
            6'd35: xpb[73] = 1024'd59702983698946847477941895282949643907535823973927027975411972859745675104957884286118592204787683157800381294129183172069478544633758084685034916433450633741411097520957441570553762796180809613733200252020480759401471276400703249945999652363966004635145930018174588613164511555879303030392406036791767230083;
            6'd36: xpb[73] = 1024'd86222122370027419971357163486282520282405104369757794171764400240162359175418508762010709082141723252769022069738658521044419271220109525444210796191958288606475263792613326225809918142946559604101902638041371036085814054342045554537452499225296637478085508701517274179561946072261581148970212746025222333523;
            6'd37: xpb[73] = 1024'd112741261041107992464772431689615396657274384765588560368116827620579043245879133237902825959495763347737662845348133870019359997806460966203386675950465943471539430064269210881066073489712309594470605024062261312770156832283387859128905346086627270321025087384859959745959380588643859267548019455258677436963;
            6'd38: xpb[73] = 1024'd15193704028063823559388772488133840287445238035683642436337399936018831979030618803779871622192129133263154213500115784415236883551592072407402430692642557402912921766353878198691989644960853863529109801695911743090138760003833390755379623264728453897144762654085587282250287031097504369007136337866538056072;
            6'd39: xpb[73] = 1024'd41712842699144396052804040691466716662314518431514408632689827316435516049491243279671988499546169228231794989109591133390177610137943513166578310451150212267977088038009762853948144991726603853897812187716802019774481537945175695346832470126059086740084341337428272848647721547479782487584943047099993159512;
            6'd40: xpb[73] = 1024'd68231981370224968546219308894799593037183798827345174829042254696852200119951867755564105376900209323200435764719066482365118336724294953925754190209657867133041254309665647509204300338492353844266514573737692296458824315886517999938285316987389719583023920020770958415045156063862060606162749756333448262952;
            6'd41: xpb[73] = 1024'd94751120041305541039634577098132469412053079223175941025394682077268884190412492231456222254254249418169076540328541831340059063310646394684930069968165521998105420581321532164460455685258103834635216959758582573143167093827860304529738163848720352425963498704113643981442590580244338724740556465566903366392;
            6'd42: xpb[73] = 1024'd121270258712386113533049845301465345786922359619006707221747109457685568260873116707348339131608289513137717315938017180314999789896997835444105949726673176863169586852977416819716611032023853825003919345779472849827509871769202609121191010710050985268903077387456329547840025096626616843318363174800358469832;
            6'd43: xpb[73] = 1024'd23722701699341944627666186099983789417093212889101789289967681773125356994024602273225384794304655298663208684089999094710876675642128941648121704468849790794543078555062084137342527187272398094062424123413123280147491799489648140747665287888152168845022752656681957084130931539080261944777480057408219088941;
            6'd44: xpb[73] = 1024'd50241840370422517121081454303316665791962493284932555486320109153542041064485226749117501671658695393631849459699474443685817402228480382407297584227357445659607244826717968792598682534038148084431126509434013556831834577430990445339118134749482801687962331340024642650528366055462540063355286766641674192381;
            6'd45: xpb[73] = 1024'd76760979041503089614496722506649542166831773680763321682672536533958725134945851225009618549012735488600490235308949792660758128814831823166473463985865100524671411098373853447854837880803898074799828895454903833516177355372332749930570981610813434530901910023367328216925800571844818181933093475875129295821;
            6'd46: xpb[73] = 1024'd103280117712583662107911990709982418541701054076594087879024963914375409205406475700901735426366775583569131010918425141635698855401183263925649343744372755389735577370029738103110993227569648065168531281475794110200520133313675054522023828472144067373841488706710013783323235088227096300510900185108584399261;
            6'd47: xpb[73] = 1024'd5732560699539493202528331508500862171871907346689169947245536229815197938557961266778781089063141369094622379070407056031575741146314370129665098486549369321109069072114405420736909382818192334227036059109444540520502061034120586148498105650245250949961163975935641319614141530680741401970017067716445018370;
            6'd48: xpb[73] = 1024'd32251699370620065695943599711833738546741187742519936143597963610231882009018585742670897966417181464063263154679882405006516467732665810888840978245057024186173235343770290075993064729583942324595738445130334817204844838975462890739950952511575883792900742659278326886011576047063019520547823776949900121810;
            6'd49: xpb[73] = 1024'd58770838041700638189358867915166614921610468138350702339950390990648566079479210218563014843771221559031903930289357753981457194319017251648016858003564679051237401615426174731249220076349692314964440831151225093889187616916805195331403799372906516635840321342621012452409010563445297639125630486183355225250;
            6'd50: xpb[73] = 1024'd85289976712781210682774136118499491296479748534181468536302818371065250149939834694455131721125261654000544705898833102956397920905368692407192737762072333916301567887082059386505375423115442305333143217172115370573530394858147499922856646234237149478779900025963698018806445079827575757703437195416810328690;
            6'd51: xpb[73] = 1024'd111809115383861783176189404321832367671349028930012234732655245751481934220400459170347248598479301748969185481508308451931338647491720133166368617520579988781365734158737944041761530769881192295701845603193005647257873172799489804514309493095567782321719478709306383585203879596209853876281243904650265432130;
            6'd52: xpb[73] = 1024'd14261558370817614270805745120350811301519882200107316800875818066921722953551944736224294261175667534494676849660290366327215533236851239370384372262756602712739225860822611359387446925129736564760350380826656077577855100519935336140783770273668965897839153978532011121494786038663498977740360787258126051239;
            6'd53: xpb[73] = 1024'd40780697041898186764221013323683687676389162595938082997228245447338407024012569212116411138529707629463317625269765715302156259823202680129560252021264257577803392132478496014643602271895486555129052766847546354262197878461277640732236617134999598740778732661874696687892220555045777096318167496491581154679;
            6'd54: xpb[73] = 1024'd67299835712978759257636281527016564051258442991768849193580672827755091094473193688008528015883747724431958400879241064277096986409554120888736131779771912442867558404134380669899757618661236545497755152868436630946540656402619945323689463996330231583718311345217382254289655071428055214895974205725036258119;
            6'd55: xpb[73] = 1024'd93818974384059331751051549730349440426127723387599615389933100208171775164933818163900644893237787819400599176488716413252037712995905561647912011538279567307931724675790265325155912965426986535866457538889326907630883434343962249915142310857660864426657890028560067820687089587810333333473780914958491361559;
            6'd56: xpb[73] = 1024'd120338113055139904244466817933682316800997003783430381586285527588588459235394442639792761770591827914369239952098191762226978439582257002407087891296787222172995890947446149980412068312192736526235159924910217184315226212285304554506595157718991497269597468711902753387084524104192611452051587624191946464999;
            6'd57: xpb[73] = 1024'd22790556042095735339083158732200760431167857053525463654506099904028247968545928205669807433288193699894731320250173676622855325327388108611103646038963836104369382649530817298037984467441280795293664702543867614635208140005750086133069434897092680845717143981128380923375430546646256553510704506799807084108;
            6'd58: xpb[73] = 1024'd49309694713176307832498426935533636806037137449356229850858527284444932039006552681561924310642233794863372095859649025597796051913739549370279525797471490969433548921186701953294139814207030785662367088564757891319550917947092390724522281758423313688656722664471066489772865063028534672088511216033262187548;
            6'd59: xpb[73] = 1024'd75828833384256880325913695138866513180906417845186996047210954664861616109467177157454041187996273889832012871469124374572736778500090990129455405555979145834497715192842586608550295160972780776031069474585648168003893695888434695315975128619753946531596301347813752056170299579410812790666317925266717290988;
            6'd60: xpb[73] = 1024'd102347972055337452819328963342199389555775698241017762243563382045278300179927801633346158065350313984800653647078599723547677505086442430888631285314486800699561881464498471263806450507738530766399771860606538444688236473829776999907427975481084579374535880031156437622567734095793090909244124634500172394428;
            6'd61: xpb[73] = 1024'd4800415042293283913945304140717833185946551511112844311783954360718088913079287199223203728046679770326145015230581637943554390831573537092647040056663414630935373166583138581432366662987075035458276638240188875008218401550222531533902252659185762950655555300382065158858640538246736010703241517108033013537;
            6'd62: xpb[73] = 1024'd31319553713373856407360572344050709560815831906943610508136381741134772983539911675115320605400719865294785790840056986918495117417924977851822919815171069495999539438239023236688522009752825025826979024261079151692561179491564836125355099520516395793595133983724750725256075054629014129281048226341488116977;
            6'd63: xpb[73] = 1024'd57838692384454428900775840547383585935685112302774376704488809121551457054000536151007437482754759960263426566449532335893435844004276418610998799573678724361063705709894907891944677356518575016195681410281969428376903957432907140716807946381847028636534712667067436291653509571011292247858854935574943220417;
        endcase
    end

    always_comb begin
        case(flag[24][16:12])
            5'd0: xpb[74] = 1024'd0;
            5'd1: xpb[74] = 1024'd84357831055535001394191108750716462310554392698605142900841236501968141124461160626899554360108800055232067342059007684868376570590627859370174679332186379226127871981550792547200832703284325006564383796302859705061246735374249445308260793243177661479474291350410121858050944087393570366436661644808398323857;
            5'd2: xpb[74] = 1024'd44648966426945261389583290096618491876410358271474601673550617938959386911613182343784037505559925801020985276660521935157689300340035384185189233648041717518565069393530367756771426215051444291818569984218479563758132620527602117651543016803125873692128679286703185685995360100858507715754633462991202163383;
            5'd3: xpb[74] = 1024'd4940101798355521384975471442520521442266323844344060446259999375950632698765204060668520651011051546809903211262036185447002030089442909000203787963897055811002266805509942966342019726818563577072756172134099422455018505680954789994825240363074085904783067222996249513939776114323445065072605281174006002909;
            5'd4: xpb[74] = 1024'd89297932853890522779166580193236983752820716542949203347101235877918773823226364687568075011119851602041970553321043870315378600680070768370378467296083435037130138787060735513542852430102888583637139968436959127516265241055204235303086033606251747384257358573406371371990720201717015431509266925982404326766;
            5'd5: xpb[74] = 1024'd49589068225300782774558761539139013318676682115818662119810617314910019610378386404452558156570977347830888487922558120604691330429478293185393021611938773329567336199040310723113445941870007868891326156352578986213151126208556907646368257166199959596911746509699435199935136215181952780827238744165208166292;
            5'd6: xpb[74] = 1024'd9880203596711042769950942885041042884532647688688120892519998751901265397530408121337041302022103093619806422524072370894004060178885818000407575927794111622004533611019885932684039453637127154145512344268198844910037011361909579989650480726148171809566134445992499027879552228646890130145210562348012005818;
            5'd7: xpb[74] = 1024'd94238034652246044164142051635757505195087040387293263793361235253869406521991568748236595662130903148851873764583080055762380630769513677370582255259980490848132405592570678479884872156921452160709896140571058549971283746736159025297911273969325833289040425796402620885930496316040460496581872207156410329675;
            5'd8: xpb[74] = 1024'd54529170023656304159534232981659534760943005960162722566070616690860652309143590465121078807582028894640791699184594306051693360518921202185596809575835829140569603004550253689455465668688571445964082328486678408668169631889511697641193497529274045501694813732695684713874912329505397845899844025339214169201;
            5'd9: xpb[74] = 1024'd14820305395066564154926414327561564326798971533032181338779998127851898096295612182005561953033154640429709633786108556341006090268328727000611363891691167433006800416529828899026059180455690731218268516402298267365055517042864369984475721089222257714349201668988748541819328342970335195217815843522018008727;
            5'd10: xpb[74] = 1024'd99178136450601565549117523078278026637353364231637324239621234629820039220756772808905116313141954695661776975845116241209382660858956586370786043223877546659134672398080621446226891883740015737782652312705157972426302252417113815292736514332399919193823493019398870399870272430363905561654477488330416332584;
            5'd11: xpb[74] = 1024'd59469271822011825544509704424180056203209329804506783012330616066811285007908794525789599458593080441450694910446630491498695390608364111185800597539732884951571869810060196655797485395507135023036838500620777831123188137570466487636018737892348131406477880955691934227814688443828842910972449306513220172110;
            5'd12: xpb[74] = 1024'd19760407193422085539901885770082085769065295377376241785039997503802530795060816242674082604044206187239612845048144741788008120357771636000815151855588223244009067222039771865368078907274254308291024688536397689820074022723819159979300961452296343619132268891984998055759104457293780260290421124696024011636;
            5'd13: xpb[74] = 1024'd104118238248957086934092994520798548079619688075981384685881234005770671919521976869573636964153006242471680187107152426656384690948399495370989831187774602470136939203590564412568911610558579314855408484839257394881320758098068605287561754695474005098606560242395119913810048544687350626727082769504422335493;
            5'd14: xpb[74] = 1024'd64409373620367346929485175866700577645475653648850843458590615442761917706673998586458120109604131988260598121708666676945697420697807020186004385503629940762574136615570139622139505122325698600109594672754877253578206643251421277630843978255422217311260948178688183741754464558152287976045054587687226175019;
            5'd15: xpb[74] = 1024'd24700508991777606924877357212602607211331619221720302231299996879753163493826020303342603255055257734049516056310180927235010150447214545001018939819485279055011334027549714831710098634092817885363780860670497112275092528404773949974126201815370429523915336114981247569698880571617225325363026405870030014545;
            5'd16: xpb[74] = 1024'd109058340047312608319068465963319069521886011920325445132141233381721304618287180930242157615164057789281583398369188612103386721037842404371193619151671658281139206009100507378910931337377142891928164656973356817336339263779023395282386995058548091003389627465391369427749824659010795691799688050678428338402;
            5'd17: xpb[74] = 1024'd69349475418722868314460647309221099087741977493194903904850614818712550405439202647126640760615183535070501332970702862392699450787249929186208173467526996573576403421080082588481524849144262177182350844888976676033225148932376067625669218618496303216044015401684433255694240672475733041117659868861232177928;
            5'd18: xpb[74] = 1024'd29640610790133128309852828655123128653597943066064362677559996255703796192591224364011123906066309280859419267572217112682012180536657454001222727783382334866013600833059657798052118360911381462436537032804596534730111034085728739968951442178444515428698403337977497083638656685940670390435631687044036017454;
            5'd19: xpb[74] = 1024'd113998441845668129704043937405839590964152335764669505578401232757671937317052384990910678266175109336091486609631224797550388751127285313371397407115568714092141472814610450345252951064195706469000920829107456239791357769459978185277212235421622176908172694688387618941689600773334240756872293331852434341311;
            5'd20: xpb[74] = 1024'd74289577217078389699436118751741620530008301337538964351110614194663183104204406707795161411626235081880404544232739047839701480876692838186411961431424052384578670226590025554823544575962825754255107017023076098488243654613330857620494458981570389120827082624680682769634016786799178106190265150035238180837;
            5'd21: xpb[74] = 1024'd34580712588488649694828300097643650095864266910408423123819995631654428891356428424679644557077360827669322478834253298129014210626100363001426515747279390677015867638569600764394138087729945039509293204938695957185129539766683529963776682541518601333481470560973746597578432800264115455508236968218042020363;
            5'd22: xpb[74] = 1024'd118938543644023651089019408848360112406418659609013566024661232133622570015817589051579198917186160882901389820893260982997390781216728222371601195079465769903143739620120393311594970791014270046073677001241555662246376275140932975272037475784696262812955761911383868455629376887657685821944898613026440344220;
            5'd23: xpb[74] = 1024'd79229679015433911084411590194262141972274625181883024797370613570613815802969610768463682062637286628690307755494775233286703510966135747186615749395321108195580937032099968521165564302781389331327863189157175520943262160294285647615319699344644475025610149847676932283573792901122623171262870431209244183746;
            5'd24: xpb[74] = 1024'd39520814386844171079803771540164171538130590754752483570079995007605061590121632485348165208088412374479225690096289483576016240715543272001630303711176446488018134444079543730736157814548508616582049377072795379640148045447638319958601922904592687238264537783969996111518208914587560520580842249392048023272;
            5'd25: xpb[74] = 1024'd123878645442379172473994880290880633848684983453357626470921231509573202714582793112247719568197212429711293032155297168444392811306171131371804983043362825714146006425630336277936990517832833623146433173375655084701394780821887765266862716147770348717738829134380117969569153001981130887017503894200446347129;
            5'd26: xpb[74] = 1024'd84169780813789432469387061636782663414540949026227085243630612946564448501734814829132202713648338175500210966756811418733705541055578656186819537359218164006583203837609911487507584029599952908400619361291274943398280665975240437610144939707718560930393217070673181797513569015446068236335475712383250186655;
            5'd27: xpb[74] = 1024'd44460916185199692464779242982684692980396914599096544016339994383555694288886836546016685859099463921289128901358325669023018270804986181001834091675073502299020401249589486697078177541367072193654805549206894802095166551128593109953427163267666773143047605006966245625457985028911005585653447530566054026181;
            5'd28: xpb[74] = 1024'd4752051556609952460171424328586722546252880171966002789049375820546940076038858262901169004550589667078046835959839919312331000554393705816848645990928840591457598661569061906648771053134191478908991737122514660792052436281945782296709386827614985355701992943259309453402401042375942934971419348748857865707;
            5'd29: xpb[74] = 1024'd89109882612144953854362533079303184856807272870571145689890612322515081200500018889800723364659389722310114178018847604180707571145021565187023325323115219817585470643119854453849603756418516485473375533425374365853299171656195227604970180070792646835176284293669431311453345129769513301408080993557256189564;
            5'd30: xpb[74] = 1024'd49401017983555213849754714425205214422663238443440604462599993759506326987652040606685206510110515468099032112620361854470020300894429090002037879638970558110022668055099429663420197268185635770727561721340994224550185056809547899948252403630740859047830672229962495139397761143234450650726052811740060029090;
            5'd31: xpb[74] = 1024'd9692153354965473845146895771107243988519204016310063235309375196497572774804062323569689655561641213887950047221876104759333030643836614817052433954825896402459865467079004872990790779952755055981747909256614083247070941962900572291534627190689071260485060166255558967342177156699388000044024629922863868616;
        endcase
    end

    always_comb begin
        case(flag[25][5:0])
            6'd0: xpb[75] = 1024'd0;
            6'd1: xpb[75] = 1024'd109058340047312608319068465963319069521886011920325445132141233381721304618287180930242157615164057789281583398369188612103386721037842404371193619151671658281139206009100507378910931337377142891928164656973356817336339263779023395282386995058548091003389627465391369427749824659010795691799688050678428338402;
            6'd2: xpb[75] = 1024'd94049984410500475239338004521823706299073596714915206136150611698465713899265222950469244015670441269120017389280883789627709601234464474187227113287012275628587737448629797420191623483237080062546131705559473788308317677337150017599795420433866732739959351516665680825393121244092958366480686274731262192473;
            6'd3: xpb[75] = 1024'd79041628773688342159607543080328343076261181509504967140159990015210123180243264970696330416176824748958451380192578967152032481431086544003260607422352892976036268888159087461472315629097017233164098754145590759280296090895276639917203845809185374476529075567939992223036417829175121041161684498784096046544;
            6'd4: xpb[75] = 1024'd64033273136876209079877081638832979853448766304094728144169368331954532461221306990923416816683208228796885371104274144676355361627708613819294101557693510323484800327688377502753007774956954403782065802731707730252274504453403262234612271184504016213098799619214303620679714414257283715842682722836929900615;
            6'd5: xpb[75] = 1024'd49024917500064076000146620197337616630636351098684489148178746648698941742199349011150503217189591708635319362015969322200678241824330683635327595693034127670933331767217667544033699920816891574400032851317824701224252918011529884552020696559822657949668523670488615018323010999339446390523680946889763754686;
            6'd6: xpb[75] = 1024'd34016561863251942920416158755842253407823935893274250152188124965443351023177391031377589617695975188473753352927664499725001122020952753451361089828374745018381863206746957585314392066676828745017999899903941672196231331569656506869429121935141299686238247721762926415966307584421609065204679170942597608757;
            6'd7: xpb[75] = 1024'd19008206226439809840685697314346890185011520687864011156197503282187760304155433051604676018202358668312187343839359677249324002217574823267394583963715362365830394646276247626595084212536765915635966948490058643168209745127783129186837547310459941422807971773037237813609604169503771739885677394995431462828;
            6'd8: xpb[75] = 1024'd3999850589627676760955235872851526962199105482453772160206881598932169585133475071831762418708742148150621334751054854773646882414196893083428078099055979713278926085805537667875776358396703086253933997076175614140188158685909751504245972685778583159377695824311549211252900754585934414566675619048265316899;
            6'd9: xpb[75] = 1024'd113058190636940285080023701836170596484085117402779217292348114980653474203420656002073920033872799937432204733120243466877033603452039297454621697250727637994418132094906045046786707695773845978182098654049532431476527422464933146786632967744326674162767323289702918639002725413596730106366363669726693655301;
            6'd10: xpb[75] = 1024'd98049835000128152000293240394675233261272702197368978296357493297397883484398698022301006434379183417270638724031938644401356483648661367270655191386068255341866663534435335088067399841633783148800065702635649402448505836023059769104041393119645315899337047340977230036646021998678892781047361893779527509372;
            6'd11: xpb[75] = 1024'd83041479363316018920562778953179870038460286991958739300366871614142292765376740042528092834885566897109072714943633821925679363845283437086688685521408872689315194973964625129348091987493720319418032751221766373420484249581186391421449818494963957635906771392251541434289318583761055455728360117832361363443;
            6'd12: xpb[75] = 1024'd68033123726503885840832317511684506815647871786548500304376249930886702046354782062755179235391950376947506705855328999450002244041905506902722179656749490036763726413493915170628784133353657490035999799807883344392462663139313013738858243870282599372476495443525852831932615168843218130409358341885195217514;
            6'd13: xpb[75] = 1024'd53024768089691752761101856070189143592835456581138261308385628247631111327332824082982265635898333856785940696767024176974325124238527576718755673792090107384212257853023205211909476279213594660653966848394000315364441076697439636056266669245601241109046219494800164229575911753925380805090356565938029071585;
            6'd14: xpb[75] = 1024'd38016412452879619681371394628693780370023041375728022312395006564375520608310866103209352036404717336624374687678719354498648004435149646534789167927430724731660789292552495253190168425073531831271933896980117286336419490255566258373675094620919882845615943546074475627219208339007543479771354789990862925656;
            6'd15: xpb[75] = 1024'd23008056816067486601640933187198417147210626170317783316404384881119929889288908123436438436911100816462808678590414532022970884631771716350822662062771342079109320732081785294470860570933469001889900945566234257308397903813692880691083519996238524582185667597348787024862504924089706154452353014043696779727;
            6'd16: xpb[75] = 1024'd7999701179255353521910471745703053924398210964907544320413763197864339170266950143663524837417484296301242669502109709547293764828393786166856156198111959426557852171611075335751552716793406172507867994152351228280376317371819503008491945371557166318755391648623098422505801509171868829133351238096530633798;
            6'd17: xpb[75] = 1024'd117058041226567961840978937709022123446284222885232989452554996579585643788554131073905682452581542085582826067871298321650680485866236190538049775349783617707697058180711582714662484054170549064436032651125708045616715581150842898290878940430105257322145019114014467850255626168182664520933039288774958972200;
            6'd18: xpb[75] = 1024'd102049685589755828761248476267526760223471807679822750456564374896330053069532173094132768853087925565421260058782993499175003366062858260354083269485124235055145589620240872755943176200030486235053999699711825016588693994708969520608287365805423899058714743165288779247898922753264827195614037512827792826271;
            6'd19: xpb[75] = 1024'd87041329952943695681518014826031397000659392474412511460573753213074462350510215114359855253594309045259694049694688676699326246259480330170116763620464852402594121059770162797223868345890423405671966748297941987560672408267096142925695791180742540795284467216563090645542219338346989870295035736880626680342;
            6'd20: xpb[75] = 1024'd72032974316131562601787553384536033777846977269002272464583131529818871631488257134586941654100692525098128040606383854223649126456102399986150257755805469750042652499299452838504560491750360576289933796884058958532650821825222765243104216556061182531854191267837402043185515923429152544976033960933460534413;
            6'd21: xpb[75] = 1024'd57024618679319429522057091943040670555034562063592033468592509846563280912466299154814028054607076004936562031518079031747972006652724469802183751891146087097491183938828742879785252637610297746907900845470175929504629235383349387560512641931379824268423915319111713440828812508511315219657032184986294388484;
            6'd22: xpb[75] = 1024'd42016263042507296442326630501545307332222146858181794472601888163307690193444341175041114455113459484774996022429774209272294886849346539618217246026486704444939715378358032921065944783470234917525867894056292900476607648941476009877921067306698466004993639370386024838472109093593477894338030409039128242555;
            6'd23: xpb[75] = 1024'd27007907405695163362596169060049944109409731652771555476611266480052099474422383195268200855619842964613430013341469386796617767045968609434250740161827321792388246817887322962346636929330172088143834942642409871448586062499602632195329492682017107741563363421660336236115405678675640569019028633091962096626;
            6'd24: xpb[75] = 1024'd11999551768883030282865707618554580886597316447361316480620644796796508755400425215495287256126226444451864004253164564320940647242590679250284234297167939139836778257416613003627329075190109258761801991228526842420564476057729254512737918057335749478133087472934647633758702263757803243700026857144795950697;
            6'd25: xpb[75] = 1024'd121057891816195638601934173581873650408483328367686761612761878178517813373687606145737444871290284233733447402622353176424327368280433083621477853448839597420975984266517120382538260412567252150689966648201883659756903739836752649795124913115883840481522714938326017061508526922768598935499714907823224289099;
            6'd26: xpb[75] = 1024'd106049536179383505522203712140378287185670913162276522616771256495262222654665648165964531271796667713571881393534048353948650248477055153437511347584180214768424515706046410423818952558427189321307933696788000630728882153394879272112533338491202482218092438989600328459151823507850761610180713131876058143170;
            6'd27: xpb[75] = 1024'd91041180542571372442473250698882923962858497956866283620780634812006631935643690186191617672303051193410315384445743531472973128673677223253544841719520832115873047145575700465099644704287126491925900745374117601700860566953005894429941763866521123954662163040874639856795120092932924284861711355928891997241;
            6'd28: xpb[75] = 1024'd76032824905759239362742789257387560740046082751456044624790013128751041216621732206418704072809434673248749375357438708997296008870299293069578335854861449463321578585104990506380336850147063662543867793960234572672838980511132516747350189241839765691231887092148951254438416678015086959542709579981725851312;
            6'd29: xpb[75] = 1024'd61024469268947106283012327815892197517233667546045805628799391445495450497599774226645790473315818153087183366269133886521618889066921362885611829990202066810770110024634280547661028996007000833161834842546351543644817394069259139064758614617158407427801611143423262652081713263097249634223707804034559705383;
            6'd30: xpb[75] = 1024'd46016113632134973203281866374396834294421252340635566632808769762239859778577816246872876873822201632925617357180829064045941769263543432701645324125542684158218641464163570588941721141866938003779801891132468514616795807627385761382167039992477049164371335194697574049725009848179412308904706028087393559454;
            6'd31: xpb[75] = 1024'd31007757995322840123551404932901471071608837135225327636818148078984269059555858267099963274328585112764051348092524241570264649460165502517678818260883301505667172903692860630222413287726875174397768939718585485588774221185512383699575465367795690900941059245971885447368306433261574983585704252140227413525;
            6'd32: xpb[75] = 1024'd15999402358510707043820943491406107848796421929815088640827526395728678340533900287327049674834968592602485339004219419094587529656787572333712312396223918853115704343222150671503105433586812345015735988304702456560752634743639006016983890743114332637510783297246196845011603018343737658266702476193061267596;
            6'd33: xpb[75] = 1024'd991046721698573964090482049910744625984006724404849644836904712473087621511942307554136075341352072440919329915914596618910409853409642149745806531564536200564235782751440712783797579446749515633703036890819427532731048301765628334392316118432974374080507348520508242654899603425900332947700700245895121667;
            6'd34: xpb[75] = 1024'd110049386769011182283158948013229814147870018644730294776978138094194392239799123237796293690505409861722502728285103208722297130891252046520939425683236194481703441791851948091694728916823892407561867693864176244869070312080789023616779311176981065377470134813911877670404724262436696024747388750924323460069;
            6'd35: xpb[75] = 1024'd95041031132199049203428486571734450925057603439320055780987516410938801520777165258023380091011793341560936719196798386246620011087874116336972919818576811829151973231381238132975421062683829578179834742450293215841048725638915645934187736552299707114039858865186189068048020847518858699428386974977157314140;
            6'd36: xpb[75] = 1024'd80032675495386916123698025130239087702245188233909816784996894727683210801755207278250466491518176821399370710108493563770942891284496186153006413953917429176600504670910528174256113208543766748797801791036410186813027139197042268251596161927618348850609582916460500465691317432601021374109385199029991168211;
            6'd37: xpb[75] = 1024'd65024319858574783043967563688743724479432773028499577789006273044427620082733249298477552892024560301237804701020188741295265771481118255969039908089258046524049036110439818215536805354403703919415768839622527157785005552755168890569004587302936990587179306967734811863334614017683184048790383423082825022282;
            6'd38: xpb[75] = 1024'd50015964221762649964237102247248361256620357823089338793015651361172029363711291318704639292530943781076238691931883918819588651677740325785073402224598663871497567549969108256817497500263641090033735888208644128756983966313295512886413012678255632323749031019009123260977910602765346723471381647135658876353;
            6'd39: xpb[75] = 1024'd35007608584950516884506640805752998033807942617679099797025029677916438644689333338931725693037327260914672682843579096343911531874362395601106896359939281218946098989498398298098189646123578260651702936794761099728962379871422135203821438053574274060318755070283434658621207187847509398152379871188492730424;
            6'd40: xpb[75] = 1024'd19999252948138383804776179364257634810995527412268860801034407994660847925667375359158812093543710740753106673755274273868234412070984465417140390495279898566394630429027688339378881791983515431269669985380878070700940793429548757521229863428892915796888479121557746056264503772929672072833378095241326584495;
            6'd41: xpb[75] = 1024'd4990897311326250725045717922762271588183112206858621805043786311405257206645417379385898494050094220591540664666969451392557292267606535233173884630620515913843161868556978380659573937843452601887637033966995041672919206987675379838638288804211557533458203172832057453907800358011834747514376319294160438566;
            6'd42: xpb[75] = 1024'd114049237358638859044114183886081341110069124127184066937185019693126561824932598309628056109214152009873124063036158063495944013305448939604367503782292174194982367877657485759570505275220595493815801690940351859009258470766698775121025283862759648536847830638223426881657625017022630439314064369972588776968;
            6'd43: xpb[75] = 1024'd99040881721826725964383722444585977887256708921773827941194398009870971105910640329855142509720535489711558053947853241020266893502071009420400997917632791542430899317186775800851197421080532664433768739526468829981236884324825397438433709238078290273417554689497738279300921602104793113995062594025422631039;
            6'd44: xpb[75] = 1024'd84032526085014592884653261003090614664444293716363588945203776326615380386888682350082228910226918969549992044859548418544589773698693079236434492052973408889879430756716065842131889566940469835051735788112585800953215297882952019755842134613396932009987278740772049676944218187186955788676060818078256485110;
            6'd45: xpb[75] = 1024'd69024170448202459804922799561595251441631878510953349949213154643359789667866724370309315310733302449388426035771243596068912653895315149052467986188314026237327962196245355883412581712800407005669702836698702771925193711441078642073250559988715573746557002792046361074587514772269118463357059042131090339181;
            6'd46: xpb[75] = 1024'd54015814811390326725192338120099888218819463305543110953222532960104198948844766390536401711239685929226860026682938773593235534091937218868501480323654643584776493635774645924693273858660344176287669885284819742897172124999205264390658985364034215483126726843320672472230811357351281138038057266183924193252;
            6'd47: xpb[75] = 1024'd39007459174578193645461876678604524996007048100132871957231911276848608229822808410763488111746069409065294017594633951117558414288559288684534974458995260932225025075303935965973966004520281346905636933870936713869150538557331886708067410739352857219696450894594983869874107942433443812719055490236758047323;
            6'd48: xpb[75] = 1024'd23999103537766060565731415237109161773194632894722632961241289593593017510800850430990574512252452888903728008506329128641881294485181358500568468594335878279673556514833226007254658150380218517523603982457053684841128952115458509025475836114671498956266174945869295267517404527515606487400053714289591901394;
            6'd49: xpb[75] = 1024'd8990747900953927486000953795613798550382217689312393965250667910337426791778892451217660912758836368742161999418024306166204174681803428316601962729676495627122087954362516048535350296240155688141571031043170655813107365673585131342884261489990140692835898997143606665160701112597769162081051938342425755465;
            6'd50: xpb[75] = 1024'd118049087948266535805069419758932868072268229609637839097391901292058731410066073381459818527922894158023745397787212918269590895719645832687795581881348153908261293963463023427446281633617298580069735688016527473149446629452608526625271256548538231696225526462534976092910525771608564853880739989020854093867;
            6'd51: xpb[75] = 1024'd103040732311454402725338958317437504849455814404227600101401279608803140691044115401686904928429277637862179388698908095793913775916267902503829076016688771255709825402992313468726973779477235750687702736602644444121425043010735148942679681923856873432795250513809287490553822356690727528561738213073687947938;
            6'd52: xpb[75] = 1024'd88032376674642269645608496875942141626643399198817361105410657925547549972022157421913991328935661117700613379610603273318236656112889972319862570152029388603158356842521603510007665925337172921305669785188761415093403456568861771260088107299175515169364974565083598888197118941772890203242736437126521802009;
            6'd53: xpb[75] = 1024'd73024021037830136565878035434446778403830983993407122109420036242291959253000199442141077729442044597539047370522298450842559536309512042135896064287370005950606888282050893551288358071197110091923636833774878386065381870126988393577496532674494156905934698616357910285840415526855052877923734661179355656080;
            6'd54: xpb[75] = 1024'd58015665401018003486147573992951415181018568787996883113429414559036368533978241462368164129948428077377481361433993628366882416506134111951929558422710623298055419721580183592569050217057047262541603882360995357037360283685115015894904958049812798642504422667632221683483712111937215552604732885232189510151;
            6'd55: xpb[75] = 1024'd43007309764205870406417112551456051958206153582586644117438792875780777814956283482595250530454811557215915352345688805891205296702756181767963052558051240645503951161109473633849742362916984433159570930947112328009338697243241638212313383425131440379074146718906533081127008697019378227285731109285023364222;
            6'd56: xpb[75] = 1024'd27998954127393737326686651109960688735393738377176405121448171192525187095934325502822336930961195037054349343257383983415528176899378251583996546693391857992952482600638763675130434508776921603777537979533229298981317110801368260529721808800450082115643870770180844478770305282101540901966729333337857218293;
            6'd57: xpb[75] = 1024'd12990598490581604246956189668465325512581323171766166125457549509269596376912367523049423331467578516892783334169079160939851057096000321400030040828732475340401014040168053716411126654636858774395505028119346269953295524359494882847130234175768723852213594821455155876413601867183703576647727557390691072364;
            6'd58: xpb[75] = 1024'd122048938537894212566024655631784395034467335092091611257598782890990900995199548453291580946631636306174366732538267773043237778133842725771223659980404133621540220049268561095322057992014001666323669685092703087289634788138518278129517229234316814855603222286846525304163426526194499268447415608069119410766;
            6'd59: xpb[75] = 1024'd107040582901082079486294194190289031811654919886681372261608161207735310276177590473518667347138019786012800723449962950567560658330464795587257154115744750968988751488797851136602750137873938836941636733678820058261613201696644900446925654609635456592172946338120836701806723111276661943128413832121953264837;
            6'd60: xpb[75] = 1024'd92032227264269946406563732748793668588842504681271133265617539524479719557155632493745753747644403265851234714361658128091883538527086865403290648251085368316437282928327141177883442283733876007559603782264937029233591615254771522764334079984954098328742670389395148099450019696358824617809412056174787118908;
            6'd61: xpb[75] = 1024'd77023871627457813326833271307298305366030089475860894269626917841224128838133674513972840148150786745689668705273353305616206418723708935219324142386425985663885814367856431219164134429593813178177570830851054000205570028812898145081742505360272740065312394440669459497093316281440987292490410280227620972979;
            6'd62: xpb[75] = 1024'd62015515990645680247102809865802942143217674270450655273636296157968538119111716534199926548657170225528102696185048483140529298920331005035357636521766603011334345807385721260444826575453750348795537879437170971177548442371024767399150930735591381801882118491943770894736612866523149967171408504280454827050;
            6'd63: xpb[75] = 1024'd47007160353833547167372348424307578920405259065040416277645674474712947400089758554427012949163553705366536687096743660664852179116953074851391130657107220358782877246915011301725518721313687519413504928023287942149526855929151389716559356110910023538451842543218082292379909451605312641852406728333288681121;
        endcase
    end

    always_comb begin
        case(flag[25][11:6])
            6'd0: xpb[76] = 1024'd0;
            6'd1: xpb[76] = 1024'd31998804717021414087641886982812215697592843859630177281655052791457356681067800574654099349669937185204970678008438838189175059313575144667424624792447837706231408686444301343006210867173624690031471976609404913121505269487278012033967781486228665275021566594492393690023206036687475316533404952386122535192;
            6'd2: xpb[76] = 1024'd63997609434042828175283773965624431395185687719260354563310105582914713362135601149308198699339874370409941356016877676378350118627150289334849249584895675412462817372888602686012421734347249380062943953218809826243010538974556024067935562972457330550043133188984787380046412073374950633066809904772245070384;
            6'd3: xpb[76] = 1024'd95996414151064242262925660948436647092778531578890531844965158374372070043203401723962298049009811555614912034025316514567525177940725434002273874377343513118694226059332904029018632601520874070094415929828214739364515808461834036101903344458685995825064699783477181070069618110062425949600214857158367605576;
            6'd4: xpb[76] = 1024'd3928523183960914951768620526434430045672948312785024998488356100852531386962063388601326184022074431376733304576261918177636396413080244114538374153460309891234960176205988034394604277177293038815690298050379806121660227728215275170892556261685211833266362963852516729986296072821268249014929982918895656437;
            6'd5: xpb[76] = 1024'd35927327900982329039410507509246645743265792172415202280143408892309888068029863963255425533692011616581703982584700756366811455726655388781962998945908147597466368862650289377400815144350917728847162274659784719243165497215493287204860337747913877108287929558344910420009502109508743565548334935305018191629;
            6'd6: xpb[76] = 1024'd67926132618003743127052394492058861440858636032045379561798461683767244749097664537909524883361948801786674660593139594555986515040230533449387623738355985303697777549094590720407026011524542418878634251269189632364670766702771299238828119234142542383309496152837304110032708146196218882081739887691140726821;
            6'd7: xpb[76] = 1024'd99924937335025157214694281474871077138451479891675556843453514475224601430165465112563624233031885986991645338601578432745161574353805678116812248530803823009929186235538892063413236878698167108910106227878594545486176036190049311272795900720371207658331062747329697800055914182883694198615144840077263262013;
            6'd8: xpb[76] = 1024'd7857046367921829903537241052868860091345896625570049996976712201705062773924126777202652368044148862753466609152523836355272792826160488229076748306920619782469920352411976068789208554354586077631380596100759612243320455456430550341785112523370423666532725927705033459972592145642536498029859965837791312874;
            6'd9: xpb[76] = 1024'd39855851084943243991179128035681075788938740485200227278631764993162419454991927351856751717714086047958437287160962674544447852139735632896501373099368457488701329038856277411795419421528210767662852572710164525364825724943708562375752894009599088941554292522197427149995798182330011814563264918223913848066;
            6'd10: xpb[76] = 1024'd71854655801964658078821015018493291486531584344830404560286817784619776136059727926510851067384023233163407965169401512733622911453310777563925997891816295194932737725300578754801630288701835457694324549319569438486330994430986574409720675495827754216575859116689820840019004219017487131096669870610036383258;
            6'd11: xpb[76] = 1024'd103853460518986072166462902001305507184124428204460581841941870576077132817127528501164950417053960418368378643177840350922797970766885922231350622684264132901164146411744880097807841155875460147725796525928974351607836263918264586443688456982056419491597425711182214530042210255704962447630074822996158918450;
            6'd12: xpb[76] = 1024'd11785569551882744855305861579303290137018844938355074995465068302557594160886190165803978552066223294130199913728785754532909189239240732343615122460380929673704880528617964103183812831531879116447070894151139418364980683184645825512677668785055635499799088891557550189958888218463804747044789948756686969311;
            6'd13: xpb[76] = 1024'd43784374268904158942947748562115505834611688797985252277120121094014950841953990740458077901736160479335170591737224592722084248552815877011039747252828767379936289215062265446190023698705503806478542870760544331486485952671923837546645450271284300774820655486049943879982094255151280063578194901142809504503;
            6'd14: xpb[76] = 1024'd75783178985925573030589635544927721532204532657615429558775173885472307523021791315112177251406097664540141269745663430911259307866391021678464372045276605086167697901506566789196234565879128496510014847369949244607991222159201849580613231757512966049842222080542337570005300291838755380111599853528932039695;
            6'd15: xpb[76] = 1024'd107781983702946987118231522527739937229797376517245606840430226676929664204089591889766276601076034849745111947754102269100434367179966166345888996837724442792399106587950868132202445433052753186541486823979354157729496491646479861614581013243741631324863788675034731260028506328526230696645004805915054574887;
            6'd16: xpb[76] = 1024'd15714092735843659807074482105737720182691793251140099993953424403410125547848253554405304736088297725506933218305047672710545585652320976458153496613841239564939840704823952137578417108709172155262761192201519224486640910912861100683570225046740847333065451855410066919945184291285072996059719931675582625748;
            6'd17: xpb[76] = 1024'd47712897452865073894716369088549935880284637110770277275608477194867482228916054129059404085758234910711903896313486510899720644965896121125578121406289077271171249391268253480584627975882796845294233168810924137608146180400139112717538006532969512608087018449902460609968390327972548312593124884061705160940;
            6'd18: xpb[76] = 1024'd79711702169886487982358256071362151577877480970400454557263529986324838909983854703713503435428172095916874574321925349088895704279471265793002746198736914977402658077712554823590838843056421535325705145420329050729651449887417124751505788019198177883108585044394854299991596364660023629126529836447827696132;
            6'd19: xpb[76] = 1024'd111710506886907902070000143054174367275470324830030631838918582777782195591051655278367602785098109281121845252330364187278070763593046410460427370991184752683634066764156856166597049710230046225357177122029733963851156719374695136785473569505426843158130151638887247990014802401347498945659934788833950231324;
            6'd20: xpb[76] = 1024'd19642615919804574758843102632172150228364741563925124992441780504262656934810316943006630920110372156883666522881309590888181982065401220572691870767301549456174800881029940171973021385886465194078451490251899030608301138641076375854462781308426059166331814819262583649931480364106341245074649914594478282185;
            6'd21: xpb[76] = 1024'd51641420636825988846484989614984365925957585423555302274096833295720013615878117517660730269780309342088637200889748429077357041378976365240116495559749387162406209567474241514979232253060089884109923466861303943729806408128354387888430562794654724441353381413754977339954686400793816561608054866980600817377;
            6'd22: xpb[76] = 1024'd83640225353847402934126876597796581623550429283185479555751886087177370296945918092314829619450246527293607878898187267266532100692551509907541120352197224868637618253918542857985443120233714574141395443470708856851311677615632399922398344280883389716374948008247371029977892437481291878141459819366723352569;
            6'd23: xpb[76] = 1024'd115639030070868817021768763580608797321143273142815656837406938878634726978013718666968928969120183712498578556906626105455707160006126654574965745144645062574869026940362844200991653987407339264172867420080113769972816947102910411956366125767112054991396514602739764720001098474168767194674864771752845887761;
            6'd24: xpb[76] = 1024'd23571139103765489710611723158606580274037689876710149990930136605115188321772380331607957104132446588260399827457571509065818378478481464687230244920761859347409761057235928206367625663063758232894141788302278836729961366369291651025355337570111270999598177783115100379917776436927609494089579897513373938622;
            6'd25: xpb[76] = 1024'd55569943820786903798253610141418795971630533736340327272585189396572545002840180906262056453802383773465370505466010347254993437792056609354654869713209697053641169743680229549373836530237382922925613764911683749851466635856569663059323119056339936274619744377607494069940982473615084810622984849899496473814;
            6'd26: xpb[76] = 1024'd87568748537808317885895497124231011669223377595970504554240242188029901683907981480916155803472320958670341183474449185444168497105631754022079494505657534759872578430124530892380047397411007612957085741521088662972971905343847675093290900542568601549641310972099887759964188510302560127156389802285619009006;
            6'd27: xpb[76] = 1024'd119567553254829731973537384107043227366816221455600681835895294979487258364975782055570255153142258143875311861482888023633343556419206898689504119298105372466103987116568832235386258264584632302988557718130493576094477174831125687127258682028797266824662877566592281449987394546990035443689794754671741544198;
            6'd28: xpb[76] = 1024'd27499662287726404662380343685041010319710638189495174989418492705967719708734443720209283288154521019637133132033833427243454774891561708801768619074222169238644721233441916240762229940241051271709832086352658642851621594097506926196247893831796482832864540746967617109904072509748877743104509880432269595059;
            6'd29: xpb[76] = 1024'd59498467004747818750022230667853226017303482049125352271073545497425076389802244294863382637824458204842103810042272265432629834205136853469193243866670006944876129919886217583768440807414675961741304062962063555973126863584784938230215675318025148107886107341460010799927278546436353059637914832818392130251;
            6'd30: xpb[76] = 1024'd91497271721769232837664117650665441714896325908755529552728598288882433070870044869517481987494395390047074488050711103621804893518711998136617868659117844651107538606330518926774651674588300651772776039571468469094632133072062950264183456804253813382907673935952404489950484583123828376171319785204514665443;
            6'd31: xpb[76] = 1024'd123496076438790646925306004633477657412489169768385706834383651080339789751937845444171581337164332575252045166059149941810979952832287142804042493451565682357338947292774820269780862541761925341804248016180873382216137402559340962298151238290482478657929240530444798179973690619811303692704724737590637200635;
            6'd32: xpb[76] = 1024'd31428185471687319614148964211475440365383586502280199987906848806820251095696507108810609472176595451013866436610095345421091171304641952916306993227682479129879681409647904275156834217418344310525522384403038448973281821825722201367140450093481694666130903710820133839890368582570145992119439863351165251496;
            6'd33: xpb[76] = 1024'd63426990188708733701790851194287656062976430361910377269561901598277607776764307683464708821846532636218837114618534183610266230618217097583731618020130316836111090096092205618163045084591969000556994361012443362094787091313000213401108231579710359941152470305312527529913574619257621308652844815737287786688;
            6'd34: xpb[76] = 1024'd95425794905730147789432738177099871760569274221540554551216954389734964457832108258118808171516469821423807792626973021799441289931792242251156242812578154542342498782536506961169255951765593690588466337621848275216292360800278225435076013065939025216174036899804921219936780655945096625186249768123410321880;
            6'd35: xpb[76] = 1024'd3357903938626820478275697755097654713463690955435047704740152116215425801590769922757836306528732697185629063177918425409552508404147052363420742588694951314883232899409590966545227627422012659309740705844013341973436780066659464504065224868938241224375700080180256879853458618703938924600964893883938372741;
            6'd36: xpb[76] = 1024'd35356708655648234565917584737909870411056534815065224986395204907672782482658570497411935656198669882390599741186357263598727567717722197030845367381142789021114641585853892309551438494595637349341212682453418255094942049553937476538033006355166906499397266674672650569876664655391414241134369846270060907933;
            6'd37: xpb[76] = 1024'd67355513372669648653559471720722086108649378674695402268050257699130139163726371072066035005868607067595570419194796101787902627031297341698269992173590626727346050272298193652557649361769262039372684659062823168216447319041215488572000787841395571774418833269165044259899870692078889557667774798656183443125;
            6'd38: xpb[76] = 1024'd99354318089691062741201358703534301806242222534325579549705310490587495844794171646720134355538544252800541097203234939977077686344872486365694616966038464433577458958742494995563860228942886729404156635672228081337952588528493500605968569327624237049440399863657437949923076728766364874201179751042305978317;
            6'd39: xpb[76] = 1024'd7286427122587735430044318281532084759136639268220072703228508217067957188552833311359162490550807128562362367754180343587188904817227296477959116742155261206118193075615579000939831904599305698125431003894393148095097007794874739674957781130623453057642063044032773609839754691525207173615894876802834029178;
            6'd40: xpb[76] = 1024'd39285231839609149517686205264344300456729483127850249984883561008525313869620633886013261840220744313767333045762619181776363964130802441145383741534603098912349601762059880343946042771772930388156902980503798061216602277282152751708925562616852118332663629638525167299862960728212682490149299829188956564370;
            6'd41: xpb[76] = 1024'd71284036556630563605328092247156516154322326987480427266538613799982670550688434460667361189890681498972303723771058019965539023444377585812808366327050936618581010448504181686952253638946555078188374957113202974338107546769430763742893344103080783607685196233017560989886166764900157806682704781575079099562;
            6'd42: xpb[76] = 1024'd103282841273651977692969979229968731851915170847110604548193666591440027231756235035321460539560618684177274401779496858154714082757952730480232991119498774324812419134948483029958464506120179768219846933722607887459612816256708775776861125589309448882706762827509954679909372801587633123216109733961201634754;
            6'd43: xpb[76] = 1024'd11214950306548650381812938807966514804809587581005097701716864317920488575514896699960488674572881559939095672330442261764825301230307540592497490895615571097353153251821567035334436181776598736941121301944772954216757235523090014845850337392308664890908426007885290339826050764346475422630824859721729685615;
            6'd44: xpb[76] = 1024'd43213755023570064469454825790778730502402431440635274983371917109377845256582697274614588024242818745144066350338881099954000360543882685259922115688063408803584561938265868378340647048950223426972593278554177867338262505010368026879818118878537330165929992602377684029849256801033950739164229812107852220807;
            6'd45: xpb[76] = 1024'd75212559740591478557096712773590946199995275300265452265026969900835201937650497849268687373912755930349037028347319938143175419857457829927346740480511246509815970624710169721346857916123848117004065255163582780459767774497646038913785900364765995440951559196870077719872462837721426055697634764493974755999;
            6'd46: xpb[76] = 1024'd107211364457612892644738599756403161897588119159895629546682022692292558618718298423922786723582693115554007706355758776332350479171032974594771365272959084216047379311154471064353068783297472807035537231772987693581273043984924050947753681850994660715973125791362471409895668874408901372231039716880097291191;
            6'd47: xpb[76] = 1024'd15143473490509565333581559334400944850482535893790122700205220418773019962476960088561814858594955991315828976906704179942461697643387784707035865049075880988588113428027555069729040458953891775756811599995152760338417463251305290016742893653993876724174788971737807069812346837167743671645754842640625342052;
            6'd48: xpb[76] = 1024'd47142278207530979421223446317213160548075379753420299981860273210230376643544760663215914208264893176520799654915143018131636756956962929374460489841523718694819522114471856412735251326127516465788283576604557673459922732738583302050710675140222541999196355566230200759835552873855218988179159795026747877244;
            6'd49: xpb[76] = 1024'd79141082924552393508865333300025376245668223613050477263515326001687733324612561237870013557934830361725770332923581856320811816270538074041885114633971556401050930800916157755741462193301141155819755553213962586581428002225861314084678456626451207274217922160722594449858758910542694304712564747412870412436;
            6'd50: xpb[76] = 1024'd111139887641573807596507220282837591943261067472680654545170378793145090005680361812524112907604767546930741010932020694509986875584113218709309739426419394107282339487360459098747673060474765845851227529823367499702933271713139326118646238112679872549239488755214988139881964947230169621245969699798992947628;
            6'd51: xpb[76] = 1024'd19071996674470480285350179860835374896155484206575147698693576519625551349439023477163141042617030422692562281482966098120098094056468028821574239202536190879823073604233543104123644736131184814572501898045532566460077690979520565187635449915679088557441151935590323799798642909989011920660684825559520998489;
            6'd52: xpb[76] = 1024'd51070801391491894372992066843647590593748328066205324980348629311082908030506824051817240392286967607897532959491404936309273153370043173488998863994984028586054482290677844447129855603304809504603973874654937479581582960466798577221603231401907753832462718530082717489821848946676487237194089777945643533681;
            6'd53: xpb[76] = 1024'd83069606108513308460633953826459806291341171925835502262003682102540264711574624626471339741956904793102503637499843774498448212683618318156423488787431866292285890977122145790136066470478434194635445851264342392703088229954076589255571012888136419107484285124575111179845054983363962553727494730331766068873;
            6'd54: xpb[76] = 1024'd115068410825534722548275840809272021988934015785465679543658734893997621392642425201125439091626841978307474315508282612687623271997193462823848113579879703998517299663566447133142277337652058884666917827873747305824593499441354601289538794374365084382505851719067504869868261020051437870260899682717888604065;
            6'd55: xpb[76] = 1024'd23000519858431395237118800387269804941828432519360172697181932620478082736401086865764467226639104854069295586059228016297734490469548272936112613355996500771058033780439531138518249013308477853388192196095912372581737918707735840358528006177364300390707514899442840529784938982810280169675614808478416654926;
            6'd56: xpb[76] = 1024'd54999324575452809324760687370082020639421276378990349978836985411935439417468887440418566576309042039274266264067666854486909549783123417603537238148444338477289442466883832481524459880482102543419664172705317285703243188195013852392495787663592965665729081493935234219808145019497755486209019760864539190118;
            6'd57: xpb[76] = 1024'd86998129292474223412402574352894236337014120238620527260492038203392796098536688015072665925978979224479236942076105692676084609096698562270961862940892176183520851153328133824530670747655727233451136149314722198824748457682291864426463569149821630940750648088427627909831351056185230802742424713250661725310;
            6'd58: xpb[76] = 1024'd118996934009495637500044461335706452034606964098250704542147090994850152779604488589726765275648916409684207620084544530865259668410273706938386487733340013889752259839772435167536881614829351923482608125924127111946253727169569876460431350636050296215772214682920021599854557092872706119275829665636784260502;
            6'd59: xpb[76] = 1024'd26929043042392310188887420913704234987501380832145197695670288721330614123363150254365793410661179285446028890635489934475370886882628517050650987509456810662292993956645519172912853290485770892203882494146292178703398146435951115529420562439049512223973877863295357259771235055631548418690544791397312311363;
            6'd60: xpb[76] = 1024'd58927847759413724276529307896516450685094224691775374977325341512787970804430950829019892760331116470650999568643928772664545946196203661718075612301904648368524402643089820515919064157659395582235354470755697091824903415923229127563388343925278177498995444457787750949794441092319023735223949743783434846555;
            6'd61: xpb[76] = 1024'd90926652476435138364171194879328666382687068551405552258980394304245327485498751403673992110001053655855970246652367610853721005509778806385500237094352486074755811329534121858925275024833020272266826447365102004946408685410507139597356125411506842774017011052280144639817647129006499051757354696169557381747;
            6'd62: xpb[76] = 1024'd122925457193456552451813081862140882080279912411035729540635447095702684166566551978328091459670990841060940924660806449042896064823353951052924861886800323780987220015978423201931485892006644962298298423974506918067913954897785151631323906897735508049038577646772538329840853165693974368290759648555679916939;
            6'd63: xpb[76] = 1024'd30857566226353225140656041440138665033174329144930222694158644822183145510325213642967119594683253716822762195211751852653007283295708761165189361662917120553527954132851507207307457567663063931019572792196671984825058374164166390700313118700734724057240240827147873989757531128452816667705474774316207967800;
        endcase
    end

    always_comb begin
        case(flag[25][16:12])
            5'd0: xpb[77] = 1024'd0;
            5'd1: xpb[77] = 1024'd62856370943374639228297928422950880730767173004560399975813697613640502191393014217621218944353190902027732873220190690842182342609283905832613986455364958259759362819295808550313668434836688621051044768806076897946563643651444402734280900186963389332261807421640267679780737165140291984238879726702330502992;
            5'd2: xpb[77] = 1024'd1646046202624537057796929441087328716835918883385115823495540162304109045476889525227366674048707494612316338982887947105300844377347477110067847894398875585828051069020399762997097678156171520791891929224913949528766437081992032503583230690697329397703711429163477329454946256351950951359069626779066521653;
            5'd3: xpb[77] = 1024'd64502417145999176286094857864038209447603091887945515799309237775944611236869903742848585618401898396640049212203078637947483186986631382942681834349763833845587413888316208313310766112992860141842936698030990847475330080733436435237864130877660718729965518850803745009235683421492242935597949353481397024645;
            5'd4: xpb[77] = 1024'd3292092405249074115593858882174657433671837766770231646991080324608218090953779050454733348097414989224632677965775894210601688754694954220135695788797751171656102138040799525994195356312343041583783858449827899057532874163984065007166461381394658795407422858326954658909892512703901902718139253558133043306;
            5'd5: xpb[77] = 1024'd66148463348623713343891787305125538164439010771330631622804777938248720282346793268075952292450605891252365551185966585052784031363978860052749682244162709431415464957336608076307863791149031662634828627255904797004096517815428467741447361568358048127669230279967222338690629677844193886957018980260463546298;
            5'd6: xpb[77] = 1024'd4938138607873611173390788323261986150507756650155347470486620486912327136430668575682100022146122483836949016948663841315902533132042431330203543683196626757484153207061199288991293034468514562375675787674741848586299311245976097510749692072091988193111134287490431988364838769055852854077208880337199564959;
            5'd7: xpb[77] = 1024'd67794509551248250401688716746212866881274929654715747446300318100552829327823682793303318966499313385864681890168854532158084875741326337162817530138561585017243516026357007839304961469305203183426720556480818746532862954897420500245030592259055377525372941709130699668145575934196144838316088607039530067951;
            5'd8: xpb[77] = 1024'd6584184810498148231187717764349314867343675533540463293982160649216436181907558100909466696194829978449265355931551788421203377509389908440271391577595502343312204276081599051988390712624686083167567716899655798115065748327968130014332922762789317590814845716653909317819785025407803805436278507116266086612;
            5'd9: xpb[77] = 1024'd69440555753872787459485646187300195598110848538100863269795858262856938373300572318530685640548020880476998229151742479263385720118673814272885378032960460603071567095377407602302059147461374704218612485705732696061629391979412532748613822949752706923076653138294176997600522190548095789675158233818596589604;
            5'd10: xpb[77] = 1024'd8230231013122685288984647205436643584179594416925579117477700811520545227384447626136833370243537473061581694914439735526504221886737385550339239471994377929140255345101998814985488390780857603959459646124569747643832185409960162517916153453486646988518557145817386647274731281759754756795348133895332608265;
            5'd11: xpb[77] = 1024'd71086601956497324517282575628387524314946767421485979093291398425161047418777461843758052314596728375089314568134630426368686564496021291382953225927359336188899618164397807365299156825617546225010504414930646645590395829061404565252197053640450036320780364567457654327055468446900046741034227860597663111257;
            5'd12: xpb[77] = 1024'd9876277215747222346781576646523972301015513300310694940973240973824654272861337151364200044292244967673898033897327682631805066264084862660407087366393253514968306414122398577982586068937029124751351575349483697172598622491952195021499384144183976386222268574980863976729677538111705708154417760674399129918;
            5'd13: xpb[77] = 1024'd72732648159121861575079505069474853031782686304871094916786938587465156464254351368985418988645435869701630907117518373473987408873368768493021073821758211774727669233418207128296254503773717745802396344155560595119162266143396597755780284331147365718484075996621131656510414703251997692393297487376729632910;
            5'd14: xpb[77] = 1024'd11522323418371759404578506087611301017851432183695810764468781136128763318338226676591566718340952462286214372880215629737105910641432339770474935260792129100796357483142798340979683747093200645543243504574397646701365059573944227525082614834881305783925980004144341306184623794463656659513487387453465651571;
            5'd15: xpb[77] = 1024'd74378694361746398632876434510562181748618605188256210740282478749769265509731240894212785662694143364313947246100406320579288253250716245603088921716157087360555720302438606891293352181929889266594288273380474544647928703225388630259363515021844695116187787425784608985965360959603948643752367114155796154563;
            5'd16: xpb[77] = 1024'd13168369620996296462375435528698629734687351067080926587964321298432872363815116201818933392389659956898530711863103576842406755018779816880542783155191004686624408552163198103976781425249372166335135433799311596230131496655936260028665845525578635181629691433307818635639570050815607610872557014232532173224;
            5'd17: xpb[77] = 1024'd76024740564370935690673363951649510465454524071641326563778018912073374555208130419440152336742850858926263585083294267684589097628063722713156769610555962946383771371459006654290449860086060787386180202605388494176695140307380662762946745712542024513891498854948086315420307215955899595111436740934862676216;
            5'd18: xpb[77] = 1024'd14814415823620833520172364969785958451523269950466042411459861460736981409292005727046300066438367451510847050845991523947707599396127293990610631049589880272452459621183597866973879103405543687127027363024225545758897933737928292532249076216275964579333402862471295965094516307167558562231626641011598694877;
            5'd19: xpb[77] = 1024'd77670786766995472748470293392736839182290442955026442387273559074377483600685019944667519010791558353538579924066182214789889942005411199823224617504954838532211822440479406417287547538242232308178072131830302443705461577389372695266529976403239353911595210284111563644875253472307850546470506367713929197869;
            5'd20: xpb[77] = 1024'd16460462026245370577969294410873287168359188833851158234955401623041090454768895252273666740487074946123163389828879471053008443773474771100678478943988755858280510690203997629970976781561715207918919292249139495287664370819920325035832306906973293977037114291634773294549462563519509513590696267790665216530;
            5'd21: xpb[77] = 1024'd79316832969620009806267222833824167899126361838411558210769099236681592646161909469894885684840265848150896263049070161895190786382758676933292465399353714118039873509499806180284645216398403828969964061055216393234228014471364727770113207093936683309298921713275040974330199728659801497829575994492995719522;
            5'd22: xpb[77] = 1024'd18106508228869907635766223851960615885195107717236274058450941785345199500245784777501033414535782440735479728811767418158309288150822248210746326838387631444108561759224397392968074459717886728710811221474053444816430807901912357539415537597670623374740825720798250624004408819871460464949765894569731738183;
            5'd23: xpb[77] = 1024'd80962879172244546864064152274911496615962280721796674034264639398985701691638798995122252358888973342763212602031958109000491630760106154043360313293752589703867924578520205943281742894554575349761855990280130342762994451553356760273696437784634012707002633142438518303785145985011752449188645621272062241175;
            5'd24: xpb[77] = 1024'd19752554431494444693563153293047944602031026600621389881946481947649308545722674302728400088584489935347796067794655365263610132528169725320814174732786507029936612828244797155965172137874058249502703150698967394345197244983904390042998768288367952772444537149961727953459355076223411416308835521348798259836;
            5'd25: xpb[77] = 1024'd82608925374869083921861081715998825332798199605181789857760179561289810737115688520349619032937680837375528941014846056105792475137453631153428161188151465289695975647540605706278840572710746870553747919505044292291760888635348792777279668475331342104706344571601995633240092241363703400547715248051128762828;
            5'd26: xpb[77] = 1024'd21398600634118981751360082734135273318866945484006505705442022109953417591199563827955766762633197429960112406777543312368910976905517202430882022627185382615764663897265196918962269816030229770294595079923881343873963682065896422546581998979065282170148248579125205282914301332575362367667905148127864781489;
            5'd27: xpb[77] = 1024'd84254971577493620979658011157086154049634118488566905681255719723593919782592578045576985706986388331987845279997734003211093319514801108263496009082550340875524026716561005469275938250866918391345639848729958241820527325717340825280862899166028671502410056000765472962695038497715654351906784874830195284481;
            5'd28: xpb[77] = 1024'd23044646836743518809157012175222602035702864367391621528937562272257526636676453353183133436681904924572428745760431259474211821282864679540949870521584258201592714966285596681959367494186401291086487009148795293402730119147888455050165229669762611567851960008288682612369247588927313319026974774906931303142;
            5'd29: xpb[77] = 1024'd85901017780118158037454940598173482766470037371952021504751259885898028828069467570804352381035095826600161618980621950316394163892148585373563856976949216461352077785581405232273035929023089912137531777954872191349293762799332857784446129856726000900113767429928950292149984754067605303265854501609261806134;
            5'd30: xpb[77] = 1024'd24690693039368055866953941616309930752538783250776737352433102434561635682153342878410500110730612419184745084743319206579512665660212156651017718415983133787420766035305996444956465172342572811878378938373709242931496556229880487553748460360459940965555671437452159941824193845279264270386044401685997824795;
            5'd31: xpb[77] = 1024'd87547063982742695095251870039260811483305956255337137328246800048202137873546357096031719055083803321212477957963509897421695008269496062483631704871348092047180128854601804995270133607179261432929423707179786140878060199881324890288029360547423330297817478859092427621604931010419556254624924128388328327787;
        endcase
    end

    always_comb begin
        case(flag[26][5:0])
            6'd0: xpb[78] = 1024'd0;
            6'd1: xpb[78] = 1024'd13168369620996296462375435528698629734687351067080926587964321298432872363815116201818933392389659956898530711863103576842406755018779816880542783155191004686624408552163198103976781425249372166335135433799311596230131496655936260028665845525578635181629691433307818635639570050815607610872557014232532173224;
            6'd2: xpb[78] = 1024'd26336739241992592924750871057397259469374702134161853175928642596865744727630232403637866784779319913797061423726207153684813510037559633761085566310382009373248817104326396207953562850498744332670270867598623192460262993311872520057331691051157270363259382866615637271279140101631215221745114028465064346448;
            6'd3: xpb[78] = 1024'd39505108862988889387126306586095889204062053201242779763892963895298617091445348605456800177168979870695592135589310730527220265056339450641628349465573014059873225656489594311930344275748116499005406301397934788690394489967808780085997536576735905544889074299923455906918710152446822832617671042697596519672;
            6'd4: xpb[78] = 1024'd52673478483985185849501742114794518938749404268323706351857285193731489455260464807275733569558639827594122847452414307369627020075119267522171132620764018746497634208652792415907125700997488665340541735197246384920525986623745040114663382102314540726518765733231274542558280203262430443490228056930128692896;
            6'd5: xpb[78] = 1024'd65841848104981482311877177643493148673436755335404632939821606492164361819075581009094666961948299784492653559315517884212033775093899084402713915775955023433122042760815990519883907126246860831675677168996557981150657483279681300143329227627893175908148457166539093178197850254078038054362785071162660866120;
            6'd6: xpb[78] = 1024'd79010217725977778774252613172191778408124106402485559527785927790597234182890697210913600354337959741391184271178621461054440530112678901283256698931146028119746451312979188623860688551496232998010812602795869577380788979935617560171995073153471811089778148599846911813837420304893645665235342085395193039344;
            6'd7: xpb[78] = 1024'd92178587346974075236628048700890408142811457469566486115750249089030106546705813412732533746727619698289714983041725037896847285131458718163799482086337032806370859865142386727837469976745605164345948036595181173610920476591553820200660918679050446271407840033154730449476990355709253276107899099627725212568;
            6'd8: xpb[78] = 1024'd105346956967970371699003484229589037877498808536647412703714570387462978910520929614551467139117279655188245694904828614739254040150238535044342265241528037492995268417305584831814251401994977330681083470394492769841051973247490080229326764204629081453037531466462549085116560406524860886980456113860257385792;
            6'd9: xpb[78] = 1024'd118515326588966668161378919758287667612186159603728339291678891685895851274336045816370400531506939612086776406767932191581660795169018351924885048396719042179619676969468782935791032827244349497016218904193804366071183469903426340257992609730207716634667222899770367720756130457340468497853013128092789559016;
            6'd10: xpb[78] = 1024'd7617000525838223224955427882171864602175083545073581751511357919351828300842023108174262709238925259542157711173542333845003709346577834250267706535579005932553410952060763702137575060976515942041156729605876115936954116338465827321679885572556902549477010918961128326289172434227443091606880315699727247909;
            6'd11: xpb[78] = 1024'd20785370146834519687330863410870494336862434612154508339475679217784700664657139309993196101628585216440688423036645910687410464365357651130810489690770010619177819504223961806114356486225888108376292163405187712167085612994402087350345731098135537731106702352268946961928742485043050702479437329932259421133;
            6'd12: xpb[78] = 1024'd33953739767830816149706298939569124071549785679235434927440000516217573028472255511812129494018245173339219134899749487529817219384137468011353272845961015305802228056387159910091137911475260274711427597204499308397217109650338347379011576623714172912736393785576765597568312535858658313351994344164791594357;
            6'd13: xpb[78] = 1024'd47122109388827112612081734468267753806237136746316361515404321814650445392287371713631062886407905130237749846762853064372223974402917284891896056001152019992426636608550358014067919336724632441046563031003810904627348606306274607407677422149292808094366085218884584233207882586674265924224551358397323767581;
            6'd14: xpb[78] = 1024'd60290479009823409074457169996966383540924487813397288103368643113083317756102487915449996278797565087136280558625956641214630729421697101772438839156343024679051045160713556118044700761974004607381698464803122500857480102962210867436343267674871443275995776652192402868847452637489873535097108372629855940805;
            6'd15: xpb[78] = 1024'd73458848630819705536832605525665013275611838880478214691332964411516190119917604117268929671187225044034811270489060218057037484440476918652981622311534029365675453712876754222021482187223376773716833898602434097087611599618147127465009113200450078457625468085500221504487022688305481145969665386862388114029;
            6'd16: xpb[78] = 1024'd86627218251816001999208041054363643010299189947559141279297285709949062483732720319087863063576885000933341982352163794899444239459256735533524405466725034052299862265039952325998263612472748940051969332401745693317743096274083387493674958726028713639255159518808040140126592739121088756842222401094920287253;
            6'd17: xpb[78] = 1024'd99795587872812298461583476583062272744986541014640067867261607008381934847547836520906796455966544957831872694215267371741850994478036552414067188621916038738924270817203150429975045037722121106387104766201057289547874592930019647522340804251607348820884850952115858775766162789936696367714779415327452460477;
            6'd18: xpb[78] = 1024'd112963957493808594923958912111760902479673892081720994455225928306814807211362952722725729848356204914730403406078370948584257749496816369294609971777107043425548679369366348533951826462971493272722240200000368885778006089585955907551006649777185984002514542385423677411405732840752303978587336429559984633701;
            6'd19: xpb[78] = 1024'd2065631430680149987535420235645099469662816023066236915058394540270784237868930014529592026088190562185784710483981090847600663674375851619992629915967007178482413351958329300298368696703659717747178025412440635643776736020995394614693925619535169917324330404614438016938774817639278572341203617166922322594;
            6'd20: xpb[78] = 1024'd15234001051676446449910855764343729204350167090147163503022715838703656601684046216348525418477850519084315422347084667690007418693155668500535413071158011865106821904121527404275150121953031884082313459211752231873908232676931654643359771145113805098954021837922256652578344868454886183213760631399454495818;
            6'd21: xpb[78] = 1024'd28402370672672742912286291293042358939037518157228090090987037137136528965499162418167458810867510475982846134210188244532414173711935485381078196226349016551731230456284725508251931547202404050417448893011063828104039729332867914672025616670692440280583713271230075288217914919270493794086317645631986669042;
            6'd22: xpb[78] = 1024'd41570740293669039374661726821740988673724869224309016678951358435569401329314278619986392203257170432881376846073291821374820928730715302261620979381540021238355639008447923612228712972451776216752584326810375424334171225988804174700691462196271075462213404704537893923857484970086101404958874659864518842266;
            6'd23: xpb[78] = 1024'd54739109914665335837037162350439618408412220291389943266915679734002273693129394821805325595646830389779907557936395398217227683749495119142163762536731025924980047560611121716205494397701148383087719760609687020564302722644740434729357307721849710643843096137845712559497055020901709015831431674097051015490;
            6'd24: xpb[78] = 1024'd67907479535661632299412597879138248143099571358470869854880001032435146056944511023624258988036490346678438269799498975059634438768274936022706545691922030611604456112774319820182275822950520549422855194408998616794434219300676694758023153247428345825472787571153531195136625071717316626703988688329583188714;
            6'd25: xpb[78] = 1024'd81075849156657928761788033407836877877786922425551796442844322330868018420759627225443192380426150303576968981662602551902041193787054752903249328847113035298228864664937517924159057248199892715757990628208310213024565715956612954786688998773006981007102479004461349830776195122532924237576545702562115361938;
            6'd26: xpb[78] = 1024'd94244218777654225224163468936535507612474273492632723030808643629300890784574743427262125772815810260475499693525706128744447948805834569783792112002304039984853273217100716028135838673449264882093126062007621809254697212612549214815354844298585616188732170437769168466415765173348531848449102716794647535162;
            6'd27: xpb[78] = 1024'd107412588398650521686538904465234137347161624559713649618772964927733763148389859629081059165205470217374030405388809705586854703824614386664334895157495044671477681769263914132112620098698637048428261495806933405484828709268485474844020689824164251370361861871076987102055335224164139459321659731027179708386;
            6'd28: xpb[78] = 1024'd120580958019646818148914339993932767081848975626794576206737286226166635512204975830899992557595130174272561117251913282429261458843394203544877678312686049358102090321427112236089401523948009214763396929606245001714960205924421734872686535349742886551991553304384805737694905274979747070194216745259711881610;
            6'd29: xpb[78] = 1024'd9682631956518373212490848117816964071837899568139818666569752459622612538710953122703854735327115821727942421657523424692604373020953685870260336451546013111035824304019093002435943757680175659788334755018316751580730852359461221936373811192092072466801341323575566343227947251866721663948083932866649570503;
            6'd30: xpb[78] = 1024'd22851001577514669674866283646515593806525250635220745254534073758055484902526069324522788127716775778626473133520627001535011128039733502750803119606737017797660232856182291106412725182929547826123470188817628347810862349015397481965039656717670707648431032756883384978867517302682329274820640947099181743727;
            6'd31: xpb[78] = 1024'd36019371198510966137241719175214223541212601702301671842498395056488357266341185526341721520106435735525003845383730578377417883058513319631345902761928022484284641408345489210389506608178919992458605622616939944040993845671333741993705502243249342830060724190191203614507087353497936885693197961331713916951;
            6'd32: xpb[78] = 1024'd49187740819507262599617154703912853275899952769382598430462716354921229630156301728160654912496095692423534557246834155219824638077293136511888685917119027170909049960508687314366288033428292158793741056416251540271125342327270002022371347768827978011690415623499022250146657404313544496565754975564246090175;
            6'd33: xpb[78] = 1024'd62356110440503559061992590232611483010587303836463525018427037653354101993971417929979588304885755649322065269109937732062231393096072953392431469072310031857533458512671885418343069458677664325128876490215563136501256838983206262051037193294406613193320107056806840885786227455129152107438311989796778263399;
            6'd34: xpb[78] = 1024'd75524480061499855524368025761310112745274654903544451606391358951786974357786534131798521697275415606220595980973041308904638148114852770272974252227501036544157867064835083522319850883927036491464011924014874732731388335639142522079703038819985248374949798490114659521425797505944759718310869004029310436623;
            6'd35: xpb[78] = 1024'd88692849682496151986743461290008742479962005970625378194355680250219846721601650333617455089665075563119126692836144885747044903133632587153517035382692041230782275616998281626296632309176408657799147357814186328961519832295078782108368884345563883556579489923422478157065367556760367329183426018261842609847;
            6'd36: xpb[78] = 1024'd101861219303492448449118896818707372214649357037706304782320001548652719085416766535436388482054735520017657404699248462589451658152412404034059818537883045917406684169161479730273413734425780824134282791613497925191651328951015042137034729871142518738209181356730296792704937607575974940055983032494374783071;
            6'd37: xpb[78] = 1024'd115029588924488744911494332347406001949336708104787231370284322847085591449231882737255321874444395476916188116562352039431858413171192220914602601693074050604031092721324677834250195159675152990469418225412809521421782825606951302165700575396721153919838872790038115428344507658391582550928540046726906956295;
            6'd38: xpb[78] = 1024'd4131262861360299975070840471290198939325632046132473830116789080541568475737860029059184052176381124371569420967962181695201327348751703239985259831934014356964826703916658600596737393407319435494356050824881271287553472041990789229387851239070339834648660809228876033877549635278557144682407234333844645188;
            6'd39: xpb[78] = 1024'd17299632482356596437446275999988828674012983113213400418081110378974440839552976230878117444566041081270100132831065758537608082367531520120528042987125019043589235256079856704573518818656691601829491484624192867517684968697927049258053696764648975016278352242536694669517119686094164755554964248566376818412;
            6'd40: xpb[78] = 1024'd30468002103352892899821711528687458408700334180294327006045431677407313203368092432697050836955701038168630844694169335380014837386311337001070826142316023730213643808243054808550300243906063768164626918423504463747816465353863309286719542290227610197908043675844513305156689736909772366427521262798908991636;
            6'd41: xpb[78] = 1024'd43636371724349189362197147057386088143387685247375253594009752975840185567183208634515984229345360995067161556557272912222421592405091153881613609297507028416838052360406252912527081669155435934499762352222816059977947962009799569315385387815806245379537735109152331940796259787725379977300078277031441164860;
            6'd42: xpb[78] = 1024'd56804741345345485824572582586084717878075036314456180181974074274273057930998324836334917621735020951965692268420376489064828347423870970762156392452698033103462460912569451016503863094404808100834897786022127656208079458665735829344051233341384880561167426542460150576435829838540987588172635291263973338084;
            6'd43: xpb[78] = 1024'd69973110966341782286948018114783347612762387381537106769938395572705930294813441038153851014124680908864222980283480065907235102442650787642699175607889037790086869464732649120480644519654180267170033219821439252438210955321672089372717078866963515742797117975767969212075399889356595199045192305496505511308;
            6'd44: xpb[78] = 1024'd83141480587338078749323453643481977347449738448618033357902716871138802658628557239972784406514340865762753692146583642749641857461430604523241958763080042476711278016895847224457425944903552433505168653620750848668342451977608349401382924392542150924426809409075787847714969940172202809917749319729037684532;
            6'd45: xpb[78] = 1024'd96309850208334375211698889172180607082137089515698959945867038169571675022443673441791717798904000822661284404009687219592048612480210421403784741918271047163335686569059045328434207370152924599840304087420062444898473948633544609430048769918120786106056500842383606483354539990987810420790306333961569857756;
            6'd46: xpb[78] = 1024'd109478219829330671674074324700879236816824440582779886533831359468004547386258789643610651191293660779559815115872790796434455367498990238284327525073462051849960095121222243432410988795402296766175439521219374041128605445289480869458714615443699421287686192275691425118994110041803418031662863348194102030980;
            6'd47: xpb[78] = 1024'd122646589450326968136449760229577866551511791649860813121795680766437419750073905845429584583683320736458345827735894373276862122517770055164870308228653056536584503673385441536387770220651668932510574955018685637358736941945417129487380460969278056469315883708999243754633680092619025642535420362426634204204;
            6'd48: xpb[78] = 1024'd11748263387198523200026268353462063541500715591206055581628146999893396776579883137233446761415306383913727132141504515540205036695329537490252966367513020289518237655977422302734312454383835377535512780430757387224507588380456616551067736811627242384125671728190004360166722069506000236289287550033571893097;
            6'd49: xpb[78] = 1024'd24916633008194819662401703882160693276188066658286982169592468298326269140394999339052380153804966340812257844004608092382611791714109354370795749522704024976142646208140620406711093879633207543870648214230068983454639085036392876579733582337205877565755363161497822995806292120321607847161844564266104066321;
            6'd50: xpb[78] = 1024'd38085002629191116124777139410859323010875417725367908757556789596759141504210115540871313546194626297710788555867711669225018546732889171251338532677895029662767054760303818510687875304882579710205783648029380579684770581692329136608399427862784512747385054594805641631445862171137215458034401578498636239545;
            6'd51: xpb[78] = 1024'd51253372250187412587152574939557952745562768792448835345521110895192013868025231742690246938584286254609319267730815246067425301751668988131881315833086034349391463312467016614664656730131951876540919081828692175914902078348265396637065273388363147929014746028113460267085432221952823068906958592731168412769;
            6'd52: xpb[78] = 1024'd64421741871183709049528010468256582480250119859529761933485432193624886231840347944509180330973946211507849979593918822909832056770448805012424098988277039036015871864630214718641438155381324042876054515628003772145033575004201656665731118913941783110644437461421278902725002272768430679779515606963700585993;
            6'd53: xpb[78] = 1024'd77590111492180005511903445996955212214937470926610688521449753492057758595655464146328113723363606168406380691457022399752238811789228621892966882143468043722640280416793412822618219580630696209211189949427315368375165071660137916694396964439520418292274128894729097538364572323584038290652072621196232759217;
            6'd54: xpb[78] = 1024'd90758481113176301974278881525653841949624821993691615109414074790490630959470580348147047115753266125304911403320125976594645566808008438773509665298659048409264688968956610926595001005880068375546325383226626964605296568316074176723062809965099053473903820328036916174004142374399645901524629635428764932441;
            6'd55: xpb[78] = 1024'd103926850734172598436654317054352471684312173060772541697378396088923503323285696549965980508142926082203442115183229553437052321826788255654052448453850053095889097521119809030571782431129440541881460817025938560835428064972010436751728655490677688655533511761344734809643712425215253512397186649661297105665;
            6'd56: xpb[78] = 1024'd117095220355168894899029752583051101418999524127853468285342717387356375687100812751784913900532586039101972827046333130279459076845568072534595231609041057782513506073283007134548563856378812708216596250825250157065559561627946696780394501016256323837163203194652553445283282476030861123269743663893829278889;
            6'd57: xpb[78] = 1024'd6196894292040449962606260706935298408988448069198710745175183620812352713606790043588776078264571686557354131451943272542801991023127554859977889747901021535447240055874987900895106090110979153241534076237321906931330208062986183844081776858605509751972991213843314050816324452917835717023610851500766967782;
            6'd58: xpb[78] = 1024'd19365263913036746424981696235633928143675799136279637333139504919245225077421906245407709470654231643455884843315046849385208746041907371740520672903092026222071648608038186004871887515360351319576669510036633503161461704718922443872747622384184144933602682647151132686455894503733443327896167865733299141006;
            6'd59: xpb[78] = 1024'd32533633534033042887357131764332557878363150203360563921103826217678097441237022447226642863043891600354415555178150426227615501060687188621063456058283030908696057160201384108848668940609723485911804943835945099391593201374858703901413467909762780115232374080458951322095464554549050938768724879965831314230;
            6'd60: xpb[78] = 1024'd45702003155029339349732567293031187613050501270441490509068147516110969805052138649045576255433551557252946267041254003070022256079467005501606239213474035595320465712364582212825450365859095652246940377635256695621724698030794963930079313435341415296862065513766769957735034605364658549641281894198363487454;
            6'd61: xpb[78] = 1024'd58870372776025635812108002821729817347737852337522417097032468814543842168867254850864509647823211514151476978904357579912429011098246822382149022368665040281944874264527780316802231791108467818582075811434568291851856194686731223958745158960920050478491756947074588593374604656180266160513838908430895660678;
            6'd62: xpb[78] = 1024'd72038742397021932274483438350428447082425203404603343684996790112976714532682371052683443040212871471050007690767461156754835766117026639262691805523856044968569282816690978420779013216357839984917211245233879888081987691342667483987411004486498685660121448380382407229014174706995873771386395922663427833902;
            6'd63: xpb[78] = 1024'd85207112018018228736858873879127076817112554471684270272961111411409586896497487254502376432602531427948538402630564733597242521135806456143234588679047049655193691368854176524755794641607212151252346679033191484312119187998603744016076850012077320841751139813690225864653744757811481382258952936895960007126;
        endcase
    end

    always_comb begin
        case(flag[26][11:6])
            6'd0: xpb[79] = 1024'd0;
            6'd1: xpb[79] = 1024'd98375481639014525199234309407825706551799905538765196860925432709842459260312603456321309824992191384847069114493668310439649276154586273023777371834238054341818099921017374628732576066856584317587482112832503080542250684654540004044742695537655956023380831246998044500293314808627088993131509951128492180350;
            6'd2: xpb[79] = 1024'd72684267593904308999669691410836980358901383951794709593719010354708023183316068002627548435326708460250988821529843186300234711467952211492394618652145067749945525272463531919834912942195962913864766617277766314720140519088183235124506821392082462779941759079879030970480101543325544969144330075631389876369;
            6'd3: xpb[79] = 1024'd46993053548794092800105073413848254166002862364824222326512587999573587106319532548933787045661225535654908528566018062160820146781318149961011865470052081158072950623909689210937249817535341510142051121723029548898030353521826466204270947246508969536502686912760017440666888278024000945157150200134287572388;
            6'd4: xpb[79] = 1024'd21301839503683876600540455416859527973104340777853735059306165644439151029322997095240025655995742611058828235602192938021405582094684088429629112287959094566200375975355846502039586692874720106419335626168292783075920187955469697284035073100935476293063614745641003910853675012722456921169970324637185268407;
            6'd5: xpb[79] = 1024'd119677321142698401799774764824685234524904246316618931920231598354281610289635600551561335480987933995905897350095861248461054858249270361453406484122197148908018475896373221130772162759731304424006817739000795863618170872610009701328777768638591432316444445992639048411146989821349545914301480275765677448757;
            6'd6: xpb[79] = 1024'd93986107097588185600210146827696508332005724729648444653025175999147174212639065097867574091322451071309817057132036124321640293562636299922023730940104162316145901247819378421874499635070683020284102243446059097796060707043652932408541894493017939073005373825520034881333776556048001890314300400268575144776;
            6'd7: xpb[79] = 1024'd68294893052477969400645528830707782139107203142677957385818753644012738135642529644173812701656968146713736764168211000182225728876002238390640977758011175724273326599265535712976836510410061616561386747891322331973950541477296163488306020347444445829566301658401021351520563290746457866327120524771472840795;
            6'd8: xpb[79] = 1024'd42603679007367753201080910833719055946208681555707470118612331288878302058645994190480051311991485222117656471204385876042811164189368176859258224575918189132400751950711693004079173385749440212838671252336585566151840375910939394568070146201870952586127229491282007821707350025444913842339940649274370536814;
            6'd9: xpb[79] = 1024'd16912464962257537001516292836730329753310159968736982851405908933743865981649458736786289922326002297521576178240560751903396599502734115327875471393825202540528177302157850295181510261088818809115955756781848800329730210344582625647834272056297459342688157324162994291894136760143369818352760773777268232833;
            6'd10: xpb[79] = 1024'd115287946601272062200750602244556036305110065507502179712331341643586325241962062193107599747318193682368645292734229062343045875657320388351652843228063256882346277223175224923914086327945403126703437869614351880871980894999122629692576967593953415366068988571161038792187451568770458811484270724905760413183;
            6'd11: xpb[79] = 1024'd89596732556161846001185984247567310112211543920531692445124919288451889164965526739413838357652710757772564999770403938203631310970686326820270090045970270290473702574621382215016423203284781722980722374059615115049870729432765860772341093448379922122629916404042025262374238303468914787497090849408658109202;
            6'd12: xpb[79] = 1024'd63905518511051629801621366250578583919313022333561205177918496933317453087968991285720076967987227833176484706806578814064216746284052265288887336863877283698601127926067539506118760078624160319258006878504878349227760563866409091852105219302806428879190844236923011732561025038167370763509910973911555805221;
            6'd13: xpb[79] = 1024'd38214304465941413602056748253589857726414500746590717910712074578183017010972455832026315578321744908580404413842753689924802181597418203757504583681784297106728553277513696797221096953963538915535291382950141583405650398300052322931869345157232935635751772069803998202747811772865826739522731098414453501240;
            6'd14: xpb[79] = 1024'd12523090420831197402492130256601131533515979159620230643505652223048580933975920378332554188656261983984324120878928565785387616910784142226121830499691310514855978628959854088323433829302917511812575887395404817583540232733695554011633471011659442392312699902684984672934598507564282715535551222917351197259;
            6'd15: xpb[79] = 1024'd110898572059845722601726439664426838085315884698385427504431084932891040194288523834653864013648453368831393235372596876225036893065370415249899202333929364856674078549977228717056009896159501829400058000227907898125790917388235558056376166549315398415693531149683029173227913316191371708667061174045843377609;
            6'd16: xpb[79] = 1024'd85207358014735506402161821667438111892417363111414940237224662577756604117291988380960102623982970444235312942408771752085622328378736353718516449151836378264801503901423386008158346771498880425677342504673171132303680751821878789136140292403741905172254458982564015643414700050889827684679881298548741073628;
            6'd17: xpb[79] = 1024'd59516143969625290202597203670449385699518841524444452970018240222622168040295452927266341234317487519639232649444946627946207763692102292187133695969743391672928929252869543299260683646838259021954627009118434366481570586255522020215904418258168411928815386815445002113601486785588283660692701423051638769647;
            6'd18: xpb[79] = 1024'd33824929924515074003032585673460659506620319937473965702811817867487731963298917473572579844652004595043152356481121503806793199005468230655750942787650405081056354604315700590363020522177637618231911513563697600659460420689165251295668544112594918685376314648325988583788273520286739636705521547554536465666;
            6'd19: xpb[79] = 1024'd8133715879404857803467967676471933313721798350503478435605395512353295886302382019878818454986521670447072063517296379667378634318834169124368189605557418489183779955761857881465357397517016214509196018008960834837350255122808482375432669967021425441937242481206975053975060254985195612718341672057434161685;
            6'd20: xpb[79] = 1024'd106509197518419383002702277084297639865521703889268675296530828222195755146614985476200128279978713055294141178010964690107027910473420442148145561439795472831001879876779232510197933464373600532096678130841463915379600939777348486420175365504677381465318073728205019554268375063612284605849851623185926342035;
            6'd21: xpb[79] = 1024'd80817983473309166803137659087308913672623182302298188029324405867061319069618450022506366890313230130698060885047139565967613345786786380616762808257702486239129305228225389801300270339712979128373962635286727149557490774210991717499939491359103888221879001561086006024455161798310740581862671747688824038054;
            6'd22: xpb[79] = 1024'd55126769428198950603573041090320187479724660715327700762117983511926882992621914568812605500647747206101980592083314441828198781100152319085380055075609499647256730579671547092402607215052357724651247139731990383735380608644634948579703617213530394978439929393966992494641948533009196557875491872191721734073;
            6'd23: xpb[79] = 1024'd29435555383088734404008423093331461286826139128357213494911561156792446915625379115118844110982264281505900299119489317688784216413518257553997301893516513055384155931117704383504944090391736320928531644177253617913270443078278179659467743067956901735000857226847978964828735267707652533888311996694619430092;
            6'd24: xpb[79] = 1024'd3744341337978518204443805096342735093927617541386726227705138801658010838628843661425082721316781356909820006155664193549369651726884196022614548711423526463511581282563861674607280965731114917205816148622516852091160277511921410739231868922383408491561785059728965435015522002406108509901132121197517126111;
            6'd25: xpb[79] = 1024'd102119822976993043403678114504168441645727523080151923088630571511500470098941447117746392546308972741756889120649332503989018927881470469046391920545661580805329681203581236303339857032587699234793298261455019932633410962166461414783974564460039364514942616306727009935308836811033197503032642072326009306461;
            6'd26: xpb[79] = 1024'd76428608931882827204113496507179715452829001493181435821424149156366034021944911664052631156643489817160808827685507379849604363194836407515009167363568594213457106555027393594442193907927077831070582765900283166811300796600104645863738690314465871271503544139607996405495623545731653479045462196828907002480;
            6'd27: xpb[79] = 1024'd50737394886772611004548878510190989259930479906210948554217726801231597944948376210358869766978006892564728534721682255710189798508202345983626414181475607621584531906473550885544530783266456427347867270345546400989190631033747876943502816168892378028064471972488982875682410280430109455058282321331804698499;
            6'd28: xpb[79] = 1024'd25046180841662394804984260513202263067031958319240461287011304446097161867951840756665108377312523967968648241757857131570775233821568284452243660999382621029711957257919708176646867658605835023625151774790809635167080465467391108023266942023318884784625399805369969345869197015128565431071102445834702394518;
            6'd29: xpb[79] = 1024'd123421662480676920004218569921027969618831863858005658147936737155939621128264444212986418202304715352815717356251525442010424509976154557476021032833620675371530057178937082805379443725462419341212633887623312715709331150121931112068009637560974840808006231052368013846162511823755654424202612396963194574868;
            6'd30: xpb[79] = 1024'd97730448435566703804653951924039243425933342271035170880730314800805185051267908759292656812639232428219637063287700317871009945289520495944638279651527688779657482530383240096481780600801797937489918392068575949887220984555574343147773763415401347564567158885249000316349298558454110400215432521466092270887;
            6'd31: xpb[79] = 1024'd72039234390456487605089333927050517233034820684064683613523892445670748974271373305598895422973749503623556770323875193731595380602886434413255526469434702187784907881829397387584117476141176533767202896513839184065110818989217574227537889269827854321128086718129986786536085293152566376228252645968989966906;
            6'd32: xpb[79] = 1024'd46348020345346271405524715930061791040136299097094196346317470090536312897274837851905134033308266579027476477360050069592180815916252372881872773287341715595912333233275554678686454351480555130044487400959102418243000653422860805307302015124254361077689014551010973256722872027851022352241072770471887662925;
            6'd33: xpb[79] = 1024'd20656806300236055205960097933073064847237777510123709079111047735401876820278302398211372643642783654431396184396224945452766251229618311350490020105248729004039758584721711969788791226819933726321771905404365652420890487856504036387066140978680867834249942383891959726909658762549478328253892894974785358944;
            6'd34: xpb[79] = 1024'd119032287939250580405194407340898771399037683048888905940036480445244336080590905854532682468634975039278465298889893255892415527384204584374267391939486783345857858505739086598521367293676518043909254018236868732963141172511044040431808836516336823857630773630890004227202973571176567321385402846103277539294;
            6'd35: xpb[79] = 1024'd93341073894140364205629789343910045206139161461918418672830058090109900003594370400838921078969492114682385005926068131753000962697570522842884638757393796753985283857185243889623704169015896640186538522682131967141031006944687271511572962370763330614191701463770990697389760305875023297398222970606175235313;
            6'd36: xpb[79] = 1024'd67649859849030148006065171346921319013240639874947931405623635734975463926597834947145159689304009190086304712962243007613586398010936461311501885575300810162112709208631401180726041044355275236463823027127395201318920841378330502591337088225189837370752629296651977167576547040573479273411043095109072931332;
            6'd37: xpb[79] = 1024'd41958645803919931806500553349932592820342118287977444138417213379841027849601299493451398299638526265490224419998417883474171833324302399780119132393207823570240134560077558471828377919694653832741107531572658435496810675811973733671101214079616344127313557129532963637763333775271935249423863219611970627351;
            6'd38: xpb[79] = 1024'd16267431758809715606935935352943866627443596701006956871210791024706591772604764039757636909973043340894144127034592759334757268637668338248736379211114836978367559911523715762930714795034032429018392036017921669674700510245616964750865339934042850883874484962413950107950120509970391225436683344114868323370;
            6'd39: xpb[79] = 1024'd114642913397824240806170244760769573179243502239772153732136223734549051032917367496078946734965234725741213241528261069774406544792254611272513751045352891320185659832541090391663290861890616746605874148850424750216951194900156968795608035471698806907255316209411994608243435318597480218568193295243360503720;
            6'd40: xpb[79] = 1024'd88951699352714024606605626763780846986344980652801666464929801379414614955920832042385185345299751801145132948564435945634991980105620549741130997863259904728313085183987247682765627737229995342883158653295687984394841029333800199875372161326125313663816244042292981078430222053295936194581013419746258199739;
            6'd41: xpb[79] = 1024'd63260485307603808407041008766792120793446459065831179197723379024280178878924296588691423955634268876549052655600610821495577415418986488209748244681166918136440510535433404973867964612569373939160443157740951218572730863767443430955136287180551820420377171875173967548617008787994392170593833544249155895758;
            6'd42: xpb[79] = 1024'd37569271262493592207476390769803394600547937478860691930516956669145742801927761134997662565968785951952972362636785697356162850732352426678365491499073931544567935886879562264970301487908752535437727662186214452750620698201086662034900413034978327176938099708054954018803795522692848146606653668752053591777;
            6'd43: xpb[79] = 1024'd11878057217383376007911772772814668407649415891890204663310534314011306724931225681303901176303303027356892069672960573216748286045718365146982738316980944952695361238325719556072638363248131131715012166631477686928510532634729893114664538889404833933499027540935940488990582257391304122619473793254951287796;
            6'd44: xpb[79] = 1024'd110253538856397901207146082180640374959449321430655401524235967023853765985243829137625211001295494412203961184166628883656397562200304638170760110151218999294513461159343094184805214430104715449302494279463980767470761217289269897159407234427060789956879858787933984989283897066018393115750983744383443468146;
            6'd45: xpb[79] = 1024'd84562324811287685007581464183651648766550799843684914257029544668719329908247293683931449611630011487607880891202803759516982997513670576639377356969126012702640886510789251475907551305444094045579778783909244001648651051722913128239171360281487296713440786620814971459470683800716849091763803868886341164165;
            6'd46: xpb[79] = 1024'd58871110766177468808016846186662922573652278256714426989823122313584893831250758230237688221964528563011800598238978635377568432827036515107994603787033026110768311862235408767009888180783472641857063288354507235826540886156556359318935486135913803470001714453695957929657470535415305067776623993389238860184;
            6'd47: xpb[79] = 1024'd33179896721067252608452228189674196380753756669743939722616699958450457754254222776543926832299045638415720305275153511238153868140402453576611850604940039518895737213681566058112225056122851238134347792799770470004430720590199590398699611990340310226562642286576944399844257270113761043789444117892136556203;
            6'd48: xpb[79] = 1024'd7488682675957036408887610192685470187855235082773452455410277603316021677257687322850165442633562713819640012311328387098739303453768392045229097422847052927023162565127723349214561931462229834411632297245033704182320555023842821478463737844766816983123570119457930870031044004812217019802264242395034252222;
            6'd49: xpb[79] = 1024'd105864164314971561608121919600511176739655140621538649316335710313158480937570290779171475267625754098666709126804996697538388579608354665069006469257085107268841262486145097977947137998318814151999114410077536784724571239678382825523206433382422773006504401366455975370324358813439306012933774193523526432572;
            6'd50: xpb[79] = 1024'd80172950269861345408557301603522450546756619034568162049129287958024044860573755325477713877960271174070628833841171573398974014921720603537623716074992120676968687837591255269049474873658192748276398914522800018902461074112026056602970559236849279763065329199336961840511145548137761988946594318026424128591;
            6'd51: xpb[79] = 1024'd54481736224751129208992683606533724353858097447597674781922865602889608783577219871783952488294788249474548540877346449259559450235086542006240962892899134085096113189037412560151811748997571344553683418968063253080350908545669287682734685091275786519626257032217948310697932282836217964959414442529321824610;
            6'd52: xpb[79] = 1024'd28790522179640913009428065609544998160959575860627187514716443247755172706580684418090191098629305324878468247913521325120144885548452480474858209710806147493223538540483569851254148624336949940830967923413326487258240742979312518762498810945702293276187184865098934780884719017534673940972234567032219520629;
            6'd53: xpb[79] = 1024'd3099308134530696809863447612556271968061054273656700247510020892620736629584148964396429708963822400282387954949696200980730320861818418943475456528713160901350963891929727142356485499676328537108252427858589721436130577412955749842262936800128800032748112697979921251071505752233129916985054691535117216648;
            6'd54: xpb[79] = 1024'd101474789773545222009097757020381978519860959812421897108435453602463195889896752420717739533956013785129457069443364511420379597016404691967252828362951215243169063812947101771089061566532912854695734540691092801978381262067495753887005632337784756056128943944977965751364820560860218910116564642663609396998;
            6'd55: xpb[79] = 1024'd75783575728435005809533139023393252326962438225451409841229031247328759812900216967023978144290530860533376776479539387280965032329770630435870075180858228651296489164393259062191398441872291450973019045136356036156271096501138984966769758192211262812689871777858952221551607295558674886129384767166507093017;
            6'd56: xpb[79] = 1024'd50092361683324789609968521026404526134063916638480922574022608892194323735903681513330216754625047935937296483515714263141550467643136568904487321998765242059423914515839416353293735317211670047250303549581619270334160930934782216046533884046637769569250799610739938691738394030257130862142204891669404789036;
            6'd57: xpb[79] = 1024'd24401147638214573410403903029415799941165395051510435306816186537059887658907146059636455364959565011341216190551889139002135902956502507373104568816672255467551339867285573644396072192551048643527588054026882504512050765368425447126298009901064276325811727443620925161925180764955586838155025016172302485055;
            6'd58: xpb[79] = 1024'd122776629277229098609638212437241506492965300590275632167741619246902346919219749515957765189951756396188285305045557449441785179111088780396881940650910309809369439788302948273128648259407632961115070166859385585054301450022965451171040705438720232349192558690618969662218495573582675831286534967300794665405;
            6'd59: xpb[79] = 1024'd97085415232118882410073594440252780300066779003305144900535196891767910842223214062264003800286273471592205012081732325302370614424454718865499187468817323217496865139749105564230985134747011557392354671304648819232191284456608682250804831293146739105753486523499956132405282308281131807299355091803692361424;
            6'd60: xpb[79] = 1024'd71394201187008666210508976443264054107168257416334657633328774536633474765226678608570242410620790546996124719117907201162956049737820657334116434286724336625624290491195262855333322010086390153669639175749912053410081118890251913330568957147573245862314414356380942602592069042979587783312175216306590057443;
            6'd61: xpb[79] = 1024'd45702987141898450010944358446275327914269735829364170366122352181499038688230143154876481020955307622400044426154082077023541485051186595802733681104631350033751715842641420146435658885425768749946923680195175287587970953323895144410333083001999752618875342189261929072778855777678043759324995340809487753462;
            6'd62: xpb[79] = 1024'd20011773096788233811379740449286601721371214242393683098915929826364602611233607701182719631289824697803964133190256952884126920364552534271350927922538363441879141194087577437537995760765147346224208184640438521765860787757538375490097208856426259375436270022142915542965642512376499735337815465312385449481;
            6'd63: xpb[79] = 1024'd118387254735802759010614049857112308273171119781158879959841362536207061871546211157504029456282016082651033247683925263323776196519138807295128299756776417783697241115104952066270571827621731663811690297472941602308111472412078379534839904394082215398817101269140960043258957321003588728469325416440877629831;
        endcase
    end

    always_comb begin
        case(flag[26][16:12])
            5'd0: xpb[80] = 1024'd0;
            5'd1: xpb[80] = 1024'd92696040690692542811049431860123582080272598194188392692634940181072625794549675703810268066616533158054952954720100139184361631832504745763745546574683431191824666466551109357372908702961110260088974801918204836486001306845721610614604030248508722155378029102021946513445744055702044704482145540943775325850;
            5'd2: xpb[80] = 1024'd61325385697260344223299936315432731415846769262641101257138025297168356251790212497605464918575392006666756501982706843789659422823789156972330968133035821449958658363531001377115578214405014798867751995449169826607641763470546448264229490813787995043936154789926834996784960037475456391845601255261956167369;
            5'd3: xpb[80] = 1024'd29954730703828145635550440770741880751420940331093809821641110413264086709030749291400661770534250855278560049245313548394957213815073568180916389691388211708092650260510893396858247725848919337646529188980134816729282220095371285913854951379067267932494280477831723480124176019248868079209056969580137008888;
            5'd4: xpb[80] = 1024'd122650771394520688446599872630865462831693538525282202514276050594336712503580424995210929837150784013333513003965413687579318845647578313944661936266071642899917316727062002754231156428810029597735503990898339653215283526941092896528458981627575990087872309579853669993569920074950912783691202510523912334738;
            5'd5: xpb[80] = 1024'd91280116401088489858850377086174612167267709593734911078779135710432442960820961789006126689109642861945316551228020392184616636638862725153247357824424033158051308624041894773973825940253934136514281184429304643336923983565917734178084442192855262976430435267758558476909136056724324471054658224842093176257;
            5'd6: xpb[80] = 1024'd59909461407656291271100881541483761502841880662187619643282220826528173418061498582801323541068501710557120098490627096789914427630147136361832779382776423416185300521021786793716495451697838675293058377960269633458564440190742571827709902758134535864988560955663446960248352038497736158418113939160274017776;
            5'd7: xpb[80] = 1024'd28538806414224092683351385996792910838416051730640328207785305942623903875302035376596520393027360559168923645753233801395212218621431547570418200941128813674319292418001678813459164963141743214071835571491234623580204896815567409477335363323413808753546686643568335443587568020271147845781569653478454859295;
            5'd8: xpb[80] = 1024'd121234847104916635494400817856916492918688649924828720900420246123696529669851711080406788459643893717223876600473333940579573850453936293334163747515812244866143958884552788170832073666102853474160810373409439460066206203661289020091939393571922530908924715745590281957033312075973192550263715194422230185145;
            5'd9: xpb[80] = 1024'd89864192111484436906651322312225642254262820993281429464923331239792260127092247874201985311602752565835680147735940645184871641445220704542749169074164635124277950781532680190574743177546758012939587566940404450187846660286113857741564854137201803797482841433495170440372528057746604237627170908740411026664;
            5'd10: xpb[80] = 1024'd58493537118052238318901826767534791589836992061734138029426416355887990584332784667997182163561611414447483694998547349790169432436505115751334590632517025382411942678512572210317412688990662551718364760471369440309487116910938695391190314702481076686040967121400058923711744039520015924990626623058591868183;
            5'd11: xpb[80] = 1024'd27122882124620039731152331222843940925411163130186846593929501471983721041573321461792379015520470263059287242261154054395467223427789526959920012190869415640545934575492464230060082200434567090497141954002334430431127573535763533040815775267760349574599092809304947407050960021293427612354082337376772709702;
            5'd12: xpb[80] = 1024'd119818922815312582542201763082967523005683761324375239286564441653056346836122997165602647082137003421114240196981254193579828855260294272723665558765552846832370601042043573587432990903395677350586116755920539266917128880381485143655419805516269071729977121911326893920496704076995472316836227878320548035552;
            5'd13: xpb[80] = 1024'd88448267821880383954452267538276672341257932392827947851067526769152077293363533959397843934095862269726043744243860898185126646251578683932250980323905237090504592939023465607175660414839581889364893949451504257038769337006309981305045266081548344618535247599231782403835920058768884004199683592638728877071;
            5'd14: xpb[80] = 1024'd57077612828448185366702771993585821676832103461280656415570611885247807750604070753193040786054721118337847291506467602790424437242863095140836401882257627348638584836003357626918329926283486428143671142982469247160409793631134818954670726646827617507093373287136670887175136040542295691563139306956909718590;
            5'd15: xpb[80] = 1024'd25706957835015986778953276448894971012406274529733364980073697001343538207844607546988237638013579966949650838769074307395722228234147506349421823440610017606772576732983249646660999437727390966922448336513434237282050250255959656604296187212106890395651498975041559370514352022315707378926595021275090560109;
            5'd16: xpb[80] = 1024'd118402998525708529590002708309018553092678872723921757672708637182416164002394283250798505704630113125004603793489174446580083860066652252113167370015293448798597243199534359004033908140688501227011423138431639073768051557101681267218900217460615612551029528077063505883960096078017752083408740562218865885959;
            5'd17: xpb[80] = 1024'd87032343532276331002253212764327702428253043792374466237211722298511894459634820044593702556588971973616407340751781151185381651057936663321752791573645839056731235096514251023776577652132405765790200331962604063889692013726506104868525678025894885439587653764968394367299312059791163770772196276537046727478;
            5'd18: xpb[80] = 1024'd55661688538844132414503717219636851763827214860827174801714807414607624916875356838388899408547830822228210888014387855790679442049221074530338213131998229314865226993494143043519247163576310304568977525493569054011332470351330942518151138591174158328145779452873282850638528041564575458135651990855227568997;
            5'd19: xpb[80] = 1024'd24291033545411933826754221674946001099401385929279883366217892530703355374115893632184096260506689670840014435276994560395977233040505485738923634690350619572999218890474035063261916675020214843347754719024534044132972926976155780167776599156453431216703905140778171333977744023337987145499107705173408410516;
            5'd20: xpb[80] = 1024'd116987074236104476637803653535069583179673984123468276058852832711775981168665569335994364327123222828894967389997094699580338864873010231502669181265034050764823885357025144420634825377981325103436729520942738880618974233821877390782380629404962153372081934242800117847423488079040031849981253246117183736366;
            5'd21: xpb[80] = 1024'd85616419242672278050054157990378732515248155191920984623355917827871711625906106129789561179082081677506770937259701404185636655864294642711254602823386441022957877254005036440377494889425229642215506714473703870740614690446702228432006089970241426260640059930705006330762704060813443537344708960435364577885;
            5'd22: xpb[80] = 1024'd54245764249240079462304662445687881850822326260373693187859002943967442083146642923584758031040940526118574484522308108790934446855579053919840024381738831281091869150984928460120164400869134180994283908004668860862255147071527066081631550535520699149198185618609894814101920042586855224708164674753545419404;
            5'd23: xpb[80] = 1024'd22875109255807880874555166900997031186396497328826401752362088060063172540387179717379954882999799374730378031784914813396232237846863465128425445940091221539225861047964820479862833912313038719773061101535633850983895603696351903731257011100799972037756311306514783297441136024360266912071620389071726260923;
            5'd24: xpb[80] = 1024'd115571149946500423685604598761120613266669095523014794444997028241135798334936855421190222949616332532785330986505014952580593869679368210892170992514774652731050527514515929837235742615274148979862035903453838687469896910542073514345861041349308694193134340408536729810886880080062311616553765930015501586773;
            5'd25: xpb[80] = 1024'd84200494953068225097855103216429762602243266591467503009500113357231528792177392214985419801575191381397134533767621657185891660670652622100756414073127042989184519411495821856978412126718053518640813096984803677591537367166898351995486501914587967081692466096441618294226096061835723303917221644333682428292;
            5'd26: xpb[80] = 1024'd52829839959636026510105607671738911937817437659920211574003198473327259249417929008780616653534050230008938081030228361791189451661937033309341835631479433247318511308475713876721081638161958057419590290515768667713177823791723189645111962479867239970250591784346506777565312043609134991280677358651863269811;
            5'd27: xpb[80] = 1024'd21459184966203827922356112127048061273391608728372920138506283589422989706658465802575813505492909078620741628292835066396487242653221444517927257189831823505452503205455605896463751149605862596198367484046733657834818280416548027294737423045146512858808717472251395260904528025382546678644133072970044111330;
            5'd28: xpb[80] = 1024'd114155225656896370733405543987171643353664206922561312831141223770495615501208141506386081572109442236675694583012935205580848874485726190281672803764515254697277169672006715253836659852566972856287342285964938494320819587262269637909341453293655235014186746574273341774350272081084591383126278613913819437180;
            5'd29: xpb[80] = 1024'd82784570663464172145656048442480792689238377991014021395644308886591345958448678300181278424068301085287498130275541910186146665477010601490258225322867644955411161568986607273579329364010877395066119479495903484442460043887094475558966913858934507902744872262178230257689488062858003070489734328232000278699;
            5'd30: xpb[80] = 1024'd51413915670031973557906552897789942024812549059466729960147394002687076415689215093976475276027159933899301677538148614791444456468295012698843646881220035213545153465966499293321998875454781933844896673026868474564100500511919313208592374424213780791302997950083118741028704044631414757853190042550181120218;
            5'd31: xpb[80] = 1024'd20043260676599774970157057353099091360386720127919438524650479118782806872929751887771672127986018782511105224800755319396742247459579423907429068439572425471679145362946391313064668386898686472623673866557833464685740957136744150858217834989493053679861123637988007224367920026404826445216645756868361961737;
        endcase
    end

    always_comb begin
        case(flag[27][5:0])
            6'd0: xpb[81] = 1024'd0;
            6'd1: xpb[81] = 1024'd118402998525708529590002708309018553092678872723921757672708637182416164002394283250798505704630113125004603793489174446580083860066652252113167370015293448798597243199534359004033908140688501227011423138431639073768051557101681267218900217460615612551029528077063505883960096078017752083408740562218865885959;
            6'd2: xpb[81] = 1024'd112739301367292317781206489213222673440659318322107831217285419299855432667479427591581940194602551940566058179520855458581103879292084169671174615014255856663503811829497500670437577089859796732712648668476038301171742263982465761472821865238001775835239152740009953737813664082106871149698791297812137287587;
            6'd3: xpb[81] = 1024'd107075604208876105972410270117426793788639763920293904761862201417294701332564571932365374684574990756127512565552536470582123898517516087229181860013218264528410380459460642336841246039031092238413874198520437528575432970863250255726743513015387939119448777402956401591667232086195990215988842033405408689215;
            6'd4: xpb[81] = 1024'd101411907050459894163614051021630914136620209518479978306438983534733969997649716273148809174547429571688966951584217482583143917742948004787189105012180672393316949089423784003244914988202387744115099728564836755979123677744034749980665160792774102403658402065902849445520800090285109282278892768998680090843;
            6'd5: xpb[81] = 1024'd95748209892043682354817831925835034484600655116666051851015765652173238662734860613932243664519868387250421337615898494584163936968379922345196350011143080258223517719386925669648583937373683249816325258609235983382814384624819244234586808570160265687868026728849297299374368094374228348568943504591951492471;
            6'd6: xpb[81] = 1024'd90084512733627470546021612830039154832581100714852125395592547769612507327820004954715678154492307202811875723647579506585183956193811839903203595010105488123130086349350067336052252886544978755517550788653635210786505091505603738488508456347546428972077651391795745153227936098463347414858994240185222894099;
            6'd7: xpb[81] = 1024'd84420815575211258737225393734243275180561546313038198940169329887051775992905149295499112644464746018373330109679260518586203975419243757461210840009067895988036654979313209002455921835716274261218776318698034438190195798386388232742430104124932592256287276054742193007081504102552466481149044975778494295727;
            6'd8: xpb[81] = 1024'd78757118416795046928429174638447395528541991911224272484746112004491044657990293636282547134437184833934784495710941530587223994644675675019218085008030303852943223609276350668859590784887569766920001848742433665593886505267172726996351751902318755540496900717688640860935072106641585547439095711371765697355;
            6'd9: xpb[81] = 1024'd73093421258378835119632955542651515876522437509410346029322894121930313323075437977065981624409623649496238881742622542588244013870107592577225330006992711717849792239239492335263259734058865272621227378786832892997577212147957221250273399679704918824706525380635088714788640110730704613729146446965037098983;
            6'd10: xpb[81] = 1024'd67429724099962623310836736446855636224502883107596419573899676239369581988160582317849416114382062465057693267774303554589264033095539510135232575005955119582756360869202634001666928683230160778322452908831232120401267919028741715504195047457091082108916150043581536568642208114819823680019197182558308500611;
            6'd11: xpb[81] = 1024'd61766026941546411502040517351059756572483328705782493118476458356808850653245726658632850604354501280619147653805984566590284052320971427693239820004917527447662929499165775668070597632401456284023678438875631347804958625909526209758116695234477245393125774706527984422495776118908942746309247918151579902239;
            6'd12: xpb[81] = 1024'd56102329783130199693244298255263876920463774303968566663053240474248119318330870999416285094326940096180602039837665578591304071546403345251247065003879935312569498129128917334474266581572751789724903968920030575208649332790310704012038343011863408677335399369474432276349344122998061812599298653744851303867;
            6'd13: xpb[81] = 1024'd50438632624713987884448079159467997268444219902154640207630022591687387983416015340199719584299378911742056425869346590592324090771835262809254310002842343177476066759092059000877935530744047295426129498964429802612340039671095198265959990789249571961545024032420880130202912127087180878889349389338122705495;
            6'd14: xpb[81] = 1024'd44774935466297776075651860063672117616424665500340713752206804709126656648501159680983154074271817727303510811901027602593344109997267180367261555001804751042382635389055200667281604479915342801127355029008829030016030746551879692519881638566635735245754648695367327984056480131176299945179400124931394107123;
            6'd15: xpb[81] = 1024'd39111238307881564266855640967876237964405111098526787296783586826565925313586304021766588564244256542864965197932708614594364129222699097925268800000767158907289204019018342333685273429086638306828580559053228257419721453432664186773803286344021898529964273358313775837910048135265419011469450860524665508751;
            6'd16: xpb[81] = 1024'd33447541149465352458059421872080358312385556696712860841360368944005193978671448362550023054216695358426419583964389626595384148448131015483276044999729566772195772648981484000088942378257933812529806089097627484823412160313448681027724934121408061814173898021260223691763616139354538077759501596117936910379;
            6'd17: xpb[81] = 1024'd27783843991049140649263202776284478660366002294898934385937151061444462643756592703333457544189134173987873969996070638596404167673562933041283289998691974637102341278944625666492611327429229318231031619142026712227102867194233175281646581898794225098383522684206671545617184143443657144049552331711208312007;
            6'd18: xpb[81] = 1024'd22120146832632928840466983680488599008346447893085007930513933178883731308841737044116892034161572989549328356027751650597424186898994850599290534997654382502008909908907767332896280276600524823932257149186425939630793574075017669535568229676180388382593147347153119399470752147532776210339603067304479713635;
            6'd19: xpb[81] = 1024'd16456449674216717031670764584692719356326893491271081475090715296322999973926881384900326524134011805110782742059432662598444206124426768157297779996616790366915478538870908999299949225771820329633482679230825167034484280955802163789489877453566551666802772010099567253324320151621895276629653802897751115263;
            6'd20: xpb[81] = 1024'd10792752515800505222874545488896839704307339089457155019667497413762268639012025725683761014106450620672237128091113674599464225349858685715305024995579198231822047168834050665703618174943115835334708209275224394438174987836586658043411525230952714951012396673046015107177888155711014342919704538491022516891;
            6'd21: xpb[81] = 1024'd5129055357384293414078326393100960052287784687643228564244279531201537304097170066467195504078889436233691514122794686600484244575290603273312269994541606096728615798797192332107287124114411341035933739319623621841865694717371152297333173008338878235222021335992462961031456159800133409209755274084293918519;
            6'd22: xpb[81] = 1024'd123532053883092823004081034702119513144966657411564986236952916713617701306491453317265701208709002561238295307611969133180568104641942855386479640009835054895325858998331551336141195264802912568047356877751262695609917251819052419516233390468954490786251549413055968844991552237817885492618495836303159804478;
            6'd23: xpb[81] = 1024'd117868356724676611195284815606323633492947103009751059781529698831056969971576597658049135698681441376799749693643650145181588123867374772944486885008797462760232427628294693002544864213974208073748582407795661923013607958699836913770155038246340654070461174076002416698845120241907004558908546571896431206106;
            6'd24: xpb[81] = 1024'd112204659566260399386488596510527753840927548607937133326106480948496238636661741998832570188653880192361204079675331157182608143092806690502494130007759870625138996258257834668948533163145503579449807937840061150417298665580621408024076686023726817354670798738948864552698688245996123625198597307489702607734;
            6'd25: xpb[81] = 1024'd106540962407844187577692377414731874188907994206123206870683263065935507301746886339616004678626319007922658465707012169183628162318238608060501375006722278490045564888220976335352202112316799085151033467884460377820989372461405902277998333801112980638880423401895312406552256250085242691488648043082974009362;
            6'd26: xpb[81] = 1024'd100877265249427975768896158318935994536888439804309280415260045183374775966832030680399439168598757823484112851738693181184648181543670525618508620005684686354952133518184118001755871061488094590852258997928859605224680079342190396531919981578499143923090048064841760260405824254174361757778698778676245410990;
            6'd27: xpb[81] = 1024'd95213568091011763960099939223140114884868885402495353959836827300814044631917175021182873658571196639045567237770374193185668200769102443176515865004647094219858702148147259668159540010659390096553484527973258832628370786222974890785841629355885307207299672727788208114259392258263480824068749514269516812618;
            6'd28: xpb[81] = 1024'd89549870932595552151303720127344235232849331000681427504413609418253313297002319361966308148543635454607021623802055205186688219994534360734523110003609502084765270778110401334563208959830685602254710058017658060032061493103759385039763277133271470491509297390734655968112960262352599890358800249862788214246;
            6'd29: xpb[81] = 1024'd83886173774179340342507501031548355580829776598867501048990391535692581962087463702749742638516074270168476009833736217187708239219966278292530355002571909949671839408073543000966877909001981107955935588062057287435752199984543879293684924910657633775718922053681103821966528266441718956648850985456059615874;
            6'd30: xpb[81] = 1024'd78222476615763128533711281935752475928810222197053574593567173653131850627172608043533177128488513085729930395865417229188728258445398195850537600001534317814578408038036684667370546858173276613657161118106456514839442906865328373547606572688043797059928546716627551675820096270530838022938901721049331017502;
            6'd31: xpb[81] = 1024'd72558779457346916724915062839956596276790667795239648138143955770571119292257752384316611618460951901291384781897098241189748277670830113408544845000496725679484976667999826333774215807344572119358386648150855742243133613746112867801528220465429960344138171379573999529673664274619957089228952456642602419130;
            6'd32: xpb[81] = 1024'd66895082298930704916118843744160716624771113393425721682720737888010387957342896725100046108433390716852839167928779253190768296896262030966552089999459133544391545297962968000177884756515867625059612178195254969646824320626897362055449868242816123628347796042520447383527232278709076155519003192235873820758;
            6'd33: xpb[81] = 1024'd61231385140514493107322624648364836972751558991611795227297520005449656622428041065883480598405829532414293553960460265191788316121693948524559334998421541409298113927926109666581553705687163130760837708239654197050515027507681856309371516020202286912557420705466895237380800282798195221809053927829145222386;
            6'd34: xpb[81] = 1024'd55567687982098281298526405552568957320732004589797868771874302122888925287513185406666915088378268347975747939992141277192808335347125866082566579997383949274204682557889251332985222654858458636462063238284053424454205734388466350563293163797588450196767045368413343091234368286887314288099104663422416624014;
            6'd35: xpb[81] = 1024'd49903990823682069489730186456773077668712450187983942316451084240328193952598329747450349578350707163537202326023822289193828354572557783640573824996346357139111251187852392999388891604029754142163288768328452651857896441269250844817214811574974613480976670031359790945087936290976433354389155399015688025642;
            6'd36: xpb[81] = 1024'd44240293665265857680933967360977198016692895786170015861027866357767462617683474088233784068323145979098656712055503301194848373797989701198581069995308765004017819817815534665792560553201049647864514298372851879261587148150035339071136459352360776765186294694306238798941504295065552420679206134608959427270;
            6'd37: xpb[81] = 1024'd38576596506849645872137748265181318364673341384356089405604648475206731282768618429017218558295584794660111098087184313195868393023421618756588314994271172868924388447778676332196229502372345153565739828417251106665277855030819833325058107129746940049395919357252686652795072299154671486969256870202230828898;
            6'd38: xpb[81] = 1024'd32912899348433434063341529169385438712653786982542162950181430592645999947853762769800653048268023610221565484118865325196888412248853536314595559993233580733830957077741817998599898451543640659266965358461650334068968561911604327578979754907133103333605544020199134506648640303243790553259307605795502230526;
            6'd39: xpb[81] = 1024'd27249202190017222254545310073589559060634232580728236494758212710085268612938907110584087538240462425783019870150546337197908431474285453872602804992195988598737525707704959665003567400714936164968190888506049561472659268792388821832901402684519266617815168683145582360502208307332909619549358341388773632154;
            6'd40: xpb[81] = 1024'd21585505031601010445749090977793679408614678178914310039334994827524537278024051451367522028212901241344474256182227349198928450699717371430610049991158396463644094337668101331407236349886231670669416418550448788876349975673173316086823050461905429902024793346092030214355776311422028685839409076982045033782;
            6'd41: xpb[81] = 1024'd15921807873184798636952871881997799756595123777100383583911776944963805943109195792150956518185340056905928642213908361199948469925149288988617294990120804328550662967631242997810905299057527176370641948594848016280040682553957810340744698239291593186234418009038478068209344315511147752129459812575316435410;
            6'd42: xpb[81] = 1024'd10258110714768586828156652786201920104575569375286457128488559062403074608194340132934391008157778872467383028245589373200968489150581206546624539989083212193457231597594384664214574248228822682071867478639247243683731389434742304594666346016677756470444042671984925922062912319600266818419510548168587837038;
            6'd43: xpb[81] = 1024'd4594413556352375019360433690406040452556014973472530673065341179842343273279484473717825498130217688028837414277270385201988508376013124104631784988045620058363800227557526330618243197400118187773093008683646471087422096315526798848587993794063919754653667334931373775916480323689385884709561283761859238666;
            6'd44: xpb[81] = 1024'd122997412082060904609363141999424593545234887697394288345773978362258507275673767724516331202760330813033441207766444831782072368442665376217799155003339068856961043427091885334652151338088619414784516147115285544855473653417208066067488211254679532305683195411994879659876576401707137968118301845980725124625;
            6'd45: xpb[81] = 1024'd117333714923644692800566922903628713893215333295580361890350760479697775940758912065299765692732769628594895593798125843783092387668097293775806400002301476721867612057055027001055820287259914920485741677159684772259164360297992560321409859032065695589892820074941327513730144405796257034408352581573996526253;
            6'd46: xpb[81] = 1024'd111670017765228480991770703807832834241195778893766435434927542597137044605844056406083200182705208444156349979829806855784112406893529211333813645001263884586774180687018168667459489236431210426186967207204083999662855067178777054575331506809451858874102444737887775367583712409885376100698403317167267927881;
            6'd47: xpb[81] = 1024'd106006320606812269182974484712036954589176224491952508979504324714576313270929200746866634672677647259717804365861487867785132426118961128891820890000226292451680749316981310333863158185602505931888192737248483227066545774059561548829253154586838022158312069400834223221437280413974495166988454052760539329509;
            6'd48: xpb[81] = 1024'd100342623448396057374178265616241074937156670090138582524081106832015581936014345087650069162650086075279258751893168879786152445344393046449828134999188700316587317946944452000266827134773801437589418267292882454470236480940346043083174802364224185442521694063780671075290848418063614233278504788353810731137;
            6'd49: xpb[81] = 1024'd94678926289979845565382046520445195285137115688324656068657888949454850601099489428433503652622524890840713137924849891787172464569824964007835379998151108181493886576907593666670496083945096943290643797337281681873927187821130537337096450141610348726731318726727118929144416422152733299568555523947082132765;
            6'd50: xpb[81] = 1024'd89015229131563633756585827424649315633117561286510729613234671066894119266184633769216938142594963706402167523956530903788192483795256881565842624997113516046400455206870735333074165033116392448991869327381680909277617894701915031591018097918996512010940943389673566782997984426241852365858606259540353534393;
            6'd51: xpb[81] = 1024'd83351531973147421947789608328853435981098006884696803157811453184333387931269778110000372632567402521963621909988211915789212503020688799123849869996075923911307023836833876999477833982287687954693094857426080136681308601582699525844939745696382675295150568052620014636851552430330971432148656995133624936021;
            6'd52: xpb[81] = 1024'd77687834814731210138993389233057556329078452482882876702388235301772656596354922450783807122539841337525076296019892927790232522246120716681857114995038331776213592466797018665881502931458983460394320387470479364084999308463484020098861393473768838579360192715566462490705120434420090498438707730726896337649;
            6'd53: xpb[81] = 1024'd72024137656314998330197170137261676677058898081068950246965017419211925261440066791567241612512280153086530682051573939791252541471552634239864359994000739641120161096760160332285171880630278966095545917514878591488690015344268514352783041251155001863569817378512910344558688438509209564728758466320167739277;
            6'd54: xpb[81] = 1024'd66360440497898786521400951041465797025039343679255023791541799536651193926525211132350676102484718968647985068083254951792272560696984551797871604992963147506026729726723301998688840829801574471796771447559277818892380722225053008606704689028541165147779442041459358198412256442598328631018809201913439140905;
            6'd55: xpb[81] = 1024'd60696743339482574712604731945669917373019789277441097336118581654090462591610355473134110592457157784209439454114935963793292579922416469355878849991925555370933298356686443665092509778972869977497996977603677046296071429105837502860626336805927328431989066704405806052265824446687447697308859937506710542533;
            6'd56: xpb[81] = 1024'd55033046181066362903808512849874037721000234875627170880695363771529731256695499813917545082429596599770893840146616975794312599147848386913886094990887963235839866986649585331496178728144165483199222507648076273699762135986621997114547984583313491716198691367352253906119392450776566763598910673099981944161;
            6'd57: xpb[81] = 1024'd49369349022650151095012293754078158068980680473813244425272145888968999921780644154700979572402035415332348226178297987795332618373280304471893339989850371100746435616612726997899847677315460988900448037692475501103452842867406491368469632360699655000408316030298701759972960454865685829888961408693253345789;
            6'd58: xpb[81] = 1024'd43705651864233939286216074658282278416961126071999317969848928006408268586865788495484414062374474230893802612209978999796352637598712222029900584988812778965653004246575868664303516626486756494601673567736874728507143549748190985622391280138085818284617940693245149613826528458954804896179012144286524747417;
            6'd59: xpb[81] = 1024'd38041954705817727477419855562486398764941571670185391514425710123847537251950932836267848552346913046455256998241660011797372656824144139587907829987775186830559572876539010330707185575658052000302899097781273955910834256628975479876312927915471981568827565356191597467680096463043923962469062879879796149045;
            6'd60: xpb[81] = 1024'd32378257547401515668623636466690519112922017268371465059002492241286805917036077177051283042319351862016711384273341023798392676049576057145915074986737594695466141506502151997110854524829347506004124627825673183314524963509759974130234575692858144853037190019138045321533664467133043028759113615473067550673;
            6'd61: xpb[81] = 1024'd26714560388985303859827417370894639460902462866557538603579274358726074582121221517834717532291790677578165770305022035799412695275007974703922319985700002560372710136465293663514523474000643011705350157870072410718215670390544468384156223470244308137246814682084493175387232471222162095049164351066338952301;
            6'd62: xpb[81] = 1024'd21050863230569092051031198275098759808882908464743612148156056476165343247206365858618152022264229493139620156336703047800432714500439892261929564984662410425279278766428435329918192423171938517406575687914471638121906377271328962638077871247630471421456439345030941029240800475311281161339215086659610353929;
            6'd63: xpb[81] = 1024'd15387166072152880242234979179302880156863354062929685692732838593604611912291510199401586512236668308701074542368384059801452733725871809819936809983624818290185847396391576996321861372343234023107801217958870865525597084152113456891999519025016634705666064007977388883094368479400400227629265822252881755557;
        endcase
    end

    always_comb begin
        case(flag[27][11:6])
            6'd0: xpb[82] = 1024'd0;
            6'd1: xpb[82] = 1024'd9723468913736668433438760083507000504843799661115759237309620711043880577376654540185021002209107124262528928400065071802472752951303727377944054982587226155092416026354718662725530321514529528809026748003270092929287791032897951145921166802402797989875688670923836736947936483489519293919316557846153157185;
            6'd2: xpb[82] = 1024'd19446937827473336866877520167014001009687599322231518474619241422087761154753309080370042004418214248525057856800130143604945505902607454755888109965174452310184832052709437325451060643029059057618053496006540185858575582065795902291842333604805595979751377341847673473895872966979038587838633115692306314370;
            6'd3: xpb[82] = 1024'd29170406741210005300316280250521001514531398983347277711928862133131641732129963620555063006627321372787586785200195215407418258853911182133832164947761678465277248079064155988176590964543588586427080244009810278787863373098693853437763500407208393969627066012771510210843809450468557881757949673538459471555;
            6'd4: xpb[82] = 1024'd38893875654946673733755040334028002019375198644463036949238482844175522309506618160740084008836428497050115713600260287209891011805214909511776219930348904620369664105418874650902121286058118115236106992013080371717151164131591804583684667209611191959502754683695346947791745933958077175677266231384612628740;
            6'd5: xpb[82] = 1024'd48617344568683342167193800417535002524218998305578796186548103555219402886883272700925105011045535621312644642000325359012363764756518636889720274912936130775462080131773593313627651607572647644045133740016350464646438955164489755729605834012013989949378443354619183684739682417447596469596582789230765785925;
            6'd6: xpb[82] = 1024'd58340813482420010600632560501042003029062797966694555423857724266263283464259927241110126013254642745575173570400390430814836517707822364267664329895523356930554496158128311976353181929087177172854160488019620557575726746197387706875527000814416787939254132025543020421687618900937115763515899347076918943110;
            6'd7: xpb[82] = 1024'd68064282396156679034071320584549003533906597627810314661167344977307164041636581781295147015463749869837702498800455502617309270659126091645608384878110583085646912184483030639078712250601706701663187236022890650505014537230285658021448167616819585929129820696466857158635555384426635057435215904923072100295;
            6'd8: xpb[82] = 1024'd77787751309893347467510080668056004038750397288926073898476965688351044619013236321480168017672856994100231427200520574419782023610429819023552439860697809240739328210837749301804242572116236230472213984026160743434302328263183609167369334419222383919005509367390693895583491867916154351354532462769225257480;
            6'd9: xpb[82] = 1024'd87511220223630015900948840751563004543594196950041833135786586399394925196389890861665189019881964118362760355600585646222254776561733546401496494843285035395831744237192467964529772893630765759281240732029430836363590119296081560313290501221625181908881198038314530632531428351405673645273849020615378414665;
            6'd10: xpb[82] = 1024'd97234689137366684334387600835070005048437996611157592373096207110438805773766545401850210022091071242625289284000650718024727529513037273779440549825872261550924160263547186627255303215145295288090267480032700929292877910328979511459211668024027979898756886709238367369479364834895192939193165578461531571850;
            6'd11: xpb[82] = 1024'd106958158051103352767826360918577005553281796272273351610405827821482686351143199942035231024300178366887818212400715789827200282464341001157384604808459487706016576289901905289980833536659824816899294228035971022222165701361877462605132834826430777888632575380162204106427301318384712233112482136307684729035;
            6'd12: xpb[82] = 1024'd116681626964840021201265121002084006058125595933389110847715448532526566928519854482220252026509285491150347140800780861629673035415644728535328659791046713861108992316256623952706363858174354345708320976039241115151453492394775413751054001628833575878508264051086040843375237801874231527031798694153837886220;
            6'd13: xpb[82] = 1024'd2338400194451948235904953680776573818270968468769185956893214178593552168587370112390201814060718305969726661743352498853081947525728121358112589757302899082510733773040125277801654988171678153207150115655271361716380433206776591931996598748006924601564049307892819550216646211435117803832425425374396559074;
            6'd14: xpb[82] = 1024'd12061869108188616669343713764283574323114768129884945194202834889637432745964024652575222816269825430232255590143417570655554700477031848736056644739890125237603149799394843940527185309686207682016176863658541454645668224239674543077917765550409722591439737978816656287164582694924637097751741983220549716259;
            6'd15: xpb[82] = 1024'd21785338021925285102782473847790574827958567791000704431512455600681313323340679192760243818478932554494784518543482642458027453428335576114000699722477351392695565825749562603252715631200737210825203611661811547574956015272572494223838932352812520581315426649740493024112519178414156391671058541066702873444;
            6'd16: xpb[82] = 1024'd31508806935661953536221233931297575332802367452116463668822076311725193900717333732945264820688039678757313446943547714260500206379639303491944754705064577547787981852104281265978245952715266739634230359665081640504243806305470445369760099155215318571191115320664329761060455661903675685590375098912856030629;
            6'd17: xpb[82] = 1024'd41232275849398621969659994014804575837646167113232222906131697022769074478093988273130285822897146803019842375343612786062972959330943030869888809687651803702880397878458999928703776274229796268443257107668351733433531597338368396515681265957618116561066803991588166498008392145393194979509691656759009187814;
            6'd18: xpb[82] = 1024'd50955744763135290403098754098311576342489966774347982143441317733812955055470642813315306825106253927282371303743677857865445712282246758247832864670239029857972813904813718591429306595744325797252283855671621826362819388371266347661602432760020914550942492662512003234956328628882714273429008214605162344999;
            6'd19: xpb[82] = 1024'd60679213676871958836537514181818576847333766435463741380750938444856835632847297353500327827315361051544900232143742929667918465233550485625776919652826256013065229931168437254154836917258855326061310603674891919292107179404164298807523599562423712540818181333435839971904265112372233567348324772451315502184;
            6'd20: xpb[82] = 1024'd70402682590608627269976274265325577352177566096579500618060559155900716210223951893685348829524468175807429160543808001470391218184854213003720974635413482168157645957523155916880367238773384854870337351678162012221394970437062249953444766364826510530693870004359676708852201595861752861267641330297468659369;
            6'd21: xpb[82] = 1024'd80126151504345295703415034348832577857021365757695259855370179866944596787600606433870369831733575300069958088943873073272863971136157940381665029618000708323250061983877874579605897560287914383679364099681432105150682761469960201099365933167229308520569558675283513445800138079351272155186957888143621816554;
            6'd22: xpb[82] = 1024'd89849620418081964136853794432339578361865165418811019092679800577988477364977260974055390833942682424332487017343938145075336724087461667759609084600587934478342478010232593242331427881802443912488390847684702198079970552502858152245287099969632106510445247346207350182748074562840791449106274445989774973739;
            6'd23: xpb[82] = 1024'd99573089331818632570292554515846578866708965079926778329989421289032357942353915514240411836151789548595015945744003216877809477038765395137553139583175160633434894036587311905056958203316973441297417595687972291009258343535756103391208266772034904500320936017131186919696011046330310743025591003835928130924;
            6'd24: xpb[82] = 1024'd109296558245555301003731314599353579371552764741042537567299042000076238519730570054425432838360896672857544874144068288680282229990069122515497194565762386788527310062942030567782488524831502970106444343691242383938546134568654054537129433574437702490196624688055023656643947529819830036944907561682081288109;
            6'd25: xpb[82] = 1024'd119020027159291969437170074682860579876396564402158296804608662711120119097107224594610453840570003797120073802544133360482754982941372849893441249548349612943619726089296749230508018846346032498915471091694512476867833925601552005683050600376840500480072313358978860393591884013309349330864224119528234445294;
            6'd26: xpb[82] = 1024'd4676800388903896471809907361553147636541936937538371913786428357187104337174740224780403628121436611939453323486704997706163895051456242716225179514605798165021467546080250555603309976343356306414300231310542723432760866413553183863993197496013849203128098615785639100433292422870235607664850850748793118148;
            6'd27: xpb[82] = 1024'd14400269302640564905248667445060148141385736598654131151096049068230984914551394764965424630330543736201982251886770069508636648002759970094169234497193024320113883572434969218328840297857885835223326979313812816362048657446451135009914364298416647193003787286709475837381228906359754901584167408594946275333;
            6'd28: xpb[82] = 1024'd24123738216377233338687427528567148646229536259769890388405669779274865491928049305150445632539650860464511180286835141311109400954063697472113289479780250475206299598789687881054370619372415364032353727317082909291336448479349086155835531100819445182879475957633312574329165389849274195503483966441099432518;
            6'd29: xpb[82] = 1024'd33847207130113901772126187612074149151073335920885649625715290490318746069304703845335466634748757984727040108686900213113582153905367424850057344462367476630298715625144406543779900940886944892841380475320353002220624239512247037301756697903222243172755164628557149311277101873338793489422800524287252589703;
            6'd30: xpb[82] = 1024'd43570676043850570205564947695581149655917135582001408863024911201362626646681358385520487636957865108989569037086965284916054906856671152228001399444954702785391131651499125206505431262401474421650407223323623095149912030545144988447677864705625041162630853299480986048225038356828312783342117082133405746888;
            6'd31: xpb[82] = 1024'd53294144957587238639003707779088150160760935243117168100334531912406507224058012925705508639166972233252097965487030356718527659807974879605945454427541928940483547677853843869230961583916003950459433971326893188079199821578042939593599031508027839152506541970404822785172974840317832077261433639979558904073;
            6'd32: xpb[82] = 1024'd63017613871323907072442467862595150665604734904232927337644152623450387801434667465890529641376079357514626893887095428521000412759278606983889509410129155095575963704208562531956491905430533479268460719330163281008487612610940890739520198310430637142382230641328659522120911323807351371180750197825712061258;
            6'd33: xpb[82] = 1024'd72741082785060575505881227946102151170448534565348686574953773334494268378811322006075550643585186481777155822287160500323473165710582334361833564392716381250668379730563281194682022226945063008077487467333433373937775403643838841885441365112833435132257919312252496259068847807296870665100066755671865218443;
            6'd34: xpb[82] = 1024'd82464551698797243939319988029609151675292334226464445812263394045538148956187976546260571645794293606039684750687225572125945918661886061739777619375303607405760795756917999857407552548459592536886514215336703466867063194676736793031362531915236233122133607983176332996016784290786389959019383313518018375628;
            6'd35: xpb[82] = 1024'd92188020612533912372758748113116152180136133887580205049573014756582029533564631086445592648003400730302213679087290643928418671613189789117721674357890833560853211783272718520133082869974122065695540963339973559796350985709634744177283698717639031112009296654100169732964720774275909252938699871364171532813;
            6'd36: xpb[82] = 1024'd101911489526270580806197508196623152684979933548695964286882635467625910110941285626630613650212507854564742607487355715730891424564493516495665729340478059715945627809627437182858613191488651594504567711343243652725638776742532695323204865520041829101884985325024006469912657257765428546858016429210324689998;
            6'd37: xpb[82] = 1024'd111634958440007249239636268280130153189823733209811723524192256178669790688317940166815634652421614978827271535887420787533364177515797243873609784323065285871038043835982155845584143513003181123313594459346513745654926567775430646469126032322444627091760673995947843206860593741254947840777332987056477847183;
            6'd38: xpb[82] = 1024'd121358427353743917673075028363637153694667532870927482761501876889713671265694594707000655654630722103089800464287485859335836930467100971251553839305652512026130459862336874508309673834517710652122621207349783838584214358808328597615047199124847425081636362666871679943808530224744467134696649544902631004368;
            6'd39: xpb[82] = 1024'd7015200583355844707714861042329721454812905406307557870679642535780656505762110337170605442182154917909179985230057496559245842577184364074337769271908697247532201319120375833404964964515034459621450346965814085149141299620329775795989796244020773804692147923678458650649938634305353411497276276123189677222;
            6'd40: xpb[82] = 1024'd16738669497092513141153621125836721959656705067423317107989263246824537083138764877355626444391262042171708913630122568361718595528488091452281824254495923402624617345475094496130495286029563988430477094969084178078429090653227726941910963046423571794567836594602295387597875117794872705416592833969342834407;
            6'd41: xpb[82] = 1024'd26462138410829181574592381209343722464500504728539076345298883957868417660515419417540647446600369166434237842030187640164191348479791818830225879237083149557717033371829813158856025607544093517239503842972354271007716881686125678087832129848826369784443525265526132124545811601284391999335909391815495991592;
            6'd42: xpb[82] = 1024'd36185607324565850008031141292850722969344304389654835582608504668912298237892073957725668448809476290696766770430252711966664101431095546208169934219670375712809449398184531821581555929058623046048530590975624363937004672719023629233753296651229167774319213936449968861493748084773911293255225949661649148777;
            6'd43: xpb[82] = 1024'd45909076238302518441469901376357723474188104050770594819918125379956178815268728497910689451018583414959295698830317783769136854382399273586113989202257601867901865424539250484307086250573152574857557338978894456866292463751921580379674463453631965764194902607373805598441684568263430587174542507507802305962;
            6'd44: xpb[82] = 1024'd55632545152039186874908661459864723979031903711886354057227746091000059392645383038095710453227690539221824627230382855571609607333703000964058044184844828022994281450893969147032616572087682103666584086982164549795580254784819531525595630256034763754070591278297642335389621051752949881093859065353955463147;
            6'd45: xpb[82] = 1024'd65356014065775855308347421543371724483875703373002113294537366802043939970022037578280731455436797663484353555630447927374082360285006728342002099167432054178086697477248687809758146893602211632475610834985434642724868045817717482671516797058437561743946279949221479072337557535242469175013175623200108620332;
            6'd46: xpb[82] = 1024'd75079482979512523741786181626878724988719503034117872531846987513087820547398692118465752457645904787746882484030512999176555113236310455719946154150019280333179113503603406472483677215116741161284637582988704735654155836850615433817437963860840359733821968620145315809285494018731988468932492181046261777517;
            6'd47: xpb[82] = 1024'd84802951893249192175224941710385725493563302695233631769156608224131701124775346658650773459855011912009411412430578070979027866187614183097890209132606506488271529529958125135209207536631270690093664330991974828583443627883513384963359130663243157723697657291069152546233430502221507762851808738892414934702;
            6'd48: xpb[82] = 1024'd94526420806985860608663701793892725998407102356349391006466228935175581702152001198835794462064119036271940340830643142781500619138917910475834264115193732643363945556312843797934737858145800218902691078995244921512731418916411336109280297465645955713573345961992989283181366985711027056771125296738568091887;
            6'd49: xpb[82] = 1024'd104249889720722529042102461877399726503250902017465150243775849646219462279528655739020815464273226160534469269230708214583973372090221637853778319097780958798456361582667562460660268179660329747711717826998515014442019209949309287255201464268048753703449034632916826020129303469200546350690441854584721249072;
            6'd50: xpb[82] = 1024'd113973358634459197475541221960906727008094701678580909481085470357263342856905310279205836466482333284796998197630773286386446125041525365231722374080368184953548777609022281123385798501174859276520744575001785107371307000982207238401122631070451551693324723303840662757077239952690065644609758412430874406257;
            6'd51: xpb[82] = 1024'd123696827548195865908979982044413727512938501339696668718395091068307223434281964819390857468691440409059527126030838358188918877992829092609666429062955411108641193635376999786111328822689388805329771323005055200300594792015105189547043797872854349683200411974764499494025176436179584938529074970277027563442;
            6'd52: xpb[82] = 1024'd9353600777807792943619814723106295273083873875076743827572856714374208674349480449560807256242873223878906646973409995412327790102912485432450359029211596330042935092160501111206619952686712612828600462621085446865521732827106367727986394992027698406256197231571278200866584845740471215329701701497586236296;
            6'd53: xpb[82] = 1024'd19077069691544461377058574806613295777927673536192503064882477425418089251726134989745828258451980348141435575373475067214800543054216212810394414011798822485135351118515219773932150274201242141637627210624355539794809523860004318873907561794430496396131885902495114937814521329229990509249018259343739393481;
            6'd54: xpb[82] = 1024'd28800538605281129810497334890120296282771473197308262302192098136461969829102789529930849260661087472403964503773540139017273296005519940188338468994386048640227767144869938436657680595715771670446653958627625632724097314892902270019828728596833294386007574573418951674762457812719509803168334817189892550666;
            6'd55: xpb[82] = 1024'd38524007519017798243936094973627296787615272858424021539501718847505850406479444070115870262870194596666493432173605210819746048956823667566282523976973274795320183171224657099383210917230301199255680706630895725653385105925800221165749895399236092375883263244342788411710394296209029097087651375036045707851;
            6'd56: xpb[82] = 1024'd48247476432754466677374855057134297292459072519539780776811339558549730983856098610300891265079301720929022360573670282622218801908127394944226578959560500950412599197579375762108741238744830728064707454634165818582672896958698172311671062201638890365758951915266625148658330779698548391006967932882198865036;
            6'd57: xpb[82] = 1024'd57970945346491135110813615140641297797302872180655540014120960269593611561232753150485912267288408845191551288973735354424691554859431122322170633942147727105505015223934094424834271560259360256873734202637435911511960687991596123457592229004041688355634640586190461885606267263188067684926284490728352022221;
            6'd58: xpb[82] = 1024'd67694414260227803544252375224148298302146671841771299251430580980637492138609407690670933269497515969454080217373800426227164307810734849700114688924734953260597431250288813087559801881773889785682760950640706004441248479024494074603513395806444486345510329257114298622554203746677586978845601048574505179406;
            6'd59: xpb[82] = 1024'd77417883173964471977691135307655298806990471502887058488740201691681372715986062230855954271706623093716609145773865498029637060762038577078058743907322179415689847276643531750285332203288419314491787698643976097370536270057392025749434562608847284335386017928038135359502140230167106272764917606420658336591;
            6'd60: xpb[82] = 1024'd87141352087701140411129895391162299311834271164002817726049822402725253293362716771040975273915730217979138074173930569832109813713342304456002798889909405570782263302998250413010862524802948843300814446647246190299824061090289976895355729411250082325261706598961972096450076713656625566684234164266811493776;
            6'd61: xpb[82] = 1024'd96864821001437808844568655474669299816678070825118576963359443113769133870739371311225996276124837342241667002573995641634582566664646031833946853872496631725874679329352969075736392846317478372109841194650516283229111852123187928041276896213652880315137395269885808833398013197146144860603550722112964650961;
            6'd62: xpb[82] = 1024'd106588289915174477278007415558176300321521870486234336200669063824813014448116025851411017278333944466504195930974060713437055319615949759211890908855083857880967095355707687738461923167832007900918867942653786376158399643156085879187198063016055678305013083940809645570345949680635664154522867279959117808146;
            6'd63: xpb[82] = 1024'd116311758828911145711446175641683300826365670147350095437978684535856895025492680391596038280543051590766724859374125785239528072567253486589834963837671084036059511382062406401187453489346537429727894690657056469087687434188983830333119229818458476294888772611733482307293886164125183448442183837805270965331;
        endcase
    end

    always_comb begin
        case(flag[27][16:12])
            5'd0: xpb[83] = 1024'd0;
            5'd1: xpb[83] = 1024'd1968532058523072746086008320375868586511042682730170547156450181923880265560196021765988068094484405586104380316697422462936984677336879412618893803927269257461252838845907726282744619343861237226723830273086715652614375000985008514061826937631825017944557868540261014135294573686069725242810569025829638185;
            5'd2: xpb[83] = 1024'd3937064117046145492172016640751737173022085365460341094312900363847760531120392043531976136188968811172208760633394844925873969354673758825237787607854538514922505677691815452565489238687722474453447660546173431305228750001970017028123653875263650035889115737080522028270589147372139450485621138051659276370;
            5'd3: xpb[83] = 1024'd5905596175569218238258024961127605759533128048190511641469350545771640796680588065297964204283453216758313140950092267388810954032010638237856681411781807772383758516537723178848233858031583711680171490819260146957843125002955025542185480812895475053833673605620783042405883721058209175728431707077488914555;
            5'd4: xpb[83] = 1024'd7874128234092290984344033281503474346044170730920682188625800727695521062240784087063952272377937622344417521266789689851747938709347517650475575215709077029845011355383630905130978477375444948906895321092346862610457500003940034056247307750527300071778231474161044056541178294744278900971242276103318552740;
            5'd5: xpb[83] = 1024'd9842660292615363730430041601879342932555213413650852735782250909619401327800980108829940340472422027930521901583487112314684923386684397063094469019636346287306264194229538631413723096719306186133619151365433578263071875004925042570309134688159125089722789342701305070676472868430348626214052845129148190925;
            5'd6: xpb[83] = 1024'd11811192351138436476516049922255211519066256096381023282938701091543281593361176130595928408566906433516626281900184534777621908064021276475713362823563615544767517033075446357696467716063167423360342981638520293915686250005910051084370961625790950107667347211241566084811767442116418351456863414154977829110;
            5'd7: xpb[83] = 1024'd13779724409661509222602058242631080105577298779111193830095151273467161858921372152361916476661390839102730662216881957240558892741358155888332256627490884802228769871921354083979212335407028660587066811911607009568300625006895059598432788563422775125611905079781827098947062015802488076699673983180807467295;
            5'd8: xpb[83] = 1024'd15748256468184581968688066563006948692088341461841364377251601455391042124481568174127904544755875244688835042533579379703495877418695035300951150431418154059690022710767261810261956954750889897813790642184693725220915000007880068112494615501054600143556462948322088113082356589488557801942484552206637105480;
            5'd9: xpb[83] = 1024'd17716788526707654714774074883382817278599384144571534924408051637314922390041764195893892612850359650274939422850276802166432862096031914713570044235345423317151275549613169536544701574094751135040514472457780440873529375008865076626556442438686425161501020816862349127217651163174627527185295121232466743665;
            5'd10: xpb[83] = 1024'd19685320585230727460860083203758685865110426827301705471564501819238802655601960217659880680944844055861043803166974224629369846773368794126188938039272692574612528388459077262827446193438612372267238302730867156526143750009850085140618269376318250179445578685402610141352945736860697252428105690258296381850;
            5'd11: xpb[83] = 1024'd21653852643753800206946091524134554451621469510031876018720952001162682921162156239425868749039328461447148183483671647092306831450705673538807831843199961832073781227304984989110190812782473609493962133003953872178758125010835093654680096313950075197390136553942871155488240310546766977670916259284126020035;
            5'd12: xpb[83] = 1024'd23622384702276872953032099844510423038132512192762046565877402183086563186722352261191856817133812867033252563800369069555243816128042552951426725647127231089535034066150892715392935432126334846720685963277040587831372500011820102168741923251581900215334694422483132169623534884232836702913726828309955658220;
            5'd13: xpb[83] = 1024'd25590916760799945699118108164886291624643554875492217113033852365010443452282548282957844885228297272619356944117066492018180800805379432364045619451054500346996286904996800441675680051470196083947409793550127303483986875012805110682803750189213725233279252291023393183758829457918906428156537397335785296405;
            5'd14: xpb[83] = 1024'd27559448819323018445204116485262160211154597558222387660190302546934323717842744304723832953322781678205461324433763914481117785482716311776664513254981769604457539743842708167958424670814057321174133623823214019136601250013790119196865577126845550251223810159563654197894124031604976153399347966361614934590;
            5'd15: xpb[83] = 1024'd29527980877846091191290124805638028797665640240952558207346752728858203983402940326489821021417266083791565704750461336944054770160053191189283407058909038861918792582688615894241169290157918558400857454096300734789215625014775127710927404064477375269168368028103915212029418605291045878642158535387444572775;
            5'd16: xpb[83] = 1024'd31496512936369163937376133126013897384176682923682728754503202910782084248963136348255809089511750489377670085067158759406991754837390070601902300862836308119380045421534523620523913909501779795627581284369387450441830000015760136224989231002109200287112925896644176226164713178977115603884969104413274210960;
            5'd17: xpb[83] = 1024'd33465044994892236683462141446389765970687725606412899301659653092705964514523332370021797157606234894963774465383856181869928739514726950014521194666763577376841298260380431346806658528845641032854305114642474166094444375016745144739051057939741025305057483765184437240300007752663185329127779673439103849145;
            5'd18: xpb[83] = 1024'd35433577053415309429548149766765634557198768289143069848816103274629844780083528391787785225700719300549878845700553604332865724192063829427140088470690846634302551099226339073089403148189502270081028944915560881747058750017730153253112884877372850323002041633724698254435302326349255054370590242464933487330;
            5'd19: xpb[83] = 1024'd37402109111938382175634158087141503143709810971873240395972553456553725045643724413553773293795203706135983226017251026795802708869400708839758982274618115891763803938072246799372147767533363507307752775188647597399673125018715161767174711815004675340946599502264959268570596900035324779613400811490763125515;
            5'd20: xpb[83] = 1024'd39370641170461454921720166407517371730220853654603410943129003638477605311203920435319761361889688111722087606333948449258739693546737588252377876078545385149225056776918154525654892386877224744534476605461734313052287500019700170281236538752636500358891157370805220282705891473721394504856211380516592763700;
            5'd21: xpb[83] = 1024'd41339173228984527667806174727893240316731896337333581490285453820401485576764116457085749429984172517308191986650645871721676678224074467664996769882472654406686309615764062251937637006221085981761200435734821028704901875020685178795298365690268325376835715239345481296841186047407464230099021949542422401885;
            5'd22: xpb[83] = 1024'd43307705287507600413892183048269108903242939020063752037441904002325365842324312478851737498078656922894296366967343294184613662901411347077615663686399923664147562454609969978220381625564947218987924266007907744357516250021670187309360192627900150394780273107885742310976480621093533955341832518568252040070;
            5'd23: xpb[83] = 1024'd45276237346030673159978191368644977489753981702793922584598354184249246107884508500617725566173141328480400747284040716647550647578748226490234557490327192921608815293455877704503126244908808456214648096280994460010130625022655195823422019565531975412724830976426003325111775194779603680584643087594081678255;
            5'd24: xpb[83] = 1024'd47244769404553745906064199689020846076265024385524093131754804366173126373444704522383713634267625734066505127600738139110487632256085105902853451294254462179070068132301785430785870864252669693441371926554081175662745000023640204337483846503163800430669388844966264339247069768465673405827453656619911316440;
            5'd25: xpb[83] = 1024'd49213301463076818652150208009396714662776067068254263678911254548097006639004900544149701702362110139652609507917435561573424616933421985315472345098181731436531320971147693157068615483596530930668095756827167891315359375024625212851545673440795625448613946713506525353382364342151743131070264225645740954625;
            5'd26: xpb[83] = 1024'd51181833521599891398236216329772583249287109750984434226067704730020886904565096565915689770456594545238713888234132984036361601610758864728091238902109000693992573809993600883351360102940392167894819587100254606967973750025610221365607500378427450466558504582046786367517658915837812856313074794671570592810;
            5'd27: xpb[83] = 1024'd53150365580122964144322224650148451835798152433714604773224154911944767170125292587681677838551078950824818268550830406499298586288095744140710132706036269951453826648839508609634104722284253405121543417373341322620588125026595229879669327316059275484503062450587047381652953489523882581555885363697400230995;
            5'd28: xpb[83] = 1024'd55118897638646036890408232970524320422309195116444775320380605093868647435685488609447665906645563356410922648867527828962235570965432623553329026509963539208915079487685416335916849341628114642348267247646428038273202500027580238393731154253691100502447620319127308395788248063209952306798695932723229869180;
            5'd29: xpb[83] = 1024'd57087429697169109636494241290900189008820237799174945867537055275792527701245684631213653974740047761997027029184225251425172555642769502965947920313890808466376332326531324062199593960971975879574991077919514753925816875028565246907792981191322925520392178187667569409923542636896022032041506501749059507365;
            5'd30: xpb[83] = 1024'd59055961755692182382580249611276057595331280481905116414693505457716407966805880652979642042834532167583131409500922673888109540320106382378566814117818077723837585165377231788482338580315837116801714908192601469578431250029550255421854808128954750538336736056207830424058837210582091757284317070774889145550;
            5'd31: xpb[83] = 1024'd61024493814215255128666257931651926181842323164635286961849955639640288232366076674745630110929016573169235789817620096351046524997443261791185707921745346981298838004223139514765083199659698354028438738465688185231045625030535263935916635066586575556281293924748091438194131784268161482527127639800718783735;
        endcase
    end

    always_comb begin
        case(flag[28][5:0])
            6'd0: xpb[84] = 1024'd0;
            6'd1: xpb[84] = 1024'd31496512936369163937376133126013897384176682923682728754503202910782084248963136348255809089511750489377670085067158759406991754837390070601902300862836308119380045421534523620523913909501779795627581284369387450441830000015760136224989231002109200287112925896644176226164713178977115603884969104413274210960;
            6'd2: xpb[84] = 1024'd62993025872738327874752266252027794768353365847365457509006405821564168497926272696511618179023500978755340170134317518813983509674780141203804601725672616238760090843069047241047827819003559591255162568738774900883660000031520272449978462004218400574225851793288352452329426357954231207769938208826548421920;
            6'd3: xpb[84] = 1024'd94489538809107491812128399378041692152530048771048186263509608732346252746889409044767427268535251468133010255201476278220975264512170211805706902588508924358140136264603570861571741728505339386882743853108162351325490000047280408674967693006327600861338777689932528678494139536931346811654907313239822632880;
            6'd4: xpb[84] = 1024'd1919356061351914350705605099241156792008304568995230889880956578151441658543406483008165143389327648067530932811141603048903178508339947852449078435014191543829507116566877144465416446489913461200127529090309955402959149842143771934978354325207351881631800172459646874552324641979829398421186591027502359509;
            6'd5: xpb[84] = 1024'd33415868997721078288081738225255054176184987492677959644384159488933525907506542831263974232901078137445201017878300362455894933345730018454351379297850499663209552538101400764989330355991693256827708813459697405844789149857903908159967585327316552168744726069103823100717037820956945002306155695440776570469;
            6'd6: xpb[84] = 1024'd64912381934090242225457871351268951560361670416360688398887362399715610156469679179519783322412828626822871102945459121862886688183120089056253680160686807782589597959635924385513244265493473052455290097829084856286619149873664044384956816329425752455857651965747999326881750999934060606191124799854050781429;
            6'd7: xpb[84] = 1024'd96408894870459406162834004477282848944538353340043417153390565310497694405432815527775592411924579116200541188012617881269878443020510159658155981023523115901969643381170448006037158174995252848082871382198472306728449149889424180609946047331534952742970577862392175553046464178911176210076093904267324992389;
            6'd8: xpb[84] = 1024'd3838712122703828701411210198482313584016609137990461779761913156302883317086812966016330286778655296135061865622283206097806357016679895704898156870028383087659014233133754288930832892979826922400255058180619910805918299684287543869956708650414703763263600344919293749104649283959658796842373182055004719018;
            6'd9: xpb[84] = 1024'd35335225059072992638787343324496210968193292061673190534265116067084967566049949314272139376290405785512731950689441965504798111854069966306800457732864691207039059654668277909454746802481606718027836342550007361247748299700047680094945939652523904050376526241563469975269362462936774400727342286468278929978;
            6'd10: xpb[84] = 1024'd66831737995442156576163476450510108352369974985355919288768318977867051815013085662527948465802156274890402035756600724911789866691460036908702758595700999326419105076202801529978660711983386513655417626919394811689578299715807816319935170654633104337489452138207646201434075641913890004612311390881553140938;
            6'd11: xpb[84] = 1024'd98328250931811320513539609576524005736546657909038648043271521888649136063976222010783757555313906764268072120823759484318781621528850107510605059458537307445799150497737325150502574621485166309282998911288782262131408299731567952544924401656742304624602378034851822427598788820891005608497280495294827351898;
            6'd12: xpb[84] = 1024'd5758068184055743052116815297723470376024913706985692669642869734454324975630219449024495430167982944202592798433424809146709535525019843557347235305042574631488521349700631433396249339469740383600382587270929866208877449526431315804935062975622055644895400517378940623656973925939488195263559773082507078527;
            6'd13: xpb[84] = 1024'd37254581120424906989492948423737367760201596630668421424146072645236409224593355797280304519679733433580262883500583568553701290362409914159249536167878882750868566771235155053920163248971520179227963871640317316650707449542191452029924293977731255932008326414023116849821687104916603799148528877495781289487;
            6'd14: xpb[84] = 1024'd68751094056794070926869081549751265144378279554351150178649275556018493473556492145536113609191483922957932968567742327960693045199799984761151837030715190870248612192769678674444077158473299974855545156009704767092537449557951588254913524979840456219121252310667293075986400283893719403033497981909055500447;
            6'd15: xpb[84] = 1024'd100247606993163234864245214675765162528554962478033878933152478466800577722519628493791922698703234412335603053634901087367684800037190055363054137893551498989628657614304202294967991067975079770483126440379092217534367449573711724479902755981949656506234178207311469302151113462870835006918467086322329711407;
            6'd16: xpb[84] = 1024'd7677424245407657402822420396964627168033218275980923559523826312605766634173625932032660573557310592270123731244566412195612714033359791409796313740056766175318028466267508577861665785959653844800510116361239821611836599368575087739913417300829407526527200689838587498209298567919317593684746364110009438036;
            6'd17: xpb[84] = 1024'd39173937181776821340198553522978524552209901199663652314027029223387850883136762280288469663069061081647793816311725171602604468870749862011698614602893074294698073887802032198385579695461433640428091400730627272053666599384335223964902648302938607813640126586482763724374011746896433197569715468523283648996;
            6'd18: xpb[84] = 1024'd70670450118145985277574686648992421936386584123346381068530232134169935132099898628544278752580811571025463901378883931009596223708139932613600915465729382414078119309336555818909493604963213436055672685100014722495496599400095360189891879305047808100753052483126939950538724925873548801454684572936557859956;
            6'd19: xpb[84] = 1024'd102166963054515149214950819775006319320563267047029109823033435044952019381063034976800087842092562060403133986446042690416587978545530003215503216328565690533458164730871079439433407514464993231683253969469402172937326599415855496414881110307157008387865978379771116176703438104850664405339653677349832070916;
            6'd20: xpb[84] = 1024'd9596780306759571753528025496205783960041522844976154449404782890757208292717032415040825716946638240337654664055708015244515892541699739262245392175070957719147535582834385722327082232449567306000637645451549777014795749210718859674891771626036759408159000862298234372761623209899146992105932955137511797545;
            6'd21: xpb[84] = 1024'd41093293243128735690904158622219681344218205768658883203907985801539292541680168763296634806458388729715324749122866774651507647379089809864147693037907265838527581004368909342850996141951347101628218929820937227456625749226478995899881002628145959695271926758942410598926336388876262595990902059550786008505;
            6'd22: xpb[84] = 1024'd72589806179497899628280291748233578728394888692341611958411188712321376790643305111552443895970139219092994834190025534058499402216479880466049993900743573957907626425903432963374910051453126897255800214190324677898455749242239132124870233630255159982384852655586586825091049567853378199875871163964060219465;
            6'd23: xpb[84] = 1024'd104086319115867063565656424874247476112571571616024340712914391623103461039606441459808252985481889708470664919257184293465491157053869951067952294763579882077287671847437956583898823960954906692883381498559712128340285749257999268349859464632364360269497778552230763051255762746830493803760840268377334430425;
            6'd24: xpb[84] = 1024'd11516136368111486104233630595446940752049827413971385339285739468908649951260438898048990860335965888405185596866849618293419071050039687114694470610085149262977042699401262866792498678939480767200765174541859732417754899052862631609870125951244111289790801034757881247313947851878976390527119546165014157054;
            6'd25: xpb[84] = 1024'd43012649304480650041609763721460838136226510337654114093788942379690734200223575246304799949847716377782855681934008377700410825887429757716596771472921457382357088120935786487316412588441260562828346458911247182859584899068622767834859356953353311576903726931402057473478661030856091994412088650578288368014;
            6'd26: xpb[84] = 1024'd74509162240849813978985896847474735520403193261336842848292145290472818449186711594560609039359466867160525767001167137107402580724819828318499072335757765501737133542470310107840326497943040358455927743280634633301414899084382904059848587955462511864016652828046233699643374209833207598297057754991562578974;
            6'd27: xpb[84] = 1024'd106005675177218977916362029973488632904579876185019571602795348201254902698149847942816418128871217356538195852068325896514394335562209898920401373198594073621117178964004833728364240407444820154083509027650022083743244899100143040284837818957571712151129578724690409925808087388810323202182026859404836789934;
            6'd28: xpb[84] = 1024'd13435492429463400454939235694688097544058131982966616229166696047060091609803845381057156003725293536472716529677991221342322249558379634967143549045099340806806549815968140011257915125429394228400892703632169687820714048895006403544848480276451463171422601207217528121866272493858805788948306137192516516563;
            6'd29: xpb[84] = 1024'd44932005365832564392315368820701994928234814906649344983669898957842175858766981729312965093237044025850386614745149980749314004395769705569045849907935648926186595237502663631781829034931174024028473988001557138262544048910766539769837711278560663458535527103861704348030985672835921392833275241605790727523;
            6'd30: xpb[84] = 1024'd76428518302201728329691501946715892312411497830332073738173101868624260107730118077568774182748794515228056699812308740156305759233159776170948150770771957045566640659037187252305742944432953819656055272370944588704374048926526675994826942280669863745648453000505880574195698851813036996718244346019064938483;
            6'd31: xpb[84] = 1024'd107925031238570892267067635072729789696588180754014802492676304779406344356693254425824583272260545004605726784879467499563297514070549846772850451633608265164946686080571710872829656853934733615283636556740332039146204048942286812219816173282779064032761378897150056800360412030790152600603213450432339149443;
            6'd32: xpb[84] = 1024'd15354848490815314805644840793929254336066436551961847119047652625211533268347251864065321147114621184540247462489132824391225428066719582819592627480113532350636056932535017155723331571919307689601020232722479643223673198737150175479826834601658815053054401379677174996418597135838635187369492728220018876072;
            6'd33: xpb[84] = 1024'd46851361427184478743020973919943151720243119475644575873550855535993617517310388212321130236626371673917917547556291583798217182904109653421494928342949840470016102354069540776247245481421087485228601517091867093665503198752910311704816065603768015340167327276321351222583310314815750791254461832633293087032;
            6'd34: xpb[84] = 1024'd78347874363553642680397107045957049104419802399327304628054058446775701766273524560576939326138122163295587632623450343205208937741499724023397229205786148589396147775604064396771159390922867280856182801461254544107333198768670447929805296605877215627280253172965527448748023493792866395139430937046567297992;
            6'd35: xpb[84] = 1024'd109844387299922806617773240171970946488596485323010033382557261357557786015236660908832748415649872652673257717690609102612200692578889794625299530068622456708776193197138588017295073300424647076483764085830641994549163198784430584154794527607986415914393179069609703674912736672769981999024400041459841508952;
            6'd36: xpb[84] = 1024'd17274204552167229156350445893170411128074741120957078008928609203362974926890658347073486290503948832607778395300274427440128606575059530672041705915127723894465564049101894300188748018409221150801147761812789598626632348579293947414805188926866166934686201552136821870970921777818464585790679319247521235581;
            6'd37: xpb[84] = 1024'd48770717488536393093726579019184308512251424044639806763431812114145059175853794695329295380015699321985448480367433186847120361412449601273944006777964032013845609470636417920712661927911000946428729046182177049068462348595054083639794419928975367221799127448780998097135634956795580189675648423660795446541;
            6'd38: xpb[84] = 1024'd80267230424905557031102712145198205896428106968322535517935015024927143424816931043585104469527449811363118565434591946254112116249839671875846307640800340133225654892170941541236575837412780742056310330551564499510292348610814219864783650931084567508912053345425174323300348135772695793560617528074069657501;
            6'd39: xpb[84] = 1024'd111763743361274720968478845271212103280604789892005264272438217935709227673780067391840913559039200300740788650501750705661103871087229742477748608503636648252605700313705465161760489746914560537683891614920951949952122348626574356089772881933193767796024979242069350549465061314749811397445586632487343868461;
            6'd40: xpb[84] = 1024'd19193560613519143507056050992411567920083045689952308898809565781514416585434064830081651433893276480675309328111416030489031785083399478524490784350141915438295071165668771444654164464899134612001275290903099554029591498421437719349783543252073518816318001724596468745523246419798293984211865910275023595090;
            6'd41: xpb[84] = 1024'd50690073549888307444432184118425465304259728613635037653312768692296500834397201178337460523405026970052979413178574789896023539920789549126393085212978223557675116587203295065178078374400914407628856575272487004471421498437197855574772774254182719103430927621240644971687959598775409588096835014688297806050;
            6'd42: xpb[84] = 1024'd82186586486257471381808317244439362688436411537317766407815971603078585083360337526593269612916777459430649498245733549303015294758179619728295386075814531677055162008737818685701992283902694203256437859641874454913251498452957991799762005256291919390543853517884821197852672777752525191981804119101572017010;
            6'd43: xpb[84] = 1024'd113683099422626635319184450370453260072613094461000495162319174513860669332323473874849078702428527948808319583312892308710007049595569690330197686938650839796435207430272342306225906193404473998884019144011261905355081498468718128024751236258401119677656779414528997424017385956729640795866773223514846227970;
            6'd44: xpb[84] = 1024'd21112916674871057857761656091652724712091350258947539788690522359665858243977471313089816577282604128742840260922557633537934963591739426376939862785156106982124578282235648589119580911389048073201402819993409509432550648263581491284761897577280870697949801897056115620075571061778123382633052501302525954599;
            6'd45: xpb[84] = 1024'd52609429611240221795137789217666622096268033182630268543193725270447942492940607661345625666794354618120510345989716392944926718429129496978842163647992415101504623703770172209643494820890827868828984104362796959874380648279341627509751128579390070985062727793700291846240284240755238986518021605715800165559;
            6'd46: xpb[84] = 1024'd84105942547609385732513922343680519480444716106312997297696928181230026741903744009601434756306105107498180431056875152351918473266519567580744464510828723220884669125304695830167408730392607664456565388732184410316210648295101763734740359581499271272175653690344468072404997419732354590402990710129074376519;
            6'd47: xpb[84] = 1024'd115602455483978549669890055469694416864621399029995726052200131092012110990866880357857243845817855596875850516124033911758910228103909638182646765373665031340264714546839219450691322639894387460084146673101571860758040648310861899959729590583608471559288579586988644298569710598709470194287959814542348587479;
            6'd48: xpb[84] = 1024'd23032272736222972208467261190893881504099654827942770678571478937817299902520877796097981720671931776810371193733699236586838142100079374229388941220170298525954085398802525733584997357878961534401530349083719464835509798105725263219740251902488222579581602069515762494627895703757952781054239092330028314108;
            6'd49: xpb[84] = 1024'd54528785672592136145843394316907778888276337751625499433074681848599384151484014144353790810183682266188041278800857995993829896937469444831291242083006606645334130820337049354108911267380741330029111633453106915277339798121485399444729482904597422866694527966159938720792608882735068384939208196743302525068;
            6'd50: xpb[84] = 1024'd86025298608961300083219527442921676272453020675308228187577884759381468400447150492609599899695432755565711363868016755400821651774859515433193542945842914764714176241871572974632825176882521125656692917822494365719169798137245535669718713906706623153807453862804114946957322061712183988824177301156576736028;
            6'd51: xpb[84] = 1024'd117521811545330464020595660568935573656629703598990956942081087670163552649410286840865408989207183244943381448935175514807813406612249586035095843808679222884094221663406096595156739086384300921284274202191881816160999798153005671894707944908815823440920379759448291173122035240689299592709146405569850946988;
            6'd52: xpb[84] = 1024'd24951628797574886559172866290135038296107959396938001568452435515968741561064284279106146864061259424877902126544840839635741320608419322081838019655184490069783592515369402878050413804368874995601657878174029420238468947947869035154718606227695574461213402241975409369180220345737782179475425683357530673617;
            6'd53: xpb[84] = 1024'd56448141733944050496548999416148935680284642320620730322955638426750825810027420627361955953573009914255572211611999599042733075445809392683740320518020798189163637936903926498574327713870654791229239162543416870680298947963629171379707837229804774748326328138619585595344933524714897783360394787770804884577;
            6'd54: xpb[84] = 1024'd87944654670313214433925132542162833064461325244303459077458841337532910058990556975617765043084760403633242296679158358449724830283199463285642621380857106308543683358438450119098241623372434586856820446912804321122128947979389307604697068231913975035439254035263761821509646703692013387245363892184079095537;
            6'd55: xpb[84] = 1024'd119441167606682378371301265668176730448638008167986187831962044248314994307953693323873574132596510893010912381746317117856716585120589533887544922243693414427923728779972973739622155532874214382484401731282191771563958947995149443829686299234023175322552179931907938047674359882669128991130332996597353306497;
            6'd56: xpb[84] = 1024'd26870984858926800909878471389376195088116263965933232458333392094120183219607690762114312007450587072945433059355982442684644499116759269934287098090198681613613099631936280022515830250858788456801785407264339375641428097790012807089696960552902926342845202414435056243732544987717611577896612274385033033126;
            6'd57: xpb[84] = 1024'd58367497795295964847254604515390092472292946889615961212836595004902267468570827110370121096962337562323103144423141202091636253954149340536189398953034989732993145053470803643039744160360568252429366691633726826083258097805772943314686191555012126629958128311079232469897258166694727181781581378798307244086;
            6'd58: xpb[84] = 1024'd89864010731665128784630737641403989856469629813298689967339797915684351717533963458625930186474088051700773229490299961498628008791539411138091699815871297852373190475005327263563658069862348048056947976003114276525088097821533079539675422557121326917071054207723408696061971345671842785666550483211581455046;
            6'd59: xpb[84] = 1024'd121360523668034292722006870767417887240646312736981418721843000826466435966497099806881739275985838541078443314557458720905619763628929481739994000678707605971753235896539850884087571979364127843684529260372501726966918097837293215764664653559230527204183980104367584922226684524648958389551519587624855666006;
            6'd60: xpb[84] = 1024'd28790340920278715260584076488617351880124568534928463348214348672271624878151097245122477150839914721012963992167124045733547677625099217786736176525212873157442606748503157166981246697348701918001912936354649331044387247632156579024675314878110278224477002586894703118284869629697440976317798865412535392635;
            6'd61: xpb[84] = 1024'd60286853856647879197960209614631249264301251458611192102717551583053709127114233593378286240351665210390634077234282805140539432462489288388638477388049181276822652170037680787505160606850481713629494220724036781486217247647916715249664545880219478511589928483538879344449582808674556580202767969825809603595;
            6'd62: xpb[84] = 1024'd91783366793017043135336342740645146648477934382293920857220754493835793376077369941634095329863415699768304162301441564547531187299879358990540778250885489396202697591572204408029074516352261509257075505093424231928047247663676851474653776882328678798702854380183055570614295987651672184087737074239083814555;
            6'd63: xpb[84] = 1024'd123279879729386207072712475866659044032654617305976649611723957404617877625040506289889904419375166189145974247368600323954522942137269429592443079113721797515582743013106728028552988425854041304884656789462811682369877247679436987699643007884437879085815780276827231796779009166628787787972706178652358025515;
        endcase
    end

    always_comb begin
        case(flag[28][11:6])
            6'd0: xpb[85] = 1024'd0;
            6'd1: xpb[85] = 1024'd30709696981630629611289681587858508672132873103923694238095305250423066536694503728130642294229242369080494924978265648782450856133439165639185254960227064701272113865070034311446663143838615379202040465444959286447346397474300350959653669203317630106108802759354349992837194271677270374738985456440037752144;
            6'd2: xpb[85] = 1024'd61419393963261259222579363175717017344265746207847388476190610500846133073389007456261284588458484738160989849956531297564901712266878331278370509920454129402544227730140068622893326287677230758404080930889918572894692794948600701919307338406635260212217605518708699985674388543354540749477970912880075504288;
            6'd3: xpb[85] = 1024'd92129090944891888833869044763575526016398619311771082714285915751269199610083511184391926882687727107241484774934796946347352568400317496917555764880681194103816341595210102934339989431515846137606121396334877859342039192422901052878961007609952890318326408278063049978511582815031811124216956369320113256432;
            6'd4: xpb[85] = 1024'd122838787926522518445158726351434034688531492415694776952381221001692266146778014912522569176916969476321979699913062595129803424533756662556741019840908258805088455460280137245786652575354461516808161861779837145789385589897201403838614676813270520424435211037417399971348777086709081498955941825760151008576;
            6'd5: xpb[85] = 1024'd29481789224028406657649480534478110615965938393882787062344671187138437346163379730638140256488537535959325217433834809333190439825975493640766149784804282572669894755778954219603076527675871174700004718837556585872371137150604981833289776333358701263724110382654691934079443284457718856576237455574594276389;
            6'd6: xpb[85] = 1024'd60191486205659036268939162122336619288098811497806481300439976437561503882857883458768782550717779905039820142412100458115641295959414659279951404745031347273942008620848988531049739671514486553902045184282515872319717534624905332792943445536676331369832913142009041926916637556134989231315222912014632028533;
            6'd7: xpb[85] = 1024'd90901183187289665880228843710195127960231684601730175538535281687984570419552387186899424844947022274120315067390366106898092152092853824919136659705258411975214122485919022842496402815353101933104085649727475158767063932099205683752597114739993961475941715901363391919753831827812259606054208368454669780677;
            6'd8: xpb[85] = 1024'd121610880168920295491518525298053636632364557705653869776630586938407636956246890915030067139176264643200809992368631755680543008226292990558321914665485476676486236350989057153943065959191717312306126115172434445214410329573506034712250783943311591582050518660717741912591026099489529980793193824894707532821;
            6'd9: xpb[85] = 1024'd28253881466426183704009279481097712559799003683841879886594037123853808155632255733145638218747832702838155509889403969883930023518511821642347044609381500444067675646487874127759489911513126970197968972230153885297395876826909612706925883463399772421339418005955033875321692297238167338413489454709150800634;
            6'd10: xpb[85] = 1024'd58963578448056813315298961068956221231931876787765574124689342374276874692326759461276280512977075071918650434867669618666380879651950987281532299569608565145339789511557908439206153055351742349400009437675113171744742274301209963666579552666717402527448220765309383868158886568915437713152474911149188552778;
            6'd11: xpb[85] = 1024'd89673275429687442926588642656814729904064749891689268362784647624699941229021263189406922807206317440999145359845935267448831735785390152920717554529835629846611903376627942750652816199190357728602049903120072458192088671775510314626233221870035032633557023524663733860996080840592708087891460367589226304922;
            6'd12: xpb[85] = 1024'd120382972411318072537878324244673238576197622995612962600879952875123007765715766917537565101435559810079640284824200916231282591918829318559902809490062694547884017241697977062099479343028973107804090368565031744639435069249810665585886891073352662739665826284018083853833275112269978462630445824029264057066;
            6'd13: xpb[85] = 1024'd27025973708823960750369078427717314503632068973800972710843403060569178965101131735653136181007127869716985802344973130434669607211048149643927939433958718315465456537196794035915903295350382765695933225622751184722420616503214243580561990593440843578954725629255375816563941310018615820250741453843707324879;
            6'd14: xpb[85] = 1024'd57735670690454590361658760015575823175764942077724666948938708310992245501795635463783778475236370238797480727323238779217120463344487315283113194394185783016737570402266828347362566439188998144897973691067710471169767013977514594540215659796758473685063528388609725809401135581695886194989726910283745077023;
            6'd15: xpb[85] = 1024'd88445367672085219972948441603434331847897815181648361187034013561415312038490139191914420769465612607877975652301504427999571319477926480922298449354412847718009684267336862658809229583027613524100014156512669757617113411451814945499869329000076103791172331147964075802238329853373156569728712366723782829167;
            6'd16: xpb[85] = 1024'd119155064653715849584238123191292840520030688285572055425129318811838378575184642920045063063694854976958470577279770076782022175611365646561483704314639912419281798132406896970255892726866228903302054621957629044064459808926115296459522998203393733897281133907318425795075524125050426944467697823163820581311;
            6'd17: xpb[85] = 1024'd25798065951221737796728877374336916447465134263760065535092768997284549774570007738160634143266423036595816094800542290985409190903584477645508834258535936186863237427905713944072316679187638561193897479015348484147445356179518874454198097723481914736570033252555717757806190322799064302087993452978263849124;
            6'd18: xpb[85] = 1024'd56507762932852367408018558962195425119598007367683759773188074247707616311264511466291276437495665405676311019778807939767860047037023643284694089218763000888135351292975748255518979823026253940395937944460307770594791753653819225413851766926799544842678836011910067750643384594476334676826978909418301601268;
            6'd19: xpb[85] = 1024'd87217459914482997019308240550053933791730880471607454011283379498130682847959015194421918731724907774756805944757073588550310903170462808923879344178990065589407465158045782566965642966864869319597978409905267057042138151128119576373505436130117174948787638771264417743480578866153605051565964365858339353412;
            6'd20: xpb[85] = 1024'd117927156896113626630597922137912442463863753575531148249378684748553749384653518922552561025954150143837300869735339237332761759303901974563064599139217130290679579023115816878412306110703484698800018875350226343489484548602419927333159105333434805054896441530618767736317773137830875426304949822298377105556;
            6'd21: xpb[85] = 1024'd24570158193619514843088676320956518391298199553719158359342134933999920584038883740668132105525718203474646387256111451536148774596120805647089729083113154058261018318614633852228730063024894356691861732407945783572470095855823505327834204853522985894185340875856059699048439335579512783925245452112820373369;
            6'd22: xpb[85] = 1024'd55279855175250144454378357908815027063431072657642852597437440184422987120733387468798774399754960572555141312234377100318599630729559971286274984043340218759533132183684668163675393206863509735893902197852905070019816493330123856287487874056840616000294143635210409691885633607256783158664230908552858125513;
            6'd23: xpb[85] = 1024'd85989552156880774065668039496673535735563945761566546835532745434846053657427891196929416693984202941635636237212642749101050486862999136925460239003567283460805246048754702475122056350702125115095942663297864356467162890804424207247141543260158246106402946394564759684722827878934053533403216364992895877657;
            6'd24: xpb[85] = 1024'd116699249138511403676957721084532044407696818865490241073628050685269120194122394925060058988213445310716131162190908397883501342996438302564645493963794348162077359913824736786568719494540740494297983128742823642914509288278724558206795212463475876212511749153919109677560022150611323908142201821432933629801;
            6'd25: xpb[85] = 1024'd23342250436017291889448475267576120335131264843678251183591500870715291393507759743175630067785013370353476679711680612086888358288657133648670623907690371929658799209323553760385143446862150152189825985800543082997494835532128136201470311983564057051800648499156401640290688348359961265762497451247376897614;
            6'd26: xpb[85] = 1024'd54051947417647921500738156855434629007264137947601945421686806121138357930202263471306272362014255739433971604689946260869339214422096299287855878867917436630930913074393588071831806590700765531391866451245502369444841233006428487161123981186881687157909451258510751633127882620037231640501482907687414649758;
            6'd27: xpb[85] = 1024'd84761644399278551112027838443293137679397011051525639659782111371561424466896767199436914656243498108514466529668211909651790070555535464927041133828144501332203026939463622383278469734539380910593906916690461655892187630480728838120777650390199317264018254017865101625965076891714502015240468364127452401902;
            6'd28: xpb[85] = 1024'd115471341380909180723317520031151646351529884155449333897877416621984491003591270927567556950472740477594961454646477558434240926688974630566226388788371566033475140804533656694725132878377996289795947382135420942339534027955029189080431319593516947370127056777219451618802271163391772389979453820567490154046;
            6'd29: xpb[85] = 1024'd22114342678415068935808274214195722278964330133637344007840866807430662202976635745683128030044308537232306972167249772637627941981193461650251518732267589801056580100032473668541556830699405947687790239193140382422519575208432767075106419113605128209415956122456743581532937361140409747599749450381933421859;
            6'd30: xpb[85] = 1024'd52824039660045698547097955802054230951097203237561038245936172057853728739671139473813770324273550906312801897145515421420078798114632627289436773692494654502328693965102507979988219974538021326889830704638099668869865972682733118034760088316922758315524758881811093574370131632817680122338734906821971174003;
            6'd31: xpb[85] = 1024'd83533736641676328158387637389912739623230076341484732484031477308276795276365643201944412618502793275393296822123781070202529654248071792928622028652721719203600807830172542291434883118376636706091871170083058955317212370157033468994413757520240388421633561641165443567207325904494950497077720363262008926147;
            6'd32: xpb[85] = 1024'd114243433623306957769677318977771248295362949445408426722126782558699861813060146930075054912732035644473791747102046718984980510381510958567807283612948783904872921695242576602881546262215252085293911635528018241764558767631333819954067426723558018527742364400519793560044520176172220871816705819702046678291;
            6'd33: xpb[85] = 1024'd20886434920812845982168073160815324222797395423596436832090232744146033012445511748190625992303603704111137264622818933188367525673729789651832413556844807672454360990741393576697970214536661743185754492585737681847544314884737397948742526243646199367031263745757085522775186373920858229437001449516489946104;
            6'd34: xpb[85] = 1024'd51596131902443475593457754748673832894930268527520131070185537994569099549140015476321268286532846073191632189601084581970818381807168955291017668517071872373726474855811427888144633358375277122387794958030696968294890712359037748908396195446963829473140066505111435515612380645598128604175986905956527698248;
            6'd35: xpb[85] = 1024'd82305828884074105204747436336532341567063141631443825308280843244992166085834519204451910580762088442272127114579350230753269237940608120930202923477298937074998588720881462199591296502213892501589835423475656254742237109833338099868049864650281459579248869264465785508449574917275398978914972362396565450392;
            6'd36: xpb[85] = 1024'd113015525865704734816037117924390850239196014735367519546376148495415232622529022932582552874991330811352622039557615879535720094074047286569388178437526001776270702585951496511037959646052507880791875888920615541189583507307638450827703533853599089685357672023820135501286769188952669353653957818836603202536;
            6'd37: xpb[85] = 1024'd19658527163210623028527872107434926166630460713555529656339598680861403821914387750698123954562898870989967557078388093739107109366266117653413308381422025543852141881450313484854383598373917538683718745978334981272569054561042028822378633373687270524646571369057427464017435386701306711274253448651046470349;
            6'd38: xpb[85] = 1024'd50368224144841252639817553695293434838763333817479223894434903931284470358608891478828766248792141240070462482056653742521557965499705283292598563341649090245124255746520347796301046742212532917885759211423294267719915452035342379782032302577004900630755374128411777456854629658378577086013238905091084222493;
            6'd39: xpb[85] = 1024'd81077921126471882251107235283151943510896206921402918132530209181707536895303395206959408543021383609150957407034919391304008821633144448931783818301876154946396369611590382107747709886051148297087799676868253554167261849509642730741685971780322530736864176887766127449691823930055847460752224361531121974637;
            6'd40: xpb[85] = 1024'd111787618108102511862396916871010452183029080025326612370625514432130603431997898935090050837250625978231452332013185040086459677766583614570969073262103219647668483476660416419194373029889763676289840142313212840614608246983943081701339640983640160842972979647120477442529018201733117835491209817971159726781;
            6'd41: xpb[85] = 1024'd18430619405608400074887671054054528110463526003514622480588964617576774631383263753205621916822194037868797849533957254289846693058802445654994203205999243415249922772159233393010796982211173334181682999370932280697593794237346659696014740503728341682261878992357769405259684399481755193111505447785602994594;
            6'd42: xpb[85] = 1024'd49140316387239029686177352641913036782596399107438316718684269867999841168077767481336264211051436406949292774512222903072297549192241611294179458166226308116522036637229267704457460126049788713383723464815891567144940191711647010655668409707045971788370681751712119398096878671159025567850490904225640746738;
            6'd43: xpb[85] = 1024'd79850013368869659297467034229771545454729272211362010956779575118422907704772271209466906505280678776029787699490488551854748405325680776933364713126453372817794150502299302015904123269888404092585763930260850853592286589185947361615322078910363601894479484511066469390934072942836295942589476360665678498882;
            6'd44: xpb[85] = 1024'd110559710350500288908756715817630054126862145315285705194874880368845974241466774937597548799509921145110282624468754200637199261459119942572549968086680437519066264367369336327350786413727019471787804395705810140039632986660247712574975748113681232000588287270420819383771267214513566317328461817105716251026;
            6'd45: xpb[85] = 1024'd17202711648006177121247470000674130054296591293473715304838330554292145440852139755713119879081489204747628141989526414840586276751338773656575098030576461286647703662868153301167210366048429129679647252763529580122618533913651290569650847633769412839877186615658111346501933412262203674948757446920159518839;
            6'd46: xpb[85] = 1024'd47912408629636806732537151588532638726429464397397409542933635804715211977546643483843762173310731573828123066967792063623037132884777939295760352990803525987919817527938187612613873509887044508881687718208488866569964931387951641529304516837087042945985989375012461339339127683939474049687742903360197270983;
            6'd47: xpb[85] = 1024'd78622105611267436343826833176391147398562337501321103781028941055138278514241147211974404467539973942908617991946057712405487989018217104934945607951030590689191931393008221924060536653725659888083728183653448153017311328862251992488958186040404673052094792134366811332176321955616744424426728359800235023127;
            6'd48: xpb[85] = 1024'd109331802592898065955116514764249656070695210605244798019124246305561345050935650940105046761769216311989112916924323361187938845151656270574130862911257655390464045258078256235507199797564275267285768649098407439464657726336552343448611855243722303158203594893721161325013516227294014799165713816240272775271;
            6'd49: xpb[85] = 1024'd15974803890403954167607268947293731998129656583432808129087696491007516250321015758220617841340784371626458434445095575391325860443875101658155992855153679158045484553577073209323623749885684925177611506156126879547643273589955921443286954763810483997492494238958453287744182425042652156786009446054716043084;
            6'd50: xpb[85] = 1024'd46684500872034583778896950535152240670262529687356502367183001741430582787015519486351260135570026740706953359423361224173776716577314267297341247815380743859317598418647107520770286893724300304379651971601086165994989671064256272402940623967128114103601296998312803280581376696719922531524994902494753795228;
            6'd51: xpb[85] = 1024'd77394197853665213390186632123010749342395402791280196605278306991853649323710023214481902429799269109787448284401626872956227572710753432936526502775607808560589712283717141832216950037562915683581692437046045452442336068538556623362594293170445744209710099757667153273418570968397192906263980358934791547372;
            6'd52: xpb[85] = 1024'd108103894835295843001476313710869258014528275895203890843373612242276715860404526942612544724028511478867943209379892521738678428844192598575711757735834873261861826148787176143663613181401531062783732902491004738889682466012856974322247962373763374315818902517021503266255765240074463281002965815374829299516;
            6'd53: xpb[85] = 1024'd14746896132801731213967067893913333941962721873391900953337062427722887059789891760728115803600079538505288726900664735942065444136411429659736887679730897029443265444285993117480037133722940720675575759548724178972668013266260552316923061893851555155107801862258795228986431437823100638623261445189272567329;
            6'd54: xpb[85] = 1024'd45456593114432360825256749481771842614095594977315595191432367678145953596484395488858758097829321907585783651878930384724516300269850595298922142639957961730715379309356027428926700277561556099877616224993683465420014410740560903276576731097169185261216604621613145221823625709500371013362246901629310319473;
            6'd55: xpb[85] = 1024'd76166290096062990436546431069630351286228468081239289429527672928569020133178899216989400392058564276666278576857196033506967156403289760938107397600185026431987493174426061740373363421400171479079656690438642751867360808214861254236230400300486815367325407380967495214660819981177641388101232358069348071617;
            6'd56: xpb[85] = 1024'd106875987077693620047836112657488859958361341185162983667622978178992086669873402945120042686287806645746773501835461682289418012536728926577292652560412091133259607039496096051820026565238786858281697155883602038314707205689161605195884069503804445473434210140321845207498014252854911762840217814509385823761;
            6'd57: xpb[85] = 1024'd13518988375199508260326866840532935885795787163350993777586428364438257869258767763235613765859374705384119019356233896492805027828947757661317782504308114900841046334994913025636450517560196516173540012941321478397692752942565183190559169023892626312723109485559137170228680450603549120460513444323829091574;
            6'd58: xpb[85] = 1024'd44228685356830137871616548428391444557928660267274688015681733614861324405953271491366256060088617074464613944334499545275255883962386923300503037464535179602113160200064947337083113661398811895375580478386280764845039150416865534150212838227210256418831912244913487163065874722280819495199498900763866843718;
            6'd59: xpb[85] = 1024'd74938382338460767482906230016249953230061533371198382253777038865284390942647775219496898354317859443545108869312765194057706740095826088939688292424762244303385274065134981648529776805237427274577620943831240051292385547891165885109866507430527886524940715004267837155903068993958089869938484357203904595862;
            6'd60: xpb[85] = 1024'd105648079320091397094195911604108461902194406475122076491872344115707457479342278947627540648547101812625603794291030842840157596229265254578873547384989309004657387930205015959976439949076042653779661409276199337739731945365466236069520176633845516631049517763622187148740263265635360244677469813643942348006;
            6'd61: xpb[85] = 1024'd12291080617597285306686665787152537829628852453310086601835794301153628678727643765743111728118669872262949311811803057043544611521484085662898677328885332772238827225703832933792863901397452311671504266333918777822717492618869814064195276153933697470338417108859479111470929463383997602297765443458385615819;
            6'd62: xpb[85] = 1024'd43000777599227914917976347375011046501761725557233780839931099551576695215422147493873754022347912241343444236790068705825995467654923251302083932289112397473510941090773867245239527045236067690873544731778878064270063890093170165023848945357251327576447219868213829104308123735061267977036750899898423367963;
            6'd63: xpb[85] = 1024'd73710474580858544529266028962869555173894598661157475078026404801999761752116651222004396316577154610423939161768334354608446323788362416941269187249339462174783054955843901556686190189074683070075585197223837350717410287567470515983502614560568957682556022627568179097145318006738538351775736356338461120107;
        endcase
    end

    always_comb begin
        case(flag[28][16:12])
            5'd0: xpb[86] = 1024'd0;
            5'd1: xpb[86] = 1024'd104420171562489174140555710550728063846027471765081169316121710052422828288811154950135038610806396979504434086746600003390897179921801582580454442209566526876055168820913935868132853332913298449277625662668796637164756685041770866943156283763886587788664825386922529089982512278415808726514721812778498872251;
            5'd2: xpb[86] = 1024'd84773647440853606882312493696641694947356516404426654504111565039868761240313170990255006006955119649565718766035706572202730519002382830605748759402802012818419663072256654398635467474309391177245053716950353427965152519862644960921333997844543726310509747359728000149858496482902984435910753798931403260171;
            5'd3: xpb[86] = 1024'd65127123319218039624069276842555326048685561043772139692101420027314694191815187030374973403103842319627003445324813141014563858082964078631043076596037498760784157323599372929138081615705483905212481771231910218765548354683519054899511711925200864832354669332533471209734480687390160145306785785084307648091;
            5'd4: xpb[86] = 1024'd45480599197582472365826059988468957150014605683117624880091275014760627143317203070494940799252564989688288124613919709826397197163545326656337393789272984703148651574942091459640695757101576633179909825513467009565944189504393148877689426005858003354199591305338942269610464891877335854702817771237212036011;
            5'd5: xpb[86] = 1024'd25834075075946905107582843134382588251343650322463110068081130002206560094819219110614908195401287659749572803903026278638230536244126574681631710982508470645513145826284809990143309898497669361147337879795023800366340024325267242855867140086515141876044513278144413329486449096364511564098849757390116423931;
            5'd6: xpb[86] = 1024'd6187550954311337849339626280296219352672694961808595256070984989652493046321235150734875591550010329810857483192132847450063875324707822706926028175743956587877640077627528520645924039893762089114765934076580591166735859146141336834044854167172280397889435250949884389362433300851687273494881743543020811851;
            5'd7: xpb[86] = 1024'd110607722516800511989895336831024283198700166726889764572192695042075321335132390100869914202356407309315291569938732850840961055246509405287380470385310483463932808898541464388778777372807060538392391596745377228331492544187912203777201137931058868186554260637872413479344945579267496000009603556321519684102;
            5'd8: xpb[86] = 1024'd90961198395164944731652119976937914300029211366235249760182550029521254286634406140989881598505129979376576249227839419652794394327090653312674787578545969406297303149884182919281391514203153266359819651026934019131888379008786297755378852011716006708399182610677884539220929783754671709405635542474424072022;
            5'd9: xpb[86] = 1024'd71314674273529377473408903122851545401358256005580734948172405016967187238136422181109848994653852649437860928516945988464627733407671901337969104771781455348661797401226901449784005655599245994327247705308490809932284213829660391733556566092373145230244104583483355599096913988241847418801667528627328459942;
            5'd10: xpb[86] = 1024'd51668150151893810215165686268765176502687300644926220136162260004413120189638438221229816390802575319499145607806052557276461072488253149363263421965016941291026291652569619980286619796995338722294675759590047600732680048650534485711734280173030283752089026556288826658972898192729023128197699514780232847862;
            5'd11: xpb[86] = 1024'd32021626030258242956922469414678807604016345284271705324152114991859053141140454261349783786951297989560430287095159126088294411568834397388557739158252427233390785903912338510789233938391431450262103813871604391533075883471408579689911994253687422273933948529094297718848882397216198837593731500933137235782;
            5'd12: xpb[86] = 1024'd12375101908622675698679252560592438705345389923617190512141969979304986092642470301469751183100020659621714966384265694900127750649415645413852056351487913175755280155255057041291848079787524178229531868153161182333471718292282673668089708334344560795778870501899768778724866601703374546989763487086041623702;
            5'd13: xpb[86] = 1024'd116795273471111849839234963111320502551372861688698359828263680031727814381453625251604789793906417639126149053130865698291024930571217227994306498561054440051810448976168992909424701412700822627507157530821957819498228403334053540611245992098231148584443695888822297868707378880119183273504485299864540495953;
            5'd14: xpb[86] = 1024'd97148749349476282580991746257234133652701906328043845016253535019173747332955641291724757190055140309187433732419972267102858269651798476019600815754289925994174943227511711439927315554096915355474585585103514610298624238154927634589423706178888287106288617861627768928583363084606358982900517286017444883873;
            5'd15: xpb[86] = 1024'd77502225227840715322748529403147764754030950967389330204243390006619680284457657331844724586203862979248718411709078835914691608732379724044895132947525411936539437478854429970429929695493008083442013639385071401099020072975801728567601420259545425628133539834433239988459347289093534692296549272170349271793;
            5'd16: xpb[86] = 1024'd57855701106205148064505312549061395855359995606734815392233244994065613235959673371964691982352585649310003090998185404726524947812960972070189450140760897878903931730197148500932543836889100811409441693666628191899415907796675822545779134340202564149978461807238711048335331493580710401692581258323253659713;
            5'd17: xpb[86] = 1024'd38209176984569580806262095694975026956689040246080300580223099981511546187461689412084659378501308319371287770287291973538358286893542220095483767333996383821268425981539867031435157978285193539376869747948184982699811742617549916523956848420859702671823383780044182108211315698067886111088613244476158047633;
            5'd18: xpb[86] = 1024'd18562652862934013548018878840888658058018084885425785768212954968957479138963705452204626774650030989432572449576398542350191625974123468120778084527231869763632920232882585561937772119681286267344297802229741773500207577438424010502134562501516841193668305752849653168087299902555061820484645230629062435553;
            5'd19: xpb[86] = 1024'd122982824425423187688574589391616721904045556650506955084334665021380307427774860402339665385456427968937006536322998545741088805895925050701232526736798396639688089053796521430070625452594584716621923464898538410664964262480194877445290846265403428982333131139772182258069812180970870546999367043407561307804;
            5'd20: xpb[86] = 1024'd103336300303787620430331372537530353005374601289852440272324520008826240379276876442459632781605150638998291215612105114552922144976506298726526843930033882582052583305139239960573239593990677444589351519180095201465360097301068971423468560346060567504178053112577653317945796385458046256395399029560465695724;
            5'd21: xpb[86] = 1024'd83689776182152053172088155683443984106703645929197925460314374996272173330778892482579600177753873309059575894901211683364755484057087546751821161123269368524417077556481958491075853735386770172556779573461651992265755932121943065401646274426717706026022975085383124377821780589945221965791431015713370083644;
            5'd22: xpb[86] = 1024'd64043252060516485913844938829357615208032690568543410648304229983718106282280908522699567573902595979120860574190318252176588823137668794777115478316504854466781571807824677021578467876782862900524207627743208783066151766942817159379823988507374844547867897058188595437697764794432397675187463001866274471564;
            5'd23: xpb[86] = 1024'd44396727938880918655601721975271246309361735207888895836294084971164039233782924562819534970051318649182145253479424820988422162218250042802409795509740340409146066059167395552081082018178955628491635682024765573866547601763691253358001702588031983069712819030994066497573748998919573384583494988019178859484;
            5'd24: xpb[86] = 1024'd24750203817245351397358505121184877410690779847234381024283939958609972185284940602939502366200041319243429932768531389800255501298831290827704112702975826351510560310510114082583696159575048356459063736306322364666943436584565347336179416668689121591557741003799537557449733203406749093979526974172083247404;
            5'd25: xpb[86] = 1024'd5103679695609784139115288267098508512019824486579866212273794946055905136786956643059469762348763989304714612057637958612088840379412538852998429896211312293875054561852832613086310300971141084426491790587879155467339271405439441314357130749346260113402662976605008617325717407893924803375558960324987635324;
            5'd26: xpb[86] = 1024'd109523851258098958279670998817826572358047296251661035528395504998478733425598111593194508373155160968809148698804237962002986020301214121433452872105777839169930223382766768481219163633884439533704117453256675792632095956447210308257513414513232847902067488363527537707308229686309733529890280773103486507575;
            5'd27: xpb[86] = 1024'd89877327136463391021427781963740203459376340891006520716385359985924666377100127633314475769303883638870433378093344530814819359381795369458747189299013325112294717634109487011721777775280532261671545507538232583432491791268084402235691128593889986423912410336333008767184213890796909239286312759256390895495;
            5'd28: xpb[86] = 1024'd70230803014827823763184565109653834560705385530352005904375214973370599328602143673434443165452606308931718057382451099626652698462376617484041506492248811054659211885452205542224391916676624989638973561819789374232887626088958496213868842674547124945757332309138479827060198095284084948682344745409295283415;
            5'd29: xpb[86] = 1024'd50584278893192256504941348255567465662034430169697491092365069960816532280104159713554410561601328978993002736671557668438486037542957865509335823685484296997023706136794924072727006058072717717606401616101346165033283460909832590192046556755204263467602254281943950886936182299771260658078376731562199671335;
            5'd30: xpb[86] = 1024'd30937754771556689246698131401481096763363474809042976280354924948262465231606175753674377957750051649054287415960664237250319376623539113534630140878719782939388200388137642603229620199468810445573829670382902955833679295730706684170224270835861401989447176254749421946812166504258436367474408717715104059255;
            5'd31: xpb[86] = 1024'd11291230649921121988454914547394727864692519448388461468344779935708398183108191793794345353898774319115572095249770806062152715704120361559924458071955268881752694639480361133732234340864903173541257724664459746634075130551580778148401984916518540511292098227554893006688150708745612076870440703868008447175;
        endcase
    end

    always_comb begin
        case(flag[29][5:0])
            6'd0: xpb[87] = 1024'd0;
            6'd1: xpb[87] = 1024'd57855701106205148064505312549061395855359995606734815392233244994065613235959673371964691982352585649310003090998185404726524947812960972070189450140760897878903931730197148500932543836889100811409441693666628191899415907796675822545779134340202564149978461807238711048335331493580710401692581258323253659713;
            6'd2: xpb[87] = 1024'd115711402212410296129010625098122791710719991213469630784466489988131226471919346743929383964705171298620006181996370809453049895625921944140378900281521795757807863460394297001865087673778201622818883387333256383798831815593351645091558268680405128299956923614477422096670662987161420803385162516646507319426;
            6'd3: xpb[87] = 1024'd49500407634490702794717010242369754821381559694468762048567879917219944370569881205879004732400082638486859865537062779600511002597662581655408225405951652703021120621020228165167392319150096712918127472612644729333886873169130694672358833337378243183115482007599075114899466406813498187959053948344166494808;
            6'd4: xpb[87] = 1024'd107356108740695850859222322791431150676741555301203577440801124911285557606529554577843696714752668287796862956535248184327035950410623553725597675546712550581925052351217376666099936156039197524327569166279272921233302780965806517218137967677580807333093943814837786163234797900394208589651635206667420154521;
            6'd5: xpb[87] = 1024'd41145114162776257524928707935678113787403123782202708704902514840374275505180089039793317482447579627663716640075940154474497057382364191240627000671142407527138309511843307829402240801411092614426813251558661266768357838541585566798938532334553922216252502207959439181463601320046285974225526638365079329903;
            6'd6: xpb[87] = 1024'd99000815268981405589434020484739509642763119388937524097135759834439888741139762411758009464800165276973719731074125559201022005195325163310816450811903305406042241242040456330334784638300193425836254945225289458667773746338261389344717666674756486366230964015198150229798932813626996375918107896688332989616;
            6'd7: xpb[87] = 1024'd32789820691061812255140405628986472753424687869936655361237149763528606639790296873707630232495076616840573414614817529348483112167065800825845775936333162351255498402666387493637089283672088515935499030504677804202828803914040438925518231331729601249389522408319803248027736233279073760491999328385992164998;
            6'd8: xpb[87] = 1024'd90645521797266960319645718178047868608784683476671470753470394757594219875749970245672322214847662266150576505613002934075008059980026772896035226077094060230159430132863535994569633120561189327344940724171305996102244711710716261471297365671932165399367984215558514296363067726859784162184580586709245824711;
            6'd9: xpb[87] = 1024'd24434527219347366985352103322294831719446251957670602017571784686682937774400504707621942982542573606017430189153694904222469166951767410411064551201523917175372687293489467157871937765933084417444184809450694341637299769286495311052097930328905280282526542608680167314591871146511861546758472018406905000093;
            6'd10: xpb[87] = 1024'd82290228325552515049857415871356227574806247564405417409805029680748551010360178079586634964895159255327433280151880308948994114764728382481254001342284815054276619023686615658804481602822185228853626503117322533536715677083171133597877064669107844432505004415918878362927202640092571948451053276730158659806;
            6'd11: xpb[87] = 1024'd16079233747632921715563801015603190685467816045404548673906419609837268909010712541536255732590070595194286963692572279096455221736469019996283326466714671999489876184312546822106786248194080318952870588396710879071770734658950183178677629326080959315663562809040531381156006059744649333024944708427817835188;
            6'd12: xpb[87] = 1024'd73934934853838069780069113564664586540827811652139364066139664603902882144970385913500947714942656244504290054690757683822980169549429992066472776607475569878393807914509695323039330085083181130362312282063339070971186642455626005724456763666283523465642024616279242429491337553325359734717525966751071494901;
            6'd13: xpb[87] = 1024'd7723940275918476445775498708911549651489380133138495330241054532991600043620920375450568482637567584371143738231449653970441276521170629581502101731905426823607065075135626486341634730455076220461556367342727416506241700031405055305257328323256638348800583009400895447720140972977437119291417398448730670283;
            6'd14: xpb[87] = 1024'd65579641382123624510280811257972945506849375739873310722474299527057213279580593747415260464990153233681146829229635058696966224334131601651691551872666324702510996805332774987274178567344177031870998061009355608405657607828080877851036462663459202498779044816639606496055472466558147520983998656771984329996;
            6'd15: xpb[87] = 1024'd123435342488328772574786123807034341362209371346608126114707544521122826515540267119379952447342738882991149920227820463423491172147092573721881002013427222581414928535529923488206722404233277843280439754675983800305073515624756700396815597003661766648757506623878317544390803960138857922676579915095237989709;
            6'd16: xpb[87] = 1024'd57224347910409179240492508951281304472870939827607257378808934450211544414190801581329573215037650222858003603768512433570952279118833211236910327137857079526628185696155854651509027049605172933379683839955372145840128573200535749977616161660634881531916065016999970562619607379790935307250471346792897165091;
            6'd17: xpb[87] = 1024'd115080049016614327304997821500342700328230935434342072771042179444277157650150474953294265197390235872168006694766697838297477226931794183307099777278617977405532117426353003152441570886494273744789125533622000337739544480997211572523395296000837445681894526824238681610954938873371645708943052605116150824804;
            6'd18: xpb[87] = 1024'd48869054438694733970704206644589663438892503915341204035143569373365875548801009415243885965085147212034860378307389808444938333903534820822129102403047834350745374586978934315743875531866168834888369618901388683274599538572990622104195860657810560565053085217360334629183742293023723093516944036813810000186;
            6'd19: xpb[87] = 1024'd106724755544899882035209519193651059294252499522076019427376814367431488784760682787208577947437732861344863469305575213171463281716495792892318552543808732229649306317176082816676419368755269646297811312568016875174015446369666444649974994998013124715031547024599045677519073786604433495209525295137063659899;
            6'd20: xpb[87] = 1024'd40513760966980288700915904337898022404914068003075150691478204296520206683411217249158198715132644201211717152846267183318924388688236430407347877668238589174862563477802013979978724014127164736397055397847405220709070503945445494230775559654986239598190105417720698695747877206256510879783416726834722835281;
            6'd21: xpb[87] = 1024'd98369462073185436765421216886959418260274063609809966083711449290585819919370890621122890697485229850521720243844452588045449336501197402477537327808999487053766495207999162480911267851016265547806497091514033412608486411742121316776554693995188803748168567224959409744083208699837221281475997985157976494994;
            6'd22: xpb[87] = 1024'd32158467495265843431127602031206381370935632090809097347812839219674537818021425083072511465180141190388573927385144558192910443472938039992566652933429343998979752368625093644213572496388160637905741176793421758143541469317900366357355258652161918631327125618081062762312012119489298666049889416855635670376;
            6'd23: xpb[87] = 1024'd90014168601470991495632914580267777226295627697543912740046084213740151053981098455037203447532726839698577018383329962919435391285899012062756103074190241877883684098822242145146116333277261449315182870460049950042957377114576188903134392992364482781305587425319773810647343613070009067742470675178889330089;
            6'd24: xpb[87] = 1024'd23803174023551398161339299724514740336957196178543044004147474142828868952631632916986824215227638179565430701924021933066896498257639649577785428198620098823096941259448173308448420978649156539414426955739438295578012434690355238483934957649337597664464145818441426828876147032722086452316362106876548505471;
            6'd25: xpb[87] = 1024'd81658875129756546225844612273576136192317191785277859396380719136894482188591306288951516197580223828875433792922207337793421446070600621647974878339380996702000872989645321809380964815538257350823868649406066487477428342487031061029714091989540161814442607625680137877211478526302796854008943365199802165184;
            6'd26: xpb[87] = 1024'd15447880551836952891550997417823099302978760266276990660482109065983200087241840750901136965275135168742287476462899307940882553042341259163004203463810853647214130150271252972683269460910152440923112734685454833012483400062810110610514656646513276697601166018801790895440281945954874238582834796897461340566;
            6'd27: xpb[87] = 1024'd73303581658042100956056309966884495158338755873011806052715354060048813323201514122865828947627720818052290567461084712667407500855302231233193653604571751526118061880468401473615813297799253252332554428352083024911899307859485933156293790986715840847579627826040501943775613439535584640275416055220715000279;
            6'd28: xpb[87] = 1024'd7092587080122507621762695111131458269000324354010937316816743989137531221852048584815449715322632157919144251001776682814868607827042868748222978729001608471331319041094332636918117943171148342431798513631471370446954365435264982737094355643688955730738186219162154962004416859187662024849307486918374175661;
            6'd29: xpb[87] = 1024'd64948288186327655686268007660192854124360319960745752709049988983203144457811721956780141697675217807229147341999962087541393555640003840818412428869762506350235250771291481137850661780060249153841240207298099562346370273231940805282873489983891519880716648026400866010339748352768372426541888745241627835374;
            6'd30: xpb[87] = 1024'd122803989292532803750773320209254249979720315567480568101283233977268757693771395328744833680027803456539150432998147492267918503452964812888601879010523404229139182501488629638783205616949349965250681900964727754245786181028616627828652624324094084030695109833639577058675079846349082828234470003564881495087;
            6'd31: xpb[87] = 1024'd56592994714613210416479705353501213090381884048479699365384623906357475592421929790694454447722714796406004116538839462415379610424705450403631204134953261174352439662114560802085510262321245055349925986244116099780841238604395677409453188981067198913853668226761230076903883266001160212808361435262540670469;
            6'd32: xpb[87] = 1024'd114448695820818358480985017902562608945741879655214514757617868900423088828381603162659146430075300445716007207537024867141904558237666422473820654275714159053256371392311709303018054099210345866759367679910744291680257146401071499955232323321269763063832130033999941125239214759581870614500942693585794330182;
            6'd33: xpb[87] = 1024'd48237701242898765146691403046809572056403448136213646021719258829511806727032137624608767197770211785582860891077716837289365665209407059988849979400144015998469628552937640466320358744582240956858611765190132637215312203976850549536032887978242877946990688427121594143468018179233947999074834125283453505564;
            6'd34: xpb[87] = 1024'd106093402349103913211196715595870967911763443742948461413952503823577419962991810996573459180122797434892863982075902242015890613022368032059039429540904913877373560283134788967252902581471341768268053458856760829114728111773526372081812022318445442096969150234360305191803349672814658400767415383606707165277;
            6'd35: xpb[87] = 1024'd39882407771184319876903100740117931022425012223947592678053893752666137861642345458523079947817708774759717665616594212163351719994108669574068754665334770822586817443760720130555207226843236858367297544136149174649783169349305421662612586975418556980127708627481958210032153092466735785341306815304366340659;
            6'd36: xpb[87] = 1024'd97738108877389467941408413289179326877785007830682408070287138746731751097602018830487771930170294424069720756614779616889876667807069641644258204806095668701490749173957868631487751063732337669776739237802777366549199077145981244208391721315621121130106170434720669258367484586047446187033888073627620000372;
            6'd37: xpb[87] = 1024'd31527114299469874607114798433426289988446576311681539334388528675820468996252553292437392697865205763936574440155471587037337774778810279159287529930525525646704006334583799794790055709104232759875983323082165712084254134721760293789192285972594236013264728827842322276596288005699523571607779505325279175754;
            6'd38: xpb[87] = 1024'd89382815405675022671620110982487685843806571918416354726621773669886082232212226664402084680217791413246577531153656991763862722591771251229476980071286423525607938064780948295722599545993333571285425016748793903983670042518436116334971420312796800163243190635081033324931619499280233973300360763648532835467;
            6'd39: xpb[87] = 1024'd23171820827755429337326496126734648954468140399415485990723163598974800130862761126351705447912702753113431214694348961911323829563511888744506305195716280470821195225406879459024904191365228661384669102028182249518725100094215165915771984969769915046401749028202686343160422918932311357874252195346192010849;
            6'd40: xpb[87] = 1024'd81027521933960577401831808675796044809828136006150301382956408593040413366822434498316397430265288402423434305692534366637848777376472860814695755336477178349725126955604027959957448028254329472794110795694810441418141007890890988461551119309972479196380210835441397391495754412513021759566833453669445670562;
            6'd41: xpb[87] = 1024'd14816527356040984067538193820043007920489704487149432647057798522129131265472968960266018197960199742290287989233226336785309884348213498329725080460907035294938384116229959123259752673626224562893354880974198786953196065466670038042351683966945594079538769228563050409724557832165099144140724885367104845944;
            6'd42: xpb[87] = 1024'd72672228462246132132043506369104403775849700093884248039291043516194744501432642332230710180312785391600291080231411741511834832161174470399914530601667933173842315846427107624192296510515325374302796574640826978852611973263345860588130818307148158229517231035801761458059889325745809545833306143690358505657;
            6'd43: xpb[87] = 1024'd6461233884326538797749891513351366886511268574883379303392433445283462400083176794180330948007696731467144763772103711659295939132915107914943855726097790119055573007053038787494601155887220464402040659920215324387667030839124910168931382964121273112675789428923414476288692745397886930407197575388017681039;
            6'd44: xpb[87] = 1024'd64316934990531686862255204062412762741871264181618194695625678439349075636042850166145022930360282380777147854770289116385820886945876079985133305866858687997959504737250187288427144992776321275811482353586843516287082938635800732714710517304323837262654251236162125524624024238978597332099778833711271340752;
            6'd45: xpb[87] = 1024'd122172636096736834926760516611474158597231259788353010087858923433414688872002523538109714912712868030087150945768474521112345834758837052055322756007619585876863436467447335789359688829665422087220924047253471708186498846432476555260489651644526401412632713043400836572959355732559307733792360092034525000465;
            6'd46: xpb[87] = 1024'd55961641518817241592466901755721121707892828269352141351960313362503406770653058000059335680407779369954004629309166491259806941730577689570352081132049442822076693628073266952661993475037317177320168132532860053721553904008255604841290216301499516295791271436522489591188159152211385118366251523732184175847;
            6'd47: xpb[87] = 1024'd113817342625022389656972214304782517563252823876086956744193558356569020006612731372024027662760365019264007720307351895986331889543538661640541531272810340700980625358270415453594537311926417988729609826199488245620969811804931427387069350641702080445769733243761200639523490645792095520058832782055437835560;
            6'd48: xpb[87] = 1024'd47606348047102796322678599449029480673914392357086088008294948285657737905263265833973648430455276359130861403848043866133792996515279299155570856397240197646193882518896346616896841957298313078828853911478876591156024869380710476967869915298675195328928291636882853657752294065444172904632724213753097010942;
            6'd49: xpb[87] = 1024'd105462049153307944387183911998090876529274387963820903400528193279723351141222939205938340412807862008440864494846229270860317944328240271225760306538001095525097814249093495117829385794187413890238295605145504783055440777177386299513649049638877759478906753444121564706087625559024883306325305472076350670655;
            6'd50: xpb[87] = 1024'd39251054575388351052890297142337839639935956444820034664629583208812069039873473667887961180502773348307718178386921241007779051299980908740789631662430952470311071409719426281131690439559308980337539690424893128590495834753165349094449614295850874362065311837243217724316428978676960690899196903774009846037;
            6'd51: xpb[87] = 1024'd97106755681593499117395609691399235495295952051554850056862828202877682275833147039852653162855358997617721269385106645734303999112941880810979081803191850349215003139916574782064234276448409791746981384091521320489911742549841171640228748636053438512043773644481928772651760472257671092591778162097263505750;
            6'd52: xpb[87] = 1024'd30895761103673905783101994835646198605957520532553981320964218131966400174483681501802273930550270337484574952925798615881765106084682518326008406927621707294428260300542505945366538921820304881846225469370909666024966800125620221221029313293026553395202332037603581790880563891909748477165669593794922681132;
            6'd53: xpb[87] = 1024'd88751462209879053847607307384707594461317516139288796713197463126032013410443354873766965912902855986794578043923984020608290053897643490396197857068382605173332192030739654446299082758709405693255667163037537857924382707922296043766808447633229117545180793844842292839215895385490458878858250852118176340845;
            6'd54: xpb[87] = 1024'd22540467631959460513313692528954557571979084620287927977298853055120731309093889335716586680597767326661431727464675990755751160869384127911227182192812462118545449191365585609601387404081300783354911248316926203459437765498075093347609012290202232428339352237963945857444698805142536263432142283815835516227;
            6'd55: xpb[87] = 1024'd80396168738164608577819005078015953427339080227022743369532098049186344545053562707681278662950352975971434818462861395482276108682345099981416632333573359997449380921562734110533931240970401594764352941983554395358853673294750915893388146630404796578317814045202656905780030298723246665124723542139089175940;
            6'd56: xpb[87] = 1024'd14185174160245015243525390222262916538000648708021874633633487978275062443704097169630899430645264315838288502003553365629737215654085737496445957458003216942662638082188665273836235886342296684863597027262942740893908730870529965474188711287377911461476372438324309924008833718375324049698614973836748351322;
            6'd57: xpb[87] = 1024'd72040875266450163308030702771324312393360644314756690025866732972340675679663770541595591412997849965148291593001738770356262163467046709566635407598764114821566569812385813774768779723231397496273038720929570932793324638667205788019967845627580475611454834245563020972344165211956034451391196232160002011035;
            6'd58: xpb[87] = 1024'd5829880688530569973737087915571275504022212795755821289968122901429393578314305003545212180692761305015145276542430740503723270438787347081664732723193971766779826973011744938071084368603292586372282806208959278328379696242984837600768410284553590494613392638684673990572968631608111835965087663857661186417;
            6'd59: xpb[87] = 1024'd63685581794735718038242400464632671359382208402490636682201367895495006814273978375509904163045346954325148367540616145230248218251748319151854182863954869645683758703208893439003628205492393397781724499875587470227795604039660660146547544624756154644591854445923385038908300125188822237657668922180914846130;
            6'd60: xpb[87] = 1024'd121541282900940866102747713013694067214742204009225452074434612889560620050233651747474596145397932603635151458538801549956773166064709291222043633004715767524587690433406041939936172042381494209191166193542215662127211511836336482692326678964958718794570316253162096087243631618769532639350250180504168505843;
            6'd61: xpb[87] = 1024'd55330288323021272768454098157941030325403772490224583338536002818649337948884186209424216913092843943502005142079493520104234273036449928737072958129145624469800947594031973103238476687753389299290410278821604007662266569412115532273127243621931833677728874646283749105472435038421610023924141612201827681225;
            6'd62: xpb[87] = 1024'd113185989429226420832959410707002426180763768096959398730769247812714951184843859581388908895445429592812008233077678924830759220849410900807262408269906522348704879324229121604171020524642490110699851972488232199561682477208791354818906377962134397827707336453522460153807766532002320425616722870525081340938;
            6'd63: xpb[87] = 1024'd46974994851306827498665795851249389291425336577958529994870637741803669083494394043338529663140340932678861916618370894978220327821151538322291733394336379293918136484855052767473325170014385200799096057767620545096737534784570404399706942619107512710865894846644113172036569951654397810190614302222740516320;
        endcase
    end

    always_comb begin
        case(flag[29][11:6])
            6'd0: xpb[88] = 1024'd0;
            6'd1: xpb[88] = 1024'd104830695957511975563171108400310785146785332184693345387103882735869282319454067415303221645492926581988865007616556299704745275634112510392481183535097277172822068215052201268405869006903486012208537751434248736996153442581246226945486076959310076860844356653882824220371901445235108211883195560545994176033;
            6'd2: xpb[88] = 1024'd85594696230899209727543289395807137548872237243651006646075910406761669301598995920591372076328178854534580607775619164830426710427004686229802242053863513411953461860533185199181498822289766303106877894481257627627946034941595680925993584235390704454868809893648590410637274816541583406647701294466393867735;
            6'd3: xpb[88] = 1024'd66358696504286443891915470391303489950959142302608667905047938077654056283743924425879522507163431127080296207934682029956108145219896862067123300572629749651084855506014169129957128637676046594005218037528266518259738627301945134906501091511471332048893263133414356600902648187848058601412207028386793559437;
            6'd4: xpb[88] = 1024'd47122696777673678056287651386799842353046047361566329164019965748546443265888852931167672937998683399626011808093744895081789580012789037904444359091395985890216249151495153060732758453062326884903558180575275408891531219662294588887008598787551959642917716373180122791168021559154533796176712762307193251139;
            6'd5: xpb[88] = 1024'd27886697051060912220659832382296194755132952420523990422991993419438830248033781436455823368833935672171727408252807760207471014805681213741765417610162222129347642796976136991508388268448607175801898323622284299523323812022644042867516106063632587236942169612945888981433394930461008990941218496227592942841;
            6'd6: xpb[88] = 1024'd8650697324448146385032013377792547157219857479481651681964021090331217230178709941743973799669187944717443008411870625333152449598573389579086476128928458368479036442457120922284018083834887466700238466669293190155116404382993496848023613339713214830966622852711655171698768301767484185705724230147992634543;
            6'd7: xpb[88] = 1024'd113481393281960121948203121778103332304005189664174997069067903826200499549632777357047195445162114526706308016028426925037897725232685899971567659664025735541301104657509322190689887090738373478908776218103541927151269846964239723793509690299023291691810979506594479392070669747002592397588919790693986810576;
            6'd8: xpb[88] = 1024'd94245393555347356112575302773599684706092094723132658328039931497092886531777705862335345875997366799252023616187489790163579160025578075808888718182791971780432498302990306121465516906124653769807116361150550817783062439324589177774017197575103919285835432746360245582336043118309067592353425524614386502278;
            6'd9: xpb[88] = 1024'd75009393828734590276947483769096037108178999782090319587011959167985273513922634367623496306832619071797739216346552655289260594818470251646209776701558208019563891948471290052241146721510934060705456504197559708414855031684938631754524704851184546879859885986126011772601416489615542787117931258534786193980;
            6'd10: xpb[88] = 1024'd55773394102121824441319664764592389510265904841047980845983986838877660496067562872911646737667871344343454816505615520414942029611362427483530835220324444258695285593952273983016776536897214351603796647244568599046647624045288085735032212127265174473884339225891777962866789860922017981882436992455185885682;
            6'd11: xpb[88] = 1024'd36537394375509058605691845760088741912352809900005642104956014509770047478212491378199797168503123616889170416664678385540623464404254603320851893739090680497826679239433257913792406352283494642502136790291577489678440216405637539715539719403345802067908792465657544153132163232228493176646942726375585577384;
            6'd12: xpb[88] = 1024'd17301394648896292770064026755585094314439714958963303363928042180662434460357419883487947599338375889434886016823741250666304899197146779158172952257856916736958072884914241844568036167669774933400476933338586380310232808765986993696047226679426429661933245705423310343397536603534968371411448460295985269086;
            6'd13: xpb[88] = 1024'd122132090606408268333235135155895879461225047143656648751031924916531716779811487298791169244831302471423751024440297550371050174831259289550654135792954193909780141099966443112973905174573260945609014684772835117306386251347233220641533303638736506522777602359306134563769438048770076583294644020841979445119;
            6'd14: xpb[88] = 1024'd102896090879795502497607316151392231863311952202614310010003952587424103761956415804079319675666554743969466624599360415496731609624151465387975194311720430148911534745447427043749534989959541236507354827819844007938178843707582674622040810914817134116802055599071900754034811420076551778059149754762379136821;
            6'd15: xpb[88] = 1024'd83660091153182736661979497146888584265398857261571971268975980258316490744101344309367470106501807016515182224758423280622413044417043641225296252830486666388042928390928410974525164805345821527405694970866852898569971436067932128602548318190897761710826508838837666944300184791383026972823655488682778828523;
            6'd16: xpb[88] = 1024'd64424091426569970826351678142384936667485762320529632527948007929208877726246272814655620537337059289060897824917486145748094479209935817062617311349252902627174322036409394905300794620732101818304035113913861789201764028428281582583055825466978389304850962078603433134565558162689502167588161222603178520225;
            6'd17: xpb[88] = 1024'd45188091699957204990723859137881289069572667379487293786920035600101264708391201319943770968172311561606613425076549010873775914002827992899938369868019138866305715681890378836076424436118382109202375256960870679833556620788631036563563332743059016898875415318369199324830931533995977362352666956523578211927;
            6'd18: xpb[88] = 1024'd25952091973344439155096040133377641471659572438444955045892063270993651690536129825231921399007563834152329025235611875999457348795720168737259428386785375105437109327371362766852054251504662400100715400007879570465349213148980490544070840019139644492899868558134965515096304905302452557117172690443977903629;
            6'd19: xpb[88] = 1024'd6716092246731673319468221128873993873746477497402616304864090941886038672681058330520071829842816106698044625394674741125138783588612344574580486905551611344568502972852346697627684066890942690999055543054888461097141805509329944524578347295220272086924321797900731705361678276608927751881678424364377595331;
            6'd20: xpb[88] = 1024'd111546788204243648882639329529184779020531809682095961691967973677755320992135125745823293475335742688686909633011231040829884059222724854967061670440648888517390571187904547966033553073794428703207593294489137198093295248090576171470064424254530348947768678451783555925733579721844035963764873984910371771364;
            6'd21: xpb[88] = 1024'd92310788477630883047011510524681131422618714741053622950940001348647707974280054251111443906170994961232625233170293905955565494015617030804382728959415124756521964833385531896809182889180708994105933437536146088725087840450925625450571931530610976541793131691549322115998953093150511158529379718830771463066;
            6'd22: xpb[88] = 1024'd73074788751018117211383691520177483824705619800011284209912029019540094956424982756399594337006247233778340833329356771081246928808509206641703787478181360995653358478866515827584812704566989285004273580583154979356880432811275079431079438806691604135817584931315088306264326464456986353293885452751171154768;
            6'd23: xpb[88] = 1024'd53838789024405351375755872515673836226792524858968945468884056690432481938569911261687744767841499506324056433488419636206928363601401382479024845996947597234784752124347499758360442519953269575902613723630163869988673025171624533411586946082772231729842038171080854496529699835763461548058391186671570846470;
            6'd24: xpb[88] = 1024'd34602789297792585540128053511170188628879429917926606727856084361324868920714839766975895198676751778869772033647482501332609798394293558316345904515713833473916145769828483689136072335339549866800953866677172760620465617531973987392094453358852859323866491410846620686795073207069936742822896920591970538172;
            6'd25: xpb[88] = 1024'd15366789571179819704500234506666541030966334976884267986828112032217255902859768272264045629512004051415487633806545366458291233187185734153666963034480069713047539415309467619911702150725830157699294009724181651252258209892323441372601960634933486917890944650612386877060446578376411937587402654512370229874;
            6'd26: xpb[88] = 1024'd120197485528691795267671342906977326177751667161577613373931994768086538222313835687567267275004930633404352641423101666163036508821298244546148146569577346885869607630361668888317571157629316169907831761158430388248411652473569668318088037594243563778735301304495211097432348023611520149470598215058364405907;
            6'd27: xpb[88] = 1024'd100961485802079029432043523902473678579838572220535274632904022438978925204458764192855417705840182905950068241582164531288717943614190420383469205088343583125001001275842652819093200973015596460806171904205439278880204244833919122298595544870324191372759754544260977287697721394917995344235103948978764097609;
            6'd28: xpb[88] = 1024'd81725486075466263596415704897970030981925477279492935891876050109871312186603692698143568136675435178495783841741227396414399378407082596220790263607109819364132394921323636749868830788401876751704512047252448169511996837194268576279103052146404818966784207784026743477963094766224470538999609682899163789311;
            6'd29: xpb[88] = 1024'd62489486348853497760787885893466383384012382338450597150848077780763699168748621203431718567510687451041499441900290261540080813199974772058111322125876055603263788566804620680644460603788157042602852190299457060143789429554618030259610559422485446560808661023792509668228468137530945733764115416819563481013;
            6'd30: xpb[88] = 1024'd43253486622240731925160066888962735786099287397408258409820105451656086150893549708719868998345939723587215042059353126665762247992866947895432380644642291842395182212285604611420090419174437333501192333346465950775582021914967484240118066698566074154833114263558275858493841508837420928528621150739963172715;
            6'd31: xpb[88] = 1024'd24017486895627966089532247884459088188186192456365919668792133122548473133038478214008019429181191996132930642218415991791443682785759123732753439163408528081526575857766588542195720234560717624399532476393474841407374614275316938220625573974646701748857567503324042048759214880143896123293126884660362864417;
            6'd32: xpb[88] = 1024'd4781487169015200253904428879955440590273097515323580927764160793440860115183406719296169860016444268678646242377478856917125117578651299570074497682174764320657969503247572472971350049946997915297872619440483732039167206635666392201133081250727329342882020743089808239024588251450371318057632618580762556119;
            6'd33: xpb[88] = 1024'd109612183126527175817075537280266225737058429700016926314868043529310142434637474134599391505509370850667511249994035156621870393212763809962555681217272041493480037718299773741377219056850483927506410370874732469035320649216912619146619158210037406203726377396972632459396489696685479529940828179126756732152;
            6'd34: xpb[88] = 1024'd90376183399914409981447718275762578139145334758974587573840071200202529416782402639887541936344623123213226850153098021747551828005655985799876739736038277732611431363780757672152848872236764218404750513921741359667113241577262073127126665486118033797750830636738398649661863067991954724705333913047156423854;
            6'd35: xpb[88] = 1024'd71140183673301644145819899271258930541232239817932248832812098871094916398927331145175692367179875395758942450312160886873233262798548161637197798254804513971742825009261741602928478687623044509303090656968750250298905833937611527107634172762198661391775283876504164839927236439298429919469839646967556115556;
            6'd36: xpb[88] = 1024'd51904183946688878310192080266755282943319144876889910091784126541987303381072259650463842798015127668304658050471223751998914697591440337474518856773570750210874218654742725533704108503009324800201430800015759140930698426297960981088141680038279288985799737116269931030192609810604905114234345380887955807258;
            6'd37: xpb[88] = 1024'd32668184220076112474564261262251635345406049935847571350756154212879690363217188155751993228850379940850373650630286617124596132384332513311839915292336986450005612300223709464479738318395605091099770943062768031562491018658310435068649187314359916579824190356035697220457983181911380308998851114808355498960;
            6'd38: xpb[88] = 1024'd13432184493463346638936442257747987747492954994805232609728181883772077345362116661040143659685632213396089250789349482250277567177224689149160973811103222689137005945704693395255368133781885381998111086109776922194283611018659889049156694590440544173848643595801463410723356553217855503763356848728755190662;
            6'd39: xpb[88] = 1024'd118262880450975322202107550658058772894278287179498577996832064619641359664816184076343365305178558795384954258405905781955022842811337199541642157346200499861959074160756894663661237140685371394206648837544025659190437053599906115994642771549750621034693000249684287631095257998452963715646552409274749366695;
            6'd40: xpb[88] = 1024'd99026880724362556366479731653555125296365192238456239255804092290533746646961112581631515736013811067930669858564968647080704277604229375378963215864966736101090467806237878594436866956071651685104988980591034549822229645960255569975150278825831248628717453489450053821360631369759438910411058143195149058397;
            6'd41: xpb[88] = 1024'd79790880997749790530851912649051477698452097297413900514776119961426133629106041086919666166849063340476385458724031512206385712397121551216284274383732972340221861451718862525212496771457931976003329123638043440454022238320605023955657786101911876222741906729215820011626004741065914105175563877115548750099;
            6'd42: xpb[88] = 1024'd60554881271137024695224093644547830100539002356371561773748147632318520611250969592207816597684315613022101058883094377332067147190013727053605332902499208579353255097199846455988126586844212266901669266685052331085814830680954477936165293377992503816766359968981586201891378112372389299940069611035948441801;
            6'd43: xpb[88] = 1024'd41318881544524258859596274640044182502625907415329223032720175303210907593395898097495967028519567885567816659042157242457748581982905902890926391421265444818484648742680830386763756402230492557800009409732061221717607423041303931916672800654073131410790813208747352392156751483678864494704575344956348133503;
            6'd44: xpb[88] = 1024'd22082881817911493023968455635540534904712812474286884291692202974103294575540826602784117459354820158113532259201220107583430016775798078728247449940031681057616042388161814317539386217616772848698349552779070112349400015401653385897180307930153759004815266448513118582422124854985339689469081078876747825205;
            6'd45: xpb[88] = 1024'd2846882091298727188340636631036887306799717533244545550664230644995681557685755108072267890190072430659247859360282972709111451568690254565568508458797917296747436033642798248315016033003053139596689695826079002981192607762002839877687815206234386598839719688278884772687498226291814884233586812797147516907;
            6'd46: xpb[88] = 1024'd107677578048810702751511745031347672453585049717937890937768113380864963877139822523375489535682999012648112866976839272413856727202802764958049691993895194469569504248694999516720885039906539151805227447260327739977346050343249066823173892165544463459684076342161708993059399671526923096116782373343141692940;
            6'd47: xpb[88] = 1024'd88441578322197936915883926026844024855671954776895552196740141051757350859284751028663639966518251285193828467135902137539538161995694940795370750512661430708700897894175983447496514855292819442703567590307336630609138642703598520803681399441625091053708529581927475183324773042833398290881288107263541384642;
            6'd48: xpb[88] = 1024'd69205578595585171080256107022340377257758859835853213455712168722649737841429679533951790397353503557739544067294965002665219596788587116632691809031427666947832291539656967378272144670679099733601907733354345521240931235063947974784188906717705718647732982821693241373590146414139873485645793841183941076344;
            6'd49: xpb[88] = 1024'd49969578868972405244628288017836729659845764894810874714684196393542124823574608039239940828188755830285259667454027867790901031581479292470012867550193903186963685185137951309047774486065380024500247876401354411872723827424297428764696413993786346241757436061459007563855519785446348680410299575104340768046;
            6'd50: xpb[88] = 1024'd30733579142359639409000469013333082061932669953768535973656224064434511805719536544528091259024008102830975267613090732916582466374371468307333926068960139426095078830618935239823404301451660315398588019448363302504516419784646882745203921269866973835781889301224773754120893156752823875174805309024740459748;
            6'd51: xpb[88] = 1024'd11497579415746873573372650008829434464019575012726197232628251735326898787864465049816241689859260375376690867772153598042263901167263644144654984587726375665226472476099919170599034116837940606296928162495372193136309012144996336725711428545947601429806342540990539944386266528059299069939311042945140151450;
            6'd52: xpb[88] = 1024'd116328275373258849136543758409140219610804907197419542619732134471196181107318532465119463335352186957365555875388709897747009176801376154537136168122823652838048540691152120439004903123741426618505465913929620930132462454726242563671197505505257678290650699194873364164758167973294407281822506603491134327483;
            6'd53: xpb[88] = 1024'd97092275646646083300915939404636572012891812256377203878704162142088568089463460970407613766187439229911271475547772762872690611594268330374457226641589889077179934336633104369780532939127706909403806056976629820764255047086592017651705012781338305884675152434639130355023541344600882476587012337411534019185;
            6'd54: xpb[88] = 1024'd77856275920033317465288120400132924414978717315334865137676189812980955071608389475695764197022691502456987075706835627998372046387160506211778285160356125316311327982114088300556162754513987200302146200023638711396047639446941471632212520057418933478699605674404896545288914715907357671351518071331933710887;
            6'd55: xpb[88] = 1024'd58620276193420551629660301395629276817065622374292526396648217483873342053753317980983914627857943775002702675865898493124053481180052682049099343679122361555442721627595072231331792569900267491200486343070647602027840231807290925612720027333499561072724058914170662735554288087213832866116023805252333402589;
            6'd56: xpb[88] = 1024'd39384276466807785794032482391125629219152527433250187655620245154765729035898246486272065058693196047548418276024961358249734915972944857886420402197888597794574115273076056162107422385286547782098826486117656492659632824167640379593227534609580188666748512153936428925819661458520308060880529539172733094291;
            6'd57: xpb[88] = 1024'd20148276740195019958404663386621981621239432492207848914592272825658116018043174991560215489528448320094133876184024223375416350765837033723741460716654834033705508918557040092883052200672828072997166629164665383291425416527989833573735041885660816260772965393702195116085034829826783255645035273093132785993;
            6'd58: xpb[88] = 1024'd912277013582254122776844382118334023326337551165510173564300496550503000188103496848365920363700592639849476343087088501097785558729209561062519235421070272836902564038024023658682016059108363895506772211674273923218008888339287554242549161741443854797418633467961306350408201133258450409541007013532477695;
            6'd59: xpb[88] = 1024'd105742972971094229685947952782429119170111669735858855560668183232419785319642170912151587565856627174628714483959643388205843061192841719953543702770518347445658970779090225292064551022962594376104044523645923010919371451469585514499728626121051520715641775287350785526722309646368366662292736567559526653728;
            6'd60: xpb[88] = 1024'd86506973244481463850320133777925471572198574794816516819640210903312172301787099417439737996691879447174430084118706253331524495985733895790864761289284583684790364424571209222840180838348874667002384666692931901551164043829934968480236133397132148309666228527116551716987683017674841857057242301479926345430;
            6'd61: xpb[88] = 1024'd67270973517868698014692314773421823974285479853774178078612238574204559283932027922727888427527131719720145684277769118457205930778626071628185819808050819923921758070052193153615810653735154957900724809739940792182956636190284422460743640673212775903690681766882317907253056388981317051821748035400326037132;
            6'd62: xpb[88] = 1024'd48034973791255932179064495768918176376372384912731839337584266245096946266076956428016038858362383992265861284436831983582887365571518247465506878326817056163053151715533177084391440469121435248799064952786949682814749228550633876441251147949293403497715135006648084097518429760287792246586253769320725728834;
            6'd63: xpb[88] = 1024'd28798974064643166343436676764414528778459289971689500596556293915989333248221884933304189289197636264811576884595894848708568800364410423302827936845583292402184545361014161015167070284507715539697405095833958573446541820910983330421758655225374031091739588246413850287783803131594267441350759503241125420536;
        endcase
    end

    always_comb begin
        case(flag[29][16:12])
            5'd0: xpb[89] = 1024'd0;
            5'd1: xpb[89] = 1024'd9562974338030400507808857759910881180546195030647161855528321586881720230366813438592339720032888537357292484754957713834250235157302599140148995364349528641315939006495144945942700099893995830595745238880967464078334413271332784402266162501454658685764041486179616478049176502900742636115265237161525112238;
            5'd2: xpb[89] = 1024'd19125948676060801015617715519821762361092390061294323711056643173763440460733626877184679440065777074714584969509915427668500470314605198280297990728699057282631878012990289891885400199787991661191490477761934928156668826542665568804532325002909317371528082972359232956098353005801485272230530474323050224476;
            5'd3: xpb[89] = 1024'd28688923014091201523426573279732643541638585091941485566584964760645160691100440315777019160098665612071877454264873141502750705471907797420446986093048585923947817019485434837828100299681987491787235716642902392235003239813998353206798487504363976057292124458538849434147529508702227908345795711484575336714;
            5'd4: xpb[89] = 1024'd38251897352121602031235431039643524722184780122588647422113286347526880921467253754369358880131554149429169939019830855337000940629210396560595981457398114565263756025980579783770800399575983322382980955523869856313337653085331137609064650005818634743056165944718465912196706011602970544461060948646100448952;
            5'd5: xpb[89] = 1024'd47814871690152002539044288799554405902730975153235809277641607934408601151834067192961698600164442686786462423774788569171251175786512995700744976821747643206579695032475724729713500499469979152978726194404837320391672066356663922011330812507273293428820207430898082390245882514503713180576326185807625561190;
            5'd6: xpb[89] = 1024'd57377846028182403046853146559465287083277170183882971133169929521290321382200880631554038320197331224143754908529746283005501410943815594840893972186097171847895634038970869675656200599363974983574471433285804784470006479627996706413596975008727952114584248917077698868295059017404455816691591422969150673428;
            5'd7: xpb[89] = 1024'd66940820366212803554662004319376168263823365214530132988698251108172041612567694070146378040230219761501047393284703996839751646101118193981042967550446700489211573045466014621598900699257970814170216672166772248548340892899329490815863137510182610800348290403257315346344235520305198452806856660130675785666;
            5'd8: xpb[89] = 1024'd76503794704243204062470862079287049444369560245177294844226572695053761842934507508738717760263108298858339878039661710674001881258420793121191962914796229130527512051961159567541600799151966644765961911047739712626675306170662275218129300011637269486112331889436931824393412023205941088922121897292200897904;
            5'd9: xpb[89] = 1024'd86066769042273604570279719839197930624915755275824456699754894281935482073301320947331057480295996836215632362794619424508252116415723392261340958279145757771843451058456304513484300899045962475361707149928707176705009719441995059620395462513091928171876373375616548302442588526106683725037387134453726010142;
            5'd10: xpb[89] = 1024'd95629743380304005078088577599108811805461950306471618555283215868817202303668134385923397200328885373572924847549577138342502351573025991401489953643495286413159390064951449459427000998939958305957452388809674640783344132713327844022661625014546586857640414861796164780491765029007426361152652371615251122380;
            5'd11: xpb[89] = 1024'd105192717718334405585897435359019692986008145337118780410811537455698922534034947824515736920361773910930217332304534852176752586730328590541638949007844815054475329071446594405369701098833954136553197627690642104861678545984660628424927787516001245543404456347975781258540941531908168997267917608776776234618;
            5'd12: xpb[89] = 1024'd114755692056364806093706293118930574166554340367765942266339859042580642764401761263108076640394662448287509817059492566011002821887631189681787944372194343695791268077941739351312401198727949967148942866571609568940012959255993412827193950017455904229168497834155397736590118034808911633383182845938301346856;
            5'd13: xpb[89] = 1024'd251970710270465202716223474027022602402108272677419993736325564485467657459435791685345145769876676201652894356956845266189216203713454266776814720212831403416532514865666959624862107104740076434490497065337186653986522306429424264481542835681113648112635906217956184532766463781021252379758256474231974763;
            5'd14: xpb[89] = 1024'd9814945048300865710525081233937903782948303303324581849264647151367187887826249230277684865802765213558945379111914559100439451361016053406925810084562360044732471521360811905567562206998735907030235735946304650732320935577762208666747705337135772333876677392397572662581942966681763888495023493635757087001;
            5'd15: xpb[89] = 1024'd19377919386331266218333938993848784963494498333971743704792968738248908118193062668870024585835653750916237863866872272934689686518318652547074805448911888686048410527855956851510262306892731737625980974827272114810655348849094993069013867838590431019640718878577189140631119469582506524610288730797282199239;
            5'd16: xpb[89] = 1024'd28940893724361666726142796753759666144040693364618905560321290325130628348559876107462364305868542288273530348621829986768939921675621251687223800813261417327364349534351101797452962406786727568221726213708239578888989762120427777471280030340045089705404760364756805618680295972483249160725553967958807311477;
            5'd17: xpb[89] = 1024'd38503868062392067233951654513670547324586888395266067415849611912012348578926689546054704025901430825630822833376787700603190156832923850827372796177610945968680288540846246743395662506680723398817471452589207042967324175391760561873546192841499748391168801850936422096729472475383991796840819205120332423715;
            5'd18: xpb[89] = 1024'd48066842400422467741760512273581428505133083425913229271377933498894068809293502984647043745934319362988115318131745414437440391990226449967521791541960474609996227547341391689338362606574719229413216691470174507045658588663093346275812355342954407076932843337116038574778648978284734432956084442281857535953;
            5'd19: xpb[89] = 1024'd57629816738452868249569370033492309685679278456560391126906255085775789039660316423239383465967207900345407802886703128271690627147529049107670786906310003251312166553836536635281062706468715060008961930351141971123993001934426130678078517844409065762696884823295655052827825481185477069071349679443382648191;
            5'd20: xpb[89] = 1024'd67192791076483268757378227793403190866225473487207552982434576672657509270027129861831723186000096437702700287641660842105940862304831648247819782270659531892628105560331681581223762806362710890604707169232109435202327415205758915080344680345863724448460926309475271530877001984086219705186614916604907760429;
            5'd21: xpb[89] = 1024'd76755765414513669265187085553314072046771668517854714837962898259539229500393943300424062906032984975059992772396618555940191097462134247387968777635009060533944044566826826527166462906256706721200452408113076899280661828477091699482610842847318383134224967795654888008926178486986962341301880153766432872667;
            5'd22: xpb[89] = 1024'd86318739752544069772995943313224953227317863548501876693491219846420949730760756739016402626065873512417285257151576269774441332619436846528117772999358589175259983573321971473109163006150702551796197646994044363358996241748424483884877005348773041819989009281834504486975354989887704977417145390927957984905;
            5'd23: xpb[89] = 1024'd95881714090574470280804801073135834407864058579149038549019541433302669961127570177608742346098762049774577741906533983608691567776739445668266768363708117816575922579817116419051863106044698382391942885875011827437330655019757268287143167850227700505753050768014120965024531492788447613532410628089483097143;
            5'd24: xpb[89] = 1024'd105444688428604870788613658833046715588410253609796200404547863020184390191494383616201082066131650587131870226661491697442941802934042044808415763728057646457891861586312261364994563205938694212987688124755979291515665068291090052689409330351682359191517092254193737443073707995689190249647675865251008209381;
            5'd25: xpb[89] = 1024'd115007662766635271296422516592957596768956448640443362260076184607066110421861197054793421786164539124489162711416449411277192038091344643948564759092407175099207800592807406310937263305832690043583433363636946755593999481562422837091675492853137017877281133740373353921122884498589932885762941102412533321619;
            5'd26: xpb[89] = 1024'd503941420540930405432446948054045204804216545354839987472651128970935314918871583370690291539753352403305788713913690532378432407426908533553629440425662806833065029731333919249724214209480152868980994130674373307973044612858848528963085671362227296225271812435912369065532927562042504759516512948463949526;
            5'd27: xpb[89] = 1024'd10066915758571330913241304707964926385350411576002001843000972715852655545285685021963030011572641889760598273468871404366628667564729507673702624804775191448149004036226478865192424314103475983464726233011641837386307457884191632931229248172816885981989313298615528847114709430462785140874781750109989061764;
            5'd28: xpb[89] = 1024'd19629890096601731421050162467875807565896606606649163698529294302734375775652498460555369731605530427117890758223829118200878902722032106813851620169124720089464943042721623811135124413997471814060471471892609301464641871155524417333495410674271544667753354784795145325163885933363527776990046987271514174002;
            5'd29: xpb[89] = 1024'd29192864434632131928859020227786688746442801637296325554057615889616096006019311899147709451638418964475183242978786832035129137879334705954000615533474248730780882049216768757077824513891467644656216710773576765542976284426857201735761573175726203353517396270974761803213062436264270413105312224433039286240;
            5'd30: xpb[89] = 1024'd38755838772662532436667877987697569926988996667943487409585937476497816236386125337740049171671307501832475727733744545869379373036637305094149610897823777372096821055711913703020524613785463475251961949654544229621310697698189986138027735677180862039281437757154378281262238939165013049220577461594564398478;
            5'd31: xpb[89] = 1024'd48318813110692932944476735747608451107535191698590649265114259063379536466752938776332388891704196039189768212488702259703629608193939904234298606262173306013412760062207058648963224713679459305847707188535511693699645110969522770540293898178635520725045479243333994759311415442065755685335842698756089510716;
        endcase
    end

    always_comb begin
        case(flag[30][5:0])
            6'd0: xpb[90] = 1024'd0;
            6'd1: xpb[90] = 1024'd28940893724361666726142796753759666144040693364618905560321290325130628348559876107462364305868542288273530348621829986768939921675621251687223800813261417327364349534351101797452962406786727568221726213708239578888989762120427777471280030340045089705404760364756805618680295972483249160725553967958807311477;
            6'd2: xpb[90] = 1024'd57881787448723333452285593507519332288081386729237811120642580650261256697119752214924728611737084576547060697243659973537879843351242503374447601626522834654728699068702203594905924813573455136443452427416479157777979524240855554942560060680090179410809520729513611237360591944966498321451107935917614622954;
            6'd3: xpb[90] = 1024'd86822681173085000178428390261278998432122080093856716680963870975391885045679628322387092917605626864820591045865489960306819765026863755061671402439784251982093048603053305392358887220360182704665178641124718736666969286361283332413840091020135269116214281094270416856040887917449747482176661903876421934431;
            6'd4: xpb[90] = 1024'd115763574897446666904571187015038664576162773458475622241285161300522513394239504429849457223474169153094121394487319947075759686702485006748895203253045669309457398137404407189811849627146910272886904854832958315555959048481711109885120121360180358821619041459027222474721183889932996642902215871835229245908;
            6'd5: xpb[90] = 1024'd20637772937683592231915056363983897975505039697358843673474596560676246405490241627296750314685037131924502335651656499265635767536885923880958879049976045703131073102184291649634572842416432119798433460153958048080587960381242114391421582016995999260203898409666970063294951788487612786509080013168442073054;
            6'd6: xpb[90] = 1024'd49578666662045258958057853117743564119545733061977749233795886885806874754050117734759114620553579420198032684273486486034575689212507175568182679863237463030495422636535393447087535249203159688020159673862197626969577722501669891862701612357041088965608658774423775681975247760970861947234633981127249384531;
            6'd7: xpb[90] = 1024'd78519560386406925684200649871503230263586426426596654794117177210937503102609993842221478926422121708471563032895316472803515610888128427255406480676498880357859772170886495244540497655989887256241885887570437205858567484622097669333981642697086178671013419139180581300655543733454111107960187949086056696008;
            6'd8: xpb[90] = 1024'd107460454110768592410343446625262896407627119791215560354438467536068131451169869949683843232290663996745093381517146459572455532563749678942630281489760297685224121705237597041993460062776614824463612101278676784747557246742525446805261673037131268376418179503937386919335839705937360268685741917044864007485;
            6'd9: xpb[90] = 1024'd12334652151005517737687315974208129806969386030098781786627902796221864462420607147131136323501531975575474322681483011762331613398150596074693957286690674078897796670017481501816183278046136671375140706599676517272186158642056451311563133693946908815003036454577134507909607604491976412292606058378076834631;
            6'd10: xpb[90] = 1024'd41275545875367184463830112727967795951010079394717687346949193121352492810980483254593500629370074263849004671303312998531271535073771847761917758099952091406262146204368583299269145684832864239596866920307916096161175920762484228782843164033991998520407796819333940126589903576975225573018160026336884146108;
            6'd11: xpb[90] = 1024'd70216439599728851189972909481727462095050772759336592907270483446483121159540359362055864935238616552122535019925142985300211456749393099449141558913213508733626495738719685096722108091619591807818593134016155675050165682882912006254123194374037088225812557184090745745270199549458474733743713994295691457585;
            6'd12: xpb[90] = 1024'd99157333324090517916115706235487128239091466123955498467591773771613749508100235469518229241107158840396065368546972972069151378425014351136365359726474926060990845273070786894175070498406319376040319347724395253939155445003339783725403224714082177931217317548847551363950495521941723894469267962254498769062;
            6'd13: xpb[90] = 1024'd4031531364327443243459575584432361638433732362838719899781209031767482519350972666965522332318026819226446309711309524259027459259415268268429035523405302454664520237850671353997793713675841222951847953045394986463784356902870788231704685370897818369802174499487298952524263420496340038076132103587711596208;
            6'd14: xpb[90] = 1024'd32972425088689109969602372338192027782474425727457625460102499356898110867910848774427886638186569107499976658333139511027967380935036519955652836336666719782028869772201773151450756120462568791173574166753634565352774119023298565702984715710942908075206934864244104571204559392979589198801686071546518907685;
            6'd15: xpb[90] = 1024'd61913318813050776695745169091951693926515119092076531020423789682028739216470724881890250944055111395773507006954969497796907302610657771642876637149928137109393219306552874948903718527249296359395300380461874144241763881143726343174264746050987997780611695229000910189884855365462838359527240039505326219162;
            6'd16: xpb[90] = 1024'd90854212537412443421887965845711360070555812456695436580745080007159367565030600989352615249923653684047037355576799484565847224286279023330100437963189554436757568840903976746356680934036023927617026594170113723130753643264154120645544776391033087486016455593757715808565151337946087520252794007464133530639;
            6'd17: xpb[90] = 1024'd119795106261774110148030762599471026214596505821314342141066370332289995913590477096814979555792195972320567704198629471334787145961900275017324238776450971764121918375255078543809643340822751495838752807878353302019743405384581898116824806731078177191421215958514521427245447310429336680978347975422940842116;
            6'd18: xpb[90] = 1024'd24669304302011035475374631948416259613938772060197563573255805592443728924841214294262272647003063951150948645362966023524663226796301192149387914573381348157795593340034963003632366556092273342750281413199353034544372317284112902623126267387893817630006072909154269015819215208983952824585212116756153669262;
            6'd19: xpb[90] = 1024'd53610198026372702201517428702175925757979465424816469133577095917574357273401090401724636952871606239424478993984796010293603148471922443836611715386642765485159942874386064801085328962879000910972007626907592613433362079404540680094406297727938907335410833273911074634499511181467201985310766084714960980739;
            6'd20: xpb[90] = 1024'd82551091750734368927660225455935591902020158789435374693898386242704985621960966509187001258740148527698009342606625997062543070147543695523835516199904182812524292408737166598538291369665728479193733840615832192322351841524968457565686328067983997040815593638667880253179807153950451146036320052673768292216;
            6'd21: xpb[90] = 1024'd111491985475096035653803022209695258046060852154054280254219676567835613970520842616649365564608690815971539691228455983831482991823164947211059317013165600139888641943088268395991253776452456047415460054324071771211341603645396235036966358408029086746220354003424685871860103126433700306761874020632575603693;
            6'd22: xpb[90] = 1024'd16366183515332960981146891558640491445403118392937501686409111827989346981771579814096658655819558794801920632392792536021359072657565864343122992810095976533562316907868152855813976991721977894326988659645071503735970515544927239543267819064844727184805210954064433460433871024988316450368738161965788430839;
            6'd23: xpb[90] = 1024'd45307077239694627707289688312400157589443811757556407246730402153119975330331455921559022961688101083075450981014622522790298994333187116030346793623357393860926666442219254653266939398508705462548714873353311082624960277665355017014547849404889816890209971318821239079114166997471565611094292129924595742316;
            6'd24: xpb[90] = 1024'd74247970964056294433432485066159823733484505122175312807051692478250603678891332029021387267556643371348981329636452509559238916008808367717570594436618811188291015976570356450719901805295433030770441087061550661513950039785782794485827879744934906595614731683578044697794462969954814771819846097883403053793;
            6'd25: xpb[90] = 1024'd103188864688417961159575281819919489877525198486794218367372982803381232027451208136483751573425185659622511678258282496328178837684429619404794395249880228515655365510921458248172864212082160598992167300769790240402939801906210571957107910084979996301019492048334850316474758942438063932545400065842210365270;
            6'd26: xpb[90] = 1024'd8063062728654886486919151168864723276867464725677439799562418063534965038701945333931044664636053638452892619422619048518054918518830536536858071046810604909329040475701342707995587427351682445903695906090789972927568713805741576463409370741795636739604348998974597905048526840992680076152264207175423192416;
            6'd27: xpb[90] = 1024'd37003956453016553213061947922624389420908158090296345359883708388665593387261821441393408970504595926726422968044449035286994840194451788224081871860072022236693390010052444505448549834138410014125422119799029551816558475926169353934689401081840726445009109363731403523728822813475929236877818175134230503893;
            6'd28: xpb[90] = 1024'd65944850177378219939204744676384055564948851454915250920204998713796221735821697548855773276373138214999953316666279022055934761870073039911305672673333439564057739544403546302901512240925137582347148333507269130705548238046597131405969431421885816150413869728488209142409118785959178397603372143093037815370;
            6'd29: xpb[90] = 1024'd94885743901739886665347541430143721708989544819534156480526289038926850084381573656318137582241680503273483665288109008824874683545694291598529473486594856891422089078754648100354474647711865150568874547215508709594538000167024908877249461761930905855818630093245014761089414758442427558328926111051845126847;
            6'd30: xpb[90] = 1024'd123826637626101553391490338183903387853030238184153062040847579364057478432941449763780501888110222791547014013909938995593814605221315543285753274299856274218786438613105749897807437054498592718790600760923748288483527762287452686348529492101975995561223390458001820379769710730925676719054480079010652438324;
            6'd31: xpb[90] = 1024'd28700835666338478718834207532848621252372504423036283473037014624211211444192186961227794979321090770377394955074275547783690686055716460417816950096786650612460113577885634357630160269768114565702129366244748021008156674186983690854830952758791635999808247408641567968343478629480292862661344220343865265470;
            6'd32: xpb[90] = 1024'd57641729390700145444977004286608287396413197787655189033358304949341839792752063068690159285189633058650925303696105534552630607731337712105040750910048067939824463112236736155083122676554842133923855579952987599897146436307411468326110983098836725705213007773398373587023774601963542023386898188302672576947;
            6'd33: xpb[90] = 1024'd86582623115061812171119801040367953540453891152274094593679595274472468141311939176152523591058175346924455652317935521321570529406958963792264551723309485267188812646587837952536085083341569702145581793661227178786136198427839245797391013438881815410617768138155179205704070574446791184112452156261479888424;
            6'd34: xpb[90] = 1024'd115523516839423478897262597794127619684494584516893000154000885599603096489871815283614887896926717635197986000939765508090510451082580215479488352536570902594553162180938939749989047490128297270367308007369466757675125960548267023268671043778926905116022528502911984824384366546930040344838006124220287199901;
            6'd35: xpb[90] = 1024'd20397714879660404224606467143072853083836850755776221586190320859756829501122552481062180988137585614028366942104102060280386531916981132611552028333501278988226837145718824209811770705397819117278836612690466490199754872447798027774972504435742545554607385453551732412958134445484656488444870265553500027047;
            6'd36: xpb[90] = 1024'd49338608604022070950749263896832519227877544120395127146511611184887457849682428588524545294006127902301897290725932047049326453592602384298775829146762696315591186680069926007264733112184546685500562826398706069088744634568225805246252534775787635260012145818308538031638430417967905649170424233512307338524;
            6'd37: xpb[90] = 1024'd78279502328383737676892060650592185371918237485014032706832901510018086198242304695986909599874670190575427639347762033818266375268223635985999629960024113642955536214421027804717695518971274253722289040106945647977734396688653582717532565115832724965416906183065343650318726390451154809895978201471114650001;
            6'd38: xpb[90] = 1024'd107220396052745404403034857404351851515958930849632938267154191835148714546802180803449273905743212478848957987969592020587206296943844887673223430773285530970319885748772129602170657925758001821944015253815185226866724158809081360188812595455877814670821666547822149268999022362934403970621532169429921961478;
            6'd39: xpb[90] = 1024'd12094594092982329730378726753297084915301197088516159699343627095302447558052918000896566996954080457679338929133928572777082377778245804805287106570215907363993560713552014061993381141027523668855543859136184959391353070708612364695114056112693455109406523498461896857572790261489020114228396310763134788624;
            6'd40: xpb[90] = 1024'd41035487817343996456521523507056751059341890453135065259664917420433075906612794108358931302822622745952869277755758559546022299453867056492510907383477324691357910247903115859446343547814251237077270072844424538280342832829040142166394086452738544814811283863218702476253086233972269274953950278721942100101;
            6'd41: xpb[90] = 1024'd69976381541705663182664320260816417203382583817753970819986207745563704255172670215821295608691165034226399626377588546314962221129488308179734708196738742018722259782254217656899305954600978805298996286552664117169332594949467919637674116792783634520216044227975508094933382206455518435679504246680749411578;
            6'd42: xpb[90] = 1024'd98917275266067329908807117014576083347423277182372876380307498070694332603732546323283659914559707322499929974999418533083902142805109559866958509010000159346086609316605319454352268361387706373520722500260903696058322357069895697108954147132828724225620804592732313713613678178938767596405058214639556723055;
            6'd43: xpb[90] = 1024'd3791473306304255236150986363521316746765543421256097812496933330848065614983283520730953005770575301330310916163755085273778223639510476999022184806930535739760284281385203914174991576657228220432251105581903428582951268969426701615255607789644364664205661543372061302187446077493383740011922355972769550201;
            6'd44: xpb[90] = 1024'd32732367030665921962293783117280982890806236785875003372818223655978693963543159628193317311639117589603841264785585072042718145315131728686245985620191953067124633815736305711627953983443955788653977319290143007471941031089854479086535638129689454369610421908128866920867742049976632900737476323931576861678;
            6'd45: xpb[90] = 1024'd61673260755027588688436579871040649034846930150493908933139513981109322312103035735655681617507659877877371613407415058811658066990752980373469786433453370394488983350087407509080916390230683356875703532998382586360930793210282256557815668469734544075015182272885672539548038022459882061463030291890384173155;
            6'd46: xpb[90] = 1024'd90614154479389255414579376624800315178887623515112814493460804306239950660662911843118045923376202166150901962029245045580597988666374232060693587246714787721853332884438509306533878797017410925097429746706622165249920555330710034029095698809779633780419942637642478158228333994943131222188584259849191484632;
            6'd47: xpb[90] = 1024'd119555048203750922140722173378559981322928316879731720053782094631370579009222787950580410229244744454424432310651075032349537910341995483747917388059976205049217682418789611103986841203804138493319155960414861744138910317451137811500375729149824723485824703002399283776908629967426380382914138227807998796109;
            6'd48: xpb[90] = 1024'd24429246243987847468066042727505214722270583118614941485971529891524312020473525148027703320455612433254813251815411584539413991176396400879981063856906581442891357383569495563809564419073660340230684565735861476663539229350668816006677189806640363924409559953039031365482397865980996526521002369141211623255;
            6'd49: xpb[90] = 1024'd53370139968349514194208839481264880866311276483233847046292820216654940369033401255490067626324154721528343600437241571308353912852017652567204864670167998770255706917920597361262526825860387908452410779444101055552528991471096593477957220146685453629814320317795836984162693838464245687246556337100018934732;
            6'd50: xpb[90] = 1024'd82311033692711180920351636235024547010351969847852752606614110541785568717593277362952431932192697009801873949059071558077293834527638904254428665483429416097620056452271699158715489232647115476674136993152340634441518753591524370949237250486730543335219080682552642602842989810947494847972110305058826246209;
            6'd51: xpb[90] = 1024'd111251927417072847646494432988784213154392663212471658166935400866916197066153153470414796238061239298075404297680901544846233756203260155941652466296690833424984405986622800956168451639433843044895863206860580213330508515711952148420517280826775633040623841047309448221523285783430744008697664273017633557686;
            6'd52: xpb[90] = 1024'd16126125457309772973838302337729446553734929451354879599124836127069930077403890667862089329272107276905785238845238097036109837037661073073716142093621209818658080951402685415991174854703364891807391812181579945855137427611483152926818741483591273479208697997949195810097053681985360152304528414350846384832;
            6'd53: xpb[90] = 1024'd45067019181671439699981099091489112697775622815973785159446126452200558425963766775324453635140649565179315587467068083805049758713282324760939942906882627146022430485753787213444137261490092460029118025889819524744127189731910930398098771823636363184613458362706001428777349654468609313030082382309653696309;
            6'd54: xpb[90] = 1024'd74007912906033106426123895845248778841816316180592690719767416777331186774523642882786817941009191853452845936088898070573989680388903576448163743720144044473386780020104889010897099668276820028250844239598059103633116951852338707869378802163681452890018218727462807047457645626951858473755636350268461007786;
            6'd55: xpb[90] = 1024'd102948806630394773152266692599008444985857009545211596280088707102461815123083518990249182246877734141726376284710728057342929602064524828135387544533405461800751129554455990808350062075063547596472570453306298682522106713972766485340658832503726542595422979092219612666137941599435107634481190318227268319263;
            6'd56: xpb[90] = 1024'd7823004670631698479610561947953678385199275784094817712278142362615548134334256187696475338088602120556757225875064609532805682898925745267451220330335838194424804519235875268172785290333069443384099058627298415046735625872297489846960293160542183034007836042859360254711709497989723778088054459560481146409;
            6'd57: xpb[90] = 1024'd36763898394993365205753358701713344529239969148713723272599432687746176482894132295158839643957144408830287574496894596301745604574546996954675021143597255521789154053586977065625747697119797011605825272335537993935725387992725267318240323500587272739412596407616165873392005470472972938813608427519288457886;
            6'd58: xpb[90] = 1024'd65704792119355031931896155455473010673280662513332628832920723012876804831454008402621203949825686697103817923118724583070685526250168248641898821956858672849153503587938078863078710103906524579827551486043777572824715150113153044789520353840632362444817356772372971492072301442956222099539162395478095769363;
            6'd59: xpb[90] = 1024'd94645685843716698658038952209232676817321355877951534393242013338007433180013884510083568255694228985377348271740554569839625447925789500329122622770120090176517853122289180660531672510693252148049277699752017151713704912233580822260800384180677452150222117137129777110752597415439471260264716363436903080840;
            6'd60: xpb[90] = 1024'd123586579568078365384181748962992342961362049242570439953563303663138061528573760617545932561562771273650878620362384556608565369601410752016346423583381507503882202656640282457984634917479979716271003913460256730602694674354008599732080414520722541855626877501886582729432893387922720420990270331395710392317;
            6'd61: xpb[90] = 1024'd28460777608315290711525618311937576360704315481453661385752738923291794539824497814993225652773639252481259561526721108798441450435811669148410099380311883897555877621420166917807358132749501563182532518781256463127323586253539604238381875177538182294211734452526330318006661286477336564597134472728923219463;
            6'd62: xpb[90] = 1024'd57401671332676957437668415065697242504745008846072566946074029248422422888384373922455589958642181540754789910148551095567381372111432920835633900193573301224920227155771268715260320539536229131404258732489496042016313348373967381709661905517583271999616494817283135936686957258960585725322688440687730530940;
            6'd63: xpb[90] = 1024'd86342565057038624163811211819456908648785702210691472506395319573553051236944250029917954264510723829028320258770381082336321293787054172522857701006834718552284576690122370512713282946322956699625984946197735620905303110494395159180941935857628361705021255182039941555367253231443834886048242408646537842417;
        endcase
    end

    always_comb begin
        case(flag[30][11:6])
            6'd0: xpb[91] = 1024'd0;
            6'd1: xpb[91] = 1024'd115283458781400290889954008573216574792826395575310378066716609898683679585504126137380318570379266117301850607392211069105261215462675424210081501820096135879648926224473472310166245353109684267847711159905975199794292872614822936652221966197673451410426015546796747174047549203927084046773796376605345153894;
            6'd2: xpb[91] = 1024'd106500221878675840381109089741618716840954364024885072005301364732390463833699113364745565926100857925160551807326928703631458590084130513865002878623861230825607177879375727282702251514702162814385224711424710553224224895008749100339465362712117453554032127679476436317988570333925535076428902926585095823457;
            6'd3: xpb[91] = 1024'd97716984975951389872264170910020858889082332474459765943886119566097248081894100592110813281822449733019253007261646338157655964705585603519924255427626325771565429534277982255238257676294641360922738262943445906654156917402675264026708759226561455697638239812156125461929591463923986106084009476564846493020;
            6'd4: xpb[91] = 1024'd88933748073226939363419252078423000937210300924034459882470874399804032330089087819476060637544041540877954207196363972683853339327040693174845632231391420717523681189180237227774263837887119907460251814462181260084088939796601427713952155741005457841244351944835814605870612593922437135739116026544597162583;
            6'd5: xpb[91] = 1024'd80150511170502488854574333246825142985338269373609153821055629233510816578284075046841307993265633348736655407131081607210050713948495782829767009035156515663481932844082492200310269999479598453997765365980916613514020962190527591401195552255449459984850464077515503749811633723920888165394222576524347832146;
            6'd6: xpb[91] = 1024'd71367274267778038345729414415227285033466237823183847759640384067217600826479062274206555348987225156595356607065799241736248088569950872484688385838921610609440184498984747172846276161072077000535278917499651966943952984584453755088438948769893462128456576210195192893752654853919339195049329126504098501709;
            6'd7: xpb[91] = 1024'd62584037365053587836884495583629427081594206272758541698225138900924385074674049501571802704708816964454057807000516876262445463191405962139609762642686705555398436153887002145382282322664555547072792469018387320373885006978379918775682345284337464272062688342874882037693675983917790224704435676483849171272;
            6'd8: xpb[91] = 1024'd53800800462329137328039576752031569129722174722333235636809893734631169322869036728937050060430408772312759006935234510788642837812861051794531139446451800501356687808789257117918288484257034093610306020537122673803817029372306082462925741798781466415668800475554571181634697113916241254359542226463599840835;
            6'd9: xpb[91] = 1024'd45017563559604686819194657920433711177850143171907929575394648568337953571064023956302297416152000580171460206869952145314840212434316141449452516250216895447314939463691512090454294645849512640147819572055858027233749051766232246150169138313225468559274912608234260325575718243914692284014648776443350510398;
            6'd10: xpb[91] = 1024'd36234326656880236310349739088835853225978111621482623513979403402044737819259011183667544771873592388030161406804669779841037587055771231104373893053981990393273191118593767062990300807441991186685333123574593380663681074160158409837412534827669470702881024740913949469516739373913143313669755326423101179961;
            6'd11: xpb[91] = 1024'd27451089754155785801504820257237995274106080071057317452564158235751522067453998411032792127595184195888862606739387414367234961677226320759295269857747085339231442773496022035526306969034469733222846675093328734093613096554084573524655931342113472846487136873593638613457760503911594343324861876402851849524;
            6'd12: xpb[91] = 1024'd18667852851431335292659901425640137322234048520632011391148913069458306315648985638398039483316776003747563806674105048893432336298681410414216646661512180285189694428398277008062313130626948279760360226612064087523545118948010737211899327856557474990093249006273327757398781633910045372979968426382602519087;
            6'd13: xpb[91] = 1024'd9884615948706884783814982594042279370362016970206705329733667903165090563843972865763286839038367811606265006608822683419629710920136500069138023465277275231147946083300531980598319292219426826297873778130799440953477141341936900899142724371001477133699361138953016901339802763908496402635074976362353188650;
            6'd14: xpb[91] = 1024'd1101379045982434274970063762444421418489985419781399268318422736871874812038960093128534194759959619464966206543540317945827085541591589724059400269042370177106197738202786953134325453811905372835387329649534794383409163735863064586386120885445479277305473271632706045280823893906947432290181526342103858213;
            6'd15: xpb[91] = 1024'd116384837827382725164924072335660996211316380995091777335035032635555554397543086230508852765139225736766816813935751387051088301004267013934140902089138506056755123962676259263300570806921589640683098489555509994177702036350686001238608087083118930687731488818429453219328373097834031479063977902947449012107;
            6'd16: xpb[91] = 1024'd107601600924658274656079153504063138259444349444666471273619787469262338645738073457874100120860817544625518013870469021577285675625722103589062278892903601002713375617578514235836576968514068187220612041074245347607634058744612164925851483597562932831337600951109142363269394227832482508719084452927199681670;
            6'd17: xpb[91] = 1024'd98818364021933824147234234672465280307572317894241165212204542302969122893933060685239347476582409352484219213805186656103483050247177193243983655696668695948671627272480769208372583130106546733758125592592980701037566081138538328613094880112006934974943713083788831507210415357830933538374191002906950351233;
            6'd18: xpb[91] = 1024'd90035127119209373638389315840867422355700286343815859150789297136675907142128047912604594832304001160342920413739904290629680424868632282898905032500433790894629878927383024180908589291699025280295639144111716054467498103532464492300338276626450937118549825216468520651151436487829384568029297552886701020796;
            6'd19: xpb[91] = 1024'd81251890216484923129544397009269564403828254793390553089374051970382691390323035139969842188025592968201621613674621925155877799490087372553826409304198885840588130582285279153444595453291503826833152695630451407897430125926390655987581673140894939262155937349148209795092457617827835597684404102866451690359;
            6'd20: xpb[91] = 1024'd72468653313760472620699478177671706451956223242965247027958806804089475638518022367335089543747184776060322813609339559682075174111542462208747786107963980786546382237187534125980601614883982373370666247149186761327362148320316819674825069655338941405762049481827898939033478747826286627339510652846202359922;
            6'd21: xpb[91] = 1024'd63685416411036022111854559346073848500084191692539940966543561637796259886713009594700336899468776583919024013544057194208272548732997551863669162911729075732504633892089789098516607776476460919908179798667922114757294170714242983362068466169782943549368161614507588082974499877824737656994617202825953029485;
            6'd22: xpb[91] = 1024'd54902179508311571603009640514475990548212160142114634905128316471503044134907996822065584255190368391777725213478774828734469923354452641518590539715494170678462885546992044071052613938068939466445693350186657468187226193108169147049311862684226945692974273747187277226915521007823188686649723752805703699048;
            6'd23: xpb[91] = 1024'd46118942605587121094164721682878132596340128591689328843713071305209828383102984049430831610911960199636426413413492463260667297975907731173511916519259265624421137201894299043588620099661418012983206901705392821617158215502095310736555259198670947836580385879866966370856542137821639716304830302785454368611;
            6'd24: xpb[91] = 1024'd37335705702862670585319802851280274644468097041264022782297826138916612631297971276796078966633552007495127613348210097786864672597362820828433293323024360570379388856796554016124626261253896559520720453224128175047090237896021474423798655713114949980186498012546655514797563267820090745959936852765205038174;
            6'd25: xpb[91] = 1024'd28552468800138220076474884019682416692596065490838716720882580972623396879492958504161326322355143815353828813282927732313062047218817910483354670126789455516337640511698808988660632422846375106058234004742863528477022260289947638111042052227558952123792610145226344658738584397818541775615043402744955707737;
            6'd26: xpb[91] = 1024'd19769231897413769567629965188084558740724033940413410659467335806330181127687945731526573678076735623212530013217645366839259421840273000138276046930554550462295892166601063961196638584438853652595747556261598881906954282683873801798285448742002954267398722277906033802679605527816992805270149952724706377300;
            6'd27: xpb[91] = 1024'd10985994994689319058785046356486700788852002389988104598052090640036965375882932958891821033798327431071231213152363001365456796461728089793197423734319645408254143821503318933732644746031332199133261107780334235336886305077799965485528845256446956411004834410585722946620626657815443834925256502704457046863;
            6'd28: xpb[91] = 1024'd2202758091964868549940127524888842836979970839562798536636845473743749624077920186257068389519919238929932413087080635891654171083183179448118800538084740354212395476405573906268650907623810745670774659299069588766818327471726129172772241770890958554610946543265412090561647787813894864580363052684207716426;
            6'd29: xpb[91] = 1024'd117486216873365159439894136098105417629806366414873176603353455372427429209582046323637386959899185356231783020479291704996915386545858603658200302358180876233861321700879046216434896260733495013518485819205044788561111200086549065824994207968564409965036962090062159264609196991740978911354159429289552870320;
            6'd30: xpb[91] = 1024'd108702979970640708931049217266507559677934334864447870541938210206134213457777033551002634315620777164090484220414009339523112761167313693313121679161945971179819573355781301188970902422325973560055999370723780141991043222480475229512237604483008412108643074222741848408550218121739429941009265979269303539883;
            6'd31: xpb[91] = 1024'd99919743067916258422204298434909701726062303314022564480522965039840997705972020778367881671342368971949185420348726974049310135788768782968043055965711066125777825010683556161506908583918452106593512922242515495420975244874401393199481000997452414252249186355421537552491239251737880970664372529249054209446;
            6'd32: xpb[91] = 1024'd91136506165191807913359379603311843774190271763597258419107719873547781954167008005733129027063960779807886620283444608575507510410223872622964432769476161071736076665585811134042914745510930653131026473761250848850907267268327556886724397511896416395855298488101226696432260381736332000319479079228804879009;
            6'd33: xpb[91] = 1024'd82353269262467357404514460771713985822318240213171952357692474707254566202361995233098376382785552587666587820218162243101704885031678962277885809573241256017694328320488066106578920907103409199668540025279986202280839289662253720573967794026340418539461410620780915840373281511734783029974585629208555548572;
            6'd34: xpb[91] = 1024'd73570032359742906895669541940116127870446208662746646296277229540961350450556982460463623738507144395525289020152879877627902259653134051932807186377006350963652579975390321079114927068695887746206053576798721555710771312056179884261211190540784420683067522753460604984314302641733234059629692179188306218135;
            6'd35: xpb[91] = 1024'd64786795457018456386824623108518269918574177112321340234861984374668134698751969687828871094228736203383990220087597512154099634274589141587728563180771445909610831630292576051650933230288366292743567128317456909140703334450106047948454587055228422826673634886140294128255323771731685089284798729168056887698;
            6'd36: xpb[91] = 1024'd56003558554294005877979704276920411966702145561896034173446739208374918946946956915194118449950328011242691420022315146680297008896044231242649939984536540855569083285194831024186939391880844839281080679836192262570635356844032211635697983569672424970279747018819983272196344901730136118939905279147807557261;
            6'd37: xpb[91] = 1024'd47220321651569555369134785445322554014830114011470728112031494042081703195141944142559365805671919819101392619957032781206494383517499320897571316788301635801527334940097085996722945553473323385818594231354927616000567379237958375322941380084116427113885859151499672416137366031728587148595011829127558226824;
            6'd38: xpb[91] = 1024'd38437084748845104860289866613724696062958082461045422050616248875788487443336931369924613161393511626960093819891750415732691758138954410552492693592066730747485586594999340969258951715065801932356107782873662969430499401631884539010184776598560429257491971284179361560078387161727038178250118379107308896387;
            6'd39: xpb[91] = 1024'd29653847846120654351444947782126838111086050910620115989201003709495271691531918597289860517115103434818795019826468050258889132760409500207414070395831825693443838249901595941794957876658280478893621334392398322860431424025810702697428173113004431401098083416859050704019408291725489207905224929087059565950;
            6'd40: xpb[91] = 1024'd20870610943396203842600028950528980159214019360194809927785758543202055939726905824655107872836695242677496219761185684785086507381864589862335447199596920639402089904803850914330964038250759025431134885911133676290363446419736866384671569627448433544704195549538739847960429421723940237560331479066810235513;
            6'd41: xpb[91] = 1024'd12087374040671753333755110118931122207341987809769503866370513376908840187921893052020355228558287050536197419695903319311283882003319679517256824003362015585360341559706105886866970199843237571968648437429869029720295468813663030071914966141892435688310307682218428991901450551722391267215438029046560905076;
            6'd42: xpb[91] = 1024'd3304137137947302824910191287333264255469956259344197804955268210615624436116880279385602584279878858394898619630620953837481256624774769172178200807127110531318593214608360859402976361435716118506161988948604383150227491207589193759158362656336437831916419814898118135842471681720842296870544579026311574639;
            6'd43: xpb[91] = 1024'd118587595919347593714864199860549839048296351834654575871671878109299304021621006416765921154659144975696749227022832022942742472087450193382259702627223246410967519439081833169569221714545400386353873148854579582944520363822412130411380328854009889242342435361694865309890020885647926343644340955631656728533;
            6'd44: xpb[91] = 1024'd109804359016623143206019281028951981096424320284229269810256632943006088269815993644131168510380736783555450426957549657468939846708905283037181079430988341356925771093984088142105227876137878932891386700373314936374452386216338294098623725368453891385948547494374554453831042015646377373299447505611407398096;
            6'd45: xpb[91] = 1024'd101021122113898692697174362197354123144552288733803963748841387776712872518010980871496415866102328591414151626892267291995137221330360372692102456234753436302884022748886343114641234037730357479428900251892050289804384408610264457785867121882897893529554659627054243597772063145644828402954554055591158067659;
            6'd46: xpb[91] = 1024'd92237885211174242188329443365756265192680257183378657687426142610419656766205968098861663221823920399272852826826984926521334595951815462347023833038518531248842274403788598087177240199322836025966413803410785643234316431004190621473110518397341895673160771759733932741713084275643279432609660605570908737222;
            6'd47: xpb[91] = 1024'd83454648308449791679484524534158407240808225632953351626010897444126441014400955326226910577545512207131554026761702561047531970573270552001945209842283626194800526058690853059713246360915314572503927354929520996664248453398116785160353914911785897816766883892413621885654105405641730462264767155550659406785;
            6'd48: xpb[91] = 1024'd74671411405725341170639605702560549288936194082528045564595652277833225262595942553592157933267104014990255226696420195573729345194725641656866586646048721140758777713593108032249252522507793119041440906448256350094180475792042948847597311426229899960372996025093311029595126535640181491919873705530410076348;
            6'd49: xpb[91] = 1024'd65888174503000890661794686870962691337064162532102739503180407111540009510790929780957405288988695822848956426631137830099926719816180731311787963449813816086717029368495363004785258684100271665578954457966991703524112498185969112534840707940673902103979108157773000173536147665638632521574980255510160745911;
            6'd50: xpb[91] = 1024'd57104937600276440152949768039364833385192130981677433441765161945246793758985917008322652644710287630707657626565855464626124094437635820966709340253578911032675281023397617977321264845692750212116468009485727056954044520579895276222084104455117904247585220290452689317477168795637083551230086805489911415474;
            6'd51: xpb[91] = 1024'd48321700697551989644104849207766975433320099431252127380349916778953578007180904235687900000431879438566358826500573099152321469059090910621630717057344005978633532678299872949857271007285228758653981561004462410383976542973821439909327500969561906391191332423132378461418189925635534580885193355469662085037;
            6'd52: xpb[91] = 1024'd39538463794827539135259930376169117481448067880826821318934671612660362255375891463053147356153471246425060026435290733678518843680546000276552093861109100924591784333202127922393277168877707305191495112523197763813908565367747603596570897484005908534797444555812067605359211055633985610540299905449412754600;
            6'd53: xpb[91] = 1024'd30755226892103088626415011544571259529576036330401515257519426446367146503570878690418394711875063054283761226370008368204716218302001089931473470664874195870550035988104382894929283330470185851729008664041933117243840587761673767283814293998449910678403556688491756749300232185632436640195406455429163424163;
            6'd54: xpb[91] = 1024'd21971989989378638117570092712973401577704004779976209196104181280073930751765865917783642067596654862142462426304726002730913592923456179586394847468639290816508287643006637867465289492062664398266522215560668470673772610155599930971057690512893912822009668821171445893241253315630887669850513005408914093726;
            6'd55: xpb[91] = 1024'd13188753086654187608725173881375543625831973229550903134688936113780714999960853145148889423318246670001163626239443637257110967544911269241316224272404385762466539297908892840001295653655142944804035767079403824103704632549526094658301087027337914965615780953851135037182274445629338699505619555388664763289;
            6'd56: xpb[91] = 1024'd4405516183929737099880255049777685673959941679125597073273690947487499248155840372514136779039838477859864826174161271783308342166366358896237601076169480708424790952811147812537301815247621491341549318598139177533636654943452258345544483541781917109221893086530824181123295575627789729160726105368415432852;
            6'd57: xpb[91] = 1024'd119688974965330027989834263622994260466786337254435975139990300846171178833659966509894455349419104595161715433566372340888569557629041783106319102896265616588073717177284620122703547168357305759189260478504114377327929527558275194997766449739455368519647908633327571355170844779554873775934522481973760586746;
            6'd58: xpb[91] = 1024'd110905738062605577480989344791396402514914305704010669078575055679877963081854953737259702705140696403020416633501089975414766932250496872761240479700030711534031968832186875095239553329949784305726774030022849730757861549952201358685009846253899370663254020766007260499111865909553324805589629031953511256309;
            6'd59: xpb[91] = 1024'd102122501159881126972144425959798544563042274153585363017159810513584747330049940964624950060862288210879117833435807609940964306871951962416161856503795806479990220487089130067775559491542262852264287581541585084187793572346127522372253242768343372806860132898686949643052887039551775835244735581933261925872;
            6'd60: xpb[91] = 1024'd93339264257156676463299507128200686611170242603160056955744565347291531578244928191990197416583880018737819033370525244467161681493407052071083233307560901425948472141991385040311565653134741398801801133060320437617725594740053686059496639282787374950466245031366638786993908169550226864899842131913012595435;
            6'd61: xpb[91] = 1024'd84556027354432225954454588296602828659298211052734750894329320180998315826439915419355444772305471826596520233305242878993359056114862141726004610111325996371906723796893640012847571814727219945339314684579055791047657617133979849746740035797231377094072357164046327930934929299548677894554948681892763264998;
            6'd62: xpb[91] = 1024'd75772790451707775445609669465004970707426179502309444832914075014705100074634902646720692128027063634455221433239960513519556430736317231380925986915091091317864975451795894985383577976319698491876828236097791144477589639527906013433983432311675379237678469296726017074875950429547128924210055231872513934561;
            6'd63: xpb[91] = 1024'd66989553548983324936764750633407112755554147951884138771498829848411884322829889874085939483748655442313922633174678148045753805357772321035847363718856186263823227106698149957919584137912177038414341787616526497907521661921832177121226828826119381381284581429405706218816971559545579953865161781852264604124;
        endcase
    end

    always_comb begin
        case(flag[30][16:12])
            5'd0: xpb[92] = 1024'd0;
            5'd1: xpb[92] = 1024'd58206316646258874427919831801809254803682116401458832710083584682118668571024877101451186839470247250172623833109395782571951179979227410690768740522621281209781478761600404930455590299504655584951855339135261851337453684315758340808470225340563383524890693562085395362757992689544030983520268331832015273687;
            5'd2: xpb[92] = 1024'd116412633292517748855839663603618509607364232802917665420167169364237337142049754202902373678940494500345247666218791565143902359958454821381537481045242562419562957523200809860911180599009311169903710678270523702674907368631516681616940450681126767049781387124170790725515985379088061967040536663664030547374;
            5'd3: xpb[92] = 1024'd50552254254651881884960568000613331666347922078640814002118898981379110375765492394338489303753067441074722091870693913136789699096461897517146096551532802695653761715229997453736531706996761033545368409018545707648000202726378249460432106338460701307852177272139128058167449994703459933442115168870451336730;
            5'd4: xpb[92] = 1024'd108758570900910756312880399802422586470030038480099646712202483663497778946790369495789676143223314691247345924980089695708740879075689308207914837074154083905435240476830402384192122006501416618497223748153807558985453887042136590268902331679024084832742870834224523420925442684247490916962383500702466610417;
            5'd5: xpb[92] = 1024'd42898191863044889342001304199417408529013727755822795294154213280639552180506107687225791768035887631976820350631992043701628218213696384343523452580444324181526044668859589977017473114488866482138881478901829563958546721136998158112393987336358019090813660982192860753576907299862888883363962005908887399773;
            5'd6: xpb[92] = 1024'd101104508509303763769921136001226663332695844157281628004237797962758220751530984788676978607506134882149444183741387826273579398192923795034292193103065605391307523430459994907473063413993522067090736818037091415296000405452756498920864212676921402615704354544278256116334899989406919866884230337740902673460;
            5'd7: xpb[92] = 1024'd35244129471437896799042040398221485391679533433004776586189527579899993985246722980113094232318707822878918609393290174266466737330930871169900808609355845667398327622489182500298414521980971930732394548785113420269093239547618066764355868334255336873775144692246593448986364605022317833285808842947323462816;
            5'd8: xpb[92] = 1024'd93450446117696771226961872200030740195361649834463609296273112262018662556271600081564281071788955073051542442502685956838417917310158281860669549131977126877179806384089587430754004821485627515684249887920375271606546923863376407572826093674818720398665838254331988811744357294566348816806077174779338736503;
            5'd9: xpb[92] = 1024'd27590067079830904256082776597025562254345339110186757878224841879160435789987338273000396696601528013781016868154588304831305256448165357996278164638267367153270610576118775023579355929473077379325907618668397276579639757958237975416317749332152654656736628402300326144395821910181746783207655679985759525859;
            5'd10: xpb[92] = 1024'd85796383726089778684002608398834817058027455511645590588308426561279104361012215374451583536071775263953640701263984087403256436427392768687046905160888648363052089337719179954034946228977732964277762957803659127917093442273996316224787974672716038181627321964385721507153814599725777766727924011817774799546;
            5'd11: xpb[92] = 1024'd19936004688223911713123512795829639117011144787368739170260156178420877594727953565887699160884348204683115126915886435396143775565399844822655520667178888639142893529748367546860297336965182827919420688551681132890186276368857884068279630330049972439698112112354058839805279215341175733129502517024195588902;
            5'd12: xpb[92] = 1024'd78142321334482786141043344597638893920693261188827571880343740860539546165752830667338886000354595454855738960025282217968094955544627255513424261189800169848924372291348772477315887636469838412871276027686942984227639960684616224876749855670613355964588805674439454202563271904885206716649770848856210862589;
            5'd13: xpb[92] = 1024'd12281942296616919170164248994633715979676950464550720462295470477681319399468568858775001625167168395585213385677184565960982294682634331649032876696090410125015176483377960070141238744457288276512933758434964989200732794779477792720241511327947290222659595822407791535214736520500604683051349354062631651945;
            5'd14: xpb[92] = 1024'd70488258942875793598084080796442970783359066866009553172379055159799987970493445960226188464637415645757837218786580348532933474661861742339801617218711691334796655244978365000596829043961943861464789097570226840538186479095236133528711736668510673747550289384493186897972729210044635666571617685894646925632;
            5'd15: xpb[92] = 1024'd4627879905009926627204985193437792842342756141732701754330784776941761204209184151662304089449988586487311644438482696525820813799868818475410232725001931610887459437007552593422180151949393725106446828318248845511279313190097701372203392325844608005621079532461524230624193825660033632973196191101067714988;
            5'd16: xpb[92] = 1024'd62834196551268801055124816995247047646024872543191534464414369459060429775234061253113490928920235836659935477547878479097771993779096229166178973247623212820668938198607957523877770451454049310058302167453510696848732997505856042180673617666407991530511773094546919593382186515204064616493464522933082988675;
            5'd17: xpb[92] = 1024'd121040513197527675483044648797056302449706988944650367174497954141179098346258938354564677768390483086832559310657274261669723173758323639856947713770244494030450416960208362454333360750958704895010157506588772548186186681821614382989143843006971375055402466656632314956140179204748095600013732854765098262362;
            5'd18: xpb[92] = 1024'd55180134159661808512165553194051124508690678220373515756449683758320871579974676546000793393203056027562033736309176609662610512896330715992556329276534734306541221152237550047158711858946154758651815237336794553159279515916475950832635498664305309313473256804600652288791643820363493566415311359971519051718;
            5'd19: xpb[92] = 1024'd113386450805920682940085384995860379312372794621832348466533268440439540150999553647451980232673303277734657569418572392234561692875558126683325069799156015516322699913837954977614302158450810343603670576472056404496733200232234291641105724004868692838363950366686047651549636509907524549935579691803534325405;
            5'd20: xpb[92] = 1024'd47526071768054815969206289392855201371356483897555497048484998057581313384715291838888095857485876218464131995070474740227449032013565202818933685305446255792413504105867142570439653266438260207245328307220078409469826034327095859484597379662202627096434740514654384984201101125522922516337158197009955114761;
            5'd21: xpb[92] = 1024'd105732388414313690397126121194664456175038600299014329758568582739699981955740168940339282696956123468636755828179870522799400211992792613509702425828067537002194982867467547500895243565942915792197183646355340260807279718642854200293067605002766010621325434076739780346959093815066953499857426528841970388448;
            5'd22: xpb[92] = 1024'd39872009376447823426247025591659278234022289574737478340520312356841755189455907131775398321768696409366230253831772870792287551130799689645311041334357777278285787059496735093720594673930365655838841377103362265780372552737715768136559260660099944879396224224708117679610558430682351466259005034048391177804;
            5'd23: xpb[92] = 1024'd98078326022706697854166857393468533037704405976196311050603897038960423760480784233226585161238943659538854086941168653364238731110027100336079781856979058488067265821097140024176184973435021240790696716238624117117826237053474108945029486000663328404286917786793513042368551120226382449779273365880406451491;
            5'd24: xpb[92] = 1024'd32217946984840830883287761790463355096688095251919459632555626656102196994196522424662700786051516600268328512593071001357126070248034176471688397363269298764158070013126327617001536081422471104432354446986646122090919071148335676788521141657997262662357707934761850375020015735841780416180851871086827240847;
            5'd25: xpb[92] = 1024'd90424263631099705311207593592272609900370211653378292342639211338220865565221399526113887625521763850440952345702466783929077250227261587162457137885890579973939548774726732547457126380927126689384209786121907973428372755464094017596991366998560646187248401496847245737778008425385811399701120202918842514534;
            5'd26: xpb[92] = 1024'd24563884593233838340328497989267431959353900929101440924590940955362638798937137717550003250334336791170426771354369131921964589365268663298065753392180820250030352966755920140282477488914576553025867516869929978401465589558955585440483022655894580445319191644815583070429473041001209366102698708125263303890;
            5'd27: xpb[92] = 1024'd82770201239492712768248329791076686763036017330560273634674525637481307369962014819001190089804584041343050604463764914493915769344496073988834493914802101459811831728356325070738067788419232137977722856005191829738919273874713926248953247996457963970209885206900978433187465730545240349622967039957278577577;
            5'd28: xpb[92] = 1024'd16909822201626845797369234188071508822019706606283422216626255254623080603677753010437305714617156982072525030115667262486803108482503150124443109421092341735902635920385512663563418896406682001619380586753213834712012107969575494092444903653791898228280675354869315765838930346160638316024545545163699366933;
            5'd29: xpb[92] = 1024'd75116138847885720225289065989880763625701823007742254926709839936741749174702630111888492554087404232245148863225063045058754288461730560815211849943713622945684114681985917594019009195911337586571235925888475686049465792285333834900915128994355281753171368916954711128596923035704669299544813876995714640620;
            5'd30: xpb[92] = 1024'd9255759810019853254409970386875585684685512283465403508661569553883522408418368303324608178899977172974623288876965393051641627599737636950820465450003863221774918874015105186844360303898787450212893656636497691022558626380195402744406784651689216011242159064923048461248387651320067265946392382202135429976;
            5'd31: xpb[92] = 1024'd67462076456278727682329802188684840488367628684924236218745154236002190979443245404775795018370224423147247121986361175623592807578965047641589205972625144431556397635615510117299950603403443035164748995771759542360012310695953743552877009992252599536132852627008443824006380340864098249466660714034150703663;
        endcase
    end

    always_comb begin
        case(flag[31][5:0])
            6'd0: xpb[93] = 1024'd0;
            6'd1: xpb[93] = 1024'd62834196551268801055124816995247047646024872543191534464414369459060429775234061253113490928920235836659935477547878479097771993779096229166178973247623212820668938198607957523877770451454049310058302167453510696848732997505856042180673617666407991530511773094546919593382186515204064616493464522933082988675;
            6'd2: xpb[93] = 1024'd1601697418412860711450706585679662547351317960647384800696883853143964213158983596211910643182797363876721547638263523616480146716972123777197821478915384707647201827644697710125301711390892898806406726519781547333105144790815311396368665649586533794203642774976781156657844956479496215868239219240571493019;
            6'd3: xpb[93] = 1024'd64435893969681661766575523580926710193376190503838919265111253312204393988393044849325401572103033200536657025186142002714252140496068352943376794726538597528316140026252655234003072162844942208864708893973292244181838142296671353577042283315994525324715415869523700750040031471683560832361703742173654481694;
            6'd4: xpb[93] = 1024'd3203394836825721422901413171359325094702635921294769601393767706287928426317967192423821286365594727753443095276527047232960293433944247554395642957830769415294403655289395420250603422781785797612813453039563094666210289581630622792737331299173067588407285549953562313315689912958992431736478438481142986038;
            6'd5: xpb[93] = 1024'd66037591388094522478026230166606372740727508464486304065808137165348358201552028445537312215285830564413378572824405526330732287213040476720574616205453982235963341853897352944128373874235835107671115620493073791514943287087486664973410948965581059118919058644500481906697876428163057048229942961414225974713;
            6'd6: xpb[93] = 1024'd4805092255238582134352119757038987642053953881942154402090651559431892639476950788635731929548392091630164642914790570849440440150916371331593464436746154122941605482934093130375905134172678696419220179559344641999315434372445934189105996948759601382610928324930343469973534869438488647604717657721714479057;
            6'd7: xpb[93] = 1024'd67639288806507383189476936752286035288078826425133688866505021018492322414711012041749222858468627928290100120462669049947212433930012600497772437684369366943610543681542050654253675585626728006477522347012855338848048431878301976369779614615167592913122701419477263063355721384642553264098182180654797467732;
            6'd8: xpb[93] = 1024'd6406789673651442845802826342718650189405271842589539202787535412575856852635934384847642572731189455506886190553054094465920586867888495108791285915661538830588807310578790840501206845563571595225626906079126189332420579163261245585474662598346135176814571099907124626631379825917984863472956876962285972076;
            6'd9: xpb[93] = 1024'd69240986224920243900927643337965697835430144385781073667201904871636286627869995637961133501651425292166821668100932573563692580646984724274970259163284751651257745509186748364378977297017620905283929073532636886181153576669117287766148280264754126707326344194454044220013566341122049479966421399895368960751;
            6'd10: xpb[93] = 1024'd8008487092064303557253532928398312736756589803236924003484419265719821065794917981059553215913986819383607738191317618082400733584860618885989107394576923538236009138223488550626508556954464494032033632598907736665525723954076556981843328247932668971018213874883905783289224782397481079341196096202857465095;
            6'd11: xpb[93] = 1024'd70842683643333104612378349923645360382781462346428458467898788724780250841028979234173044144834222656043543215739196097180172727363956848052168080642200136358904947336831446074504279008408513804090335800052418433514258721459932599162516945914340660501529986969430825376671411297601545695834660619135940453770;
            6'd12: xpb[93] = 1024'd9610184510477164268704239514077975284107907763884308804181303118863785278953901577271463859096784183260329285829581141698880880301832742663186928873492308245883210965868186260751810268345357392838440359118689283998630868744891868378211993897519202765221856649860686939947069738876977295209435315443428958114;
            6'd13: xpb[93] = 1024'd72444381061745965323829056509325022930132780307075843268595672577924215054187962830384954788017020019920264763377459620796652874080928971829365902121115521066552149164476143784629580719799406702896742526572199980847363866250747910558885611563927194295733629744407606533329256254081041911702899838376511946789;
            6'd14: xpb[93] = 1024'd11211881928890024980154946099757637831459225724531693604878186972007749492112885173483374502279581547137050833467844665315361027018804866440384750352407692953530412793512883970877111979736250291644847085638470831331736013535707179774580659547105736559425499424837468096604914695356473511077674534684000451133;
            6'd15: xpb[93] = 1024'd74046078480158826035279763095004685477484098267723228069292556431068179267346946426596865431199817383796986311015723144413133020797901095606563723600030905774199350992120841494754882431190299601703149253091981528180469011041563221955254277213513728089937272519384387689987101210560538127571139057617083439808;
            6'd16: xpb[93] = 1024'd12813579347302885691605652685437300378810543685179078405575070825151713705271868769695285145462378911013772381106108188931841173735776990217582571831323077661177614621157581681002413691127143190451253812158252378664841158326522491170949325196692270353629142199814249253262759651835969726945913753924571944152;
            6'd17: xpb[93] = 1024'd75647775898571686746730469680684348024835416228370612869989440284212143480505930022808776074382614747673707858653986668029613167514873219383761545078946290481846552819765539204880184142581192500509555979611763075513574155832378533351622942863100261884140915294361168846644946167040034343439378276857654932827;
            6'd18: xpb[93] = 1024'd14415276765715746403056359271116962926161861645826463206271954678295677918430852365907195788645176274890493928744371712548321320452749113994780393310238462368824816448802279391127715402518036089257660538678033925997946303117337802567317990846278804147832784974791030409920604608315465942814152973165143437171;
            6'd19: xpb[93] = 1024'd77249473316984547458181176266364010572186734189017997670686324137356107693664913619020686717565412111550429406292250191646093314231845343160959366557861675189493754647410236915005485853972085399315962706131544622846679300623193844747991608512686795678344558069337950003302791123519530559307617496098226425846;
            6'd20: xpb[93] = 1024'd16016974184128607114507065856796625473513179606473848006968838531439642131589835962119106431827973638767215476382635236164801467169721237771978214789153847076472018276446977101253017113908928988064067265197815473331051447908153113963686656495865337942036427749767811566578449564794962158682392192405714930190;
            6'd21: xpb[93] = 1024'd78851170735397408169631882852043673119538052149665382471383207990500071906823897215232597360748209475427150953930513715262573460948817466938157188036777059897140956475054934625130787565362978298122369432651326170179784445414009156144360274162273329472548200844314731159960636079999026775175856715338797918865;
            6'd22: xpb[93] = 1024'd17618671602541467825957772442476288020864497567121232807665722384583606344748819558331017075010771002643937024020898759781281613886693361549176036268069231784119220104091674811378318825299821886870473991717597020664156592698968425360055322145451871736240070524744592723236294521274458374550631411646286423209;
            6'd23: xpb[93] = 1024'd80452868153810268881082589437723335666889370110312767272080091843644036119982880811444508003931006839303872501568777238879053607665789590715355009515692444604788158302699632335256089276753871196928776159171107717512889590204824467540728939811859863266751843619291512316618481036478522991044095934579369411884;
            6'd24: xpb[93] = 1024'd19220369020954328537408479028155950568215815527768617608362606237727570557907803154542927718193568366520658571659162283397761760603665485326373857746984616491766421931736372521503620536690714785676880718237378567997261737489783736756423987795038405530443713299721373879894139477753954590418870630886857916228;
            6'd25: xpb[93] = 1024'd82054565572223129592533296023402998214240688070960152072776975696788000333141864407656418647113804203180594049207040762495533754382761714492552830994607829312435360130344330045381390988144764095735182885690889264845994734995639778937097605461446397060955486394268293473276325992958019206912335153819940904903;
            6'd26: xpb[93] = 1024'd20822066439367189248859185613835613115567133488416002409059490090871534771066786750754838361376365730397380119297425807014241907320637609103571679225900001199413623759381070231628922248081607684483287444757160115330366882280599048152792653444624939324647356074698155036551984434233450806287109850127429409247;
            6'd27: xpb[93] = 1024'd83656262990635990303984002609082660761592006031607536873473859549931964546300848003868329290296601567057315596845304286112013901099733838269750652473523214020082561957989027755506692699535656994541589612210670812179099879786455090333466271111032930855159129169245074629934170949437515422780574373060512397922;
            6'd28: xpb[93] = 1024'd22423763857780049960309892199515275662918451449063387209756373944015498984225770346966749004559163094274101666935689330630722054037609732880769500704815385907060825587025767941754223959472500583289694171276941662663472027071414359549161319094211473118850998849674936193209829390712947022155349069368000902266;
            6'd29: xpb[93] = 1024'd85257960409048851015434709194762323308943323992254921674170743403075928759459831600080239933479398930934037144483567809728494047816705962046948473952438598727729763785633725465631994410926549893347996338730452359512205024577270401729834936760619464649362771944221855786592015905917011638648813592301083890941;
            6'd30: xpb[93] = 1024'd24025461276192910671760598785194938210269769409710772010453257797159463197384753943178659647741960458150823214573952854247202200754581856657967322183730770614708027414670465651879525670863393482096100897796723209996577171862229670945529984743798006913054641624651717349867674347192443238023588288608572395285;
            6'd31: xpb[93] = 1024'd86859657827461711726885415780441985856294641952902306474867627256219892972618815196292150576662196294810758692121831333344974194533678085824146295431353983435376965613278423175757296122317442792154403065250233906845310169368085713126203602410205998443566414719198636943249860862396507854517052811541655383960;
            6'd32: xpb[93] = 1024'd25627158694605771383211305370874600757621087370358156811150141650303427410543737539390570290924757822027544762212216377863682347471553980435165143662646155322355229242315163362004827382254286380902507624316504757329682316653044982341898650393384540707258284399628498506525519303671939453891827507849143888304;
            6'd33: xpb[93] = 1024'd88461355245874572438336122366121648403645959913549691275564511109363857185777798792504061219844993658687480239760094856961454341250650209601344116910269368143024167440923120885882597833708335690960809791770015454178415314158901024522572268059792532237770057494175418099907705818876004070385292030782226876979;
            6'd34: xpb[93] = 1024'd27228856113018632094662011956554263304972405331005541611847025503447391623702721135602480934107555185904266309850479901480162494188526104212362965141561540030002431069959861072130129093645179279708914350836286304662787461443860293738267316042971074501461927174605279663183364260151435669760066727089715381323;
            6'd35: xpb[93] = 1024'd90063052664287433149786828951801310950997277874197076076261394962507821398936782388715971863027791022564201787398358380577934487967622333378541938389184752850671369268567818596007899545099228589767216518289797001511520458949716335918940933709379066031973700269152199256565550775355500286253531250022798369998;
            6'd36: xpb[93] = 1024'd28830553531431492806112718542233925852323723291652926412543909356591355836861704731814391577290352549780987857488743425096642640905498227989560786620476924737649632897604558782255430805036072178515321077356067851995892606234675605134635981692557608295665569949582060819841209216630931885628305946330286874342;
            6'd37: xpb[93] = 1024'd91664750082700293861237535537480973498348595834844460876958278815651785612095765984927882506210588386440923335036621904194414634684594457155739759868100137558318571096212516306133201256490121488573623244809578548844625603740531647315309599358965599826177343044128980413223395731834996502121770469263369863017;
            6'd38: xpb[93] = 1024'd30432250949844353517563425127913588399675041252300311213240793209735320050020688328026302220473149913657709405127006948713122787622470351766758608099392309445296834725249256492380732516426965077321727803875849399328997751025490916531004647342144142089869212724558841976499054173110428101496545165570858367361;
            6'd39: xpb[93] = 1024'd93266447501113154572688242123160636045699913795491845677655162668795749825254749581139793149393385750317644882674885427810894781401566580932937581347015522265965772923857214016258502967881014387380029971329360096177730748531346958711678265008552133620380985819105761569881240688314492717990009688503941356036;
            6'd40: xpb[93] = 1024'd32033948368257214229014131713593250947026359212947696013937677062879284263179671924238212863655947277534430952765270472329602934339442475543956429578307694152944036552893954202506034227817857976128134530395630946662102895816306227927373312991730675884072855499535623133156899129589924317364784384811429860380;
            6'd41: xpb[93] = 1024'd94868144919526015284138948708840298593051231756139230478352046521939714038413733177351703792576183114194366430313148951427374928118538704710135402825930906973612974751501911726383804679271907286186436697849141643510835893322162270108046930658138667414584628594082542726539085644793988933858248907744512849055;
            6'd42: xpb[93] = 1024'd33635645786670074940464838299272913494377677173595080814634560916023248476338655520450123506838744641411152500403533995946083081056414599321154251057223078860591238380538651912631335939208750874934541256915412493995208040607121539323741978641317209678276498274512404289814744086069420533233023604052001353399;
            6'd43: xpb[93] = 1024'd96469842337938875995589655294519961140402549716786615279048930375083678251572716773563614435758980478071087977951412475043855074835510828487333224304846291681260176579146609436509106390662800184992843424368923190843941038112977581504415596307725201208788271369059323883196930601273485149726488126985084342074;
            6'd44: xpb[93] = 1024'd35237343205082935651915544884952576041728995134242465615331444769167212689497639116662034150021542005287874048041797519562563227773386723098352072536138463568238440208183349622756637650599643773740947983435194041328313185397936850720110644290903743472480141049489185446472589042548916749101262823292572846418;
            6'd45: xpb[93] = 1024'd98071539756351736707040361880199623687753867677434000079745814228227642464731700369775525078941777841947809525589675998660335221552482952264531045783761676388907378406791307146634408102053693083799250150888704738177046182903792892900784261957311735002991914144036105039854775557752981365594727346225655835093;
            6'd46: xpb[93] = 1024'd36839040623495796363366251470632238589080313094889850416028328622311176902656622712873944793204339369164595595680061043179043374490358846875549894015053848275885642035828047332881939361990536672547354709954975588661418330188752162116479309940490277266683783824465966603130433999028412964969502042533144339437;
            6'd47: xpb[93] = 1024'd99673237174764597418491068465879286235105185638081384880442698081371606677890683965987435722124575205824531073227939522276815368269455076041728867262677061096554580234436004856759709813444585982605656877408486285510151327694608204297152927606898268797195556919012886196512620514232477581462966565466227328112;
            6'd48: xpb[93] = 1024'd38440738041908657074816958056311901136431631055537235216725212475455141115815606309085855436387136733041317143318324566795523521207330970652747715493969232983532843863472745043007241073381429571353761436474757135994523474979567473512847975590076811060887426599442747759788278955507909180837741261773715832456;
            6'd49: xpb[93] = 1024'd101274934593177458129941775051558948782456503598728769681139581934515570891049667562199346365307372569701252620866203045893295514986427199818926688741592445804201782062080702566885011524835478881412063603928267832843256472485423515693521593256484802591399199693989667353170465470711973797331205784706798821131;
            6'd50: xpb[93] = 1024'd40042435460321517786267664641991563683782949016184620017422096328599105328974589905297766079569934096918038690956588090412003667924303094429945536972884617691180045691117442753132542784772322470160168162994538683327628619770382784909216641239663344855091069374419528916446123911987405396705980481014287325475;
            6'd51: xpb[93] = 1024'd102876632011590318841392481637238611329807821559376154481836465787659535104208651158411257008490169933577974168504466569509775661703399323596124510220507830511848983889725400277010313236226371780218470330448049380176361617276238827089890258906071336385602842468966448509828310427191470013199445003947370314150;
            6'd52: xpb[93] = 1024'd41644132878734378497718371227671226231134266976832004818118980181743069542133573501509676722752731460794760238594851614028483814641275218207143358451800002398827247518762140463257844496163215368966574889514320230660733764561198096305585306889249878649294712149396310073103968868466901612574219700254858818494;
            6'd53: xpb[93] = 1024'd104478329430003179552843188222918273877159139520023539282533349640803499317367634754623167651672967297454695716142730093126255808420371447373322331699423215219496185717370097987135614947617264679024877056967830927509466762067054138486258924555657870179806485243943229666486155383670966229067684223187941807169;
            6'd54: xpb[93] = 1024'd43245830297147239209169077813350888778485584937479389618815864034887033755292557097721587365935528824671481786233115137644963961358247341984341179930715387106474449346406838173383146207554108267772981616034101777993838909352013407701953972538836412443498354924373091229761813824946397828442458919495430311513;
            6'd55: xpb[93] = 1024'd106080026848416040264293894808597936424510457480670924083230233493947463530526618350835078294855764661331417263780993616742735955137343571150520153178338599927143387545014795697260916659008157577831283783487612474842571906857869449882627590205244403974010128018920010823144000340150462444935923442428513300188;
            6'd56: xpb[93] = 1024'd44847527715560099920619784399030551325836902898126774419512747888030997968451540693933498009118326188548203333871378661261444108075219465761539001409630771814121651174051535883508447918945001166579388342553883325326944054142828719098322638188422946237701997699349872386419658781425894044310698138736001804532;
            6'd57: xpb[93] = 1024'd107681724266828900975744601394277598971861775441318308883927117347091427743685601947046988938038562025208138811419257140359216101854315694927717974657253984634790589372659493407386218370399050476637690510007394022175677051648684761278996255854830937768213770793896791979801845296629958660804162661669084793207;
            6'd58: xpb[93] = 1024'd46449225133972960632070490984710213873188220858774159220209631741174962181610524290145408652301123552424924881509642184877924254792191589538736822888546156521768853001696233593633749630335894065385795069073664872660049198933644030494691303838009480031905640474326653543077503737905390260178937357976573297551;
            6'd59: xpb[93] = 1024'd109283421685241761687195307979957261519213093401965693684624001200235391956844585543258899581221359389084860359057520663975696248571287818704915796136169369342437791200304191117511520081789943375444097236527175569508782196439500072675364921504417471562417413568873573136459690253109454876672401880909656286226;
            6'd60: xpb[93] = 1024'd48050922552385821343521197570389876420539538819421544020906515594318926394769507886357319295483920916301646429147905708494404401509163713315934644367461541229416054829340931303759051341726786964192201795593446419993154343724459341891059969487596013826109283249303434699735348694384886476047176577217144790570;
            6'd61: xpb[93] = 1024'd110885119103654622398646014565636924066564411362613078485320885053379356170003569139470810224404156752961581906695784187592176395288259942482113617615084754050084993027948888827636821793180836274250503963046957116841887341230315384071733587154004005356621056343850354293117535209588951092540641100150227779245;
            6'd62: xpb[93] = 1024'd49652619970798682054971904156069538967890856780068928821603399447462890607928491482569229938666718280178367976786169232110884548226135837093132465846376925937063256656985629013884353053117679862998608522113227967326259488515274653287428635137182547620312926024280215856393193650864382691915415796457716283589;
            6'd63: xpb[93] = 1024'd112486816522067483110096721151316586613915729323260463286017768906523320383162552735682720867586954116838303454334047711208656542005232066259311439094000138757732194855593586537762123504571729173056910689566738664174992486021130695468102252803590539150824699118827135449775380166068447308408880319390799272264;
        endcase
    end

    always_comb begin
        case(flag[31][11:6])
            6'd0: xpb[94] = 1024'd0;
            6'd1: xpb[94] = 1024'd51254317389211542766422610741749201515242174740716313622300283300606854821087475078781140581849515644055089524424432755727364694943107960870330287325292310644710458484630326724009654764508572761805015248633009514659364633306089964683797300786769081414516568799256997013051038607343878907783655015698287776608;
            6'd2: xpb[94] = 1024'd102508634778423085532845221483498403030484349481432627244600566601213709642174950157562281163699031288110179048848865511454729389886215921740660574650584621289420916969260653448019309529017145523610030497266019029318729266612179929367594601573538162829033137598513994026102077214687757815567310031396575553216;
            6'd3: xpb[94] = 1024'd29696256483509886900468904820433171801028097096413256738768994836843669125953286326328350530890872622722119165815804832603030243988103548055830736959545891000440700884319762834398725102008512564104848137511788697613733049697373121086413332677077794976729802983653933009046587748103003706232275220469268845493;
            6'd4: xpb[94] = 1024'd80950573872721429666891515562182373316270271837129570361069278137450523947040761405109491112740388266777208690240237588330394938931211508926161024284838201645151159368950089558408379866517085325909863386144798212273097683003463085770210633463846876391246371782910930022097626355446882614015930236167556622101;
            6'd5: xpb[94] = 1024'd8138195577808231034515198899117142086814019452110199855237706373080483430819097573875560479932229601389148807207176909478695793033099135241331186593799471356170943284009198944787795439508452366404681026390567880568101466088656277489029364567386508538943037168050869005042136888862128504680895425240249914378;
            6'd6: xpb[94] = 1024'd59392512967019773800937809640866343602056194192826513477537989673687338251906572652656701061781745245444238331631609665206060487976207096111661473919091782000881401768639525668797450204017025128209696275023577395227466099394746242172826665354155589953459605967307866018093175496206007412464550440938537690986;
            6'd7: xpb[94] = 1024'd110646830356231316567360420382615545117298368933542827099838272974294193072994047731437841643631260889499327856056042420933425182919315056981991761244384092645591860253269852392807104968525597890014711523656586909886830732700836206856623966140924671367976174766564863031144214103549886320248205456636825467594;
            6'd8: xpb[94] = 1024'd37834452061318117934984103719550313887842116548523456594006701209924152556772383900203911010823102224111267973022981742081726037021202683297161923553345362356611644168328961779186520541516964930509529163902356578181834515786029398575442697244464303515672840151704802014088724636965132210913170645709518759871;
            6'd9: xpb[94] = 1024'd89088769450529660701406714461299515403084291289239770216306984510531007377859858978985051592672617868166357497447414497809090731964310644167492210878637673001322102652959288503196175306025537692314544412535366092841199149092119363259239998031233384930189408950961799027139763244309011118696825661407806536479;
            6'd10: xpb[94] = 1024'd16276391155616462069030397798234284173628038904220399710475412746160966861638195147751120959864459202778297614414353818957391586066198270482662373187598942712341886568018397889575590879016904732809362052781135761136202932177312554978058729134773017077886074336101738010084273777724257009361790850480499828756;
            6'd11: xpb[94] = 1024'd67530708544828004835453008539983485688870213644936713332775696046767821682725670226532261541713974846833387138838786574684756281009306231352992660512891253357052345052648724613585245643525477494614377301414145275795567565483402519661856029921542098492402643135358735023135312385068135917145445866178787605364;
            6'd12: xpb[94] = 1024'd118785025934039547601875619281732687204112388385653026955075979347374676503813145305313402123563490490888476663263219330412120975952414192223322947838183564001762803537279051337594900408034050256419392550047154790454932198789492484345653330708311179906919211934615732036186350992412014824929100881877075381972;
            6'd13: xpb[94] = 1024'd45972647639126348969499302618667455974656136000633656449244407583004635987591481474079471490755331825500416780230158651560421830054301818538493110147144833712782587452338160723974315981025417296914210190292924458749935981874685676064472061811850812054615877319755671019130861525827260715594066070949768674249;
            6'd14: xpb[94] = 1024'd97226965028337891735921913360416657489898310741349970071544690883611490808678956552860612072604847469555506304654591407287786524997409779408823397472437144357493045936968487447983970745533990058719225438925933973409300615180775640748269362598619893469132446119012668032181900133171139623377721086648056450857;
            6'd15: xpb[94] = 1024'd24414586733424693103545596697351426260442058356330599565713119119241450292457292721626681439796688804167446421621530728436087379099297405723993559781398414068512829852027596834363386318525357099214043079171703641704304398265968832467088093702159525616829111504152607015126410666586385514042686275720749743134;
            6'd16: xpb[94] = 1024'd75668904122636235869968207439100627775684233097046913188013402419848305113544767800407822021646204448222535946045963484163452074042405366594323847106690724713223288336657923558373041083033929861019058327804713156363669031572058797150885394488928607031345680303409604028177449273930264421826341291419037519742;
            6'd17: xpb[94] = 1024'd2856525827723037237591890776035396546227980712027542682181830655478264597323103969173891388838045782834476063012902805311752928144292992909494009415651994424243072251717032944752456656025296901513875968050482824658672814657251988869704125592468239179042345688549543011121959807345510312491306480491730812019;
            6'd18: xpb[94] = 1024'd54110843216934580004014501517784598061470155452743856304482113956085119418410579047955031970687561426889565587437335561039117623087400953779824296740944305068953530736347359668762111420533869663318891216683492339318037447963341953553501426379237320593558914487806540024172998414689389220274961496190018588627;
            6'd19: xpb[94] = 1024'd105365160606146122770437112259533799576712330193460169926782397256691974239498054126736172552537077070944655111861768316766482318030508914650154584066236615713663989220977686392771766185042442425123906465316501853977402081269431918237298727166006402008075483287063537037224037022033268128058616511888306365235;
            6'd20: xpb[94] = 1024'd32552782311232924138060795596468568347256077808440799420950825492321933723276390295502241919728918405556595228828707637914783172132396540965324746375197885424683773136036795779151181758033809465618724105562271522272405864354625109956117458269546034155772148672203476020168547555448514018723581700960999657512;
            6'd21: xpb[94] = 1024'd83807099700444466904483406338217769862498252549157113043251108792928788544363865374283382501578434049611684753253140393642147867075504501835655033700490196069394231620667122503160836522542382227423739354195281036931770497660715074639914759056315115570288717471460473033219586162792392926507236716659287434120;
            6'd22: xpb[94] = 1024'd10994721405531268272107089675152538633042000164137742537419537028558748028142201543049451868770275384223624870220079714790448721177392128150825196009451465780414015535726231889540252095533749267918556994441050705226774280745908266358733490159854747717985382856600412016164096696207638817172201905731980726397;
            6'd23: xpb[94] = 1024'd62249038794742811038529700416901740148284174904854056159719820329165602849229676621830592450619791028278714394644512470517813416120500089021155483334743776425124474020356558613549906860042322029723572243074060219886138914051998231042530790946623829132501951655857409029215135303551517724955856921430268503005;
            6'd24: xpb[94] = 1024'd113503356183954353804952311158650941663526349645570369782020103629772457670317151700611733032469306672333803919068945226245178111063608049891485770660036087069834932504986885337559561624550894791528587491707069734545503547358088195726328091733392910547018520455114406042266173910895396632739511937128556279613;
            6'd25: xpb[94] = 1024'd40690977889041155172575994495585710434070097260550999276188531865402417154095487869377802399661148006945744036035884547393478965165495676206655932968997356780854716420045994723938977197542261832023405131952839402840507330443281387445146822836932542694715185840254345025210684444310642523404477126201249571890;
            6'd26: xpb[94] = 1024'd91945295278252697938998605237334911949312272001267312898488815166009271975182962948158942981510663651000833560460317303120843660108603637076986220294289667425565174904676321447948631962050834593828420380585848917499871963749371352128944123623701624109231754639511342038261723051654521431188132141899537348498;
            6'd27: xpb[94] = 1024'd19132916983339499306622288574269680719856019616247942392657243401639231458961299116925012348702504985612773677427256624269144514210491263392156382603250937136584958819735430834328047535042201634323238020831618585794875746834564543847762854727241256256928420024651281021206233585069767321853097330972230640775;
            6'd28: xpb[94] = 1024'd70387234372551042073044899316018882235098194356964256014957526702246086280048774195706152930552020629667863201851689379996509209153599224262486669928543247781295417304365757558337702299550774396128253269464628100454240380140654508531560155514010337671444988823908278034257272192413646229636752346670518417383;
            6'd29: xpb[94] = 1024'd121641551761762584839467510057768083750340369097680569637257810002852941101136249274487293512401536273722952726276122135723873904096707185132816957253835558426005875788996084282347357064059347157933268518097637615113605013446744473215357456300779419085961557623165275047308310799757525137420407362368806193991;
            6'd30: xpb[94] = 1024'd48829173466849386207091193394702852520884116712661199131426238238482900584914585443253362879593377608334892843243061456872174758198594811447987119562796828137025659704055193668726772637050714198428086158343407283408608796531937664934176187404319051233658223008305214030252821333172771028085372551441499486268;
            6'd31: xpb[94] = 1024'd100083490856060928973513804136452054036126291453377512753726521539089755406002060522034503461442893252389982367667494212599539453141702772318317406888089138781736118188685520392736427401559286960233101406976416798067973429838027629617973488191088132648174791807562211043303859940516649935869027567139787262876;
            6'd32: xpb[94] = 1024'd27271112561147730341137487473386822806670039068358142247894949774719714889780396690800572828634734587001922484634433533747840307243590398633487569197050408492755902103744629779115842974550654000727919047222186466362977212923220821336792219294627764795871457192702150026248370473931895826533992756212480555153;
            6'd33: xpb[94] = 1024'd78525429950359273107560098215136024321912213809074455870195233075326569710867871769581713410484250231057012009058866289475205002186698359503817856522342719137466360588374956503125497739059226762532934295855195981022341846229310786020589520081396846210388025991959147039299409081275774734317647771910768331761;
            6'd34: xpb[94] = 1024'd5713051655446074475183781552070793092455961424055085364363661310956529194646207938347782777676091565668952126025805610623505856288585985818988018831303988848486144503434065889504913312050593803027751936100965649317345629314503977739408251184936478358084691377099086022243919614691020624982612960983461624038;
            6'd35: xpb[94] = 1024'd56967369044657617241606392293819994607698136164771398986663944611563384015733683017128923359525607209724041650450238366350870551231693946689318306156596299493196602988064392613514568076559166564832767184733975163976710262620593942423205551971705559772601260176356083035294958222034899532766267976681749400646;
            6'd36: xpb[94] = 1024'd108221686433869160008029003035569196122940310905487712608964227912170238836821158095910063941375122853779131174874671122078235246174801907559648593481888610137907061472694719337524222841067739326637782433366984678636074895926683907107002852758474641187117828975613080048345996829378778440549922992380037177254;
            6'd37: xpb[94] = 1024'd35409308138955961375652686372503964893484058520468342103132656147800198320599494264676133308566964188391071291841610443226536100276689533874818755790849879848926845387753828723903638414059106367132600073612754346931078679011877098825821583862014273334814494360753019031290507362794024331214888181452730469531;
            6'd38: xpb[94] = 1024'd86663625528167504142075297114253166408726233261184655725432939448407053141686969343457273890416479832446160816266043198953900795219797494745149043116142190493637303872384155447913293178567679128937615322245763861590443312317967063509618884648783354749331063160010016044341545970137903238998543197151018246139;
            6'd39: xpb[94] = 1024'd13851247233254305509698980451187935179269980876165285219601367684037012625465305512223343257608321167058100933232982520102201649321685121060319205425103460204657087787443264834292708751559046169432432962491533529885447095403160255228437615752322986897027728545149955027286056503553149129663508386223711538416;
            6'd40: xpb[94] = 1024'd65105564622465848276121591192937136694512155616881598841901650984643867446552780591004483839457836811113190457657415275829566344264793081930649492750395770849367546272073591558302363516067618931237448211124543044544811728709250219912234916539092068311544297344406952040337095110897028037447163401921999315024;
            6'd41: xpb[94] = 1024'd116359882011677391042544201934686338209754330357597912464201934285250722267640255669785624421307352455168279982081848031556931039207901042800979780075688081494078004756703918282312018280576191693042463459757552559204176362015340184596032217325861149726060866143663949053388133718240906945230818417620287091632;
            6'd42: xpb[94] = 1024'd43547503716764192410167885271621106980298077972578541958370362520880681751418591838551693788499193789780220099048787352705231893309788669116149942384649351205097788671763027668691433853567558733537281100003322227499180145100533376314850948429400781873757531528803888036332644251656152835895783606692980383909;
            6'd43: xpb[94] = 1024'd94801821105975735176590496013370308495540252713294855580670645821487536572506066917332834370348709433835309623473220108432596588252896629986480229709941661849808247156393354392701088618076131495342296348636331742158544778406623340998648249216169863288274100328060885049383682859000031743679438622391268160517;
            6'd44: xpb[94] = 1024'd21989442811062536544214179350305077266084000328275485074839074057117496056284403086098903737540550768447249740440159429580897442354784256301650392018902931560828031071452463779080504191067498535837113988882101410453548561491816532717466980319709495435970765713200824032328193392415277634344403811463961452794;
            6'd45: xpb[94] = 1024'd73243760200274079310636790092054278781326175068991798697139357357724350877371878164880044319390066412502339264864592185308262137297892217171980679344195242205538489556082790503090158955576071297642129237515110925112913194797906497401264281106478576850487334512457821045379231999759156542128058827162249229402;
            6'd46: xpb[94] = 1024'd431381905360880678260473428989047551869922683972428191307785593354310361150214333646113686581907747114279381831531506456562991399779843487150841653156511916558273471141899889469574528567438338136946877760880593407916977883099689120083012210018208998183999897597760028323742533174402432793024016234942521679;
            6'd47: xpb[94] = 1024'd51685699294572423444683084170738249067112097424688741813608068893961165182237689412427254268431423391169368906255964262183927686342887804357481128978448822561268731955772226613479229293076011099941962126393890108067281611189189653803880312996787290412700568696854757041374781140518281340576679031933230298287;
            6'd48: xpb[94] = 1024'd102940016683783966211105694912487450582354272165405055435908352194568020003325164491208394850280939035224458430680397017911292381285995765227811416303741133205979190440402553337488884057584583861746977375026899622726646244495279618487677613783556371827217137496111754054425819747862160248360334047631518074895;
            6'd49: xpb[94] = 1024'd30127638388870767578729378249422219352898019780385684930076780430197979487103500659974464217472780369836398547647336339059593235387883391542981578612702402916998974355461662723868299630575950902241795015272669291021650027580472810206496344887096003974913802881251693037370330281277406139025299236704211367172;
            6'd50: xpb[94] = 1024'd81381955778082310345151988991171420868140194521101998552377063730804834308190975738755604799322296013891488072071769094786957930330991352413311865937994713561709432840091989447877954395084523664046810263905678805681014660886562774890293645673865085389430371680508690050421368888621285046808954252402499143780;
            6'd51: xpb[94] = 1024'd8569577483169111712775672328106189638683942136082628046545491966434793791969311907521674166514137348503428189038708415935258784432878978728482028246955983272729216755151098834257369968075890704541627904151448473976018443971755966609112376777404717537127037065648629033365879422036530937473919441475192436057;
            6'd52: xpb[94] = 1024'd59823894872380654479198283069855391153926116876798941668845775267041648613056786986302814748363652992558517713463141171662623479375986939598812315572248293917439675239781425558267024732584463466346643152784457988635383077277845931292909677564173798951643605864905626046416918029380409845257574457173480212665;
            6'd53: xpb[94] = 1024'd111078212261592197245620893811604592669168291617515255291146058567648503434144262065083955330213168636613607237887573927389988174319094900469142602897540604562150133724411752282276679497093036228151658401417467503294747710583935895976706978350942880366160174664162623059467956636724288753041229472871767989273;
            6'd54: xpb[94] = 1024'd38265833966678998613244577148539361439712039232495884785314486803278462917922598233850024697405009971225547354854513248538289028420982526784312765206501874273169917639470861668656095070084403268646476041663237171589751493669129087695525709454482512513856840049302562042412467170139534643706194661944461281550;
            6'd55: xpb[94] = 1024'd89520151355890541379667187890288562954954213973212198407614770103885317739010073312631165279254525615280636879278946004265653723364090487654643052531794184917880376124101188392665749834592976030451491290296246686249116126975219052379323010241251593928373408848559559055463505777483413551489849677642749058158;
            6'd56: xpb[94] = 1024'd16707773060977342747290871227223331725497961588192827901783198339515277222788409481397234646446366949892576996245885325413954577465978113969813214840755454628900160039160297779045165407584343070946308930542016354544119910060412244098141741344791226076070074233699498038408016310898659442154814866715442350435;
            6'd57: xpb[94] = 1024'd67962090450188885513713481968972533240740136328909141524083481640122132043875884560178375228295882593947666520670318081141319272409086074840143502166047765273610618523790624503054820172092915832751324179175025869203484543366502208781939042131560307490586643032956495051459054918242538349938469882413730127043;
            6'd58: xpb[94] = 1024'd119216407839400428280136092710721734755982311069625455146383764940728986864963359638959515810145398238002756045094750836868683967352194035710473789491340075918321077008420951227064474936601488594556339427808035383862849176672592173465736342918329388905103211832213492064510093525586417257722124898112017903651;
            6'd59: xpb[94] = 1024'd46404029544487229647759776047656503526526058684606084640552193176358946348741695807725585177337239572614696162061690158016984821454081662025643951800301345629340860923480060613443890509592855635051157068053805052157852959757785365184555074021869021052799877217353431047454604059001663148387090087184711195928;
            6'd60: xpb[94] = 1024'd97658346933698772414182386789405705041768233425322398262852476476965801169829170886506725759186755216669785686486122913744349516397189622895974239125593656274051319408110387337453545274101428396856172316686814566817217593063875329868352374808638102467316446016610428060505642666345542056170745102882998972536;
            6'd61: xpb[94] = 1024'd24845968638785573781806070126340473812311981040303027757020904712595760653607507055272795126378596551281725803453062234892650370499077249211144401434554925985071103323169496723832960847092795437350989956932584235112221376149068521587171105912177734615013111401750367043450153199760787946835710291955692264813;
            6'd62: xpb[94] = 1024'd76100286027997116548228680868089675327554155781019341379321188013202615474694982134053935708228112195336815327877494990620015065442185210081474688759847236629781561807799823447842615611601368199156005205565593749771586009455158486270968406698946816029529680201007364056501191807104666854619365307653980041421;
            6'd63: xpb[94] = 1024'd3287907733083917915852364205024444098097903395999970873489616248832574958473318302820005075419953529948755444844434311768315919544072836396644851068808506340801345722858932834222031184592735239650822845811363418066589792540351677989787137802486448177226345586147303039445702340519912745284330496726673333698;
        endcase
    end

    always_comb begin
        case(flag[31][16:12])
            5'd0: xpb[95] = 1024'd0;
            5'd1: xpb[95] = 1024'd54542225122295460682274974946773645613340078136716284495789899549439429779560793381601145657269469174003844969268867067495680614487180797266975138394100816985511804207489259558231685949101308001455838094444372932725954425846441642673584438589255529591742914385404300052496740947863791653067985512424961110306;
            5'd2: xpb[95] = 1024'd109084450244590921364549949893547291226680156273432568991579799098878859559121586763202291314538938348007689938537734134991361228974361594533950276788201633971023608414978519116463371898202616002911676188888745865451908851692883285347168877178511059183485828770808600104993481895727583306135971024849922220612;
            5'd3: xpb[95] = 1024'd39559979682761640648025997435506504095321807284413169359237843583341394001373241234788365757150733212568385500349107767907978002620322057245765290165971410022844738052896561337064818655786718283057316674945878951813502427318428155055774746084537139508408839742095842127383694769662741942085266710649288846587;
            5'd4: xpb[95] = 1024'd94102204805057101330300972382280149708661885421129453855027743132780823780934034616389511414420202386572230469617974835403658617107502854512740428560072227008356542260385820895296504604888026284513154769390251884539456853164869797729359184673792669100151754127500142179880435717526533595153252223074249956893;
            5'd5: xpb[95] = 1024'd24577734243227820613777019924239362577303536432110054222685787617243358223185689087975585857031997251132926031429348468320275390753463317224555441937842003060177671898303863115897951362472128564658795255447384970901050428790414667437965053579818749425074765098787384202270648591461692231102547908873616582868;
            5'd6: xpb[95] = 1024'd79119959365523281296051994871013008190643614568826338718475687166682788002746482469576731514301466425136771000698215535815956005240644114491530580331942820045689476105793122674129637311573436566114633349891757903627004854636856310111549492169074279016817679484191684254767389539325483884170533421298577693174;
            5'd7: xpb[95] = 1024'd9595488803694000579528042412972221059285265579806939086133731651145322444998136941162805956913261289697466562509589168732572778886604577203345593709712596097510605743711164894731084069157538846260273835948890989988598430262401179820155361075100359341740690455478926277157602413260642520119829107097944319149;
            5'd8: xpb[95] = 1024'd64137713925989461261803017359745866672625343716523223581923631200584752224558930322763951614182730463701311531778456236228253393373785374470320732103813413083022409951200424452962770018258846847716111930393263922714552856108842822493739799664355888933483604840883226329654343361124434173187814619522905429455;
            5'd9: xpb[95] = 1024'd118679939048284921944077992306519512285965421853239508077713530750024182004119723704365097271452199637705156501047323303723934007860966171737295870497914230068534214158689684011194455967360154849171950024837636855440507281955284465167324238253611418525226519226287526382151084308988225826255800131947866539761;
            5'd10: xpb[95] = 1024'd49155468486455641227554039848478725154607072864220108445371575234486716446371378175951171714063994502265852062858696936640550781506926634449110883875684006120355343796607726231795902724944257129317590510894769941802100857580829334875930107159637498850149530197574768404541297182923384462205095817747233165736;
            5'd11: xpb[95] = 1024'd103697693608751101909829014795252370767947151000936392941161474783926146225932171557552317371333463676269697032127564004136231395994107431716086022269784823105867148004096985790027588674045565130773428605339142874528055283427270977549514545748893028441892444582979068457038038130787176115273081330172194276042;
            5'd12: xpb[95] = 1024'd34173223046921821193305062337211583636588802011916993308819519268388680668183826029138391813945258540830392593938937637052848169640067894427901035647554599157688277642015028010629035431629667410919069091396275960889648859052815847258120414654919108766815455554266310479428251004722334751222377015971560902017;
            5'd13: xpb[95] = 1024'd88715448169217281875580037283985229249928880148633277804609418817828110447744619410739537471214727714834237563207804704548528784127248691694876174041655416143200081849504287568860721380730975412374907185840648893615603284899257489931704853244174638358558369939670610531924991952586126404290362528396522012323;
            5'd14: xpb[95] = 1024'd19190977607388001159056084825944442118570531159613878172267463302290644889996273882325611913826522579394933125019178337465145557773209154406691187419425192195021211487422329789462168138315077692520547671897781979977196860524802359640310722150200718683481380910957852554315204826521285040239658214195888638298;
            5'd15: xpb[95] = 1024'd73733202729683461841331059772718087731910609296330162668057362851730074669557067263926757571095991753398778094288045404960826172260389951673666325813526009180533015694911589347693854087416385693976385766342154912703151286371244002313895160739456248275224295296362152606811945774385076693307643726620849748604;
            5'd16: xpb[95] = 1024'd4208732167854181124807107314677300600552260307310763035715407336192609111808721735512832013707786617959473656099419037877442945906350414385481339191295785232354145332829631568295300845000487974122026252399287999064744861996788872022501029645482328600147306267649394629202158648320235329256939412420216374579;
            5'd17: xpb[95] = 1024'd58750957290149641807082082261450946213892338444027047531505306885632038891369515117113977670977255791963318625368286105373123560393531211652456477585396602217865949540318891126526986794101795975577864346843660931790699287843230514696085468234737858191890220653053694681698899596184026982324924924845177484885;
            5'd18: xpb[95] = 1024'd113293182412445102489357057208224591827232416580743332027295206435071468670930308498715123328246724965967163594637153172868804174880712008919431615979497419203377753747808150684758672743203103977033702441288033864516653713689672157369669906823993387783633135038457994734195640544047818635392910437270138595191;
            5'd19: xpb[95] = 1024'd43768711850615821772833104750183804695874067591723932394953250919534003113181962970301197770858519830527859156448526805785420948526672471631246629357267195255198883385726192905360119500787206257179342927345166950878247289315217027078275775730019468108556146009745236756585853417982977271342206123069505221166;
            5'd20: xpb[95] = 1024'd98310936972911282455108079696957450309214145728440216890743150468973432892742756351902343428127989004531704125717393873281101563013853268898221767751368012240710687593215452463591805449888514258635181021789539883604201715161658669751860214319274997700299060395149536809082594365846768924410191635494466331472;
            5'd21: xpb[95] = 1024'd28786466411082001738584127238916663177855796739420817258401194953435967334994410823488417870739783869092399687528767506197718336659813731610036781129137788292531817231133494684193252207472616538780821507846672969965795290787203539460466083225301078025222071366436778831472807239781927560359487321293832957447;
            5'd22: xpb[95] = 1024'd83328691533377462420859102185690308791195874876137101754191094502875397114555204205089563528009253043096244656797634573693398951146994528877011919523238605278043621438622754242424938156573924540236659602291045902691749716633645182134050521814556607616964985751841078883969548187645719213427472833718794067753;
            5'd23: xpb[95] = 1024'd13804220971548181704335149727649521659837525887117702121849138987337931556806858676675637970621047907656940218609008206610015724792954991588826932901008381329864751076540796463026384914158026820382300088348178989053343292259190051842656390720582687941887996723128320906359761061580877849376768519518160693728;
            5'd24: xpb[95] = 1024'd68346446093843642386610124674423167273177604023833986617639038536777361336367652058276783627890517081660785187877875274105696339280135788855802071295109198315376555284030056021258070863259334821838138182792551921779297718105631694516240829309838217533630911108532620958856502009444669502444754031943121804034;
            5'd25: xpb[95] = 1024'd122888671216139103068885099621196812886517682160550271113428938086216791115928445439877929285159986255664630157146742341601376953767316586122777209689210015300888359491519315579489756812360642823293976277236924854505252143952073337189825267899093747125373825493936921011353242957308461155512739544368082914340;
            5'd26: xpb[95] = 1024'd53364200654309822352361147163156025755159333171530871481086982570679325558180099911464003727771781120225325718958115974517993727413277048834592223066979791352709489129437357800091203569944745103439616763294057940866845719577618206898431136805119827450296836465224163033743455831243619791462035230167449540315;
            5'd27: xpb[95] = 1024'd107906425776605283034636122109929671368499411308247155976876882120118755337740893293065149385041250294229170688226983042013674341900457846101567361461080608338221293336926617358322889519046053104895454857738430873592800145424059849572015575394375357042039750850628463086240196779107411444530020742592410650621;
            5'd28: xpb[95] = 1024'd38381955214776002318112169651888884237141062319227756344534926604581289779992547764651223827653045158789866250038356674930291115546418308813382374838850384390042422974844659578924336276630155385041095343795563959954393721049604719280621444300401437366962761821915705108630409653042570080479316428391777276596;
            5'd29: xpb[95] = 1024'd92924180337071463000387144598662529850481140455944040840324826154020719559553341146252369484922514332793711219307223742425971730033599106080357513232951201375554227182333919137156022225731463386496933438239936892680348146896046361954205882889656966958705676207320005161127150600906361733547301940816738386902;
            5'd30: xpb[95] = 1024'd23399709775242182283863192140621742719122791466924641207982870638483254001804995617838443927534309197354406781118597375342588503679559568792172526610720977427375356820251961357757468983315565666642573924297069979041941722521591231662811751795683047283628687178607247183517363474841520369496597626616105012877;
            5'd31: xpb[95] = 1024'd77941934897537642966138167087395388332462869603640925703772770187922683781365788999439589584803778371358251750387464442838269118166740366059147665004821794412887161027741220915989154932416873668098412018741442911767896148368032874336396190384938576875371601564011547236014104422705312022564583139041066123183;
        endcase
    end

    always_comb begin
        case(flag[32][5:0])
            6'd0: xpb[96] = 1024'd0;
            6'd1: xpb[96] = 1024'd4208732167854181124807107314677300600552260307310763035715407336192609111808721735512832013707786617959473656099419037877442945906350414385481339191295785232354145332829631568295300845000487974122026252399287999064744861996788872022501029645482328600147306267649394629202158648320235329256939412420216374579;
            6'd2: xpb[96] = 1024'd8417464335708362249614214629354601201104520614621526071430814672385218223617443471025664027415573235918947312198838075754885891812700828770962678382591570464708290665659263136590601690000975948244052504798575998129489723993577744045002059290964657200294612535298789258404317296640470658513878824840432749158;
            6'd3: xpb[96] = 1024'd12626196503562543374421321944031901801656780921932289107146222008577827335426165206538496041123359853878420968298257113632328837719051243156444017573887355697062435998488894704885902535001463922366078757197863997194234585990366616067503088936446985800441918802948183887606475944960705987770818237260649123737;
            6'd4: xpb[96] = 1024'd16834928671416724499228429258709202402209041229243052142861629344770436447234886942051328054831146471837894624397676151509771783625401657541925356765183140929416581331318526273181203380001951896488105009597151996258979447987155488090004118581929314400589225070597578516808634593280941317027757649680865498316;
            6'd5: xpb[96] = 1024'd21043660839270905624035536573386503002761301536553815178577036680963045559043608677564160068538933089797368280497095189387214729531752071927406695956478926161770726664148157841476504225002439870610131261996439995323724309983944360112505148227411643000736531338246973146010793241601176646284697062101081872895;
            6'd6: xpb[96] = 1024'd25252393007125086748842643888063803603313561843864578214292444017155654670852330413076992082246719707756841936596514227264657675438102486312888035147774711394124871996977789409771805070002927844732157514395727994388469171980733232135006177872893971600883837605896367775212951889921411975541636474521298247474;
            6'd7: xpb[96] = 1024'd29461125174979267873649751202741104203865822151175341250007851353348263782661052148589824095954506325716315592695933265142100621344452900698369374339070496626479017329807420978067105915003415818854183766795015993453214033977522104157507207518376300201031143873545762404415110538241647304798575886941514622053;
            6'd8: xpb[96] = 1024'd33669857342833448998456858517418404804418082458486104285723258689540872894469773884102656109662292943675789248795352303019543567250803315083850713530366281858833162662637052546362406760003903792976210019194303992517958895974310976180008237163858628801178450141195157033617269186561882634055515299361730996632;
            6'd9: xpb[96] = 1024'd37878589510687630123263965832095705404970342765796867321438666025733482006278495619615488123370079561635262904894771340896986513157153729469332052721662067091187307995466684114657707605004391767098236271593591991582703757971099848202509266809340957401325756408844551662819427834882117963312454711781947371211;
            6'd10: xpb[96] = 1024'd42087321678541811248071073146773006005522603073107630357154073361926091118087217355128320137077866179594736560994190378774429459063504143854813391912957852323541453328296315682953008450004879741220262523992879990647448619967888720225010296454823286001473062676493946292021586483202353292569394124202163745790;
            6'd11: xpb[96] = 1024'd46296053846395992372878180461450306606074863380418393392869480698118700229895939090641152150785652797554210217093609416651872404969854558240294731104253637555895598661125947251248309295005367715342288776392167989712193481964677592247511326100305614601620368944143340921223745131522588621826333536622380120369;
            6'd12: xpb[96] = 1024'd50504786014250173497685287776127607206627123687729156428584888034311309341704660826153984164493439415513683873193028454529315350876204972625776070295549422788249743993955578819543610140005855689464315028791455988776938343961466464270012355745787943201767675211792735550425903779842823951083272949042596494948;
            6'd13: xpb[96] = 1024'd54713518182104354622492395090804907807179383995039919464300295370503918453513382561666816178201226033473157529292447492406758296782555387011257409486845208020603889326785210387838910985006343663586341281190743987841683205958255336292513385391270271801914981479442130179628062428163059280340212361462812869527;
            6'd14: xpb[96] = 1024'd58922250349958535747299502405482208407731644302350682500015702706696527565322104297179648191909012651432631185391866530284201242688905801396738748678140993252958034659614841956134211830006831637708367533590031986906428067955044208315014415036752600402062287747091524808830221076483294609597151773883029244106;
            6'd15: xpb[96] = 1024'd63130982517812716872106609720159509008283904609661445535731110042889136677130826032692480205616799269392104841491285568161644188595256215782220087869436778485312179992444473524429512675007319611830393785989319985971172929951833080337515444682234929002209594014740919438032379724803529938854091186303245618685;
            6'd16: xpb[96] = 1024'd67339714685666897996913717034836809608836164916972208571446517379081745788939547768205312219324585887351578497590704606039087134501606630167701427060732563717666325325274105092724813520007807585952420038388607985035917791948621952360016474327717257602356900282390314067234538373123765268111030598723461993264;
            6'd17: xpb[96] = 1024'd71548446853521079121720824349514110209388425224282971607161924715274354900748269503718144233032372505311052153690123643916530080407957044553182766252028348950020470658103736661020114365008295560074446290787895984100662653945410824382517503973199586202504206550039708696436697021444000597367970011143678367843;
            6'd18: xpb[96] = 1024'd75757179021375260246527931664191410809940685531593734642877332051466964012556991239230976246740159123270525809789542681793973026314307458938664105443324134182374615990933368229315415210008783534196472543187183983165407515942199696405018533618681914802651512817689103325638855669764235926624909423563894742422;
            6'd19: xpb[96] = 1024'd79965911189229441371335038978868711410492945838904497678592739387659573124365712974743808260447945741229999465888961719671415972220657873324145444634619919414728761323762999797610716055009271508318498795586471982230152377938988568427519563264164243402798819085338497954841014318084471255881848835984111117001;
            6'd20: xpb[96] = 1024'd84174643357083622496142146293546012011045206146215260714308146723852182236174434710256640274155732359189473121988380757548858918127008287709626783825915704647082906656592631365906016900009759482440525047985759981294897239935777440450020592909646572002946125352987892584043172966404706585138788248404327491580;
            6'd21: xpb[96] = 1024'd88383375524937803620949253608223312611597466453526023750023554060044791347983156445769472287863518977148946778087799795426301864033358702095108123017211489879437051989422262934201317745010247456562551300385047980359642101932566312472521622555128900603093431620637287213245331614724941914395727660824543866159;
            6'd22: xpb[96] = 1024'd92592107692791984745756360922900613212149726760836786785738961396237400459791878181282304301571305595108420434187218833303744809939709116480589462208507275111791197322251894502496618590010735430684577552784335979424386963929355184495022652200611229203240737888286681842447490263045177243652667073244760240738;
            6'd23: xpb[96] = 1024'd96800839860646165870563468237577913812701987068147549821454368732430009571600599916795136315279092213067894090286637871181187755846059530866070801399803060344145342655081526070791919435011223404806603805183623978489131825926144056517523681846093557803388044155936076471649648911365412572909606485664976615317;
            6'd24: xpb[96] = 1024'd101009572028500346995370575552255214413254247375458312857169776068622618683409321652307968328986878831027367746386056909058630701752409945251552140591098845576499487987911157639087220280011711378928630057582911977553876687922932928540024711491575886403535350423585471100851807559685647902166545898085192989896;
            6'd25: xpb[96] = 1024'd105218304196354528120177682866932515013806507682769075892885183404815227795218043387820800342694665448986841402485475946936073647658760359637033479782394630808853633320740789207382521125012199353050656309982199976618621549919721800562525741137058215003682656691234865730053966208005883231423485310505409364475;
            6'd26: xpb[96] = 1024'd109427036364208709244984790181609815614358767990079838928600590741007836907026765123333632356402452066946315058584894984813516593565110774022514818973690416041207778653570420775677821970012687327172682562381487975683366411916510672585026770782540543603829962958884260359256124856326118560680424722925625739054;
            6'd27: xpb[96] = 1024'd113635768532062890369791897496287116214911028297390601964315998077200446018835486858846464370110238684905788714684314022690959539471461188407996158164986201273561923986400052343973122815013175301294708814780775974748111273913299544607527800428022872203977269226533654988458283504646353889937364135345842113633;
            6'd28: xpb[96] = 1024'd117844500699917071494599004810964416815463288604701365000031405413393055130644208594359296383818025302865262370783733060568402485377811602793477497356281986505916069319229683912268423660013663275416735067180063973812856135910088416630028830073505200804124575494183049617660442152966589219194303547766058488212;
            6'd29: xpb[96] = 1024'd122053232867771252619406112125641717416015548912012128035746812749585664242452930329872128397525811920824736026883152098445845431284162017178958836547577771738270214652059315480563724505014151249538761319579351972877600997906877288652529859718987529404271881761832444246862600801286824548451242960186274862791;
            6'd30: xpb[96] = 1024'd2195269351500692345414292035504585271869382093587206943330365020801378016952513155369889196575924229341060275525077701744224536349292097009280050722542516036933685415317729711228786158497433502350589963591400125577985009682769387710052319681240408737599284615364780845958231375678426860589492545980896753039;
            6'd31: xpb[96] = 1024'd6404001519354873470221399350181885872421642400897969979045772356993987128761234890882721210283710847300533931624496739621667482255642511394761389913838301269287830748147361279524087003497921476472616215990688124642729871679558259732553349326722737337746590883014175475160390023998662189846431958401113127618;
            6'd32: xpb[96] = 1024'd10612733687209054595028506664859186472973902708208733014761179693186596240569956626395553223991497465260007587723915777499110428161992925780242729105134086501641976080976992847819387848498409450594642468389976123707474733676347131755054378972205065937893897150663570104362548672318897519103371370821329502197;
            6'd33: xpb[96] = 1024'd14821465855063235719835613979536487073526163015519496050476587029379205352378678361908385237699284083219481243823334815376553374068343340165724068296429871733996121413806624416114688693498897424716668720789264122772219595673136003777555408617687394538041203418312964733564707320639132848360310783241545876776;
            6'd34: xpb[96] = 1024'd19030198022917416844642721294213787674078423322830259086191994365571814464187400097421217251407070701178954899922753853253996319974693754551205407487725656966350266746636255984409989538499385398838694973188552121836964457669924875800056438263169723138188509685962359362766865968959368177617250195661762251355;
            6'd35: xpb[96] = 1024'd23238930190771597969449828608891088274630683630141022121907401701764423575996121832934049265114857319138428556022172891131439265881044168936686746679021442198704412079465887552705290383499873372960721225587840120901709319666713747822557467908652051738335815953611753991969024617279603506874189608081978625934;
            6'd36: xpb[96] = 1024'd27447662358625779094256935923568388875182943937451785157622809037957032687804843568446881278822643937097902212121591929008882211787394583322168085870317227431058557412295519121000591228500361347082747477987128119966454181663502619845058497554134380338483122221261148621171183265599838836131129020502195000513;
            6'd37: xpb[96] = 1024'd31656394526479960219064043238245689475735204244762548193338216374149641799613565303959713292530430555057375868221010966886325157693744997707649425061613012663412702745125150689295892073500849321204773730386416119031199043660291491867559527199616708938630428488910543250373341913920074165388068432922411375092;
            6'd38: xpb[96] = 1024'd35865126694334141343871150552922990076287464552073311229053623710342250911422287039472545306238217173016849524320430004763768103600095412093130764252908797895766848077954782257591192918501337295326799982785704118095943905657080363890060556845099037538777734756559937879575500562240309494645007845342627749671;
            6'd39: xpb[96] = 1024'd40073858862188322468678257867600290676839724859384074264769031046534860023231008774985377319946003790976323180419849042641211049506445826478612103444204583128120993410784413825886493763501825269448826235184992117160688767653869235912561586490581366138925041024209332508777659210560544823901947257762844124250;
            6'd40: xpb[96] = 1024'd44282591030042503593485365182277591277391985166694837300484438382727469135039730510498209333653790408935796836519268080518653995412796240864093442635500368360475138743614045394181794608502313243570852487584280116225433629650658107935062616136063694739072347291858727137979817858880780153158886670183060498829;
            6'd41: xpb[96] = 1024'd48491323197896684718292472496954891877944245474005600336199845718920078246848452246011041347361577026895270492618687118396096941319146655249574781826796153592829284076443676962477095453502801217692878739983568115290178491647446979957563645781546023339219653559508121767181976507201015482415826082603276873408;
            6'd42: xpb[96] = 1024'd52700055365750865843099579811632192478496505781316363371915253055112687358657173981523873361069363644854744148718106156273539887225497069635056121018091938825183429409273308530772396298503289191814904992382856114354923353644235851980064675427028351939366959827157516396384135155521250811672765495023493247987;
            6'd43: xpb[96] = 1024'd56908787533605046967906687126309493079048766088627126407630660391305296470465895717036705374777150262814217804817525194150982833131847484020537460209387724057537574742102940099067697143503777165936931244782144113419668215641024724002565705072510680539514266094806911025586293803841486140929704907443709622566;
            6'd44: xpb[96] = 1024'd61117519701459228092713794440986793679601026395937889443346067727497905582274617452549537388484936880773691460916944232028425779038197898406018799400683509289891720074932571667362997988504265140058957497181432112484413077637813596025066734717993009139661572362456305654788452452161721470186644319863925997145;
            6'd45: xpb[96] = 1024'd65326251869313409217520901755664094280153286703248652479061475063690514694083339188062369402192723498733165117016363269905868724944548312791500138591979294522245865407762203235658298833504753114180983749580720111549157939634602468047567764363475337739808878630105700283990611100481956799443583732284142371724;
            6'd46: xpb[96] = 1024'd69534984037167590342328009070341394880705547010559415514776882399883123805892060923575201415900510116692638773115782307783311670850898727176981477783275079754600010740591834803953599678505241088303010001980008110613902801631391340070068794008957666339956184897755094913192769748802192128700523144704358746303;
            6'd47: xpb[96] = 1024'd73743716205021771467135116385018695481257807317870178550492289736075732917700782659088033429608296734652112429215201345660754616757249141562462816974570864986954156073421466372248900523505729062425036254379296109678647663628180212092569823654439994940103491165404489542394928397122427457957462557124575120882;
            6'd48: xpb[96] = 1024'd77952448372875952591942223699695996081810067625180941586207697072268342029509504394600865443316083352611586085314620383538197562663599555947944156165866650219308301406251097940544201368506217036547062506778584108743392525624969084115070853299922323540250797433053884171597087045442662787214401969544791495461;
            6'd49: xpb[96] = 1024'd82161180540730133716749331014373296682362327932491704621923104408460951141318226130113697457023869970571059741414039421415640508569949970333425495357162435451662446739080729508839502213506705010669088759177872107808137387621757956137571882945404652140398103700703278800799245693762898116471341381965007870040;
            6'd50: xpb[96] = 1024'd86369912708584314841556438329050597282914588239802467657638511744653560253126947865626529470731656588530533397513458459293083454476300384718906834548458220684016592071910361077134803058507192984791115011577160106872882249618546828160072912590886980740545409968352673430001404342083133445728280794385224244619;
            6'd51: xpb[96] = 1024'd90578644876438495966363545643727897883466848547113230693353919080846169364935669601139361484439443206490007053612877497170526400382650799104388173739754005916370737404739992645430103903507680958913141263976448105937627111615335700182573942236369309340692716236002068059203562990403368774985220206805440619198;
            6'd52: xpb[96] = 1024'd94787377044292677091170652958405198484019108854423993729069326417038778476744391336652193498147229824449480709712296535047969346289001213489869512931049791148724882737569624213725404748508168933035167516375736105002371973612124572205074971881851637940840022503651462688405721638723604104242159619225656993777;
            6'd53: xpb[96] = 1024'd98996109212146858215977760273082499084571369161734756764784733753231387588553113072165025511855016442408954365811715572925412292195351627875350852122345576381079028070399255782020705593508656907157193768775024104067116835608913444227576001527333966540987328771300857317607880287043839433499099031645873368356;
            6'd54: xpb[96] = 1024'd103204841380001039340784867587759799685123629469045519800500141089423996700361834807677857525562803060368428021911134610802855238101702042260832191313641361613433173403228887350316006438509144881279220021174312103131861697605702316250077031172816295141134635038950251946810038935364074762756038444066089742935;
            6'd55: xpb[96] = 1024'd107413573547855220465591974902437100285675889776356282836215548425616605812170556543190689539270589678327901678010553648680298184008052456646313530504937146845787318736058518918611307283509632855401246273573600102196606559602491188272578060818298623741281941306599646576012197583684310092012977856486306117514;
            6'd56: xpb[96] = 1024'd111622305715709401590399082217114400886228150083667045871930955761809214923979278278703521552978376296287375334109972686557741129914402871031794869696232932078141464068888150486906608128510120829523272525972888101261351421599280060295079090463780952341429247574249041205214356232004545421269917268906522492093;
            6'd57: xpb[96] = 1024'd115831037883563582715206189531791701486780410390977808907646363098001824035788000014216353566686162914246848990209391724435184075820753285417276208887528717310495609401717782055201908973510608803645298778372176100326096283596068932317580120109263280941576553841898435834416514880324780750526856681326738866672;
            6'd58: xpb[96] = 1024'd120039770051417763840013296846469002087332670698288571943361770434194433147596721749729185580393949532206322646308810762312627021727103699802757548078824502542849754734547413623497209818511096777767325030771464099390841145592857804340081149754745609541723860109547830463618673528645016079783796093746955241251;
            6'd59: xpb[96] = 1024'd181806535147203566021476756331869943186503879863650850945322705410146922096304575226946379444061840722646894950736365611006126792233779633078762253789246841513225497805827854162271471994379030579153674783512252091225157368749903397603609716998488875051262963080167062714304103036618391922045679541577131499;
            6'd60: xpb[96] = 1024'd4390538703001384690828584071009170543738764187174413886660730041602756033905026310739778393151848458682120551050155403488449072698584194018560101445085032073867370830635459422457572316994867004701179927182800251155970019365538775420104639362480817475198569230729561691916462751356853721178985091961793506078;
            6'd61: xpb[96] = 1024'd8599270870855565815635691385686471144291024494485176922376137377795365145713748046252610406859635076641594207149574441365892018604934608404041440636380817306221516163465090990752873161995354978823206179582088250220714881362327647442605669007963146075345875498378956321118621399677089050435924504382009880657;
            6'd62: xpb[96] = 1024'd12808003038709746940442798700363771744843284801795939958091544713987974257522469781765442420567421694601067863248993479243334964511285022789522779827676602538575661496294722559048174006995842952945232431981376249285459743359116519465106698653445474675493181766028350950320780047997324379692863916802226255236;
            6'd63: xpb[96] = 1024'd17016735206563928065249906015041072345395545109106702993806952050180583369331191517278274434275208312560541519348412517120777910417635437175004119018972387770929806829124354127343474851996330927067258684380664248350204605355905391487607728298927803275640488033677745579522938696317559708949803329222442629815;
        endcase
    end

    always_comb begin
        case(flag[32][11:6])
            6'd0: xpb[97] = 1024'd0;
            6'd1: xpb[97] = 1024'd21225467374418109190057013329718372945947805416417466029522359386373192481139913252791106447982994930520015175447831554998220856323985851560485458210268173003283952161953985695638775696996818901189284936779952247414949467352694263510108757944410131875787794301327140208725097344637795038206742741642659004394;
            6'd2: xpb[97] = 1024'd42450934748836218380114026659436745891895610832834932059044718772746384962279826505582212895965989861040030350895663109996441712647971703120970916420536346006567904323907971391277551393993637802378569873559904494829898934705388527020217515888820263751575588602654280417450194689275590076413485483285318008788;
            6'd3: xpb[97] = 1024'd63676402123254327570171039989155118837843416249252398088567078159119577443419739758373319343948984791560045526343494664994662568971957554681456374630804519009851856485861957086916327090990456703567854810339856742244848402058082790530326273833230395627363382903981420626175292033913385114620228224927977013182;
            6'd4: xpb[97] = 1024'd84901869497672436760228053318873491783791221665669864118089437545492769924559653011164425791931979722080060701791326219992883425295943406241941832841072692013135808647815942782555102787987275604757139747119808989659797869410777054040435031777640527503151177205308560834900389378551180152826970966570636017576;
            6'd5: xpb[97] = 1024'd106127336872090545950285066648591864729739027082087330147611796931865962405699566263955532239914974652600075877239157774991104281619929257802427291051340865016419760809769928478193878484984094505946424683899761237074747336763471317550543789722050659378938971506635701043625486723188975191033713708213295021970;
            6'd6: xpb[97] = 1024'd3286108562383913741543152573495804930988405372769112049002301253262259549530340606731567473240295273676941645229495895410261297102694774807752624245277997086013038402152696836202414990463707685825512012292473638125335953895268808095673977983231341987906862393845783222244055993898137212121766623230359542033;
            6'd7: xpb[97] = 1024'd24511575936802022931600165903214177876936210789186578078524660639635452030670253859522673921223290204196956820677327450408482153426680626368238082455546170089296990564106682531841190687460526587014796949072425885540285421247963071605782735927641473863694656695172923430969153338535932250328509364873018546427;
            6'd8: xpb[97] = 1024'd45737043311220132121657179232932550822884016205604044108047020026008644511810167112313780369206285134716971996125159005406703009750666477928723540665814343092580942726060668227479966384457345488204081885852378132955234888600657335115891493872051605739482450996500063639694250683173727288535252106515677550821;
            6'd9: xpb[97] = 1024'd66962510685638241311714192562650923768831821622021510137569379412381836992950080365104886817189280065236987171572990560404923866074652329489208998876082516095864894888014653923118742081454164389393366822632330380370184355953351598626000251816461737615270245297827203848419348027811522326741994848158336555215;
            6'd10: xpb[97] = 1024'd88187978060056350501771205892369296714779627038438976167091738798755029474089993617895993265172274995757002347020822115403144722398638181049694457086350689099148847049968639618757517778450983290582651759412282627785133823306045862136109009760871869491058039599154344057144445372449317364948737589800995559609;
            6'd11: xpb[97] = 1024'd109413445434474459691828219222087669660727432454856442196614098185128221955229906870687099713155269926277017522468653670401365578722624032610179915296618862102432799211922625314396293475447802191771936696192234875200083290658740125646217767705282001366845833900481484265869542717087112403155480331443654564003;
            6'd12: xpb[97] = 1024'd6572217124767827483086305146991609861976810745538224098004602506524519099060681213463134946480590547353883290458991790820522594205389549615505248490555994172026076804305393672404829980927415371651024024584947276250671907790537616191347955966462683975813724787691566444488111987796274424243533246460719084066;
            6'd13: xpb[97] = 1024'd27797684499185936673143318476709982807924616161955690127526961892897711580200594466254241394463585477873898465906823345818743450529375401175990706700824167175310028966259379368043605677924234272840308961364899523665621375143231879701456713910872815851601519089018706653213209332434069462450275988103378088460;
            6'd14: xpb[97] = 1024'd49023151873604045863200331806428355753872421578373156157049321279270904061340507719045347842446580408393913641354654900816964306853361252736476164911092340178593981128213365063682381374921053174029593898144851771080570842495926143211565471855282947727389313390345846861938306677071864500657018729746037092854;
            6'd15: xpb[97] = 1024'd70248619248022155053257345136146728699820226994790622186571680665644096542480420971836454290429575338913928816802486455815185163177347104296961623121360513181877933290167350759321157071917872075218878834924804018495520309848620406721674229799693079603177107691672987070663404021709659538863761471388696097248;
            6'd16: xpb[97] = 1024'd91474086622440264243314358465865101645768032411208088216094040052017289023620334224627560738412570269433943992250318010813406019501332955857447081331628686185161885452121336454959932768914690976408163771704756265910469777201314670231782987744103211478964901993000127279388501366347454577070504213031355101642;
            6'd17: xpb[97] = 1024'd112699553996858373433371371795583474591715837827625554245616399438390481504760247477418667186395565199953959167698149565811626875825318807417932539541896859188445837614075322150598708465911509877597448708484708513325419244554008933741891745688513343354752696294327267488113598710985249615277246954674014106036;
            6'd18: xpb[97] = 1024'd9858325687151741224629457720487414792965216118307336147006903759786778648591021820194702419720885821030824935688487686230783891308084324423257872735833991258039115206458090508607244971391123057476536036877420914376007861685806424287021933949694025963720587181537349666732167981694411636365299869691078626099;
            6'd19: xpb[97] = 1024'd31083793061569850414686471050205787738913021534724802176529263146159971129730935072985808867703880751550840111136319241229004747632070175983743330946102164261323067368412076204246020668387941958665820973657373161790957329038500687797130691894104157839508381482864489875457265326332206674572042611333737630493;
            6'd20: xpb[97] = 1024'd52309260435987959604743484379924160684860826951142268206051622532533163610870848325776915315686875682070855286584150796227225603956056027544228789156370337264607019530366061899884796365384760859855105910437325409205906796391194951307239449838514289715296175784191630084182362670970001712778785352976396634887;
            6'd21: xpb[97] = 1024'd73534727810406068794800497709642533630808632367559734235573981918906356092010761578568021763669870612590870462031982351225446460280041879104714247366638510267890971692320047595523572062381579761044390847217277656620856263743889214817348207782924421591083970085518770292907460015607796750985528094619055639281;
            6'd22: xpb[97] = 1024'd94760195184824177984857511039360906576756437783977200265096341305279548573150674831359128211652865543110885637479813906223667316604027730665199705576906683271174923854274033291162347759378398662233675783997229904035805731096583478327456965727334553466871764386845910501632557360245591789192270836261714643675;
            6'd23: xpb[97] = 1024'd115985662559242287174914524369079279522704243200394666294618700691652741054290588084150234659635860473630900812927645461221888172928013582225685163787174856274458876016228018986801123456375217563422960720777182151450755198449277741837565723671744685342659558688173050710357654704883386827399013577904373648069;
            6'd24: xpb[97] = 1024'd13144434249535654966172610293983219723953621491076448196009205013049038198121362426926269892961181094707766580917983581641045188410779099231010496981111988344052153608610787344809659961854830743302048049169894552501343815581075232382695911932925367951627449575383132888976223975592548848487066492921438168132;
            6'd25: xpb[97] = 1024'd34369901623953764156229623623701592669901426907493914225531564399422230679261275679717376340944176025227781756365815136639266044734764950791495955191380161347336105770564773040448435658851649644491332985949846799916293282933769495892804669877335499827415243876710273097701321320230343886693809234564097172526;
            6'd26: xpb[97] = 1024'd55595368998371873346286636953419965615849232323911380255053923785795423160401188932508482788927170955747796931813646691637486901058750802351981413401648334350620057932518758736087211355848468545680617922729799047331242750286463759402913427821745631703203038178037413306426418664868138924900551976206756176920;
            6'd27: xpb[97] = 1024'd76820836372789982536343650283138338561797037740328846284576283172168615641541102185299589236910165886267812107261478246635707757382736653912466871611916507353904010094472744431725987052845287446869902859509751294746192217639158022913022185766155763578990832479364553515151516009505933963107294717849415181314;
            6'd28: xpb[97] = 1024'd98046303747208091726400663612856711507744843156746312314098642558541808122681015438090695684893160816787827282709309801633928613706722505472952329822184680357187962256426730127364762749842106348059187796289703542161141684991852286423130943710565895454778626780691693723876613354143729001314037459492074185708;
            6'd29: xpb[97] = 1024'd119271771121626200916457676942575084453692648573163778343621001944915000603820928690881802132876155747307842458157141356632149470030708357033437788032452853360471914418380715823003538446838925249248472733069655789576091152344546549933239701654976027330566421082018833932601710698781524039520780201134733190102;
            6'd30: xpb[97] = 1024'd16430542811919568707715762867479024654942026863845560245011506266311297747651703033657837366201476368384708226147479477051306485513473874038763121226389985430065192010763484181012074952318538429127560061462368190626679769476344040478369889916156709939534311969228916111220279969490686060608833116151797710165;
            6'd31: xpb[97] = 1024'd37656010186337677897772776197197397600889832280263026274533865652684490228791616286448943814184471298904723401595311032049527341837459725599248579436658158433349144172717469876650850649315357330316844998242320438041629236829038303988478647860566841815322106270556056319945377314128481098815575857794456714559;
            6'd32: xpb[97] = 1024'd58881477560755787087829789526915770546837637696680492304056225039057682709931529539240050262167466229424738577043142587047748198161445577159734037646926331436633096334671455572289626346312176231506129935022272685456578704181732567498587405804976973691109900571883196528670474658766276137022318599437115718953;
            6'd33: xpb[97] = 1024'd80106944935173896277886802856634143492785443113097958333578584425430875191071442792031156710150461159944753752490974142045969054485431428720219495857194504439917048496625441267928402043308995132695414871802224932871528171534426831008696163749387105566897694873210336737395572003404071175229061341079774723347;
            6'd34: xpb[97] = 1024'd101332412309592005467943816186352516438733248529515424363100943811804067672211356044822263158133456090464768927938805697044189910809417280280704954067462677443201000658579426963567177740305814033884699808582177180286477638887121094518804921693797237442685489174537476946120669348041866213435804082722433727741;
            6'd35: xpb[97] = 1024'd122557879684010114658000829516070889384681053945932890392623303198177260153351269297613369606116451020984784103386637252042410767133403131841190412277730850446484952820533412659205953437302632935073984745362129427701427106239815358028913679638207369318473283475864617154845766692679661251642546824365092732135;
            6'd36: xpb[97] = 1024'd19716651374303482449258915440974829585930432236614672294013807519573557297182043640389404839441771642061649871376975372461567782616168648846515745471667982516078230412916181017214489942782246114953072073754841828752015723371612848574043867899388051927441174363074699333464335963388823272730599739382157252198;
            6'd37: xpb[97] = 1024'd40942118748721591639315928770693202531878237653032138323536166905946749778321956893180511287424766572581665046824806927459788638940154500407001203681936155519362182574870166712853265639779065016142357010534794076166965190724307112084152625843798183803228968664401839542189433308026618310937342481024816256592;
            6'd38: xpb[97] = 1024'd62167586123139700829372942100411575477826043069449604353058526292319942259461870145971617735407761503101680222272638482458009495264140351967486661892204328522646134736824152408492041336775883917331641947314746323581914658077001375594261383788208315679016762965728979750914530652664413349144085222667475260986;
            6'd39: xpb[97] = 1024'd83393053497557810019429955430129948423773848485867070382580885678693134740601783398762724183390756433621695397720470037456230351588126203527972120102472501525930086898778138104130817033772702818520926884094698570996864125429695639104370141732618447554804557267056119959639627997302208387350827964310134265380;
            6'd40: xpb[97] = 1024'd104618520871975919209486968759848321369721653902284536412103245065066327221741696651553830631373751364141710573168301592454451207912112055088457578312740674529214039060732123799769592730769521719710211820874650818411813592782389902614478899677028579430592351568383260168364725341940003425557570705952793269774;
            6'd41: xpb[97] = 1024'd1777292562269287000745054684752261570971032192966318313493749386462624365572470994329865864699071985218576341158639712873608223394877572093782911506677806598807316653114892157778129236249134899589299149267363219462402209914187393159609087938209262039560242455593342346983294612649165446645623620969857789837;
            6'd42: xpb[97] = 1024'd23002759936687396190802068014470634516918837609383784343016108772835816846712384247120972312682066915738591516606471267871829079718863423654268369716945979602091268815068877853416904933245953800778584086047315466877351677266881656669717845882619393915348036756920482555708391957286960484852366362612516794231;
            6'd43: xpb[97] = 1024'd44228227311105505380859081344189007462866643025801250372538468159209009327852297499912078760665061846258606692054302822870049936042849275214753827927214152605375220977022863549055680630242772701967869022827267714292301144619575920179826603827029525791135831058247622764433489301924755523059109104255175798625;
            6'd44: xpb[97] = 1024'd65453694685523614570916094673907380408814448442218716402060827545582201808992210752703185208648056776778621867502134377868270792366835126775239286137482325608659173138976849244694456327239591603157153959607219961707250611972270183689935361771439657666923625359574762973158586646562550561265851845897834803019;
            6'd45: xpb[97] = 1024'd86679162059941723760973108003625753354762253858636182431583186931955394290132124005494291656631051707298637042949965932866491648690820978335724744347750498611943125300930834940333232024236410504346438896387172209122200079324964447200044119715849789542711419660901903181883683991200345599472594587540493807413;
            6'd46: xpb[97] = 1024'd107904629434359832951030121333344126300710059275053648461105546318328586771272037258285398104614046637818652218397797487864712505014806829896210202558018671615227077462884820635972007721233229405535723833167124456537149546677658710710152877660259921418499213962229043390608781335838140637679337329183152811807;
            6'd47: xpb[97] = 1024'd5063401124653200742288207258248066501959437565735430362496050639724883915102811601061433337939367258895517986388135608283869520497572346901535535751955803684820355055267588993980544226712842585414811161559836857587738163809456201255283065921440604027467104849439125569227350606547302658767390244200217331870;
            6'd48: xpb[97] = 1024'd26288868499071309932345220587966439447907242982152896392018410026098076396242724853852539785922362189415533161835967163282090376821558198462020993962223976688104307217221574689619319923709661486604096098339789105002687631162150464765391823865850735903254899150766265777952447951185097696974132985842876336264;
            6'd49: xpb[97] = 1024'd47514335873489419122402233917684812393855048398570362421540769412471268877382638106643646233905357119935548337283798718280311233145544050022506452172492149691388259379175560385258095620706480387793381035119741352417637098514844728275500581810260867779042693452093405986677545295822892735180875727485535340658;
            6'd50: xpb[97] = 1024'd68739803247907528312459247247403185339802853814987828451063128798844461358522551359434752681888352050455563512731630273278532089469529901582991910382760322694672211541129546080896871317703299288982665971899693599832586565867538991785609339754670999654830487753420546195402642640460687773387618469128194345052;
            6'd51: xpb[97] = 1024'd89965270622325637502516260577121558285750659231405294480585488185217653839662464612225859129871346980975578688179461828276752945793515753143477368593028495697956163703083531776535647014700118190171950908679645847247536033220233255295718097699081131530618282054747686404127739985098482811594361210770853349446;
            6'd52: xpb[97] = 1024'd111190737996743746692573273906839931231698464647822760510107847571590846320802377865016965577854341911495593863627293383274973802117501604703962826803296668701240115865037517472174422711696937091361235845459598094662485500572927518805826855643491263406406076356074826612852837329736277849801103952413512353840;
            6'd53: xpb[97] = 1024'd8349509687037114483831359831743871432947842938504542411498351892987143464633152207793000811179662532572459631617631503694130817600267121709288159997233800770833393457420285830182959217176550271240323173852310495713074117704725009350957043904671946015373967243284908791471406600445439870889156867430576873903;
            6'd54: xpb[97] = 1024'd29574977061455223673888373161462244378895648354922008441020711279360335945773065460584107259162657463092474807065463058692351673924252973269773618207501973774117345619374271525821734914173369172429608110632262743128023585057419272861065801849082077891161761544612049000196503945083234909095899609073235878297;
            6'd55: xpb[97] = 1024'd50800444435873332863945386491180617324843453771339474470543070665733528426912978713375213707145652393612489982513294613690572530248238824830259076417770146777401297781328257221460510611170188073618893047412214990542973052410113536371174559793492209766949555845939189208921601289721029947302642350715894882691;
            6'd56: xpb[97] = 1024'd72025911810291442054002399820898990270791259187756940500065430052106720908052891966166320155128647324132505157961126168688793386572224676390744534628038319780685249943282242917099286308167006974808177984192167237957922519762807799881283317737902341642737350147266329417646698634358824985509385092358553887085;
            6'd57: xpb[97] = 1024'd93251379184709551244059413150617363216739064604174406529587789438479913389192805218957426603111642254652520333408957723687014242896210527951229992838306492783969202105236228612738062005163825875997462920972119485372871987115502063391392075682312473518525144448593469626371795978996620023716127834001212891479;
            6'd58: xpb[97] = 1024'd114476846559127660434116426480335736162686870020591872559110148824853105870332718471748533051094637185172535508856789278685235099220196379511715451048574665787253154267190214308376837702160644777186747857752071732787821454468196326901500833626722605394312938749920609835096893323634415061922870575643871895873;
            6'd59: xpb[97] = 1024'd11635618249421028225374512405239676363936248311273654460500653146249403014163492814524568284419957806249401276847127399104392114702961896517040784242511797856846431859572982666385374207640257957065835186144784133838410071599993817446631021887903288003280829637130692013715462594343577083010923490660936415936;
            6'd60: xpb[97] = 1024'd32861085623839137415431525734958049309884053727691120490023012532622595495303406067315674732402952736769416452294958954102612971026947748077526242452779970860130384021526968362024149904637076858255120122924736381253359538952688080956739779832313419879068623938457832222440559938981372121217666232303595420330;
            6'd61: xpb[97] = 1024'd54086552998257246605488539064676422255831859144108586519545371918995787976443319320106781180385947667289431627742790509100833827350933599638011700663048143863414336183480954057662925601633895759444405059704688628668309006305382344466848537776723551754856418239784972431165657283619167159424408973946254424724;
            6'd62: xpb[97] = 1024'd75312020372675355795545552394394795201779664560526052549067731305368980457583232572897887628368942597809446803190622064099054683674919451198497158873316316866698288345434939753301701298630714660633689996484640876083258473658076607976957295721133683630644212541112112639890754628256962197631151715588913429118;
            6'd63: xpb[97] = 1024'd96537487747093464985602565724113168147727469976943518578590090691742172938723145825688994076351937528329461978638453619097275539998905302758982617083584489869982240507388925448940476995627533561822974933264593123498207941010770871487066053665543815506432006842439252848615851972894757235837894457231572433512;
        endcase
    end

    always_comb begin
        case(flag[32][16:12])
            5'd0: xpb[98] = 1024'd0;
            5'd1: xpb[98] = 1024'd117762955121511574175659579053831541093675275393360984608112450078115365419863059078480100524334932458849477154086285174095496396322891154319468075293852662873266192669342911144579252692624352463012259870044545370913157408363465134997174811609953947382219801143766393057340949317532552274044637198874231437906;
            5'd2: xpb[98] = 1024'd111459214558898406952520230702848649442652123660986285088093045091253835502416979246945129834012190608255804900715076913611928951804561974083776025571374284812841710769114604951528266193731499204714322131701850895461953966506033497029371053536678445497619698873415728084575370561136471530970584571122868391481;
            5'd3: xpb[98] = 1024'd105155473996285239729380882351865757791628971928611585568073640104392305584970899415410159143689448757662132647343868653128361507286232793848083975848895906752417228868886298758477279694838645946416384393359156420010750524648601859061567295463402943613019596603065063111809791804740390787896531943371505345056;
            5'd4: xpb[98] = 1024'd98851733433672072506241534000882866140605820196236886048054235117530775667524819583875188453366706907068460393972660392644794062767903613612391926126417528691992746968657992565426293195945792688118446655016461944559547082791170221093763537390127441728419494332714398139044213048344310044822479315620142298631;
            5'd5: xpb[98] = 1024'd92547992871058905283102185649899974489582668463862186528034830130669245750078739752340217763043965056474788140601452132161226618249574433376699876403939150631568265068429686372375306697052939429820508916673767469108343640933738583125959779316851939843819392062363733166278634291948229301748426687868779252206;
            5'd6: xpb[98] = 1024'd86244252308445738059962837298917082838559516731487487008015425143807715832632659920805247072721223205881115887230243871677659173731245253141007826681460772571143783168201380179324320198160086171522571178331072993657140199076306945158156021243576437959219289792013068193513055535552148558674374060117416205781;
            5'd7: xpb[98] = 1024'd79940511745832570836823488947934191187536364999112787487996020156946185915186580089270276382398481355287443633859035611194091729212916072905315776958982394510719301267973073986273333699267232913224633439988378518205936757218875307190352263170300936074619187521662403220747476779156067815600321432366053159356;
            5'd8: xpb[98] = 1024'd73636771183219403613684140596951299536513213266738087967976615170084655997740500257735305692075739504693771380487827350710524284694586892669623727236504016450294819367744767793222347200374379654926695701645684042754733315361443669222548505097025434190019085251311738247981898022759987072526268804614690112931;
            5'd9: xpb[98] = 1024'd67333030620606236390544792245968407885490061534363388447957210183223126080294420426200335001752997654100099127116619090226956840176257712433931677514025638389870337467516461600171360701481526396628757963302989567303529873504012031254744747023749932305418982980961073275216319266363906329452216176863327066506;
            5'd10: xpb[98] = 1024'd61029290057993069167405443894985516234466909801988688927937805196361596162848340594665364311430255803506426873745410829743389395657928532198239627791547260329445855567288155407120374202588673138330820224960295091852326431646580393286940988950474430420818880710610408302450740509967825586378163549111964020081;
            5'd11: xpb[98] = 1024'd54725549495379901944266095544002624583443758069613989407918400209500066245402260763130393621107513952912754620374202569259821951139599351962547578069068882269021373667059849214069387703695819880032882486617600616401122989789148755319137230877198928536218778440259743329685161753571744843304110921360600973656;
            5'd12: xpb[98] = 1024'd48421808932766734721126747193019732932420606337239289887898995222638536327956180931595422930784772102319082367002994308776254506621270171726855528346590504208596891766831543021018401204802966621734944748274906140949919547931717117351333472803923426651618676169909078356919582997175664100230058293609237927231;
            5'd13: xpb[98] = 1024'd42118068370153567497987398842036841281397454604864590367879590235777006410510101100060452240462030251725410113631786048292687062102940991491163478624112126148172409866603236827967414705910113363437007009932211665498716106074285479383529714730647924767018573899558413384154004240779583357156005665857874880806;
            5'd14: xpb[98] = 1024'd35814327807540400274848050491053949630374302872489890847860185248915476493064021268525481550139288401131737860260577787809119617584611811255471428901633748087747927966374930634916428207017260105139069271589517190047512664216853841415725956657372422882418471629207748411388425484383502614081953038106511834381;
            5'd15: xpb[98] = 1024'd29510587244927233051708702140071057979351151140115191327840780262053946575617941436990510859816546550538065606889369527325552173066282631019779379179155370027323446066146624441865441708124406846841131533246822714596309222359422203447922198584096920997818369358857083438622846727987421871007900410355148787956;
            5'd16: xpb[98] = 1024'd23206846682314065828569353789088166328327999407740491807821375275192416658171861605455540169493804699944393353518161266841984728547953450784087329456676991966898964165918318248814455209231553588543193794904128239145105780501990565480118440510821419113218267088506418465857267971591341127933847782603785741531;
            5'd17: xpb[98] = 1024'd16903106119700898605430005438105274677304847675365792287801970288330886740725781773920569479171062849350721100146953006358417284029624270548395279734198613906474482265690012055763468710338700330245256056561433763693902338644558927512314682437545917228618164818155753493091689215195260384859795154852422695106;
            5'd18: xpb[98] = 1024'd10599365557087731382290657087122383026281695942991092767782565301469356823279701942385598788848320998757048846775744745874849839511295090312703230011720235846050000365461705862712482211445847071947318318218739288242698896787127289544510924364270415344018062547805088520326110458799179641785742527101059648681;
            5'd19: xpb[98] = 1024'd4295624994474564159151308736139491375258544210616393247763160314607826905833622110850628098525579148163376593404536485391282394992965910077011180289241857785625518465233399669661495712552993813649380579876044812791495454929695651576707166290994913459417960277454423547560531702403098898711689899349696602256;
            5'd20: xpb[98] = 1024'd122058580115986138334810887789971032468933819603977377855875610392723192325696681189330728622860511607012853747490821659486778791315857064396479255583094520658891711134576310814240748405177346276661640449920590183704652863293160786573881977900948860841637761421220816604901481019935651172756327098223928040162;
            5'd21: xpb[98] = 1024'd115754839553372971111671539438988140817910667871602678335856205405861662408250601357795757932537769756419181494119613399003211346797527884160787205860616142598467229234348004621189761906284493018363702711577895708253449421435729148606078219827673358957037659150870151632135902263539570429682274470472564993737;
            5'd22: xpb[98] = 1024'd109451098990759803888532191088005249166887516139227978815836800419000132490804521526260787242215027905825509240748405138519643902279198703925095156138137764538042747334119698428138775407391639760065764973235201232802245979578297510638274461754397857072437556880519486659370323507143489686608221842721201947312;
            5'd23: xpb[98] = 1024'd103147358428146636665392842737022357515864364406853279295817395432138602573358441694725816551892286055231836987377196878036076457760869523689403106415659386477618265433891392235087788908498786501767827234892506757351042537720865872670470703681122355187837454610168821686604744750747408943534169214969838900887;
            5'd24: xpb[98] = 1024'd96843617865533469442253494386039465864841212674478579775797990445277072655912361863190845861569544204638164734005988617552509013242540343453711056693181008417193783533663086042036802409605933243469889496549812281899839095863434234702666945607846853303237352339818156713839165994351328200460116587218475854462;
            5'd25: xpb[98] = 1024'd90539877302920302219114146035056574213818060942103880255778585458415542738466282031655875171246802354044492480634780357068941568724211163218019006970702630356769301633434779848985815910713079985171951758207117806448635654006002596734863187534571351418637250069467491741073587237955247457386063959467112808037;
            5'd26: xpb[98] = 1024'd84236136740307134995974797684073682562794909209729180735759180471554012821020202200120904480924060503450820227263572096585374124205881982982326957248224252296344819733206473655934829411820226726874014019864423330997432212148570958767059429461295849534037147799116826768308008481559166714312011331715749761612;
            5'd27: xpb[98] = 1024'd77932396177693967772835449333090790911771757477354481215739775484692482903574122368585933790601318652857147973892363836101806679687552802746634907525745874235920337832978167462883842912927373468576076281521728855546228770291139320799255671388020347649437045528766161795542429725163085971237958703964386715187;
            5'd28: xpb[98] = 1024'd71628655615080800549696100982107899260748605744979781695720370497830952986128042537050963100278576802263475720521155575618239235169223622510942857803267496175495855932749861269832856414034520210278138543179034380095025328433707682831451913314744845764836943258415496822776850968767005228163906076213023668762;
            5'd29: xpb[98] = 1024'd65324915052467633326556752631125007609725454012605082175700965510969423068681962705515992409955834951669803467149947315134671790650894442275250808080789118115071374032521555076781869915141666951980200804836339904643821886576276044863648155241469343880236840988064831850011272212370924485089853448461660622337;
            5'd30: xpb[98] = 1024'd59021174489854466103417404280142115958702302280230382655681560524107893151235882873981021719633093101076131213778739054651104346132565262039558758358310740054646892132293248883730883416248813693682263066493645429192618444718844406895844397168193841995636738717714166877245693455974843742015800820710297575912;
            5'd31: xpb[98] = 1024'd52717433927241298880278055929159224307679150547855683135662155537246363233789803042446051029310351250482458960407530794167536901614236081803866708635832361994222410232064942690679896917355960435384325328150950953741415002861412768928040639094918340111036636447363501904480114699578762998941748192958934529487;
        endcase
    end

    always_comb begin
        case(flag[33][5:0])
            6'd0: xpb[99] = 1024'd0;
            6'd1: xpb[99] = 1024'd23206846682314065828569353789088166328327999407740491807821375275192416658171861605455540169493804699944393353518161266841984728547953450784087329456676991966898964165918318248814455209231553588543193794904128239145105780501990565480118440510821419113218267088506418465857267971591341127933847782603785741531;
            6'd2: xpb[99] = 1024'd46413693364628131657138707578176332656655998815480983615642750550384833316343723210911080338987609399888786707036322533683969457095906901568174658913353983933797928331836636497628910418463107177086387589808256478290211561003981130960236881021642838226436534177012836931714535943182682255867695565207571483062;
            6'd3: xpb[99] = 1024'd69620540046942197485708061367264498984983998223221475423464125825577249974515584816366620508481414099833180060554483800525954185643860352352261988370030975900696892497754954746443365627694660765629581384712384717435317341505971696440355321532464257339654801265519255397571803914774023383801543347811357224593;
            6'd4: xpb[99] = 1024'd92827386729256263314277415156352665313311997630961967231285501100769666632687446421822160677975218799777573414072645067367938914191813803136349317826707967867595856663673272995257820836926214354172775179616512956580423122007962261920473762043285676452873068354025673863429071886365364511735391130415142966124;
            6'd5: xpb[99] = 1024'd116034233411570329142846768945440831641639997038702459039106876375962083290859308027277700847469023499721966767590806334209923642739767253920436647283384959834494820829591591244072276046157767942715968974520641195725528902509952827400592202554107095566091335442532092329286339857956705639669238913018928707655;
            6'd6: xpb[99] = 1024'd15174384409759653572617195329714565225269569320707266718796396586177604611722030722718169802305153890223210713651474166472844530446500370149363851723730910867703110425938692155256492063872115809948965161037529588506273832791046619915732073381699065412489699116921452765037079755619413750484396868997119964855;
            6'd7: xpb[99] = 1024'd38381231092073719401186549118802731553597568728447758526617771861370021269893892328173709971798958590167604067169635433314829258994453820933451181180407902834602074591857010404070947273103669398492158955941657827651379613293037185395850513892520484525707966205427871230894347727210754878418244651600905706386;
            6'd8: xpb[99] = 1024'd61588077774387785229755902907890897881925568136188250334439147136562437928065753933629250141292763290111997420687796700156813987542407271717538510637084894801501038757775328652885402482335222987035352750845786066796485393795027750875968954403341903638926233293934289696751615698802096006352092434204691447917;
            6'd9: xpb[99] = 1024'd84794924456701851058325256696979064210253567543928742142260522411754854586237615539084790310786567990056390774205957966998798716090360722501625840093761886768400002923693646901699857691566776575578546545749914305941591174297018316356087394914163322752144500382440708162608883670393437134285940216808477189448;
            6'd10: xpb[99] = 1024'd108001771139015916886894610486067230538581566951669233950081897686947271244409477144540330480280372690000784127724119233840783444638314173285713169550438878735298967089611965150514312900798330164121740340654042545086696954799008881836205835424984741865362767470947126628466151641984778262219787999412262930979;
            6'd11: xpb[99] = 1024'd7141922137205241316665036870340964122211139233674041629771417897162792565272199839980799435116503080502028073784787066103704332345047289514640373990784829768507256685959066061698528918512678031354736527170930937867441885080102674351345706252576711711761131145336487064216891539647486373034945955390454188179;
            6'd12: xpb[99] = 1024'd30348768819519307145234390659429130450539138641414533437592793172355209223444061445436339604610307780446421427302948332945689060893000740298727703447461821735406220851877384310512984127744231619897930322075059177012547665582093239831464146763398130824979398233842905530074159511238827500968793737994239929710;
            6'd13: xpb[99] = 1024'd53555615501833372973803744448517296778867138049155025245414168447547625881615923050891879774104112480390814780821109599787673789440954191082815032904138813702305185017795702559327439336975785208441124116979187416157653446084083805311582587274219549938197665322349323995931427482830168628902641520598025671241;
            6'd14: xpb[99] = 1024'd76762462184147438802373098237605463107195137456895517053235543722740042539787784656347419943597917180335208134339270866629658517988907641866902362360815805669204149183714020808141894546207338796984317911883315655302759226586074370791701027785040969051415932410855742461788695454421509756836489303201811412772;
            6'd15: xpb[99] = 1024'd99969308866461504630942452026693629435523136864636008861056918997932459197959646261802960113091721880279601487857432133471643246536861092650989691817492797636103113349632339056956349755438892385527511706787443894447865007088064936271819468295862388164634199499362160927645963426012850884770337085805597154303;
            6'd16: xpb[99] = 1024'd123176155548775570459511805815781795763851136272376500668878294273124875856131507867258500282585526580223994841375593400313627975084814543435077021274169789603002077515550657305770804964670445974070705501691572133592970787590055501751937908806683807277852466587868579393503231397604192012704184868409382895834;
            6'd17: xpb[99] = 1024'd22316306546964894889282232200055529347480708554381308348567814483340397176994230562698969237421656970725238787436261232576548862791547659664004225714515740636210367111897758216955020982384793841303701688208460526373715717871149294267077779634275777124250830262257939829253971295266900123519342824387574153034;
            6'd18: xpb[99] = 1024'd45523153229278960717851585989143695675808707962121800156389189758532813835166092168154509406915461670669632140954422499418533591339501110448091555171192732603109331277816076465769476191616347429846895483112588765518821498373139859747196220145097196237469097350764358295111239266858241251453190606991359894565;
            6'd19: xpb[99] = 1024'd68729999911593026546420939778231862004136707369862291964210565033725230493337953773610049576409266370614025494472583766260518319887454561232178884627869724570008295443734394714583931400847901018390089278016717004663927278875130425227314660655918615350687364439270776760968507238449582379387038389595145636096;
            6'd20: xpb[99] = 1024'd91936846593907092374990293567320028332464706777602783772031940308917647151509815379065589745903071070558418847990745033102503048435408012016266214084546716536907259609652712963398386610079454606933283072920845243809033059377120990707433101166740034463905631527777195226825775210040923507320886172198931377627;
            6'd21: xpb[99] = 1024'd115143693276221158203559647356408194660792706185343275579853315584110063809681676984521129915396875770502812201508906299944487776983361462800353543541223708503806223775571031212212841819311008195476476867824973482954138839879111556187551541677561453577123898616283613692683043181632264635254733954802717119158;
            6'd22: xpb[99] = 1024'd14283844274410482633330073740681928244422278467348083259542835794325585130544399679961598870233006161004056147569574132207408664690094579029280747981569659537014513371918132123397057837025356062709473054341861875734883770160205348702691412505153423423522262290672974128433783079294972746069891910780908376358;
            6'd23: xpb[99] = 1024'd37490690956724548461899427529770094572750277875088575067364211069518001788716261285417139039726810860948449501087735399049393393238048029813368077438246651503913477537836450372211513046256909651252666849245990114879989550662195914182809853015974842536740529379179392594291051050886313874003739693384694117889;
            6'd24: xpb[99] = 1024'd60697537639038614290468781318858260901078277282829066875185586344710418446888122890872679209220615560892842854605896665891378121786001480597455406894923643470812441703754768621025968255488463239795860644150118354025095331164186479662928293526796261649958796467685811060148319022477655001937587475988479859420;
            6'd25: xpb[99] = 1024'd83904384321352680119038135107946427229406276690569558683006961619902835105059984496328219378714420260837236208124057932733362850333954931381542736351600635437711405869673086869840423464720016828339054439054246593170201111666177045143046734037617680763177063556192229526005586994068996129871435258592265600951;
            6'd26: xpb[99] = 1024'd107111231003666745947607488897034593557734276098310050490828336895095251763231846101783759548208224960781629561642219199575347578881908382165630065808277627404610370035591405118654878673951570416882248233958374832315306892168167610623165174548439099876395330644698647991862854965660337257805283041196051342482;
            6'd27: xpb[99] = 1024'd6251382001856070377377915281308327141363848380314858170517857105310773084094568797224228503044355351282873507702887031838268466588641498394557270248623578437818659631938506029839094691665918284115244420475263225096051822449261403138305045376031069722793694319088008427613594863323045368620440997174242599682;
            6'd28: xpb[99] = 1024'd29458228684170136205947269070396493469691847788055349978339232380503189742266430402679768672538160051227266861221048298680253195136594949178644599705300570404717623797856824278653549900897471872658438215379391464241157602951251968618423485886852488836011961407594426893470862834914386496554288779778028341213;
            6'd29: xpb[99] = 1024'd52665075366484202034516622859484659798019847195795841786160607655695606400438292008135308842031964751171660214739209565522237923684548399962731929161977562371616587963775142527468005110129025461201632010283519703386263383453242534098541926397673907949230228496100845359328130806505727624488136562381814082744;
            6'd30: xpb[99] = 1024'd75871922048798267863085976648572826126347846603536333593981982930888023058610153613590849011525769451116053568257370832364222652232501850746819258618654554338515552129693460776282460319360579049744825805187647942531369163955233099578660366908495327062448495584607263825185398778097068752421984344985599824275;
            6'd31: xpb[99] = 1024'd99078768731112333691655330437660992454675846011276825401803358206080439716782015219046389181019574151060446921775532099206207380780455301530906588075331546305414516295611779025096915528592132638288019600091776181676474944457223665058778807419316746175666762673113682291042666749688409880355832127589385565806;
            6'd32: xpb[99] = 1024'd122285615413426399520224684226749158783003845419017317209624733481272856374953876824501929350513378851004840275293693366048192109328408752314993917532008538272313480461530097273911370737823686226831213394995904420821580724959214230538897247930138165288885029761620100756899934721279751008289679910193171307337;
            6'd33: xpb[99] = 1024'd21425766411615723949995110611022892366633417701022124889314253691488377695816599519942398305349509241506084221354361198311112997035141868543921121972354489305521770057877198185095586755538034094064209581512792813602325655240308023054037118757730135135283393436009461192650674618942459119104837866171362564537;
            6'd34: xpb[99] = 1024'd44632613093929789778564464400111058694961417108762616697135628966680794353988461125397938474843313941450477574872522465153097725583095319328008451429031481272420734223795516433910041964769587682607403376416921052747431435742298588534155559268551554248501660524515879658507942590533800247038685648775148306068;
            6'd35: xpb[99] = 1024'd67839459776243855607133818189199225023289416516503108504957004241873211012160322730853478644337118641394870928390683731995082454131048770112095780885708473239319698389713834682724497174001141271150597171321049291892537216244289154014273999779372973361719927613022298124365210562125141374972533431378934047599;
            6'd36: xpb[99] = 1024'd91046306458557921435703171978287391351617415924243600312778379517065627670332184336309018813830923341339264281908844998837067182679002220896183110342385465206218662555632152931538952383232694859693790966225177531037642996746279719494392440290194392474938194701528716590222478533716482502906381213982719789130;
            6'd37: xpb[99] = 1024'd114253153140871987264272525767375557679945415331984092120599754792258044328504045941764558983324728041283657635427006265679051911226955671680270439799062457173117626721550471180353407592464248448236984761129305770182748777248270284974510880801015811588156461790035135056079746505307823630840228996586505530661;
            6'd38: xpb[99] = 1024'd13393304139061311694042952151649291263574987613988899800289275002473565649366768637205027938160858431784901581487674097941972798933688787909197644239408408206325916317897572091537623610178596315469980947646194162963493707529364077489650751628607781434554825464424495491830486402970531741655386952564696787861;
            6'd39: xpb[99] = 1024'd36600150821375377522612305940737457591902987021729391608110650277665982307538630242660568107654663131729294935005835364783957527481642238693284973696085400173224880483815890340352078819410149904013174742550322402108599488031354642969769192139429200547773092552930913957687754374561872869589234735168482529392;
            6'd40: xpb[99] = 1024'd59806997503689443351181659729825623920230986429469883415932025552858398965710491848116108277148467831673688288523996631625942256029595689477372303152762392140123844649734208589166534028641703492556368537454450641253705268533345208449887632650250619660991359641437332423545022346153213997523082517772268270923;
            6'd41: xpb[99] = 1024'd83013844186003509179751013518913790248558985837210375223753400828050815623882353453571648446642272531618081642042157898467926984577549140261459632609439384107022808815652526837980989237873257081099562332358578880398811049035335773930006073161072038774209626729943750889402290317744555125456930300376054012454;
            6'd42: xpb[99] = 1024'd106220690868317575008320367308001956576886985244950867031574776103243232282054215059027188616136077231562474995560319165309911713125502591045546962066116376073921772981570845086795444447104810669642756127262707119543916829537326339410124513671893457887427893818450169355259558289335896253390778082979839753985;
            6'd43: xpb[99] = 1024'd5360841866506899438090793692275690160516557526955674711264296313458753602916937754467657570972207622063718941620986997572832600832235707274474166506462327107130062577917945997979660464819158536875752313779595512324661759818420131925264384499485427733826257492839529791010298186998604364205936038958031011185;
            6'd44: xpb[99] = 1024'd28567688548820965266660147481363856488844556934696166519085671588651170261088799359923197740466012322008112295139148264414817329380189158058561495963139319074029026743836264246794115674050712125418946108683723751469767540320410697405382825010306846847044524581345948256867566158589945492139783821561816752716;
            6'd45: xpb[99] = 1024'd51774535231135031095229501270452022817172556342436658326907046863843586919260660965378737909959817021952505648657309531256802057928142608842648825419816311040927990909754582495608570883282265713962139903587851990614873320822401262885501265521128265960262791669852366722724834130181286620073631604165602494247;
            6'd46: xpb[99] = 1024'd74981381913449096923798855059540189145500555750177150134728422139036003577432522570834278079453621721896899002175470798098786786476096059626736154876493303007826955075672900744423026092513819302505333698491980229759979101324391828365619706031949685073481058758358785188582102101772627748007479386769388235778;
            6'd47: xpb[99] = 1024'd98188228595763162752368208848628355473828555157917641942549797414228420235604384176289818248947426421841292355693632064940771515024049510410823484333170294974725919241591218993237481301745372891048527493396108468905084881826382393845738146542771104186699325846865203654439370073363968875941327169373173977309;
            6'd48: xpb[99] = 1024'd121395075278077228580937562637716521802156554565658133750371172689420836893776245781745358418441231121785685709211793331782756243572002961194910813789847286941624883407509537242051936510976926479591721288300236708050190662328372959325856587053592523299917592935371622120296638044955310003875174951976959718840;
            6'd49: xpb[99] = 1024'd20535226276266553010707989021990255385786126847662941430060692899636358214638968477185827373277361512286929655272461164045677131278736077423838018230193237974833173003856638153236152528691274346824717474817125100830935592609466751840996457881184493146315956609760982556047377942618018114690332907955150976040;
            6'd50: xpb[99] = 1024'd43742072958580618839277342811078421714114126255403433237882068174828774872810830082641367542771166212231323008790622430887661859826689528207925347686870229941732137169774956402050607737922827935367911269721253339976041373111457317321114898392005912259534223698267401021904645914209359242624180690558936717571;
            6'd51: xpb[99] = 1024'd66948919640894684667846696600166588042442125663143925045703443450021191530982691688096907712264970912175716362308783697729646588374642978992012677143547221908631101335693274650865062947154381523911105064625381579121147153613447882801233338902827331372752490786773819487761913885800700370558028473162722459102;
            6'd52: xpb[99] = 1024'd90155766323208750496416050389254754370770125070884416853524818725213608189154553293552447881758775612120109715826944964571631316922596429776100006600224213875530065501611592899679518156385935112454298859529509818266252934115438448281351779413648750485970757875280237953619181857392041498491876255766508200633;
            6'd53: xpb[99] = 1024'd113362613005522816324985404178342920699098124478624908661346194000406024847326414899007988051252580312064503069345106231413616045470549880560187336056901205842429029667529911148493973365617488700997492654433638057411358714617429013761470219924470169599189024963786656419476449828983382626425724038370293942164;
            6'd54: xpb[99] = 1024'd12502764003712140754755830562616654282727696760629716341035714210621546168189137594448457006088710702565747015405774063676536933177282996789114540497247156875637319263877012059678189383331836568230488840950526450192103644898522806276610090752062139445587388638176016855227189726646090737240881994348485199364;
            6'd55: xpb[99] = 1024'd35709610686026206583325184351704820611055696168370208148857089485813962826360999199903997175582515402510140368923935330518521661725236447573201869953924148842536283429795330308492644592563390156773682635854654689337209425400513371756728531262883558558805655726682435321084457698237431865174729776952270940895;
            6'd56: xpb[99] = 1024'd58916457368340272411894538140792986939383695576110699956678464761006379484532860805359537345076320102454533722442096597360506390273189898357289199410601140809435247595713648557307099801794943745316876430758782928482315205902503937236846971773704977672023922815188853786941725669828772993108577559556056682426;
            6'd57: xpb[99] = 1024'd82123304050654338240463891929881153267711694983851191764499840036198796142704722410815077514570124802398927075960257864202491118821143349141376528867278132776334211761631966806121555011026497333860070225662911167627420986404494502716965412284526396785242189903695272252798993641420114121042425342159842423957;
            6'd58: xpb[99] = 1024'd105330150732968404069033245718969319596039694391591683572321215311391212800876584016270617684063929502343320429478419131044475847369096799925463858323955124743233175927550285054936010220258050922403264020567039406772526766906485068197083852795347815898460456992201690718656261613011455248976273124763628165488;
            6'd59: xpb[99] = 1024'd4470301731157728498803672103243053179669266673596491252010735521606734121739306711711086638900059892844564375539086963307396735075829916154391062764301075776441465523897385966120226237972398789636260207083927799553271697187578860712223723622939785744858820666591051154407001510674163359791431080741819422688;
            6'd60: xpb[99] = 1024'd27677148413471794327373025892331219507997266081336983059832110796799150779911168317166626808393864592788957729057248230149381463623783366938478392220978067743340429689815704214934681447203952378179454001988056038698377477689569426192342164133761204858077087755097469620264269482265504487725278863345605164219;
            6'd61: xpb[99] = 1024'd50883995095785860155942379681419385836325265489077474867653486071991567438083029922622166977887669292733351082575409496991366192171736817722565721677655059710239393855734022463749136656435505966722647796892184277843483258191559991672460604644582623971295354843603888086121537453856845615659126645949390905750;
            6'd62: xpb[99] = 1024'd74090841778099925984511733470507552164653264896817966675474861347183984096254891528077707147381473992677744436093570763833350920719690268506653051134332051677138358021652340712563591865667059555265841591796312516988589038693550557152579045155404043084513621932110306551978805425448186743592974428553176647281;
            6'd63: xpb[99] = 1024'd97297688460413991813081087259595718492981264304558458483296236622376400754426753133533247316875278692622137789611732030675335649267643719290740380591009043644037322187570658961378047074898613143809035386700440756133694819195541122632697485666225462197731889020616725017836073397039527871526822211156962388812;
        endcase
    end

    always_comb begin
        case(flag[33][11:6])
            6'd0: xpb[100] = 1024'd0;
            6'd1: xpb[100] = 1024'd120504535142728057641650441048683884821309263712298950291117611897568817412598614738988787486369083392566531143129893297517320377815597170074827710047686035610936286353488977210192502284130166732352229181604568995278800599697531688112815926177046881310950156109123143483693341368630868999460669993760748130343;
            6'd2: xpb[100] = 1024'd116942374601331373884501954692553336897920100298862216454103368730160739487888090567962503758080492475689912878802293160455576914789974005594495295079041030288181898137406737082754765376743127743394260754821898144193240349174166603260653282670864313355080408804129228937280154663333104981802650160895901776355;
            6'd3: xpb[100] = 1024'd113380214059934690127353468336422788974530936885425482617089125562752661563177566396936220029791901558813294614474693023393833451764350841114162880110396024965427509921324496955317028469356088754436292328039227293107680098650801518408490639164681745399210661499135314390866967958035340964144630328031055422367;
            6'd4: xpb[100] = 1024'd109818053518538006370204981980292241051141773471988748780074882395344583638467042225909936301503310641936676350147092886332089988738727676633830465141751019642673121705242256827879291561969049765478323901256556442022119848127436433556327995658499177443340914194141399844453781252737576946486610495166209068379;
            6'd5: xpb[100] = 1024'd106255892977141322613056495624161693127752610058552014943060639227936505713756518054883652573214719725060058085819492749270346525713104512153498050173106014319918733489160016700441554654582010776520355474473885590936559597604071348704165352152316609487471166889147485298040594547439812928828590662301362714391;
            6'd6: xpb[100] = 1024'd102693732435744638855908009268031145204363446645115281106046396060528427789045993883857368844926128808183439821491892612208603062687481347673165635204461008997164345273077776573003817747194971787562387047691214739850999347080706263852002708646134041531601419584153570751627407842142048911170570829436516360403;
            6'd7: xpb[100] = 1024'd99131571894347955098759522911900597280974283231678547269032152893120349864335469712831085116637537891306821557164292475146859599661858183192833220235816003674409957056995536445566080839807932798604418620908543888765439096557341178999840065139951473575731672279159656205214221136844284893512550996571670006415;
            6'd8: xpb[100] = 1024'd95569411352951271341611036555770049357585119818241813432017909725712271939624945541804801388348946974430203292836692338085116136636235018712500805267170998351655568840913296318128343932420893809646450194125873037679878846033976094147677421633768905619861924974165741658801034431546520875854531163706823652427;
            6'd9: xpb[100] = 1024'd92007250811554587584462550199639501434195956404805079595003666558304194014914421370778517660060356057553585028509092201023372673610611854232168390298525993028901180624831056190690607025033854820688481767343202186594318595510611009295514778127586337663992177669171827112387847726248756858196511330841977298439;
            6'd10: xpb[100] = 1024'd88445090270157903827314063843508953510806792991368345757989423390896116090203897199752233931771765140676966764181492063961629210584988689751835975329880987706146792408748816063252870117646815831730513340560531335508758344987245924443352134621403769708122430364177912565974661020950992840538491497977130944451;
            6'd11: xpb[100] = 1024'd84882929728761220070165577487378405587417629577931611920975180223488038165493373028725950203483174223800348499853891926899885747559365525271503560361235982383392404192666575935815133210259776842772544913777860484423198094463880839591189491115221201752252683059183998019561474315653228822880471665112284590463;
            6'd12: xpb[100] = 1024'd81320769187364536313017091131247857664028466164494878083960937056079960240782848857699666475194583306923730235526291789838142284533742360791171145392590977060638015976584335808377396302872737853814576486995189633337637843940515754739026847609038633796382935754190083473148287610355464805222451832247438236475;
            6'd13: xpb[100] = 1024'd77758608645967852555868604775117309740639302751058144246946693888671882316072324686673382746905992390047111971198691652776398821508119196310838730423945971737883627760502095680939659395485698864856608060212518782252077593417150669886864204102856065840513188449196168926735100905057700787564431999382591882487;
            6'd14: xpb[100] = 1024'd74196448104571168798720118418986761817250139337621410409932450721263804391361800515647099018617401473170493706871091515714655358482496031830506315455300966415129239544419855553501922488098659875898639633429847931166517342893785585034701560596673497884643441144202254380321914199759936769906412166517745528499;
            6'd15: xpb[100] = 1024'd70634287563174485041571632062856213893860975924184676572918207553855726466651276344620815290328810556293875442543491378652911895456872867350173900486655961092374851328337615426064185580711620886940671206647177080080957092370420500182538917090490929928773693839208339833908727494462172752248392333652899174511;
            6'd16: xpb[100] = 1024'd67072127021777801284423145706725665970471812510747942735903964386447648541940752173594531562040219639417257178215891241591168432431249702869841485518010955769620463112255375298626448673324581897982702779864506228995396841847055415330376273584308361972903946534214425287495540789164408734590372500788052820523;
            6'd17: xpb[100] = 1024'd63509966480381117527274659350595118047082649097311208898889721219039570617230228002568247833751628722540638913888291104529424969405626538389509070549365950446866074896173135171188711765937542909024734353081835377909836591323690330478213630078125794017034199229220510741082354083866644716932352667923206466535;
            6'd18: xpb[100] = 1024'd59947805938984433770126172994464570123693485683874475061875478051631492692519703831541964105463037805664020649560690967467681506380003373909176655580720945124111686680090895043750974858550503920066765926299164526824276340800325245626050986571943226061164451924226596194669167378568880699274332835058360112547;
            6'd19: xpb[100] = 1024'd56385645397587750012977686638334022200304322270437741224861234884223414767809179660515680377174446888787402385233090830405938043354380209428844240612075939801357298464008654916313237951163464931108797499516493675738716090276960160773888343065760658105294704619232681648255980673271116681616313002193513758559;
            6'd20: xpb[100] = 1024'd52823484856191066255829200282203474276915158857001007387846991716815336843098655489489396648885855971910784120905490693344194580328757044948511825643430934478602910247926414788875501043776425942150829072733822824653155839753595075921725699559578090149424957314238767101842793967973352663958293169328667404571;
            6'd21: xpb[100] = 1024'd49261324314794382498680713926072926353525995443564273550832748549407258918388131318463112920597265055034165856577890556282451117303133880468179410674785929155848522031844174661437764136389386953192860645951151973567595589230229991069563056053395522193555210009244852555429607262675588646300273336463821050583;
            6'd22: xpb[100] = 1024'd45699163773397698741532227569942378430136832030127539713818505381999180993677607147436829192308674138157547592250290419220707654277510715987846995706140923833094133815761934534000027229002347964234892219168481122482035338706864906217400412547212954237685462704250938009016420557377824628642253503598974696595;
            6'd23: xpb[100] = 1024'd42137003232001014984383741213811830506747668616690805876804262214591103068967082976410545464020083221280929327922690282158964191251887551507514580737495918510339745599679694406562290321615308975276923792385810271396475088183499821365237769041030386281815715399257023462603233852080060610984233670734128342607;
            6'd24: xpb[100] = 1024'd38574842690604331227235254857681282583358505203254072039790019047183025144256558805384261735731492304404311063595090145097220728226264387027182165768850913187585357383597454279124553414228269986318955365603139420310914837660134736513075125534847818325945968094263108916190047146782296593326213837869281988619;
            6'd25: xpb[100] = 1024'd35012682149207647470086768501550734659969341789817338202775775879774947219546034634357978007442901387527692799267490008035477265200641222546849750800205907864830969167515214151686816506841230997360986938820468569225354587136769651660912482028665250370076220789269194369776860441484532575668194005004435634631;
            6'd26: xpb[100] = 1024'd31450521607810963712938282145420186736580178376380604365761532712366869294835510463331694279154310470651074534939889870973733802175018058066517335831560902542076580951432974024249079599454192008403018512037797718139794336613404566808749838522482682414206473484275279823363673736186768558010174172139589280643;
            6'd27: xpb[100] = 1024'd27888361066414279955789795789289638813191014962943870528747289544958791370124986292305410550865719553774456270612289733911990339149394893586184920862915897219322192735350733896811342692067153019445050085255126867054234086090039481956587195016300114458336726179281365276950487030889004540352154339274742926655;
            6'd28: xpb[100] = 1024'd24326200525017596198641309433159090889801851549507136691733046377550713445414462121279126822577128636897838006284689596850246876123771729105852505894270891896567804519268493769373605784680114030487081658472456015968673835566674397104424551510117546502466978874287450730537300325591240522694134506409896572667;
            6'd29: xpb[100] = 1024'd20764039983620912441492823077028542966412688136070402854718803210142635520703937950252843094288537720021219741957089459788503413098148564625520090925625886573813416303186253641935868877293075041529113231689785164883113585043309312252261908003934978546597231569293536184124113620293476505036114673545050218679;
            6'd30: xpb[100] = 1024'd17201879442224228684344336720897995043023524722633669017704560042734557595993413779226559365999946803144601477629489322726759950072525400145187675956980881251059028087104013514498131969906036052571144804907114313797553334519944227400099264497752410590727484264299621637710926914995712487378094840680203864691;
            6'd31: xpb[100] = 1024'd13639718900827544927195850364767447119634361309196935180690316875326479671282889608200275637711355886267983213301889185665016487046902235664855260988335875928304639871021773387060395062518997063613176378124443462711993083996579142547936620991569842634857736959305707091297740209697948469720075007815357510703;
            6'd32: xpb[100] = 1024'd10077558359430861170047364008636899196245197895760201343676073707918401746572365437173991909422764969391364948974289048603273024021279071184522846019690870605550251654939533259622658155131958074655207951341772611626432833473214057695773977485387274678987989654311792544884553504400184452062055174950511156715;
            6'd33: xpb[100] = 1024'd6515397818034177412898877652506351272856034482323467506661830540510323821861841266147708181134174052514746684646688911541529560995655906704190431051045865282795863438857293132184921247744919085697239524559101760540872582949848972843611333979204706723118242349317877998471366799102420434404035342085664802727;
            6'd34: xpb[100] = 1024'd2953237276637493655750391296375803349466871068886733669647587373102245897151317095121424452845583135638128420319088774479786097970032742223858016082400859960041475222775053004747184340357880096739271097776430909455312332426483887991448690473022138767248495044323963452058180093804656416746015509220818448739;
            6'd35: xpb[100] = 1024'd123457772419365551297400832345059688170776134781185683960765199270671063309749931834110211939214666528204659563448982071997106475785629912298685726130086895570977761576264030214939686624488046829091500279380999904734112932124015576104264616650069020078198651153447106935751521462435525416206685502981566579082;
            6'd36: xpb[100] = 1024'd119895611877968867540252345988929140247386971367748950123750956103262985385039407663083928210926075611328041299121381934935363012760006747818353311161441890248223373360181790087501949717101007840133531852598329053648552681600650491252101973143886452122328903848453192389338334757137761398548665670116720225094;
            6'd37: xpb[100] = 1024'd116333451336572183783103859632798592323997807954312216286736712935854907460328883492057644482637484694451423034793781797873619549734383583338020896192796884925468985144099549960064212809713968851175563425815658202562992431077285406399939329637703884166459156543459277842925148051839997380890645837251873871106;
            6'd38: xpb[100] = 1024'd112771290795175500025955373276668044400608644540875482449722469768446829535618359321031360754348893777574804770466181660811876086708760418857688481224151879602714596928017309832626475902326929862217594999032987351477432180553920321547776686131521316210589409238465363296511961346542233363232626004387027517118;
            6'd39: xpb[100] = 1024'd109209130253778816268806886920537496477219481127438748612708226601038751610907835150005077026060302860698186506138581523750132623683137254377356066255506874279960208711935069705188738994939890873259626572250316500391871930030555236695614042625338748254719661933471448750098774641244469345574606171522181163130;
            6'd40: xpb[100] = 1024'd105646969712382132511658400564406948553830317714002014775693983433630673686197310978978793297771711943821568241810981386688389160657514089897023651286861868957205820495852829577751002087552851884301658145467645649306311679507190151843451399119156180298849914628477534203685587935946705327916586338657334809142;
            6'd41: xpb[100] = 1024'd102084809170985448754509914208276400630441154300565280938679740266222595761486786807952509569483121026944949977483381249626645697631890925416691236318216863634451432279770589450313265180165812895343689718684974798220751428983825066991288755612973612342980167323483619657272401230648941310258566505792488455154;
            6'd42: xpb[100] = 1024'd98522648629588764997361427852145852707051990887128547101665497098814517836776262636926225841194530110068331713155781112564902234606267760936358821349571858311697044063688349322875528272778773906385721291902303947135191178460459982139126112106791044387110420018489705110859214525351177292600546672927642101166;
            6'd43: xpb[100] = 1024'd94960488088192081240212941496015304783662827473691813264651253931406439912065738465899942112905939193191713448828180975503158771580644596456026406380926852988942655847606109195437791365391734917427752865119633096049630927937094897286963468600608476431240672713495790564446027820053413274942526840062795747178;
            6'd44: xpb[100] = 1024'd91398327546795397483064455139884756860273664060255079427637010763998361987355214294873658384617348276315095184500580838441415308555021431975693991412281847666188267631523869068000054458004695928469784438336962244964070677413729812434800825094425908475370925408501876018032841114755649257284507007197949393190;
            6'd45: xpb[100] = 1024'd87836167005398713725915968783754208936884500646818345590622767596590284062644690123847374656328757359438476920172980701379671845529398267495361576443636842343433879415441628940562317550617656939511816011554291393878510426890364727582638181588243340519501178103507961471619654409457885239626487174333103039202;
            6'd46: xpb[100] = 1024'd84274006464002029968767482427623661013495337233381611753608524429182206137934165952821090928040166442561858655845380564317928382503775103015029161474991837020679491199359388813124580643230617950553847584771620542792950176366999642730475538082060772563631430798514046925206467704160121221968467341468256685214;
            6'd47: xpb[100] = 1024'd80711845922605346211618996071493113090106173819944877916594281261774128213223641781794807199751575525685240391517780427256184919478151938534696746506346831697925102983277148685686843735843578961595879157988949691707389925843634557878312894575878204607761683493520132378793280998862357204310447508603410331226;
            6'd48: xpb[100] = 1024'd77149685381208662454470509715362565166717010406508144079580038094366050288513117610768523471462984608808622127190180290194441456452528774054364331537701826375170714767194908558249106828456539972637910731206278840621829675320269473026150251069695636651891936188526217832380094293564593186652427675738563977238;
            6'd49: xpb[100] = 1024'd73587524839811978697322023359232017243327846993071410242565794926957972363802593439742239743174393691932003862862580153132697993426905609574031916569056821052416326551112668430811369921069500983679942304423607989536269424796904388173987607563513068696022188883532303285966907588266829168994407842873717623250;
            6'd50: xpb[100] = 1024'd70025364298415294940173537003101469319938683579634676405551551759549894439092069268715956014885802775055385598534980016070954530401282445093699501600411815729661938335030428303373633013682461994721973877640937138450709174273539303321824964057330500740152441578538388739553720882969065151336388010008871269262;
            6'd51: xpb[100] = 1024'd66463203757018611183025050646970921396549520166197942568537308592141816514381545097689672286597211858178767334207379879009211067375659280613367086631766810406907550118948188175935896106295423005764005450858266287365148923750174218469662320551147932784282694273544474193140534177671301133678368177144024915274;
            6'd52: xpb[100] = 1024'd62901043215621927425876564290840373473160356752761208731523065424733738589671020926663388558308620941302149069879779741947467604350036116133034671663121805084153161902865948048498159198908384016806037024075595436279588673226809133617499677044965364828412946968550559646727347472373537116020348344279178561286;
            6'd53: xpb[100] = 1024'd59338882674225243668728077934709825549771193339324474894508822257325660664960496755637104830020030024425530805552179604885724141324412951652702256694476799761398773686783707921060422291521345027848068597292924585194028422703444048765337033538782796872543199663556645100314160767075773098362328511414332207298;
            6'd54: xpb[100] = 1024'd55776722132828559911579591578579277626382029925887741057494579089917582740249972584610821101731439107548912541224579467823980678298789787172369841725831794438644385470701467793622685384134306038890100170510253734108468172180078963913174390032600228916673452358562730553900974061778009080704308678549485853310;
            6'd55: xpb[100] = 1024'd52214561591431876154431105222448729702992866512451007220480335922509504815539448413584537373442848190672294276896979330762237215273166622692037426757186789115889997254619227666184948476747267049932131743727582883022907921656713879061011746526417660960803705053568816007487787356480245063046288845684639499322;
            6'd56: xpb[100] = 1024'd48652401050035192397282618866318181779603703099014273383466092755101426890828924242558253645154257273795676012569379193700493752247543458211705011788541783793135609038536987538747211569360228060974163316944912031937347671133348794208849103020235093004933957748574901461074600651182481045388269012819793145334;
            6'd57: xpb[100] = 1024'd45090240508638508640134132510187633856214539685577539546451849587693348966118400071531969916865666356919057748241779056638750289221920293731372596819896778470381220822454747411309474661973189072016194890162241180851787420609983709356686459514052525049064210443580986914661413945884717027730249179954946791346;
            6'd58: xpb[100] = 1024'd41528079967241824882985646154057085932825376272140805709437606420285271041407875900505686188577075440042439483914178919577006826196297129251040181851251773147626832606372507283871737754586150083058226463379570329766227170086618624504523816007869957093194463138587072368248227240586953010072229347090100437358;
            6'd59: xpb[100] = 1024'd37965919425845141125837159797926538009436212858704071872423363252877193116697351729479402460288484523165821219586578782515263363170673964770707766882606767824872444390290267156434000847199111094100258036596899478680666919563253539652361172501687389137324715833593157821835040535289188992414209514225254083370;
            6'd60: xpb[100] = 1024'd34403758884448457368688673441795990086047049445267338035409120085469115191986827558453118731999893606289202955258978645453519900145050800290375351913961762502118056174208027028996263939812072105142289609814228627595106669039888454800198528995504821181454968528599243275421853829991424974756189681360407729382;
            6'd61: xpb[100] = 1024'd30841598343051773611540187085665442162657886031830604198394876918061037267276303387426835003711302689412584690931378508391776437119427635810042936945316757179363667958125786901558527032425033116184321183031557776509546418516523369948035885489322253225585221223605328729008667124693660957098169848495561375394;
            6'd62: xpb[100] = 1024'd27279437801655089854391700729534894239268722618393870361380633750652959342565779216400551275422711772535966426603778371330032974093804471329710521976671751856609279742043546774120790125037994127226352756248886925423986167993158285095873241983139685269715473918611414182595480419395896939440150015630715021406;
            6'd63: xpb[100] = 1024'd23717277260258406097243214373404346315879559204957136524366390583244881417855255045374267547134120855659348162276178234268289511068181306849378107008026746533854891525961306646683053217650955138268384329466216074338425917469793200243710598476957117313845726613617499636182293714098132921782130182765868667418;
        endcase
    end

    always_comb begin
        case(flag[33][16:12])
            5'd0: xpb[101] = 1024'd0;
            5'd1: xpb[101] = 1024'd20155116718861722340094728017273798392490395791520402687352147415836803493144730874347983818845529938782729897948578097206546048042558142369045692039381741211100503309879066519245316310263916149310415902683545223252865666946428115391547954970774549357975979308623585089769107008800368904124110349901022313430;
            5'd2: xpb[101] = 1024'd40310233437723444680189456034547596784980791583040805374704294831673606986289461748695967637691059877565459795897156194413092096085116284738091384078763482422201006619758133038490632620527832298620831805367090446505731333892856230783095909941549098715951958617247170179538214017600737808248220699802044626860;
            5'd3: xpb[101] = 1024'd60465350156585167020284184051821395177471187374561208062056442247510410479434192623043951456536589816348189693845734291619638144127674427107137076118145223633301509929637199557735948930791748447931247708050635669758597000839284346174643864912323648073927937925870755269307321026401106712372331049703066940290;
            5'd4: xpb[101] = 1024'd80620466875446889360378912069095193569961583166081610749408589663347213972578923497391935275382119755130919591794312388826184192170232569476182768157526964844402013239516266076981265241055664597241663610734180893011462667785712461566191819883098197431903917234494340359076428035201475616496441399604089253720;
            5'd5: xpb[101] = 1024'd100775583594308611700473640086368991962451978957602013436760737079184017465723654371739919094227649693913649489742890486032730240212790711845228460196908706055502516549395332596226581551319580746552079513417726116264328334732140576957739774853872746789879896543117925448845535044001844520620551749505111567150;
            5'd6: xpb[101] = 1024'd120930700313170334040568368103642790354942374749122416124112884495020820958868385246087902913073179632696379387691468583239276288255348854214274152236290447266603019859274399115471897861583496895862495416101271339517194001678568692349287729824647296147855875851741510538614642052802213424744662099406133880580;
            5'd7: xpb[101] = 1024'd17019121347907314981864168716102156002734343414907134683333176845880729114703977210420815517261035262035959878182553245866758495456686662028159719259341147544012848599582248297086974980330207323862713710397576716405698818404100034775857115112192396239011951746248037598277220987673949311750082622681561709679;
            5'd8: xpb[101] = 1024'd37174238066769037321958896733375954395224739206427537370685324261717532607848708084768799336106565200818689776131131343073304543499244804397205411298722888755113351909461314816332291290594123473173129613081121939658564485350528150167405070082966945596987931054871622688046327996474318215874192972582584023109;
            5'd9: xpb[101] = 1024'd57329354785630759662053624750649752787715134997947940058037471677554336100993438959116783154952095139601419674079709440279850591541802946766251103338104629966213855219340381335577607600858039622483545515764667162911430152296956265558953025053741494954963910363495207777815435005274687119998303322483606336539;
            5'd10: xpb[101] = 1024'd77484471504492482002148352767923551180205530789468342745389619093391139594138169833464766973797625078384149572028287537486396639584361089135296795377486371177314358529219447854822923911121955771793961418448212386164295819243384380950500980024516044312939889672118792867584542014075056024122413672384628649969;
            5'd11: xpb[101] = 1024'd97639588223354204342243080785197349572695926580988745432741766509227943087282900707812750792643155017166879469976865634692942687626919231504342487416868112388414861839098514374068240221385871921104377321131757609417161486189812496342048934995290593670915868980742377957353649022875424928246524022285650963399;
            5'd12: xpb[101] = 1024'd117794704942215926682337808802471147965186322372509148120093913925064746580427631582160734611488684955949609367925443731899488735669477373873388179456249853599515365148977580893313556531649788070414793223815302832670027153136240611733596889966065143028891848289365963047122756031675793832370634372186673276829;
            5'd13: xpb[101] = 1024'd13883125976952907623633609414930513612978291038293866679314206275924654736263223546493647215676540585289189858416528394526970942870815181687273746479300553876925193889285430074928633650396498498415011518111608209558531969861771954160166275253610243120047924183872490106785334966547529719376054895462101105928;
            5'd14: xpb[101] = 1024'd34038242695814629963728337432204312005468686829814269366666353691761458229407954420841631034522070524071919756365106491733516990913373324056319438518682295088025697199164496594173949960660414647725427420795153432811397636808200069551714230224384792478023903492496075196554441975347898623500165245363123419358;
            5'd15: xpb[101] = 1024'd54193359414676352303823065449478110397959082621334672054018501107598261722552685295189614853367600462854649654313684588940063038955931466425365130558064036299126200509043563113419266270924330797035843323478698656064263303754628184943262185195159341835999882801119660286323548984148267527624275595264145732788;
            5'd16: xpb[101] = 1024'd74348476133538074643917793466751908790449478412855074741370648523435065215697416169537598672213130401637379552262262686146609086998489608794410822597445777510226703818922629632664582581188246946346259226162243879317128970701056300334810140165933891193975862109743245376092655992948636431748385945165168046218;
            5'd17: xpb[101] = 1024'd94503592852399796984012521484025707182939874204375477428722795939271868708842147043885582491058660340420109450210840783353155135041047751163456514636827518721327207128801696151909898891452163095656675128845789102569994637647484415726358095136708440551951841418366830465861763001749005335872496295066190359648;
            5'd18: xpb[101] = 1024'd114658709571261519324107249501299505575430269995895880116074943355108672201986877918233566309904190279202839348159418880559701183083605893532502206676209259932427710438680762671155215201716079244967091031529334325822860304593912531117906050107482989909927820726990415555630870010549374239996606644967212673078;
            5'd19: xpb[101] = 1024'd10747130605998500265403050113758871223222238661680598675295235705968580357822469882566478914092045908542419838650503543187183390284943701346387773699259960209837539178988611852770292320462789672967309325825639702711365121319443873544475435395028090001083896621496942615293448945421110127002027168242640502177;
            5'd20: xpb[101] = 1024'd30902247324860222605497778131032669615712634453201001362647383121805383850967200756914462732937575847325149736599081640393729438327501843715433465738641701420938042488867678372015608630726705822277725228509184925964230788265871988936023390365802639359059875930120527705062555954221479031126137518143662815607;
            5'd21: xpb[101] = 1024'd51057364043721944945592506148306468008203030244721404049999530537642187344111931631262446551783105786107879634547659737600275486370059986084479157778023442632038545798746744891260924940990621971588141131192730149217096455212300104327571345336577188717035855238744112794831662963021847935250247868044685129037;
            5'd22: xpb[101] = 1024'd71212480762583667285687234165580266400693426036241806737351677953478990837256662505610430370628635724890609532496237834806821534412618128453524849817405183843139049108625811410506241251254538120898557033876275372469962122158728219719119300307351738075011834547367697884600769971822216839374358217945707442467;
            5'd23: xpb[101] = 1024'd91367597481445389625781962182854064793183821827762209424703825369315794330401393379958414189474165663673339430444815932013367582455176270822570541856786925054239552418504877929751557561518454270208972936559820595722827789105156335110667255278126287432987813855991282974369876980622585743498468567846729755897;
            5'd24: xpb[101] = 1024'd111522714200307111965876690200127863185674217619282612112055972785152597823546124254306398008319695602456069328393394029219913630497734413191616233896168666265340055728383944448996873871782370419519388839243365818975693456051584450502215210248900836790963793164614868064138983989422954647622578917747752069327;
            5'd25: xpb[101] = 1024'd7611135235044092907172490812587228833466186285067330671276265136012505979381716218639310612507551231795649818884478691847395837699072221005501800919219366542749884468691793630611950990529080847519607133539671195864198272777115792928784595536445936882119869059121395123801562924294690534627999441023179898426;
            5'd26: xpb[101] = 1024'd27766251953905815247267218829861027225956582076587733358628412551849309472526447092987294431353081170578379716833056789053941885741630363374547492958601107753850387778570860149857267300792996996830023036223216419117063939723543908320332550507220486240095848367744980213570669933095059438752109790924202211856;
            5'd27: xpb[101] = 1024'd47921368672767537587361946847134825618446977868108136045980559967686112965671177967335278250198611109361109614781634886260487933784188505743593184997982848964950891088449926669102583611056913146140438938906761642369929606669972023711880505477995035598071827676368565303339776941895428342876220140825224525286;
            5'd28: xpb[101] = 1024'd68076485391629259927456674864408624010937373659628538733332707383522916458815908841683262069044141048143839512730212983467033981826746648112638877037364590176051394398328993188347899921320829295450854841590306865622795273616400139103428460448769584956047806984992150393108883950695797247000330490726246838716;
            5'd29: xpb[101] = 1024'd88231602110490982267551402881682422403427769451148941420684854799359719951960639716031245887889670986926569410678791080673580029869304790481684569076746331387151897708208059707593216231584745444761270744273852088875660940562828254494976415419544134314023786293615735482877990959496166151124440840627269152146;
            5'd30: xpb[101] = 1024'd108386718829352704607646130898956220795918165242669344108037002215196523445105370590379229706735200925709299308627369177880126077911862932850730261116128072598252401018087126226838532541848661594071686646957397312128526607509256369886524370390318683671999765602239320572647097968296535055248551190528291465576;
            5'd31: xpb[101] = 1024'd4475139864089685548941931511415586443710133908454062667257294566056431600940962554712142310923056555048879799118453840507608285113200740664615828139178772875662229758394975408453609660595372022071904941253702689017031424234787712313093755677863783763155841496745847632309676903168270942253971713803719294675;
        endcase
    end

    always_comb begin
        case(flag[34][5:0])
            6'd0: xpb[102] = 1024'd0;
            6'd1: xpb[102] = 1024'd74348476133538074643917793466751908790449478412855074741370648523435065215697416169537598672213130401637379552262262686146609086998489608794410822597445777510226703818922629632664582581188246946346259226162243879317128970701056300334810140165933891193975862109743245376092655992948636431748385945165168046218;
            6'd2: xpb[102] = 1024'd24630256582951407889036659528689384836200529699974465354609441981893235094085693429060126129768586493831609697067031937714154333155758883033661520178560514086762733068274041927698925970859288171382320843937247912269897091181215827704641710648638333121131820805369432722078783911968639846378082063704741608105;
            6'd3: xpb[102] = 1024'd98978732716489482532954452995441293626650008112829540095980090505328300309783109598597724801981716895468989249329294623860763420154248491828072342776006291596989436887196671560363508552047535117728580070099491791587026061882272128039451850814572224315107682915112678098171439904917276278126468008869909654323;
            6'd4: xpb[102] = 1024'd49260513165902815778073319057378769672401059399948930709218883963786470188171386858120252259537172987663219394134063875428308666311517766067323040357121028173525466136548083855397851941718576342764641687874495824539794182362431655409283421297276666242263641610738865444157567823937279692756164127409483216210;
            6'd5: xpb[102] = 1024'd123608989299440890421991112524130678462850537812804005450589532487221535403868803027657850931750303389300598946396326561574917753310007374861733862954566805683752169955470713488062434522906823289110900914036739703856923153063487955744093561463210557436239503720482110820250223816885916124504550072574651262428;
            6'd6: xpb[102] = 1024'd73890769748854223667109978586068154508601589099923396063828325945679705282257080287180378389305759481494829091201095813142462999467276649100984560535681542260288199204822125783096777912577864514146962531811743736809691273543647483113925131945914999363395462416108298166236351735905919539134246191114224824315;
            6'd7: xpb[102] = 1024'd24172550198267556912228844648005630554352640387042786677067119404137875160645357546702905846861215573689059236005865064710008245624545923340235258116796278836824228454173538078131121302248905739183024149586747769762459394023807010483756702428619441290551421111734485512222479654925922953763942309653798386202;
            6'd8: xpb[102] = 1024'd98521026331805631556146638114757539344802118799897861418437767927572940376342773716240504519074345975326438788268127750856617332623035532134646080714242056347050932273096167710795703883437152685529283375748991649079588364724863310818566842594553332484527283221477730888315135647874559385512328254818966432420;
            6'd9: xpb[102] = 1024'd48802806781218964801265504176695015390553170087017252031676561386031110254731050975763031976629802067520668933072897002424162578780304806373896778295356792923586961522447580005830047273108193910565344993523995682032356485205022838188398413077257774411683241917103918234301263566894562800142024373358539994307;
            6'd10: xpb[102] = 1024'd123151282914757039445183297643446924181002648499872326773047209909466175470428467145300630648842932469158048485335159688570771665778794415168307600892802570433813665341370209638494629854296440856911604219686239561349485455906079138523208553243191665605659104026847163610393919559843199231890410318523708040525;
            6'd11: xpb[102] = 1024'd73433063364170372690302163705384400226753699786991717386286003367924345348816744404823158106398388561352278630139928940138316911936063689407558298473917307010349694590721621933528973243967482081947665837461243594302253576386238665893040123725896107532815062722473350956380047478863202646520106437063281602412;
            6'd12: xpb[102] = 1024'd23714843813583705935421029767321876272504751074111107999524796826382515227205021664345685563953844653546508774944698191705862158093332963646808996055032043586885723840073034228563316633638523306983727455236247627255021696866398193262871694208600549459971021418099538302366175397883206061149802555602855164299;
            6'd13: xpb[102] = 1024'd98063319947121780579338823234073785062954229486966182740895445349817580442902437833883284236166975055183888327206960877852471245091822572441219818652477821097112427658995663861227899214826770253329986681398491506572150667567454493597681834374534440653946883527842783678458831390831842492898188500768023210517;
            6'd14: xpb[102] = 1024'd48345100396535113824457689296011261108705280774085573354134238808275750321290715093405811693722431147378118472011730129420016491249091846680470516233592557673648456908347076156262242604497811478366048299173495539524918788047614020967513404857238882581102842223468971024444959309851845907527884619307596772404;
            6'd15: xpb[102] = 1024'd122693576530073188468375482762763169899154759186940648095504887331710815536988131262943410365935561549015498024273992815566625578247581455474881338831038335183875160727269705788926825185686058424712307525335739418842047758748670321302323545023172773775078704333212216400537615302800482339276270564472764818622;
            6'd16: xpb[102] = 1024'd72975356979486521713494348824700645944905810474060038708743680790168985415376408522465937823491017641209728169078762067134170824404850729714132036412153071760411189976621118083961168575357099649748369143110743451794815879228829848672155115505877215702234663028838403746523743221820485753905966683012338380509;
            6'd17: xpb[102] = 1024'd23257137428899854958613214886638121990656861761179429321982474248627155293764685781988465281046473733403958313883531318701716070562120003953382733993267808336947219225972530378995511965028140874784430760885747484747583999708989376041986685988581657629390621724464591092509871140840489168535662801551911942396;
            6'd18: xpb[102] = 1024'd97605613562437929602531008353390030781106340174034504063353122772062220509462101951526063953259604135041337866145794004848325157560609612747793556590713585847173923044895160011660094546216387821130689987047991364064712970410045676376796826154515548823366483834207836468602527133789125600284048746717079988614;
            6'd19: xpb[102] = 1024'd47887394011851262847649874415327506826857391461153894676591916230520390387850379211048591410815060227235568010950563256415870403717878886987044254171828322423709952294246572306694437935887429046166751604822995397017481090890205203746628396637219990750522442529834023814588655052809129014913744865256653550501;
            6'd20: xpb[102] = 1024'd122235870145389337491567667882079415617306869874008969417962564753955455603547795380586190083028190628872947563212825942562479490716368495781455076769274099933936656113169201939359020517075675992513010830985239276334610061591261504081438536803153881944498304639577269190681311045757765446662130810421821596719;
            6'd21: xpb[102] = 1024'd72517650594802670736686533944016891663057921161128360031201358212413625481936072640108717540583646721067177708017595194130024736873637770020705774350388836510472685362520614234393363906746717217549072448760243309287378182071421031451270107285858323871654263335203456536667438964777768861291826928961395158606;
            6'd22: xpb[102] = 1024'd22799431044216003981805400005954367708808972448247750644440151670871795360324349899631244998139102813261407852822364445697569983030907044259956471931503573087008714611872026529427707296417758442585134066535247342240146302551580558821101677768562765798810222030829643882653566883797772275921523047500968720493;
            6'd23: xpb[102] = 1024'd97147907177754078625723193472706276499258450861102825385810800194306860576021766069168843670352233214898787405084627131844179070029396653054367294528949350597235418430794656162092289877606005388931393292697491221557275273252636859155911817934496656992786084140572889258746222876746408707669908992666136766711;
            6'd24: xpb[102] = 1024'd47429687627167411870842059534643752545009502148222215999049593652765030454410043328691371127907689307093017549889396383411724316186665927293617992110064087173771447680146068457126633267277046613967454910472495254510043393732796386525743388417201098919942042836199076604732350795766412122299605111205710328598;
            6'd25: xpb[102] = 1024'd121778163760705486514759853001395661335458980561077290740420242176200095670107459498228969800120819708730397102151659069558333403185155536088028814707509864683998151499068698089791215848465293560313714136634739133827172364433852686860553528583134990113917904945942321980825006788715048554047991056370878374816;
            6'd26: xpb[102] = 1024'd72059944210118819759878719063333137381210031848196681353659035634658265548495736757751497257676275800924627246956428321125878649342424810327279512288624601260534180748420110384825559238136334785349775754409743166779940484914012214230385099065839432041073863641568509326811134707735051968677687174910451936703;
            6'd27: xpb[102] = 1024'd22341724659532153004997585125270613426961083135316071966897829093116435426884014017274024715231731893118857391761197572693423895499694084566530209869739337837070209997771522679859902627807376010385837372184747199732708605394171741600216669548543873968229822337194696672797262626755055383307383293450025498590;
            6'd28: xpb[102] = 1024'd96690200793070227648915378592022522217410561548171146708268477616551500642581430186811623387444862294756236944023460258840032982498183693360941032467185115347296913816694152312524485208995622956732096598346991079049837576095228041935026809714477765162205684446937942048889918619703691815055769238615193544808;
            6'd29: xpb[102] = 1024'd46971981242483560894034244653959998263161612835290537321507271075009670520969707446334150845000318386950467088828229510407578228655452967600191730048299851923832943066045564607558828598666664181768158216121995112002605696575387569304858380197182207089361643142564129394876046538723695229685465357154767106695;
            6'd30: xpb[102] = 1024'd121320457376021635537952038120711907053611091248145612062877919598444735736667123615871749517213448788587846641090492196554187315653942576394602552645745629434059646884968194240223411179854911128114417442284238991319734667276443869639668520363116098283337505252307374770968702531672331661433851302319935152913;
            6'd31: xpb[102] = 1024'd71602237825434968783070904182649383099362142535265002676116713056902905615055400875394276974768904880782076785895261448121732561811211850633853250226860366010595676134319606535257754569525952353150479060059243024272502787756603397009500090845820540210493463947933562116954830450692335076063547420859508714800;
            6'd32: xpb[102] = 1024'd21884018274848302028189770244586859145113193822384393289355506515361075493443678134916804432324360972976306930700030699689277807968481124873103947807975102587131705383671018830292097959196993578186540677834247057225270908236762924379331661328524982137649422643559749462940958369712338490693243539399082276687;
            6'd33: xpb[102] = 1024'd96232494408386376672107563711338767935562672235239468030726155038796140709141094304454403104537491374613686482962293385835886894966970733667514770405420880097358409202593648462956680540385240524532799903996490936542399878937819224714141801494458873331625284753302994839033614362660974922441629484564250322905;
            6'd34: xpb[102] = 1024'd46514274857799709917226429773276243981313723522358858643964948497254310587529371563976930562092947466807916627767062637403432141124240007906765467986535616673894438451945060757991023930056281749568861521771494969495167999417978752083973371977163315258781243448929182185019742281680978337071325603103823884792;
            6'd35: xpb[102] = 1024'd120862750991337784561144223240028152771763201935213933385335597020689375803226787733514529234306077868445296180029325323550041228122729616701176290583981394184121142270867690390655606511244528695915120747933738848812296970119035052418783512143097206452757105558672427561112398274629614768819711548268991931010;
            6'd36: xpb[102] = 1024'd71144531440751117806263089301965628817514253222333323998574390479147545681615064993037056691861533960639526324834094575117586474279998890940426988165096130760657171520219102685689949900915569920951182365708742881765065090599194579788615082625801648379913064254298614907098526193649618183449407666808565492897;
            6'd37: xpb[102] = 1024'd21426311890164451051381955363903104863265304509452714611813183937605715560003342252559584149416990052833756469638863826685131720437268165179677685746210867337193200769570514980724293290586611145987243983483746914717833211079354107158446653108506090307069022949924802253084654112669621598079103785348139054784;
            6'd38: xpb[102] = 1024'd95774788023702525695299748830655013653714782922307789353183832461040780775700758422097182821630120454471136021901126512831740807435757773974088508343656644847419904588493144613388875871774858092333503209645990794034962181780410407493256793274439981501044885059668047629177310105618258029827489730513307101002;
            6'd39: xpb[102] = 1024'd46056568473115858940418614892592489699465834209427179966422625919498950654089035681619710279185576546665366166705895764399286053593027048213339205924771381423955933837844556908423219261445899317369564827420994826987730302260569934863088363757144423428200843755294234975163438024638261444457185849052880662889;
            6'd40: xpb[102] = 1024'd120405044606653933584336408359344398489915312622282254707793274442934015869786451851157308951398706948302745718968158450545895140591516657007750028522217158934182637656767186541087801842634146263715824053583238706304859272961626235197898503923078314622176705865037480351256094017586897876205571794218048709107;
            6'd41: xpb[102] = 1024'd70686825056067266829455274421281874535666363909401645321032067901392185748174729110679836408954163040496975863772927702113440386748785931247000726103331895510718666906118598836122145232305187488751885671358242739257627393441785762567730074405782756549332664560663667697242221936606901290835267912757622270994;
            6'd42: xpb[102] = 1024'd20968605505480600074574140483219350581417415196521035934270861359850355626563006370202363866509619132691206008577696953680985632906055205486251423684446632087254696155470011131156488621976228713787947289133246772210395513921945289937561644888487198476488623256289855043228349855626904705464964031297195832881;
            6'd43: xpb[102] = 1024'd95317081639018674718491933949971259371866893609376110675641509883285420842260422539739962538722749534328585560839959639827594719904544814280662246281892409597481399974392640763821071203164475660134206515295490651527524484623001590272371785054421089670464485366033100419321005848575541137213349976462363879099;
            6'd44: xpb[102] = 1024'd45598862088432007963610800011908735417617944896495501288880303341743590720648699799262489996278205626522815705644728891395139966061814088519912943863007146174017429223744053058855414592835516885170268133070494684480292605103161117642203355537125531597620444061659287765307133767595544551843046095001937440986;
            6'd45: xpb[102] = 1024'd119947338221970082607528593478660644208067423309350576030250951865178655936346115968800088668491336028160195257906991577541749053060303697314323766460452923684244133042666682691519997174023763831516527359232738563797421575804217417977013495703059422791596306171402533141399789760544180983591432040167105487204;
            6'd46: xpb[102] = 1024'd70229118671383415852647459540598120253818474596469966643489745323636825814734393228322616126046792120354425402711760829109294299217572971553574464041567660260780162292018094986554340563694805056552588977007742596750189696284376945346845066185763864718752264867028720487385917679564184398221128158706679049091;
            6'd47: xpb[102] = 1024'd20510899120796749097766325602535596299569525883589357256728538782094995693122670487845143583602248212548655547516530080676839545374842245792825161622682396837316191541369507281588683953365846281588650594782746629702957816764536472716676636668468306645908223562654907833372045598584187812850824277246252610978;
            6'd48: xpb[102] = 1024'd94859375254334823741684119069287505090019004296444431998099187305530060908820086657382742255815378614186035099778792766823448632373331854587235984220128174347542895360292136914253266534554093227934909820944990509020086787465592773051486776834402197839884085672398153209464701591532824244599210222411420657196;
            6'd49: xpb[102] = 1024'd45141155703748156986802985131224981135770055583563822611337980763988230787208363916905269713370834706380265244583562018390993878530601128826486681801242910924078924609643549209287609924225134452970971438719994541972854907945752300421318347317106639767040044368024340555450829510552827659228906340950994219083;
            6'd50: xpb[102] = 1024'd119489631837286231630720778597976889926219533996418897352708629287423296002905780086442868385583965108017644796845824704537602965529090737620897504398688688434305628428566178841952192505413381399317230664882238421289983878646808600756128487483040530961015906477767585931543485503501464090977292286116162265301;
            6'd51: xpb[102] = 1024'd69771412286699564875839644659914365971970585283538287965947422745881465881294057345965395843139421200211874941650593956105148211686360011860148201979803425010841657677917591136986535895084422624353292282657242454242751999126968128125960057965744972888171865173393773277529613422521467505606988404655735827188;
            6'd52: xpb[102] = 1024'd20053192736112898120958510721851842017721636570657678579186216204339635759682334605487923300694877292406105086455363207672693457843629286099398899560918161587377686927269003432020879284755463849389353900432246487195520119607127655495791628448449414815327823869019960623515741341541470920236684523195309389075;
            6'd53: xpb[102] = 1024'd94401668869650972764876304188603750808171114983512753320556864727774700975379750775025521972908007694043484638717625893819302544842118894893809722158363939097604390746191633064685461865943710795735613126594490366512649090308183955830601768614383306009303685978763205999608397334490107351985070468360477435293;
            6'd54: xpb[102] = 1024'd44683449319064306009995170250541226853922166270632143933795658186232870853768028034548049430463463786237714783522395145386847790999388169133060419739478675674140419995543045359719805255614752020771674744369494399465417210788343483200433339097087747936459644674389393345594525253510110766614766586900050997180;
            6'd55: xpb[102] = 1024'd119031925452602380653912963717293135644371644683487218675166306709667936069465444204085648102676594187875094335784657831533456877997877777927471242336924453184367123814465674992384387836802998967117933970531738278782546181489399783535243479263021639130435506784132638721687181246458747198363152532065219043398;
            6'd56: xpb[102] = 1024'd69313705902015713899031829779230611690122695970606609288405100168126105947853721463608175560232050280069324480589427083101002124155147052166721939918039189760903153063817087287418731226474040192153995588306742311735314301969559310905075049745726081057591465479758826067673309165478750612992848650604792605285;
            6'd57: xpb[102] = 1024'd19595486351429047144150695841168087735873747257725999901643893626584275826241998723130703017787506372263554625394196334668547370312416326405972637499153926337439182313168499582453074616145081417190057206081746344688082422449718838274906620228430522984747424175385013413659437084498754027622544769144366167172;
            6'd58: xpb[102] = 1024'd93943962484967121788068489307919996526323225670581074643014542150019341041939414892668301690000636773900934177656459020815156457310905935200383460096599703847665886132091129215117657197333328363536316432243990224005211393150775138609716760394364414178723286285128258789752093077447390459370930714309534213390;
            6'd59: xpb[102] = 1024'd44225742934380455033187355369857472572074276957700465256253335608477510920327692152190829147556092866095164322461228272382701703468175209439634157677714440424201915381442541510152000587004369588572378050018994256957979513630934665979548330877068856105879244980754446135738220996467393874000626832849107775277;
            6'd60: xpb[102] = 1024'd118574219067918529677105148836609381362523755370555539997623984131912576136025108321728427819769223267732543874723490958529310790466664818234044980275160217934428619200365171142816583168192616534918637276181238136275108484331990966314358471043002747299855107090497691511830876989416030305749012778014275821495;
            6'd61: xpb[102] = 1024'd68855999517331862922224014898546857408274806657674930610862777590370746014413385581250955277324679359926774019528260210096856036623934092473295677856274954510964648449716583437850926557863657759954698893956242169227876604812150493684190041525707189227011065786123878857817004908436033720378708896553849383382;
            6'd62: xpb[102] = 1024'd19137779966745196167342880960484333454025857944794321224101571048828915892801662840773482734880135452121004164333029461664401282781203366712546375437389691087500677699067995732885269947534698984990760511731246202180644725292310021054021612008411631154167024481750066203803132827456037135008405015093422945269;
            6'd63: xpb[102] = 1024'd93486256100283270811260674427236242244475336357649395965472219572263981108499079010311081407093265853758383716595292147811010369779692975506957198034835468597727381517990625365549852528722945931337019737893490081497773695993366321388831752174345522348142886591493311579895788820404673566756790960258590991487;
        endcase
    end

    always_comb begin
        case(flag[34][11:6])
            6'd0: xpb[103] = 1024'd0;
            6'd1: xpb[103] = 1024'd43768036549696604056379540489173718290226387644768786578711013030722150986887356269833608864648721945952613861400061399378555615936962249746207895615950205174263410767342037660584195918393987156373081355668494114450541816473525848758663322657049964275298845287119498925881916739424676981386487078798164553374;
            6'd2: xpb[103] = 1024'd87536073099393208112759080978347436580452775289537573157422026061444301973774712539667217729297443891905227722800122798757111231873924499492415791231900410348526821534684075321168391836787974312746162711336988228901083632947051697517326645314099928550597690574238997851763833478849353962772974157596329106748;
            6'd3: xpb[103] = 1024'd7237413964965070770339694062706722125980735808570675608001184027189557623352929899485755379288491528414692176742690763556603006969666414683463561831519574589099557732454895644122348563664755747809046458618242496987264599199680773311011398287920443559076632447241438747539222144345397927040771409768899175791;
            6'd4: xpb[103] = 1024'd51005450514661674826719234551880440416207123453339462186712197057911708610240286169319364243937213474367306038142752162935158622906628664429671457447469779763362968499796933304706544482058742904182127814286736611437806415673206622069674720944970407834375477734360937673421138883770074908427258488567063729165;
            6'd5: xpb[103] = 1024'd94773487064358278883098775041054158706433511098108248765423210088633859597127642439152973108585935420319919899542813562313714238843590914175879353063419984937626379267138970965290740400452730060555209169955230725888348232146732470828338043602020372109674323021480436599303055623194751889813745567365228282539;
            6'd6: xpb[103] = 1024'd14474827929930141540679388125413444251961471617141351216002368054379115246705859798971510758576983056829384353485381527113206013939332829366927123663039149178199115464909791288244697127329511495618092917236484993974529198399361546622022796575840887118153264894482877495078444288690795854081542819537798351582;
            6'd7: xpb[103] = 1024'd58242864479626745597058928614587162542187859261910137794713381085101266233593216068805119623225705002781998214885442926491761629876295079113135019278989354352462526232251828948828893045723498651991174272904979108425071014872887395380686119232890851393452110181602376420960361028115472835468029898335962904956;
            6'd8: xpb[103] = 1024'd102010901029323349653438469103760880832414246906678924373424394115823417220480572338638728487874426948734612076285504325870317245813257328859342914894939559526725936999593866609413088964117485808364255628573473222875612831346413244139349441889940815668750955468721875346842277767540149816854516977134127458330;
            6'd9: xpb[103] = 1024'd21712241894895212311019082188120166377942207425712026824003552081568672870058789698457266137865474585244076530228072290669809020908999244050390685494558723767298673197364686932367045690994267243427139375854727490961793797599042319933034194863761330677229897341724316242617666433036193781122314229306697527373;
            6'd10: xpb[103] = 1024'd65480278444591816367398622677293884668168595070480813402714565112290823856946145968290875002514196531196690391628133690048364636845961493796598581110508928941562083964706724592951241609388254399800220731523221605412335614072568168691697517520811294952528742628843815168499583172460870762508801308104862080747;
            6'd11: xpb[103] = 1024'd109248314994288420423778163166467602958394982715249599981425578143012974843833502238124483867162918477149304253028195089426920252782923743542806476726459134115825494732048762253535437527782241556173302087191715719862877430546094017450360840177861259227827587915963314094381499911885547743895288386903026634121;
            6'd12: xpb[103] = 1024'd28949655859860283081358776250826888503922943234282702432004736108758230493411719597943021517153966113658768706970763054226412027878665658733854247326078298356398230929819582576489394254659022991236185834472969987949058396798723093244045593151681774236306529788965754990156888577381591708163085639075596703164;
            6'd13: xpb[103] = 1024'd72717692409556887137738316740000606794149330879051489010715749139480381480299075867776630381802688059611382568370824453604967643815627908480062142942028503530661641697161620237073590173053010147609267190141464102399600213272248942002708915808731738511605375076085253916038805316806268689549572717873761256538;
            6'd14: xpb[103] = 1024'd116485728959253491194117857229174325084375718523820275589426762170202532467186432137610239246451410005563996429770885852983523259752590158226270038557978708704925052464503657897657786091446997303982348545809958216850142029745774790761372238465781702786904220363204752841920722056230945670936059796671925809912;
            6'd15: xpb[103] = 1024'd36187069824825353851698470313533610629903679042853378040005920135947788116764649497428776896442457642073460883713453817783015034848332073417317809157597872945497788662274478220611742818323778739045232293091212484936322995998403866555056991439602217795383162236207193737696110721726989635203857048844495878955;
            6'd16: xpb[103] = 1024'd79955106374521957908078010802707328920130066687622164618716933166669939103652005767262385761091179588026074745113515217161570650785294323163525704773548078119761199429616515881195938736717765895418313648759706599386864812471929715313720314096652182070682007523326692663578027461151666616590344127642660432329;
            6'd17: xpb[103] = 1024'd123723142924218561964457551291881047210356454332390951197427946197392090090539362037095994625739901533978688606513576616540126266722256572909733600389498283294024610196958553541780134655111753051791395004428200713837406628945455564072383636753702146345980852810446191589459944200576343597976831206440824985703;
            6'd18: xpb[103] = 1024'd43424483789790424622038164376240332755884414851424053648007104163137345740117579396914532275730949170488153060456144581339618041817998488100781370989117447534597346394729373864734091381988534486854278751709454981923587595198084639866068389727522661354459794683448632485235332866072387562244628458613395054746;
            6'd19: xpb[103] = 1024'd87192520339487028678417704865414051046110802496192840226718117193859496727004935666748141140379671116440766921856205980718173657754960737846989266605067652708860757162071411525318287300382521643227360107377949096374129411671610488624731712384572625629758639970568131411117249605497064543631115537411559608120;
            6'd20: xpb[103] = 1024'd6893861205058891335998317949773336591638763015225942677297275159604752376583153026566678790370718752950231375798773945517665432850702653038037037204686816949433493359842231848272244027259303078290243854659203364460310377924239564418416465358393140638237581843570572306892638270993108507898912789584129677163;
            6'd21: xpb[103] = 1024'd50661897754755495392377858438947054881865150659994729256008288190326903363470509296400287655019440698902845237198835344896221048787664902784244932820637022123696904127184269508856439945653290234663325210327697478910852194397765413177079788015443104913536427130690071232774555010417785489285399868382294230537;
            6'd22: xpb[103] = 1024'd94429934304452099448757398928120773172091538304763515834719301221049054350357865566233896519668162644855459098598896744274776664724627152530452828436587227297960314894526307169440635864047277391036406565996191593361394010871291261935743110672493069188835272417809570158656471749842462470671886947180458783911;
            6'd23: xpb[103] = 1024'd14131275170023962106338012012480058717619498823796618285298459186794309999936082926052434169659210281364923552541464709074268439820369067721500599036206391538533051092297127492394592590924058826099290313277445861447574977123920337729427863646313584197314214290812011054431860415338506434939684199353028852954;
            6'd24: xpb[103] = 1024'd57899311719720566162717552501653777007845886468565404864009472217516460986823439195886043034307932227317537413941526108452824055757331317467708494652156596712796461859639165152978788509318045982472371668945939975898116793597446186488091186303363548472613059577931509980313777154763183416326171278151193406328;
            6'd25: xpb[103] = 1024'd101667348269417170219097092990827495298072274113334191442720485248238611973710795465719651898956654173270151275341587507831379671694293567213916390268106801887059872626981202813562984427712033138845453024614434090348658610070972035246754508960413512747911904865051008906195693894187860397712658356949357959702;
            6'd26: xpb[103] = 1024'd21368689134989032876677706075186780843600234632367293893299643213983867623289012825538189548947701809779615729284155472630871446790035482404964160867725966127632608824752023136516941154588814573908336771895688358434839576323601111040439261934234027756390846738053449801971082559683904361980455609121928028745;
            6'd27: xpb[103] = 1024'd65136725684685636933057246564360499133826622277136080472010656244706018610176369095371798413596423755732229590684216872009427062726997732151172056483676171301896019592094060797101137072982801730281418127564182472885381392797126959799102584591283992031689692025172948727852999299108581343366942687920092582119;
            6'd28: xpb[103] = 1024'd108904762234382240989436787053534217424053009921904867050721669275428169597063725365205407278245145701684843452084278271387982678663959981897379952099626376476159430359436098457685332991376788886654499483232676587335923209270652808557765907248333956306988537312292447653734916038533258324753429766718257135493;
            6'd29: xpb[103] = 1024'd28606103099954103647017400137893502969580970440937969501300827241173425246641942725023944928236193338194307906026846236187474453759701897088427722699245540716732166557206918780639289718253570321717383230513930855422104175523281884351450660222154471315467479185294888549510304704029302289021227018890827204536;
            6'd30: xpb[103] = 1024'd72374139649650707703396940627067221259807358085706756080011840271895576233529298994857553792884915284146921767426907635566030069696664146834635618315195745890995577324548956441223485636647557478090464586182424969872645991996807733110113982879204435590766324472414387475392221443453979270407714097688991757910;
            6'd31: xpb[103] = 1024'd116142176199347311759776481116240939550033745730475542658722853302617727220416655264691162657533637230099535628826969034944585685633626396580843513931145951065258988091890994101807681555041544634463545941850919084323187808470333581868777305536254399866065169759533886401274138182878656251794201176487156311284;
            6'd32: xpb[103] = 1024'd35843517064919174417357094200600225095561706249508645109302011268362982869994872624509700307524684866609000082769536999744077460729368311771891284530765115305831724289661814424761638281918326069526429689132173352409368774722962657662462058510074914874544111632536327297049526848374700216061998428659726380327;
            6'd33: xpb[103] = 1024'd79611553614615778473736634689773943385788093894277431688013024299085133856882228894343309172173406812561613944169598399122633076666330561518099180146715320480095135057003852085345834200312313225899511044800667466859910591196488506421125381167124879149842956919655826222931443587799377197448485507457890933701;
            6'd34: xpb[103] = 1024'd123379590164312382530116175178947661676014481539046218266724037329807284843769585164176918036822128758514227805569659798501188692603292811264307075762665525654358545824345889745930030118706300382272592400469161581310452407670014355179788703824174843425141802206775325148813360327224054178834972586256055487075;
            6'd35: xpb[103] = 1024'd43080931029884245187696788263306947221542442058079320717303195295552540493347802523995455686813176395023692259512227763300680467699034726455354846362284689894931282022116710068883986845583081817335476147750415849396633373922643430973473456797995358433620744079777766044588748992720098143102769838428625556118;
            6'd36: xpb[103] = 1024'd86848967579580849244076328752480665511768829702848107296014208326274691480235158793829064551461898340976306120912289162679236083635996976201562741978234895069194692789458747729468182763977068973708557503418909963847175190396169279732136779455045322708919589366897264970470665732144775124489256917226790109492;
            6'd37: xpb[103] = 1024'd6550308445152711901656941836839951057296790221881209746593366292019947129813376153647602201452945977485770574854857127478727858731738891392610512577854059309767428987229568052422139490853850408771441250700164231933356156648798355525821532428865837717398531239899705866246054397640819088757054169399360178535;
            6'd38: xpb[103] = 1024'd50318344994849315958036482326013669347523177866649996325304379322742098116700732423481211066101667923438384436254918526857283474668701141138818408193804264484030839754571605713006335409247837565144522606368658346383897973122324204284484855085915801992697376527019204792127971137065496070143541248197524731909;
            6'd39: xpb[103] = 1024'd94086381544545920014416022815187387637749565511418782904015392353464249103588088693314819930750389869390998297654979926235839090605663390885026303809754469658294250521913643373590531327641824721517603962037152460834439789595850053043148177742965766267996221814138703718009887876490173051530028326995689285283;
            6'd40: xpb[103] = 1024'd13787722410117782671996635899546673183277526030451885354594550319209504753166306053133357580741437505900462751597547891035330865701405306076074074409373633898866986719684463696544488054518606156580487709318406728920620755848479128836832930716786281276475163687141144613785276541986217015797825579168259354326;
            6'd41: xpb[103] = 1024'd57555758959814386728376176388720391473503913675220671933305563349931655740053662322966966445390159451853076612997609290413886481638367555822281970025323839073130397487026501357128683972912593312953569064986900843371162572322004977595496253373836245551774008974260643539667193281410893997184312657966423907700;
            6'd42: xpb[103] = 1024'd101323795509510990784755716877894109763730301319989458512016576380653806726941018592800575310038881397805690474397670689792442097575329805568489865641274044247393808254368539017712879891306580469326650420655394957821704388795530826354159576030886209827072854261380142465549110020835570978570799736764588461074;
            6'd43: xpb[103] = 1024'd21025136375082853442336329962253395309258261839022560962595734346399062376519235952619112960029929034315154928340238654591933872671071720759537636240893208487966544452139359340666836618183361904389534167936649225907885355048159902147844329004706724835551796134382583361324498686331614942838596988937158530117;
            6'd44: xpb[103] = 1024'd64793172924779457498715870451427113599484649483791347541306747377121213363406592222452721824678650980267768789740300053970489488608033970505745531856843413662229955219481397001251032536577349060762615523605143340358427171521685750906507651661756689110850641421502082287206415425756291924225084067735323083491;
            6'd45: xpb[103] = 1024'd108561209474476061555095410940600831889711037128560134120017760407843364350293948492286330689327372926220382651140361453349045104544996220251953427472793618836493365986823434661835228454971336217135696879273637454808968987995211599665170974318806653386149486708621581213088332165180968905611571146533487636865;
            6'd46: xpb[103] = 1024'd28262550340047924212676024024960117435238997647593236570596918373588619999872165852104868339318420562729847105082929418148536879640738135443001198072412783077066102184594254984789185181848117652198580626554891722895149954247840675458855727292627168394628428581624022108863720830677012869879368398706057705908;
            6'd47: xpb[103] = 1024'd72030586889744528269055564514133835725465385292362023149307931404310770986759522121938477203967142508682460966482990817527092495577700385189209093688362988251329512951936292645373381100242104808571661982223385837345691770721366524217519049949677132669927273868743521034745637570101689851265855477504222259282;
            6'd48: xpb[103] = 1024'd115798623439441132325435105003307554015691772937130809728018944435032921973646878391772086068615864454635074827883052216905648111514662634935416989304313193425592923719278330305957577018636091964944743337891879951796233587194892372976182372606727096945226119155863019960627554309526366832652342556302386812656;
            6'd49: xpb[103] = 1024'd35499964305012994983015718087666839561219733456163912178598102400778177623225095751590623718606912091144539281825620181705139886610404550126464759903932357666165659917049150628911533745512873400007627085173134219882414553447521448769867125580547611953705061028865460856402942975022410796920139808474956881699;
            6'd50: xpb[103] = 1024'd79268000854709599039395258576840557851446121100932698757309115431500328610112452021424232583255634037097153143225681581083695502547366799872672655519882562840429070684391188289495729663906860556380708440841628334332956369921047297528530448237597576229003906315984959782284859714447087778306626887273121435073;
            6'd51: xpb[103] = 1024'd123036037404406203095774799066014276141672508745701485336020128462222479596999808291257841447904355983049767004625742980462251118484329049618880551135832768014692481451733225950079925582300847712753789796510122448783498186394573146287193770894647540504302751603104458708166776453871764759693113966071285988447;
            6'd52: xpb[103] = 1024'd42737378269978065753355412150373561687200469264734587786599286427967735246578025651076379097895403619559231458568310945261742893580070964809928321735451932255265217649504046273033882309177629147816673543791376716869679152647202222080878523868468055512781693476106899603942165119367808723960911218243856057490;
            6'd53: xpb[103] = 1024'd86505414819674669809734952639547279977426856909503374365310299458689886233465381920909987962544125565511845319968372344640298509517033214556136217351402137429528628416846083933618078227571616304189754899459870831320220969120728070839541846525518019788080538763226398529824081858792485705347398297042020610864;
            6'd54: xpb[103] = 1024'd6206755685246532467315565723906565522954817428536476815889457424435141883043599280728525612535173202021309773910940309439790284612775129747183987951021301670101364614616904256572034954448397739252638646741125099406401935373357146633226599499338534796559480636228839425599470524288529669615195549214590679907;
            6'd55: xpb[103] = 1024'd49974792234943136523695106213080283813181205073305263394600470455157292869930955550562134477183895147973923635311001708818345900549737379493391883566971506844364775381958941917156230872842384895625720002409619213856943751846882995391889922156388499071858325923348338351481387263713206651001682628012755233281;
            6'd56: xpb[103] = 1024'd93742828784639740580074646702254002103407592718074049973311483485879443856818311820395743341832617093926537496711063108196901516486699629239599779182921712018628186149300979577740426791236372051998801358078113328307485568320408844150553244813438463347157171210467837277363304003137883632388169706810919786655;
            6'd57: xpb[103] = 1024'd13444169650211603237655259786613287648935553237107152423890641451624699506396529180214280991823664730436001950653631072996393291582441544430647549782540876259200922347071799900694383518113153487061685105359367596393666534573037919944237997787258978355636113083470278173138692668633927596655966958983489855698;
            6'd58: xpb[103] = 1024'd57212206199908207294034800275787005939161940881875939002601654482346850493283885450047889856472386676388615812053692472374948907519403794176855445398491081433464333114413837561278579436507140643434766461027861710844208351046563768702901320444308942630934958370589777099020609408058604578042454037781654409072;
            6'd59: xpb[103] = 1024'd100980242749604811350414340764960724229388328526644725581312667513069001480171241719881498721121108622341229673453753871753504523456366043923063341014441286607727743881755875221862775354901127799807847816696355825294750167520089617461564643101358906906233803657709276024902526147483281559428941116579818962446;
            6'd60: xpb[103] = 1024'd20681583615176674007994953849320009774916289045677828031891825478814257129749459079700036371112156258850694127396321836552996298552107959114111111614060450848300480079526695544816732081777909234870731563977610093380931133772718693255249396075179421914712745530711716920677914812979325523696738368752389031489;
            6'd61: xpb[103] = 1024'd64449620164873278064374494338493728065142676690446614610602838509536408116636815349533645235760878204803307988796383235931551914489070208860319007230010656022563890846868733205400928000171896391243812919646104207831472950246244542013912718732229386190011590817831215846559831552404002505083225447550553584863;
            6'd62: xpb[103] = 1024'd108217656714569882120754034827667446355369064335215401189313851540258559103524171619367254100409600150755921850196444635310107530426032458606526902845960861196827301614210770865985123918565883547616894275314598322282014766719770390772576041389279350465310436104950714772441748291828679486469712526348718138237;
            6'd63: xpb[103] = 1024'd27918997580141744778334647912026731900897024854248503639893009506003814753102388979185791750400647787265386304139012600109599305521774373797574673445580025437400037811981591188939080645442664982679778022595852590368195732972399466566260794363099865473789377977953155668217136957324723450737509778521288207280;
        endcase
    end

    always_comb begin
        case(flag[34][16:12])
            5'd0: xpb[104] = 1024'd0;
            5'd1: xpb[104] = 1024'd71687034129838348834714188401200450191123412499017290218604022536725965739989745249019400615049369733218000165539073999488154921458736623543782569061530230611663448579323628849523276563836652139052859378264346704818737549445925315324924117020149829749088223265072654594099053696749400432123996857319452760654;
            5'd2: xpb[104] = 1024'd19307372575551956270629449397586467637548397872298896309076190008475036142670351588023730015441065156992850923620654564397246002076252912532405013106729420289636222589076040361416313936156098556795521148141453563273114248670953857684869664357070210231356543116028251158091579319570167847129303888013311036977;
            5'd3: xpb[104] = 1024'd90994406705390305105343637798786917828671810371316186527680212545201001882660096837043130630490434890210851089159728563885400923534989536076187582168259650901299671168399669210939590499992750695848380526405800268091851798116879173009793781377220039980444766381100905752190633016319568279253300745332763797631;
            5'd4: xpb[104] = 1024'd38614745151103912541258898795172935275096795744597792618152380016950072285340703176047460030882130313985701847241309128794492004152505825064810026213458840579272445178152080722832627872312197113591042296282907126546228497341907715369739328714140420462713086232056502316183158639140335694258607776026622073954;
            5'd5: xpb[104] = 1024'd110301779280942261375973087196373385466220208243615082836756402553676038025330448425066860645931500047203702012780383128282646925611242448608592595274989071190935893757475709572355904436148849252643901674547253831364966046787833030694663445734290250211801309497129156910282212335889736126382604633346074834608;
            5'd6: xpb[104] = 1024'd57922117726655868811888348192759402912645193616896688927228570025425108428011054764071190046323195470978552770861963693191738006228758737597215039320188260868908667767228121084248941808468295670386563444424360689819342746012861573054608993071210630694069629348084753474274737958710503541387911664039933110931;
            5'd7: xpb[104] = 1024'd5542456172369476247803609189145420359070178990178295017700737497174178830691661103075519446714890894753403528943544258100829086846275026585837483365387450546881441776980532596141979180787742088129225214301467548273719445237890115414554540408131011176337949199040350038267263581531270956393218694733791387254;
            5'd8: xpb[104] = 1024'd77229490302207825082517797590345870550193591489195585236304760033900144570681406352094920061764260627971403694482618257588984008305011650129620052426917681158544890356304161445665255744624394227182084592565814253092456994683815430739478657428280840925426172464113004632366317278280671388517215552053244147908;
            5'd9: xpb[104] = 1024'd24849828747921432518433058586731887996618576862477191326776927505649214973362012691099249462155956051746254452564198822498075088922527939118242496472116870836517664366056572957558293116943840644924746362442921111546833693908843973099424204765201221407694492315068601196358842901101438803522522582747102424231;
            5'd10: xpb[104] = 1024'd96536862877759781353147246987932338187741989361494481545380950042375180713351757940118650077205325784964254618103272821986230010381264562662025065533647101448181112945380201807081569680780492783977605740707267816365571243354769288424348321785351051156782715580141255790457896597850839235646519440066555184885;
            5'd11: xpb[104] = 1024'd44157201323473388789062507984318355634166974734776087635853117514124251116032364279122979477597021208739105376184853386895321090998780851650647509578846291126153886955132613318974607053099939201720267510584374674819947942579797830784293869122271431639051035431096852354450422220671606650651826470760413461208;
            5'd12: xpb[104] = 1024'd115844235453311737623776696385518805825290387233793377854457140050850216856022109528142380092646390941957105541723927386383476012457517475194430078640376521737817335534456242168497883616936591340773126888848721379638685492025723146109217986142421261388139258696169506948549475917421007082775823328079866221862;
            5'd13: xpb[104] = 1024'd63464573899025345059691957381904823271715372607074983944929307522599287258702715867146709493038086365731956299805507951292567093075033764183052522685575711415790109544208653680390920989256037758515788658725828238093062191250751688469163533479341641870407578547125103512542001540241774497781130358773724498185;
            5'd14: xpb[104] = 1024'd11084912344738952495607218378290840718140357980356590035401474994348357661383322206151038893429781789506807057887088516201658173692550053171674966730774901093762883553961065192283958361575484176258450428602935096547438890475780230829109080816262022352675898398080700076534527163062541912786437389467582774508;
            5'd15: xpb[104] = 1024'd82771946474577301330321406779491290909263770479373880254005497531074323401373067455170439508479151522724807223426162515689813095151286676715457535792305131705426332133284694041807234925412136315311309806867281801366176439921705546154033197836411852101764121663153354670633580859811942344910434246787035535162;
            5'd16: xpb[104] = 1024'd30392284920290908766236667775877308355688755852655486344477665002823393804053673794174768908870846946499657981507743080598904175768802965704079979837504321383399106143037105553700272297731582733053971576744388659820553139146734088513978745173332232584032441514108951234626106482632709759915741277480893811485;
            5'd17: xpb[104] = 1024'd102079319050129257600950856177077758546812168351672776563081687539549359544043419043194169523920216679717658147046817080087059097227539589247862548899034551995062554722360734403223548861568234872106830955008735364639290688592659403838902862193482062333120664779181605828725160179382110192039738134800346572139;
            5'd18: xpb[104] = 1024'd49699657495842865036866117173463775993237153724954382653553855011298429946724025382198498924311912103492508905128397644996150177845055878236484992944233741673035328732113145915116586233887681289849492724885842223093667387817687946198848409530402442815388984630137202392717685802202877607045045165494204848462;
            5'd19: xpb[104] = 1024'd121386691625681213871580305574664226184360566223971672872157877548024395686713770631217899539361281836710509070667471644484305099303792501780267562005763972284698777311436774764639862797724333428902352103150188927912404937263613261523772526550552272564477207895209856986816739498952278039169042022813657609116;
            5'd20: xpb[104] = 1024'd69007030071394821307495566571050243630785551597253278962630045019773466089394376970222228939752977260485359828749052209393396179921308790768890006050963161962671551321189186276532900170043779846645013873027295786366781636488641803883718073887472653046745527746165453550809265121773045454174349053507515885439;
            5'd21: xpb[104] = 1024'd16627368517108428743410827567436261077210536970534885053102212491522536492074983309226558340144672684260210586830632774302487260538825079757512450096162351640644325330941597788425937542363226264387675642904402644821158335713670346243663621224393033529013847597121050114801790744593812869179656084201374161762;
            5'd22: xpb[104] = 1024'd88314402646946777578125015968636711268333949469552175271706235028248502232064728558245958955194042417478210752369706773790642181997561703301295019157692582252307773910265226637949214106199878403440535021168749349639895885159595661568587738244542863278102070862193704708900844441343213301303652941520826922416;
            5'd23: xpb[104] = 1024'd35934741092660385014040276965022728714758934842833781362178402499997572634745334897250288355585737841253061510451287338699733262615077992289917463202891771930280547920017638149842251478519324821183196791045856208094272584384624203928533285581463243760370390713149301272893370064163980716308959972214685198739;
            5'd24: xpb[104] = 1024'd107621775222498733848754465366223178905882347341851071580782425036723538374735080146269688970635107574471061675990361338187888184073814615833700032264422002541943996499341266999365528042355976960236056169310202912913010133830549519253457402601613073509458613978221955866992423760913381148432956829534137959393;
            5'd25: xpb[104] = 1024'd55242113668212341284669726362609196352307332715132677671254592508472608777415686485274018371026802998245912434071941903096979264691330904822322476309621192219916770509093678511258565414675423377978717939187309771367386833055578061613402949938533453991726933829177552430984949383734148563438263860227996235716;
            5'd26: xpb[104] = 1024'd2862452113925948720584987358995213798732318088414283761726759980221679180096292824278347771418498422020763192153522468006070345308847193810944920354820381897889544518846090023151602786994869795721379709064416629821763532280606603973348497275453834473995253680133148994977475006554915978443570890921854512039;
            5'd27: xpb[104] = 1024'd74549486243764297555299175760195663989855730587431573980330782516947644920086038073297748386467868155238763357692596467494225266767583817354727489416350612509552993098169718872674879350831521934774239087328763334640501081726531919298272614295603664223083476945205803589076528703304316410567567748241307272693;
            5'd28: xpb[104] = 1024'd22169824689477904991214436756581681436280715960713180070802949988696715322766644412302077786859563579013614115774177032403316347385100106343349933461549802187525767107922130384567916723150968352516900857205870193094877780951560461658218161632524044705351796796161400153069054326125083825572874778935165549016;
            5'd29: xpb[104] = 1024'd93856858819316253825928625157782131627404128459730470289406972525422681062756389661321478401908933312231614281313251031891471268843836729887132502523080032799189215687245759234091193286987620491569760235470216897913615330397485776983142278652673874454440020061234054747168108022874484257696871636254618309670;
            5'd30: xpb[104] = 1024'd41477197265029861261843886154168149073829113833012076379879139997171751465436996000325807802300628736006465039394831596800562349461353018875754946568279222477161989696998170745984230659307066909312422005347323756367992029622514319343087825989594254936708339912189651311160633645695251672702178666948476585993;
            5'd31: xpb[104] = 1024'd113164231394868210096558074555368599264952526332029366598483162533897717205426741249345208417349998469224465204933905596288717270920089642419537515629809453088825438276321799595507507223143719048365281383611670461186729579068439634668011943009744084685796563177262305905259687342444652104826175524267929346647;
        endcase
    end

    always_comb begin
        case(flag[35][5:0])
            6'd0: xpb[105] = 1024'd0;
            6'd1: xpb[105] = 1024'd30392284920290908766236667775877308355688755852655486344477665002823393804053673794174768908870846946499657981507743080598904175768802965704079979837504321383399106143037105553700272297731582733053971576744388659820553139146734088513978745173332232584032441514108951234626106482632709759915741277480893811485;
            6'd2: xpb[105] = 1024'd60784569840581817532473335551754616711377511705310972688955330005646787608107347588349537817741693892999315963015486161197808351537605931408159959675008642766798212286074211107400544595463165466107943153488777319641106278293468177027957490346664465168064883028217902469252212965265419519831482554961787622970;
            6'd3: xpb[105] = 1024'd91176854760872726298710003327631925067066267557966459033432995008470181412161021382524306726612540839498973944523229241796712527306408897112239939512512964150197318429111316661100816893194748199161914730233165979461659417440202265541936235519996697752097324542326853703878319447898129279747223832442681434455;
            6'd4: xpb[105] = 1024'd121569139681163635064946671103509233422755023410621945377910660011293575216214695176699075635483387785998631926030972322395616703075211862816319919350017285533596424572148422214801089190926330932215886306977554639282212556586936354055914980693328930336129766056435804938504425930530839039662965109923575245940;
            6'd5: xpb[105] = 1024'd27894728917329802432384411474572109033745352137541747594256469949140073682959230060858773329696560423055140500081221968415457038002794493965239774171190565983304856145614310430871122297140707943959660275334703452738404845512773669604915156183431713653342304156427698143024004339234915782460016560778874573094;
            6'd6: xpb[105] = 1024'd58287013837620711198621079250449417389434107990197233938734134951963467487012903855033542238567407369554798481588965049014361213771597459669319754008694887366703962288651415984571394594872290677013631852079092112558957984659507758118893901356763946237374745670536649377650110821867625542375757838259768384579;
            6'd7: xpb[105] = 1024'd88679298757911619964857747026326725745122863842852720283211799954786861291066577649208311147438254316054456463096708129613265389540400425373399733846199208750103068431688521538271666892603873410067603428823480772379511123806241846632872646530096178821407187184645600612276217304500335302291499115740662196064;
            6'd8: xpb[105] = 1024'd119071583678202528731094414802204034100811619695508206627689464957610255095120251443383080056309101262554114444604451210212169565309203391077479713683703530133502174574725627091971939190335456143121575005567869432200064262952975935146851391703428411405439628698754551846902323787133045062207240393221556007549;
            6'd9: xpb[105] = 1024'd25397172914368696098532155173266909711801948422428008844035274895456753561864786327542777750522273899610623018654700856232009900236786022226399568504876810583210606148191515308041972296549833154865348973925018245656256551878813250695851567193531194722652166798746445051421902195837121805004291844076855334703;
            6'd10: xpb[105] = 1024'd55789457834659604864768822949144218067490704275083495188512939898280147365918460121717546659393120846110281000162443936830914076005588987930479548342381131966609712291228620861742244594281415887919320550669406905476809691025547339209830312366863427306684608312855396286048008678469831564920033121557749146188;
            6'd11: xpb[105] = 1024'd86181742754950513631005490725021526423179460127738981532990604901103541169972133915892315568263967792609938981670187017429818251774391953634559528179885453350008818434265726415442516892012998620973292127413795565297362830172281427723809057540195659890717049826964347520674115161102541324835774399038642957673;
            6'd12: xpb[105] = 1024'd116574027675241422397242158500898834778868215980394467877468269903926934974025807710067084477134814739109596963177930098028722427543194919338639508017389774733407924577302831969142789189744581354027263704158184225117915969319015516237787802713527892474749491341073298755300221643735251084751515676519536769158;
            6'd13: xpb[105] = 1024'd22899616911407589764679898871961710389858544707314270093814079841773433440770342594226782171347987376166105537228179744048562762470777550487559362838563055183116356150768720185212822295958958365771037672515333038574108258244852831786787978203630675791962029441065191959819800052439327827548567127374836096312;
            6'd14: xpb[105] = 1024'd53291901831698498530916566647839018745547300559969756438291744844596827244824016388401551080218834322665763518735922824647466938239580516191639342676067376566515462293805825738913094593690541098825009249259721698394661397391586920300766723376962908375994470955174143194445906535072037587464308404855729907797;
            6'd15: xpb[105] = 1024'd83684186751989407297153234423716327101236056412625242782769409847420221048877690182576319989089681269165421500243665905246371114008383481895719322513571697949914568436842931292613366891422123831878980826004110358215214536538321008814745468550295140960026912469283094429072013017704747347380049682336623719282;
            6'd16: xpb[105] = 1024'd114076471672280316063389902199593635456924812265280729127247074850243614852931363976751088897960528215665079481751408985845275289777186447599799302351076019333313674579880036846313639189153706564932952402748499018035767675685055097328724213723627373544059353983392045663698119500337457107295790959817517530767;
            6'd17: xpb[105] = 1024'd20402060908446483430827642570656511067915140992200531343592884788090113319675898860910786592173700852721588055801658631865115624704769078748719157172249299783022106153345925062383672295368083576676726371105647831491959964610892412877724389213730156861271892083383938868217697909041533850092842410672816857921;
            6'd18: xpb[105] = 1024'd50794345828737392197064310346533819423603896844856017688070549790913507123729572655085555501044547799221246037309401712464019800473572044452799137009753621166421212296383030616083944593099666309730697947850036491312513103757626501391703134387062389445304333597492890102843804391674243610008583688153710669406;
            6'd19: xpb[105] = 1024'd81186630749028300963300978122411127779292652697511504032548214793736900927783246449260324409915394745720904018817144793062923976242375010156879116847257942549820318439420136169784216890831249042784669524594425151133066242904360589905681879560394622029336775111601841337469910874306953369924324965634604480891;
            6'd20: xpb[105] = 1024'd111578915669319209729537645898288436134981408550166990377025879796560294731836920243435093318786241692220562000324887873661828152011177975860959096684762263933219424582457241723484489188562831775838641101338813810953619382051094678419660624733726854613369216625710792572096017356939663129840066243115498292376;
            6'd21: xpb[105] = 1024'd17904504905485377096975386269351311745971737277086792593371689734406793198581455127594791012999414329277070574375137519681668486938760607009878951505935544382927856155923129939554522294777208787582415069695962624409811670976931993968660800223829637930581754725702685776615595765643739872637117693970797619530;
            6'd22: xpb[105] = 1024'd48296789825776285863212054045228620101660493129742278937849354737230187002635128921769559921870261275776728555882880600280572662707563572713958931343439865766326962298960235493254794592508791520636386646440351284230364810123666082482639545397161870514614196239811637011241702248276449632552858971451691431015;
            6'd23: xpb[105] = 1024'd78689074746067194629448721821105928457349248982397765282327019740053580806688802715944328830741108222276386537390623680879476838476366538418038911180944187149726068441997341046955066890240374253690358223184739944050917949270400170996618290570494103098646637753920588245867808730909159392468600248932585242500;
            6'd24: xpb[105] = 1024'd109081359666358103395685389596983236813038004835053251626804684742876974610742476510119097739611955168776044518898366761478381014245169504122118891018448508533125174585034446600655339187971956986744329799929128603871471088417134259510597035743826335682679079268029539480493915213541869152384341526413479053985;
            6'd25: xpb[105] = 1024'd15406948902524270763123129968046112424028333561973053843150494680723473077487011394278795433825127805832553092948616407498221349172752135271038745839621788982833606158500334816725372294186333998488103768286277417327663377342971575059597211233929118999891617368021432685013493622245945895181392977268778381139;
            6'd26: xpb[105] = 1024'd45799233822815179529359797743923420779717089414628540187628159683546866881540685188453564342695974752332211074456359488097125524941555100975118725677126110366232712301537440370425644591917916731542075345030666077148216516489705663573575956407261351583924058882130383919639600104878655655097134254749672192624;
            6'd27: xpb[105] = 1024'd76191518743106088295596465519800729135405845267284026532105824686370260685594358982628333251566821698831869055964102568696029700710358066679198705514630431749631818444574545924125916889649499464596046921775054736968769655636439752087554701580593584167956500396239335154265706587511365415012875532230566004109;
            6'd28: xpb[105] = 1024'd106583803663396997061833133295678037491094601119939512876583489689193654489648032776803102160437668645331527037471845649294933876479161032383278685352134753133030924587611651477826189187381082197650018498519443396789322794783173840601533446753925816751988941910348286388891813070144075174928616809711459815594;
            6'd29: xpb[105] = 1024'd12909392899563164429270873666740913102084929846859315092929299627040152956392567660962799854650841282388035611522095295314774211406743663532198540173308033582739356161077539693896222293595459209393792466876592210245515083709011156150533622244028600069201480010340179593411391478848151917725668260566759142748;
            6'd30: xpb[105] = 1024'd43301677819854073195507541442618221457773685699514801437406964629863546760446241455137568763521688228887693593029838375913678387175546629236278520010812354966138462304114645247596494591327041942447764043620980870066068222855745244664512367417360832653233921524449130828037497961480861677641409538047652954233;
            6'd31: xpb[105] = 1024'd73693962740144981961744209218495529813462441552170287781884629632686940564499915249312337672392535175387351574537581456512582562944349594940358499848316676349537568447151750801296766889058624675501735620365369529886621362002479333178491112590693065237266363038558082062663604444113571437557150815528546765718;
            6'd32: xpb[105] = 1024'd104086247660435890727980876994372838169151197404825774126362294635510334368553589043487106581263382121887009556045324537111486738713152560644438479685820997732936674590188856354997039186790207408555707197109758189707174501149213421692469857764025297821298804552667033297289710926746281197472892093009440577203;
            6'd33: xpb[105] = 1024'd10411836896602058095418617365435713780141526131745576342708104573356832835298123927646804275476554758943518130095574183131327073640735191793358334506994278182645106163654744571067072293004584420299481165466907003163366790075050737241470033254128081138511342652658926501809289335450357940269943543864739904357;
            6'd34: xpb[105] = 1024'd40804121816892966861655285141313022135830281984401062687185769576180226639351797721821573184347401705443176111603317263730231249409538157497438314344498599566044212306691850124767344590736167153353452742211295662983919929221784825755448778427460313722543784166767877736435395818083067700185684821345633715842;
            6'd35: xpb[105] = 1024'd71196406737183875627891952917190330491519037837056549031663434579003620443405471515996342093218248651942834093111060344329135425178341123201518294182002920949443318449728955678467616888467749886407424318955684322804473068368518914269427523600792546306576225680876828971061502300715777460101426098826527527327;
            6'd36: xpb[105] = 1024'd101588691657474784394128620693067638847207793689712035376141099581827014247459145310171111002089095598442492074618803424928039600947144088905598274019507242332842424592766061232167889186199332619461395895700072982625026207515253002783406268774124778890608667194985780205687608783348487220017167376307421338812;
            6'd37: xpb[105] = 1024'd7914280893640951761566361064130514458198122416631837592486909519673512714203680194330808696302268235499000648669053070947879935874726720054518128840680522782550856166231949448237922292413709631205169864057221796081218496441090318332406444264227562207821205294977673410207187192052563962814218827162720665966;
            6'd38: xpb[105] = 1024'd38306565813931860527803028840007822813886878269287323936964574522496906518257353988505577605173115181998658630176796151546784111643529685758598108678184844165949962309269055001938194590145292364259141440801610455901771635587824406846385189437559794791853646809086624644833293674685273722729960104643614477451;
            6'd39: xpb[105] = 1024'd68698850734222769294039696615885131169575634121942810281442239525320300322311027782680346514043962128498316611684539232145688287412332651462678088515689165549349068452306160555638466887876875097313113017545999115722324774734558495360363934610892027375886088323195575879459400157317983482645701382124508288936;
            6'd40: xpb[105] = 1024'd99091135654513678060276364391762439525264389974598296625919904528143694126364701576855115422914809074997974593192282312744592463181135617166758068353193486932748174595343266109338739185608457830367084594290387775542877913881292583874342679784224259959918529837304527114085506639950693242561442659605402100421;
            6'd41: xpb[105] = 1024'd5416724890679845427714104762825315136254718701518098842265714465990192593109236461014813117127981712054483167242531958764432798108718248315677923174366767382456606168809154325408772291822834842110858562647536588999070202807129899423342855274327043277131067937296420318605085048654769985358494110460701427575;
            6'd42: xpb[105] = 1024'd35809009810970754193950772538702623491943474554173585186743379468813586397162910255189582025998828658554141148750275039363336973877521214019757903011871088765855712311846259879109044589554417575164830139391925248819623341953863987937321600447659275861163509451405371553231191531287479745274235387941595239060;
            6'd43: xpb[105] = 1024'd66201294731261662960187440314579931847632230406829071531221044471636980201216584049364350934869675605053799130258018119962241149646324179723837882849375410149254818454883365432809316887286000308218801716136313908640176481100598076451300345620991508445195950965514322787857298013920189505189976665422489050545;
            6'd44: xpb[105] = 1024'd96593579651552571726424108090457240203320986259484557875698709474460374005270257843539119843740522551553457111765761200561145325415127145427917862686879731532653924597920470986509589185017583041272773292880702568460729620247332164965279090794323741029228392479623274022483404496552899265105717942903382862030;
            6'd45: xpb[105] = 1024'd2919168887718739093861848461520115814311314986404360092044519412306872472014792727698817537953695188609965685816010846580985660342709776576837717508053011982362356171386359202579622291231960053016547261237851381916921909173169480514279266284426524346440930579615167227002982905256976007902769393758682189184;
            6'd46: xpb[105] = 1024'd33311453808009647860098516237397424170000070839059846436522184415130266276068466521873586446824542135109623667323753927179889836111512742280917697345557333365761462314423464756279894588963542786070518837982240041737475048319903569028258011457758756930473372093724118461629089387889685767818510671239576000669;
            6'd47: xpb[105] = 1024'd63703738728300556626335184013274732525688826691715332780999849417953660080122140316048355355695389081609281648831497007778794011880315707984997677183061654749160568457460570309980166886695125519124490414726628701558028187466637657542236756631090989514505813607833069696255195870522395527734251948720469812154;
            6'd48: xpb[105] = 1024'd94096023648591465392571851789152040881377582544370819125477514420777053884175814110223124264566236028108939630339240088377698187649118673689077657020565976132559674600497675863680439184426708252178461991471017361378581326613371746056215501804423222098538255121942020930881302353155105287649993226201363623639;
            6'd49: xpb[105] = 1024'd421612884757632760009592160214916492367911271290621341823324358623552350920348994382821958779408665165448204389489734397538522576701304837997511841739256582268106173963564079750472290641085263922235959828166174834773615539209061605215677294526005415750793221933914135400880761859182030447044677056662950793;
            6'd50: xpb[105] = 1024'd30813897805048541526246259936092224848056667123946107686300989361446946154974022788557590867650255611665106185897232814996442698345504270542077491679243577965667212317000669633450744588372667996976207536572554834655326754685943150119194422467858237999783234736042865370026987244491891790362785954537556762278;
            6'd51: xpb[105] = 1024'd61206182725339450292482927711969533203745422976601594030778654364270339959027696582732359776521102558164764167404975895595346874114307236246157471516747899349066318460037775187151016886104250730030179113316943494475879893832677238633173167641190470583815676250151816604653093727124601550278527232018450573763;
            6'd52: xpb[105] = 1024'd91598467645630359058719595487846841559434178829257080375256319367093733763081370376907128685391949504664422148912718976194251049883110201950237451354252220732465424603074880740851289183835833463084150690061332154296433032979411327147151912814522703167848117764260767839279200209757311310194268509499344385248;
            6'd53: xpb[105] = 1024'd121990752565921267824956263263724149915122934681912566719733984369917127567135044171081897594262796451164080130420462056793155225651913167654317431191756542115864530746111986294551561481567416196138122266805720814116986172126145415661130657987854935751880559278369719073905306692390021070110009786980238196733;
            6'd54: xpb[105] = 1024'd28316341802087435192394003634787025526113263408832368936079794307763626033879579055241595288475969088220588704470711702812995560579495798803237286012929822565572962319577874510621594587781793207881896235162869627573178461051982731210130833477957719069093097378361612278424885101094097812907061237835537523887;
            6'd55: xpb[105] = 1024'd58708626722378343958630671410664333881802019261487855280557459310587019837933252849416364197346816034720246685978454783411899736348298764507317265850434143948972068462614980064321866885513375940935867811907258287393731600198716819724109578651289951653125538892470563513050991583726807572822802515316431335372;
            6'd56: xpb[105] = 1024'd89100911642669252724867339186541642237490775114143341625035124313410413641986926643591133106217662981219904667486197864010803912117101730211397245687938465332371174605652085618022139183244958673989839388651646947214284739345450908238088323824622184237157980406579514747677098066359517332738543792797325146857;
            6'd57: xpb[105] = 1024'd119493196562960161491104006962418950593179530966798827969512789316233807446040600437765902015088509927719562648993940944609708087885904695915477225525442786715770280748689191171722411480976541407043810965396035607034837878492184996752067068997954416821190421920688465982303204548992227092654285070278218958342;
            6'd58: xpb[105] = 1024'd25818785799126328858541747333481826204169859693718630185858599254080305912785135321925599709301682564776071223044190590629548422813487327064397080346616067165478712322155079387792444587190918418787584933753184420491030167418022312301067244488057200138402960020680359186822782957696303835451336521133518285496;
            6'd59: xpb[105] = 1024'd56211070719417237624778415109359134559858615546374116530336264256903699716838809116100368618172529511275729204551933671228452598582290292768477060184120388548877818465192184941492716884922501151841556510497573080311583306564756400815045989661389432722435401534789310421448889440329013595367077798614412096981;
            6'd60: xpb[105] = 1024'd86603355639708146391015082885236442915547371399029602874813929259727093520892482910275137527043376457775387186059676751827356774351093258472557040021624709932276924608229290495192989182654083884895528087241961740132136445711490489329024734834721665306467843048898261656074995922961723355282819076095305908466;
            6'd61: xpb[105] = 1024'd116995640559999055157251750661113751271236127251685089219291594262550487324946156704449906435914223404275045167567419832426260950119896224176637019859129031315676030751266396048893261480385666617949499663986350399952689584858224577843003480008053897890500284563007212890701102405594433115198560353576199719951;
            6'd62: xpb[105] = 1024'd23321229796165222524689491032176626882226455978604891435637404200396985791690691588609604130127396041331553741617669478446101285047478855325556874680302311765384462324732284264963294586600043629693273632343499213408881873784061893392003655498156681207712822662999106095220680814298509857995611804431499047105;
            6'd63: xpb[105] = 1024'd53713514716456131290926158808053935237915211831260377780115069203220379595744365382784373038998242987831211723125412559045005460816281821029636854517806633148783568467769389818663566884331626362747245209087887873229435012930795981905982400671488913791745264177108057329846787296931219617911353081912392858590;
        endcase
    end

    always_comb begin
        case(flag[35][11:6])
            6'd0: xpb[106] = 1024'd0;
            6'd1: xpb[106] = 1024'd84105799636747040057162826583931243593603967683915864124592734206043773399798039176959141947869089934330869704633155639643909636585084786733716834355310954532182674610806495372363839182063209095801216785832276533049988152077530070419961145844821146375777705691217008564472893779563929377827094359393286670075;
            6'd2: xpb[106] = 1024'd44144903589369338715526725763048054442509508242096044121053613347110651462286939443903212681080505559218590001808817844708755432328949238912273543694290868130674674652041773407097439172609212470292235963277313219735615453934163367874943722006412843484735507968316959098839259485199225738535498892160978855819;
            6'd3: xpb[106] = 1024'd4184007541991637373890624942164865291415048800276224117514492488177529524775839710847283414291921184106310298984480049773601228072813691090830253033270781729166674693277051441831039163155215844783255140722349906421242755790796665329926298168004540593693310245416909633205625190834522099243903424928671041563;
            6'd4: xpb[106] = 1024'd88289807178738677431053451526096108885019016484192088242107226694221302924573878887806425362161011118437180003617635689417510864657898477824547087388581736261349349304083546814194878345218424940584471926554626439471230907868326735749887444012825686969471015936633918197678518970398451477070997784321957711638;
            6'd5: xpb[106] = 1024'd48328911131360976089417350705212919733924557042372268238568105835288180987062779154750496095372426743324900300793297894482356660401762930003103796727561649859841349345318824848928478335764428315075491103999663126156858209724960033204870020174417384078428818213733868732044884676033747837779402317089649897382;
            6'd6: xpb[106] = 1024'd8368015083983274747781249884329730582830097600552448235028984976355059049551679421694566828583842368212620597968960099547202456145627382181660506066541563458333349386554102883662078326310431689566510281444699812842485511581593330659852596336009081187386620490833819266411250381669044198487806849857342083126;
            6'd7: xpb[106] = 1024'd92473814720730314804944076468260974176434065284468312359621719182398832449349718598653708776452932302543490302602115739191112092730712168915377340421852517990516023997360598256025917508373640785367727067276976345892473663659123401079813742180830227563164326182050827830884144161232973576314901209250628753201;
            6'd8: xpb[106] = 1024'd52512918673352613463307975647377785025339605842648492356082598323465710511838618865597779509664347927431210599777777944255957888474576621093934049760832431589008024038595876290759517498919644159858746244722013032578100965515756698534796318342421924672122128459150778365250509866868269937023305742018320938945;
            6'd9: xpb[106] = 1024'd12552022625974912121671874826494595874245146400828672352543477464532588574327519132541850242875763552318930896953440149320803684218441073272490759099812345187500024079831154325493117489465647534349765422167049719263728267372389995989778894504013621781079930736250728899616875572503566297731710274786013124689;
            6'd10: xpb[106] = 1024'd96657822262721952178834701410425839467849114084744536477136211670576361974125558309500992190744853486649800601586595788964713320803525860006207593455123299719682698690637649697856956671528856630150982207999326252313716419449920066409740040348834768156857636427467737464089769352067495675558804634179299794764;
            6'd11: xpb[106] = 1024'd56696926215344250837198600589542650316754654642924716473597090811643240036614458576445062923956269111537520898762257994029559116547390312184764302794103213318174698731872927732590556662074860004642001385444362938999343721306553363864722616510426465265815438704567687998456135057702792036267209166946991980508;
            6'd12: xpb[106] = 1024'd16736030167966549495562499768659461165660195201104896470057969952710118099103358843389133657167684736425241195937920199094404912291254764363321012133083126916666698773108205767324156652620863379133020562889399625684971023163186661319705192672018162374773240981667638532822500763338088396975613699714684166252;
            6'd13: xpb[106] = 1024'd100841829804713589552725326352590704759264162885020760594650704158753891498901398020348275605036774670756110900571075838738314548876339551097037846488394081448849373383914701139687995834684072474934237348721676158734959175240716731739666338516839308750550946672884647097295394542902017774802708059107970836327;
            6'd14: xpb[106] = 1024'd60880933757335888211089225531707515608169703443200940591111583299820769561390298287292346338248190295643831197746738043803160344620204003275594555827373995047341373425149979174421595825230075849425256526166712845420586477097350029194648914678431005859508748949984597631661760248537314135511112591875663022071;
            6'd15: xpb[106] = 1024'd20920037709958186869453124710824326457075244001381120587572462440887647623879198554236417071459605920531551494922400248868006140364068455454151265166353908645833373466385257209155195815776079223916275703611749532106213778953983326649631490840022702968466551227084548166028125954172610496219517124643355207815;
            6'd16: xpb[106] = 1024'd105025837346705226926615951294755570050679211685296984712165196646931421023677237731195559019328695854862421199555555888511915776949153242187868099521664863178016048077191752581519034997839288319717492489444026065156201931031513397069592636684843849344244256918301556730501019733736539874046611484036641877890;
            6'd17: xpb[106] = 1024'd65064941299327525584979850473872380899584752243477164708626075787998299086166137998139629752540111479750141496731218093576761572693017694366424808860644776776508048118427030616252634988385291694208511666889062751841829232888146694524575212846435546453202059195401507264867385439371836234755016016804334063634;
            6'd18: xpb[106] = 1024'd25104045251949824243343749652989191748490292801657344705086954929065177148655038265083700485751527104637861793906880298641607368436882146544981518199624690375000048159662308650986234978931295068699530844334099438527456534744779991979557789008027243562159861472501457799233751145007132595463420549572026249378;
            6'd19: xpb[106] = 1024'd109209844888696864300506576236920435342094260485573208829679689135108950548453077442042842433620617038968731498540035938285517005021966933278698352554935644907182722770468804023350074160994504164500747630166375971577444686822310062399518934852848389937937567163718466363706644924571061973290514908965312919453;
            6'd20: xpb[106] = 1024'd69248948841319162958870475416037246190999801043753388826140568276175828610941977708986913166832032663856451795715698143350362800765831385457255061893915558505674722811704082058083674151540507538991766807611412658263071988678943359854501511014440087046895369440818416898073010630206358333998919441733005105197;
            6'd21: xpb[106] = 1024'd29288052793941461617234374595154057039905341601933568822601447417242706673430877975930983900043448288744172092891360348415208596509695837635811771232895472104166722852939360092817274142086510913482785985056449344948699290535576657309484087176031784155853171717918367432439376335841654694707323974500697290941;
            6'd22: xpb[106] = 1024'd113393852430688501674397201179085300633509309285849432947194181623286480073228917152890125847912538223075041797524515988059118233094780624369528605588206426636349397463745855465181113324149720009284002770888725877998687442613106727729445233020852930531630877409135375996912270115405584072534418333893983961016;
            6'd23: xpb[106] = 1024'd73432956383310800332761100358202111482414849844029612943655060764353358135717817419834196581123953847962762094700178193123964028838645076548085314927186340234841397504981133499914713314695723383775021948333762564684314744469740025184427809182444627640588679686235326531278635821040880433242822866661676146760;
            6'd24: xpb[106] = 1024'd33472060335933098991124999537318922331320390402209792940115939905420236198206717686778267314335369472850482391875840398188809824582509528726642024266166253833333397546216411534648313305241726758266041125778799251369942046326373322639410385344036324749546481963335277065645001526676176793951227399429368332504;
            6'd25: xpb[106] = 1024'd117577859972680139048287826121250165924924358086125657064708674111464009598004756863737409262204459407181352096508996037832719461167594315460358858621477208365516072157022906907012152487304935854067257911611075784419930198403903393059371531188857471125324187654552285630117895306240106171778321758822655002579;
            6'd26: xpb[106] = 1024'd77616963925302437706651725300366976773829898644305837061169553252530887660493657130681479995415875032069072393684658242897565256911458767638915567960457121964008072198258184941745752477850939228558277089056112471105557500260536690514354107350449168234281989931652236164484261011875402532486726291590347188323;
            6'd27: xpb[106] = 1024'd37656067877924736365015624479483787622735439202486017057630432393597765722982557397625550728627290656956792690860320447962411052655323219817472277299437035562500072239493462976479352468396942603049296266501149157791184802117169987969336683512040865343239792208752186698850626717510698893195130824358039374067;
            6'd28: xpb[106] = 1024'd121761867514671776422178451063415031216339406886401881182223166599641539122780596574584692676496380591287662395493476087606320689240408006551189111654747990094682746850299958348843191650460151698850513052333425690841172954194700058389297829356862011719017497899969195263323520497074628271022225183751326044142;
            6'd29: xpb[106] = 1024'd81800971467294075080542350242531842065244947444582061178684045740708417185269496841528763409707796216175382692669138292671166484984272458729745820993727903693174746891535236383576791641006155073341532229778462377526800256051333355844280405518453708827975300177069145797689886202709924631730629716519018229886;
            6'd30: xpb[106] = 1024'd41840075419916373738906249421648652914150488002762241175144924881775295247758397108472834142919211841063102989844800497736012280728136910908302530332707817291666746932770514418310391631552158447832551407223499064212427557907966653299262981680045405936933102454169096332056251908345220992439034249286710415630;
            6'd31: xpb[106] = 1024'd1879179372538672397270148600765463763056028560942421171605804022842173310247297375416904876130627465950823287020462702800858076472001363086859239671687730890158746974005792453043991622098161822323570584668535750898054859764599950754245557841637103045890904731269046866422617613980517353147438782054402601374;
            6'd32: xpb[106] = 1024'd85984979009285712454432975184696707356659996244858285296198538228885946710045336552376046823999717400281692991653618342444767713057086149820576074026998685422341421584812287825407830804161370918124787370500812283948043011842130021174206703686458249421668610422486055430895511393544446730974533141447689271449;
            6'd33: xpb[106] = 1024'd46024082961908011112796874363813518205565536803038465292659417369952824772534236819320117557211133025169413288829280547509613508800950601999132783365978599020833421626047565860141430794707374292615806547945848970633670313698763318629189279848049946530626412699586005965261877099179743091682937674215381457193;
            6'd34: xpb[106] = 1024'd6063186914530309771160773542930329054471077361218645289120296511019702835023137086264188290422548650057133586004942752574459304544815054177689492704958512619325421667282843894875030785253377667106825725390885657319297615555396616084171856009641643639584214976685956499628242804815039452391342206983073642937;
            6'd35: xpb[106] = 1024'd90168986551277349828323600126861572648075045045134509413713030717063476234821176263223330238291638584388003290638098392218368941129899840911406327060269467151508096278089339267238869967316586762908042511223162190369285767632926686504133001854462790015361920667902965064101136584378968830218436566376360313012;
            6'd36: xpb[106] = 1024'd50208090503899648486687499305978383496980585603314689410173909858130354297310076530167400971503054209275723587813760597283214736873764293089963036399249380750000096319324617301972469957862590137399061688668198877054913069489559983959115578016054487124319722945002915598467502290014265190926841099144052498756;
            6'd37: xpb[106] = 1024'd10247194456521947145051398485095194345886126161494869406634788999197232359798976797111471704714469834163443884989422802348060532617628745268519745738229294348492096360559895336706069948408593511890080866113235563740540371346193281414098154177646184233277525222102866132833867995649561551635245631911744684500;
            6'd38: xpb[106] = 1024'd94352994093268987202214225069026437939490093845410733531227523205241005759597015974070613652583559768494313589622578441991970169202713532002236580093540248880674770971366390709069909130471802607691297651945512096790528523423723351834059300022467330609055230913319874697306761775213490929462339991305031354575;
            6'd39: xpb[106] = 1024'd54392098045891285860578124248143248788395634403590913527688402346307883822085916241014684385794975393382033886798240647056815964946577984180793289432520162479166771012601668743803509121017805982182316829390548783476155825280356649289041876184059027718013033190419825231673127480848787290170744524072723540319;
            6'd40: xpb[106] = 1024'd14431201998513584518942023427260059637301174961771093524149281487374761884574816507958755119006391018269754183973902852121661760690442436359349998771500076077658771053836946778537109111563809356673336006835585470161783127136989946744024452345650724826970835467519775766039493186484083650879149056840415726063;
            6'd41: xpb[106] = 1024'd98537001635260624576104850011191303230905142645686957648742015693418535284372855684917897066875480952600623888607058491765571397275527223093066833126811030609841445664643442150900948293627018452474552792667862003211771279214520017163985598190471871202748541158736784330512386966048013028706243416233702396138;
            6'd42: xpb[106] = 1024'd58576105587882923234468749190308114079810683203867137645202894834485413346861755951861967800086896577488344185782720696830417193019391675271623542465790944208333445705878720185634548284173021826965571970112898689897398581071153314618968174352063568311706343435836734864878752671683309389414647949001394581882;
            6'd43: xpb[106] = 1024'd18615209540505221892832648369424924928716223762047317641663773975552291409350656218806038533298312202376064482958382901895262988763256127450180251804770857806825445747113998220368148274719025201456591147557935376583025882927786612073950750513655265420664145712936685399245118377318605750123052481769086767626;
            6'd44: xpb[106] = 1024'd102721009177252261949995474953356168522320191445963181766256508181596064809148695395765180481167402136706934187591538541539172625348340914183897086160081812339008120357920493592731987456782234297257807933390211909633014035005316682493911896358476411796441851404153693963718012156882535127950146841162373437701;
            6'd45: xpb[106] = 1024'd62760113129874560608359374132472979371225732004143361762717387322662942871637595662709251214378817761594654484767200746604018421092205366362453795499061725937500120399155771627465587447328237671748827110835248596318641336861949979948894472520068108905399653681253644498084377862517831488658551373930065623445;
            6'd46: xpb[106] = 1024'd22799217082496859266723273311589790220131272562323541759178266463729820934126495929653321947590233386482374781942862951668864216836069818541010504838041639535992120440391049662199187437874241046239846288280285283004268638718583277403877048681659806014357455958353595032450743568153127849366955906697757809189;
            6'd47: xpb[106] = 1024'd106905016719243899323886099895521033813735240246239405883771000669773594333924535106612463895459323320813244486576018591312773853421154605274727339193352594068174795051197545034563026619937450142041063074112561816054256790796113347823838194526480952390135161649570603596923637347717057227194050266091044479264;
            6'd48: xpb[106] = 1024'd66944120671866197982249999074637844662640780804419585880231879810840472396413435373556534628670738945700964783751680796377619649165019057453284048532332507666666795092432823069296626610483453516532082251557598502739884092652746645278820770688072649499092963926670554131290003053352353587902454798858736665008;
            6'd49: xpb[106] = 1024'd26983224624488496640613898253754655511546321362599765876692758951907350458902335640500605361882154570588685080927343001442465444908883509631840757871312421265158795133668101104030226601029456891023101429002635189425511394509379942733803346849664346608050766203770504665656368758987649948610859331626428850752;
            6'd50: xpb[106] = 1024'd111089024261235536697776724837685899105150289046515630001285493157951123858700374817459747309751244504919554785560498641086375081493968296365557592226623375797341469744474596476394065783092665986824318214834911722475499546586910013153764492694485492983828471894987513230129262538551579326437953691019715520827;
            6'd51: xpb[106] = 1024'd71128128213857835356140624016802709954055829604695809997746372299018001921189275084403818042962660129807275082736160846151220877237832748544114301565603289395833469785709874511127665773638669361315337392279948409161126848443543310608747068856077190092786274172087463764495628244186875687146358223787407706571;
            6'd52: xpb[106] = 1024'd31167232166480134014504523195919520802961370162875989994207251440084879983678175351347888776174075754694995379911823051216066672981697200722671010904583202994325469826945152545861265764184672735806356569724985095846754150300176608063729645017668887201744076449187414298861993949822172047854762756555099892315;
            6'd53: xpb[106] = 1024'd115273031803227174071667349779850764396565337846791854118799985646128653383476214528307030724043165689025865084544978690859976309566781987456387845259894157526508144437751647918225104946247881831607573355557261628896742302377706678483690790862490033577521782140404422863334887729386101425681857115948386562390;
            6'd54: xpb[106] = 1024'd75312135755849472730031248958967575245470878404972034115260864787195531445965114795251101457254581313913585381720640895924822105310646439634944554598874071125000144478986925952958704936793885206098592533002298315582369604234339975938673367024081730686479584417504373397701253435021397786390261648716078748134;
            6'd55: xpb[106] = 1024'd35351239708471771388395148138084386094376418963152214111721743928262409508454015062195172190465996938801305678896303100989667901054510891813501263937853984723492144520222203987692304927339888580589611710447335002267996906090973273393655943185673427795437386694604323932067619140656694147098666181483770933878;
            6'd56: xpb[106] = 1024'd119457039345218811445557974722015629687980386647068078236314478134306182908252054239154314138335086873132175383529458740633577537639595678547218098293164939255674819131028699360056144109403097676390828496279611535317985058168503343813617089030494574171215092385821332496540512920220623524925760540877057603953;
            6'd57: xpb[106] = 1024'd79496143297841110103921873901132440536885927205248258232775357275373060970740954506098384871546502498019895680705120945698423333383460130725774807632144852854166819172263977394789744099949101050881847673724648222003612360025136641268599665192086271280172894662921283030906878625855919885634165073644749789697;
            6'd58: xpb[106] = 1024'd39535247250463408762285773080249251385791467763428438229236236416439939033229854773042455604757918122907615977880783150763269129127324582904331516971124766452658819213499255429523344090495104425372866851169684908689239661881769938723582241353677968389130696940021233565273244331491216246342569606412441975441;
            6'd59: xpb[106] = 1024'd123641046887210448819448599664180494979395435447344302353828970622483712433027893950001597552627008057238485682513938790407178765712409369638048351326435720984841493824305750801887183272558313521174083637001961441739227813959300009143543387198499114764908402631238242129746138111055145624169663965805728645516;
            6'd60: xpb[106] = 1024'd83680150839832747477812498843297305828300976005524482350289849763550590495516794216945668285838423682126205979689600995472024561456273821816605060665415634583333493865541028836620783263104316895665102814446998128424855115815933306598525963360090811873866204908338192664112503816690441984878068498573420831260;
            6'd61: xpb[106] = 1024'd43719254792455046136176398022414116677206516563704662346750728904617468558005694483889739019049839307013926276865263200536870357200138273995161770004395548181825493906776306871354383253650320270156121991892034815110482417672566604053508539521682508982824007185438143198478869522325738345586473031341113017004;
            6'd62: xpb[106] = 1024'd3758358745077344794540297201530927526112057121884842343211608045684346620494594750833809752261254931901646574040925405601716152944002726173718479343375461780317493948011584906087983244196323644647141169337071501796109719529199901508491115683274206091781809462538093732845235227961034706294877564108805202748;
            6'd63: xpb[106] = 1024'd87864158381824384851703123785462171119716024805800706467804342251728120020292633927792951700130344866232516278674081045245625789529087512907435313698686416312500168558818080278451822426259532740448357955169348034846097871606729971928452261528095352467559515153755102297318129007524964084121971923502091872823;
        endcase
    end

    always_comb begin
        case(flag[35][16:12])
            5'd0: xpb[107] = 1024'd0;
            5'd1: xpb[107] = 1024'd47903262334446683510067022964578981968621565363980886464265221392794998082781534194737022433341760491120236575849743250310471585272951965085992023037666329910992168600053358313185422416805536114939377132614384721531725173463363269383434837689687049576517317430855052831684494713160260444830376456269784058567;
            5'd2: xpb[107] = 1024'd95806524668893367020134045929157963937243130727961772928530442785589996165563068389474044866683520982240473151699486500620943170545903930171984046075332659821984337200106716626370844833611072229878754265228769443063450346926726538766869675379374099153034634861710105663368989426320520889660752912539568117134;
            5'd3: xpb[107] = 1024'd19643091319215309131402141488922513161166268966206975264663809113408098911035463674195996085367607163917560320091736316352350914977635560702815944096667948799285831230588857601926028058899402623507933789455914318230814670169193035185325943385831699462732048878448100464946956065552148317372439542183757691370;
            5'd4: xpb[107] = 1024'd67546353653661992641469164453501495129787834330187861728929030506203096993816997868933018518709367655037796895941479566662822500250587525788807967134334278710277999830642215915111450475704938738447310922070299039762539843632556304568760781075518749039249366309303153296631450778712408762202815998453541749937;
            5'd5: xpb[107] = 1024'd115449615988108676151536187418080477098409399694168748193194251898998095076598532063670040952051128146158033471791222816973294085523539490874799990172000608621270168430695574228296872892510474853386688054684683761294265017095919573952195618765205798615766683740158206128315945491872669207033192454723325808504;
            5'd6: xpb[107] = 1024'd39286182638430618262804282977845026322332537932413950529327618226816197822070927348391992170735214327835120640183472632704701829955271121405631888193335897598571662461177715203852056117798805247015867578911828636461629340338386070370651886771663398925464097756896200929893912131104296634744879084367515382740;
            5'd7: xpb[107] = 1024'd87189444972877301772871305942424008290954103296394836993592839619611195904852461543129014604076974818955357216033215883015173415228223086491623911231002227509563831061231073517037478534604341361955244711526213357993354513801749339754086724461350448501981415187751253761578406844264557079575255540637299441307;
            5'd8: xpb[107] = 1024'd11026011623199243884139401502188557514877241534640039329726205947429298650324856827850965822761061000632444384425465698746581159659954717022455809252337516486865325091713214492592661759892671755584424235753358233160718837044215836172542992467808048811678829204489248563156373483496184507286942170281489015543;
            5'd9: xpb[107] = 1024'd58929273957645927394206424466767539483498806898620925793991427340224296733106391022587988256102821491752680960275208949057052744932906682108447832290003846397857493691766572805778084176698207870523801368367742954692444010507579105555977830157495098388196146635344301394840868196656444952117318626551273074110;
            5'd10: xpb[107] = 1024'd106832536292092610904273447431346521452120372262601812258256648733019294815887925217325010689444581982872917536124952199367524330205858647194439855327670176308849662291819931118963506593503743985463178500982127676224169183970942374939412667847182147964713464066199354226525362909816705396947695082821057132677;
            5'd11: xpb[107] = 1024'd30669102942414553015541542991111070676043510500847014594390015060837397561360320502046961908128668164550004704517202015098932074637590277725271753349005465286151156322302072094518689818792074379092358025209272551391533507213408871357868935853639748274410878082937349028103329549048332824659381712465246706913;
            5'd12: xpb[107] = 1024'd78572365276861236525608565955690052644665075864827901058655236453632395644141854696783984341470428655670241280366945265409403659910542242811263776386671795197143324922355430407704112235597610494031735157823657272923258680676772140741303773543326797850928195513792401859787824262208593269489758168735030765480;
            5'd13: xpb[107] = 1024'd2408931927183178636876661515454601868588214103073103394788602781450498389614249981505935560154514837347328448759195081140811404342273873342095674408007084174444818952837571383259295460885940887660914682050802148090623003919238637159760041549784398160625609530530396661365790901440220697201444798379220339716;
            5'd14: xpb[107] = 1024'd50312194261629862146943684480033583837209779467053989859053824174245496472395784176242957993496275328467565024608938331451282989615225838428087697445673414085436987552890929696444717877691477002600291814665186869622348177382601906543194879239471447737142926961385449493050285614600481142031821254649004398283;
            5'd15: xpb[107] = 1024'd98215456596076545657010707444612565805831344831034876323319045567040494555177318370979980426838035819587801600458681581761754574888177803514079720483339743996429156152944288009630140294497013117539668947279571591154073350845965175926629716929158497313660244392240502324734780327760741586862197710918788456850;
            5'd16: xpb[107] = 1024'd22052023246398487768278803004377115029754483069280078659452411894858597300649713655701931645522122001264888768850931397493162319319909434044911618504675032973730650183426428985185323519785343511168848471506716466321437674088431672345085984935616097623357658408978497126312746966992369014573884340562978031086;
            5'd17: xpb[107] = 1024'd69955285580845171278345825968956096998376048433260965123717633287653595383431247850438954078863882492385125344700674647803633904592861399130903641542341362884722818783479787298370745936590879626108225604121101187853162847551794941728520822625303147199874975839833549957997241680152629459404260796832762089653;
            5'd18: xpb[107] = 1024'd117858547915291854788412848933535078966997613797241851587982854680448593466212782045175976512205642983505361920550417898114105489865813364216895664580007692795714987383533145611556168353396415741047602736735485909384888021015158211111955660314990196776392293270688602789681736393312889904234637253102546148220;
            5'd19: xpb[107] = 1024'd41695114565613796899680944493299628190920752035487053924116221008266696211685177329897927730889729165182449088942667713845513234297544994747727562601342981773016481414015286587111351578684746134676782260962630784552252344257624707530411928321447797086089707287426597591259703032544517331946323882746735722456;
            5'd20: xpb[107] = 1024'd89598376900060480409747967457878610159542317399467940388381442401061694294466711524634950164231489656302685664792410964155984819570496959833719585639009311684008650014068644900296773995490282249616159393577015506083977517720987976913846766011134846662607024718281650422944197745704777776776700339016519781023;
            5'd21: xpb[107] = 1024'd13434943550382422521016063017643159383465455637713142724514808728879797039939106809356901382915575837979772833184660779887392564002228590364551483660344600661310144044550785875851957220778612643245338917804160381251341840963454473332303034017592446972304438735019645224522164384936405204488386968660709355259;
            5'd22: xpb[107] = 1024'd61338205884829106031083085982222141352087021001694029188780030121674795122720641004093923816257336329100009409034404030197864149275180555450543506698010930572302312644604144189037379637584148758184716050418545102783067014426817742715737871707279496548821756165874698056206659098096665649318763424930493413826;
            5'd23: xpb[107] = 1024'd109241468219275789541150108946801123320708586365674915653045251514469793205502175198830946249599096820220245984884147280508335734548132520536535529735677260483294481244657502502222802054389684873124093183032929824314792187890181012099172709396966546125339073596729750887891153811256926094149139881200277472393;
            5'd24: xpb[107] = 1024'd33078034869597731652418204506565672544631724603920117989178617842287895950974570483552897468283183001897333153276397096239743478979864151067367427757012549460595975275139643477777985279678015266753272707260074699482156511132647508517628977403424146435036487613467745689469120450488553521860826510844467046629;
            5'd25: xpb[107] = 1024'd80981297204044415162485227471144654513253289967901004453443839235082894033756104678289919901624943493017569729126140346550215064252816116153359450794678879371588143875193001790963407696483551381692649839874459421013881684596010777901063815093111196011553805044322798521153615163648813966691202967114251105196;
            5'd26: xpb[107] = 1024'd4817863854366357273753323030909203737176428206146206789577205562900996779228499963011871120309029674694656897518390162281622808684547746684191348816014168348889637905675142766518590921771881775321829364101604296181246007838477274319520083099568796321251219061060793322731581802880441394402889596758440679432;
            5'd27: xpb[107] = 1024'd52721126188813040783820345995488185705797993570127093253842426955695994862010034157748893553650790165814893473368133412592094393957499711770183371853680498259881806505728501079704013338577417890261206496715989017712971181301840543702954920789255845897768536491915846154416076516040701839233266053028224737999;
            5'd28: xpb[107] = 1024'd100624388523259724293887368960067167674419558934107979718107648348490992944791568352485915986992550656935130049217876662902565979230451676856175394891346828170873975105781859392889435755382954005200583629330373739244696354765203813086389758478942895474285853922770898986100571229200962284063642509298008796566;
            5'd29: xpb[107] = 1024'd24460955173581666405155464519831716898342697172353182054241014676309095690263963637207867205676636838612217217610126478633973723662183307387007292912682117148175469136264000368444618980671284398829763153557518614412060678007670309504846026485400495783983267939508893787678537868432589711775329138942198370802;
            5'd30: xpb[107] = 1024'd72364217508028349915222487484410698866964262536334068518506236069104093773045497831944889639018397329732453793459869728944445308935135272472999315950348447059167637736317358681630041397476820513769140286171903335943785851471033578888280864175087545360500585370363946619363032581592850156605705595211982429369;
            5'd31: xpb[107] = 1024'd120267479842475033425289510448989680835585827900314954982771457461899091855827032026681912072360157820852690369309612979254916894208087237558991338988014776970159806336370716994815463814282356628708517418786288057475511024934396848271715701864774594937017902801218999451047527294753110601436082051481766487936;
        endcase
    end

    always_comb begin
        case(flag[36][5:0])
            6'd0: xpb[108] = 1024'd0;
            6'd1: xpb[108] = 1024'd22052023246398487768278803004377115029754483069280078659452411894858597300649713655701931645522122001264888768850931397493162319319909434044911618504675032973730650183426428985185323519785343511168848471506716466321437674088431672345085984935616097623357658408978497126312746966992369014573884340562978031086;
            6'd2: xpb[108] = 1024'd44104046492796975536557606008754230059508966138560157318904823789717194601299427311403863291044244002529777537701862794986324638639818868089823237009350065947461300366852857970370647039570687022337696943013432932642875348176863344690171969871232195246715316817956994252625493933984738029147768681125956062172;
            6'd3: xpb[108] = 1024'd66156069739195463304836409013131345089263449207840235978357235684575791901949140967105794936566366003794666306552794192479486957959728302134734855514025098921191950550279286955555970559356030533506545414520149398964313022265295017035257954806848292870072975226935491378938240900977107043721653021688934093258;
            6'd4: xpb[108] = 1024'd88208092985593951073115212017508460119017932277120314637809647579434389202598854622807726582088488005059555075403725589972649277279637736179646474018700131894922600733705715940741294079141374044675393886026865865285750696353726689380343939742464390493430633635913988505250987867969476058295537362251912124344;
            6'd5: xpb[108] = 1024'd110260116231992438841394015021885575148772415346400393297262059474292986503248568278509658227610610006324443844254656987465811596599547170224558092523375164868653250917132144925926617598926717555844242357533582331607188370442158361725429924678080488116788292044892485631563734834961845072869421702814890155430;
            6'd6: xpb[108] = 1024'd8245443794266185210873890621448257433828471289944787828582616304174688466589143024196518658475057698146183205648094950379910075078236269714309586011719156908693226530987356573481701927194855345702893220653058951564265194309693261105537339930467136473326047039753924727769953728025581070324616216752273702185;
            6'd7: xpb[108] = 1024'd30297467040664672979152693625825372463582954359224866488035028199033285767238856679898450303997179699411071974499026347873072394398145703759221204516394189882423876714413785558667025446980198856871741692159775417885702868398124933450623324866083234096683705448732421854082700695017950084898500557315251733271;
            6'd8: xpb[108] = 1024'd52349490287063160747431496630202487493337437428504945147487440093891883067888570335600381949519301700675960743349957745366234713718055137804132823021069222856154526897840214543852348966765542368040590163666491884207140542486556605795709309801699331720041363857710918980395447662010319099472384897878229764357;
            6'd9: xpb[108] = 1024'd74401513533461648515710299634579602523091920497785023806939851988750480368538283991302313595041423701940849512200889142859397033037964571849044441525744255829885177081266643529037672486550885879209438635173208350528578216574988278140795294737315429343399022266689416106708194629002688114046269238441207795443;
            6'd10: xpb[108] = 1024'd96453536779860136283989102638956717552846403567065102466392263883609077669187997647004245240563545703205738281051820540352559352357874005893956060030419288803615827264693072514222996006336229390378287106679924816850015890663419950485881279672931526966756680675667913233020941595995057128620153579004185826529;
            6'd11: xpb[108] = 1024'd118505560026258624052267905643333832582600886636345181125844675778467674969837711302706176886085667704470627049902751937845721671677783439938867678535094321777346477448119501499408319526121572901547135578186641283171453564751851622830967264608547624590114339084646410359333688562987426143194037919567163857615;
            6'd12: xpb[108] = 1024'd16490887588532370421747781242896514867656942579889575657165232608349376933178286048393037316950115396292366411296189900759820150156472539428619172023438313817386453061974713146963403854389710691405786441306117903128530388619386522211074679860934272946652094079507849455539907456051162140649232433504547404370;
            6'd13: xpb[108] = 1024'd38542910834930858190026584247273629897411425649169654316617644503207974233827999704094968962472237397557255180147121298252982469476381973473530790528113346791117103245401142132148727374175054202574634912812834369449968062707818194556160664796550370570009752488486346581852654423043531155223116774067525435456;
            6'd14: xpb[108] = 1024'd60594934081329345958305387251650744927165908718449732976070056398066571534477713359796900607994359398822143948998052695746144788796291407518442409032788379764847753428827571117334050893960397713743483384319550835771405736796249866901246649732166468193367410897464843708165401390035900169797001114630503466542;
            6'd15: xpb[108] = 1024'd82646957327727833726584190256027859956920391787729811635522468292925168835127427015498832253516481400087032717848984093239307108116200841563354027537463412738578403612254000102519374413745741224912331855826267302092843410884681539246332634667782565816725069306443340834478148357028269184370885455193481497628;
            6'd16: xpb[108] = 1024'd104698980574126321494862993260404974986674874857009890294974880187783766135777140671200763899038603401351921486699915490732469427436110275608265646042138445712309053795680429087704697933531084736081180327332983768414281084973113211591418619603398663440082727715421837960790895324020638198944769795756459528714;
            6'd17: xpb[108] = 1024'd2684308136400067864342868859967657271730930800554284826295437017665468099117715416887624329903051093173660848093353453646567905914799375098017139530482437752349029409535640735259782261799222525939831190452460388371357908840648110971526034855785311796620482710283277056997114217084374196399964309693843075469;
            6'd18: xpb[108] = 1024'd24736331382798555632621671864344772301485413869834363485747848912524065399767429072589555975425173094438549616944284851139730225234708809142928758035157470726079679592962069720445105781584566037108679661959176854692795582929079783316612019791401409419978141119261774183309861184076743210973848650256821106555;
            6'd19: xpb[108] = 1024'd46788354629197043400900474868721887331239896939114442145200260807382662700417142728291487620947295095703438385795216248632892544554618243187840376539832503699810329776388498705630429301369909548277528133465893321014233257017511455661698004727017507043335799528240271309622608151069112225547732990819799137641;
            6'd20: xpb[108] = 1024'd68840377875595531169179277873099002360994380008394520804652672702241260001066856383993419266469417096968327154646147646126054863874527677232751995044507536673540979959814927690815752821155253059446376604972609787335670931105943128006783989662633604666693457937218768435935355118061481240121617331382777168727;
            6'd21: xpb[108] = 1024'd90892401121994018937458080877476117390748863077674599464105084597099857301716570039695350911991539098233215923497079043619217183194437111277663613549182569647271630143241356676001076340940596570615225076479326253657108605194374800351869974598249702290051116346197265562248102085053850254695501671945755199813;
            6'd22: xpb[108] = 1024'd112944424368392506705736883881853232420503346146954678123557496491958454602366283695397282557513661099498104692348010441112379502514346545322575232053857602621002280326667785661186399860725940081784073547986042719978546279282806472696955959533865799913408774755175762688560849052046219269269386012508733230899;
            6'd23: xpb[108] = 1024'd10929751930666253075216759481415914705559402090499072654878053321840156565706858441084142988378108791319844053741448404026477980993035644812326725542201594661042255940522997308741484188994077871642724411105519339935623103150341372077063374786252448269946529750037201784767067945109955266724580526446116777654;
            6'd24: xpb[108] = 1024'd32981775177064740843495562485793029735313885159779151314330465216698753866356572096786074633900230792584732822592379801519640300312945078857238344046876627634772906123949426293926807708779421382811572882612235806257060777238773044422149359721868545893304188159015698911079814912102324281298464867009094808740;
            6'd25: xpb[108] = 1024'd55033798423463228611774365490170144765068368229059229973782877111557351167006285752488006279422352793849621591443311199012802619632854512902149962551551660608503556307375855279112131228564764893980421354118952272578498451327204716767235344657484643516661846567994196037392561879094693295872349207572072839826;
            6'd26: xpb[108] = 1024'd77085821669861716380053168494547259794822851298339308633235289006415948467655999408189937924944474795114510360294242596505964938952763946947061581056226693582234206490802284264297454748350108405149269825625668738899936125415636389112321329593100741140019504976972693163705308846087062310446233548135050870912;
            6'd27: xpb[108] = 1024'd99137844916260204148331971498924374824577334367619387292687700901274545768305713063891869570466596796379399129145173993999127258272673380991973199560901726555964856674228713249482778268135451916318118297132385205221373799504068061457407314528716838763377163385951190290018055813079431325020117888698028901998;
            6'd28: xpb[108] = 1024'd121189868162658691916610774503301489854331817436899465952140112796133143068955426719593801215988718797644287897996105391492289577592582815036884818065576759529695506857655142234668101787920795427486966768639101671542811473592499733802493299464332936386734821794929687416330802780071800339594002229261006933084;
            6'd29: xpb[108] = 1024'd19175195724932438286090650102864172139387873380443860483460669626014845032296001465280661646853166489466027259389543354406388056071271914526636311553920751569735482471510353882223186116188933217345617631758578291499888297460034633182600714716719584743272576789791126512537021673135536337049196743198390479839;
            6'd30: xpb[108] = 1024'd41227218971330926054369453107241287169142356449723939142913081520873442332945715120982593292375288490730916028240474751899550375391181348571547930058595784543466132654936782867408509635974276728514466103265294757821325971548466305527686699652335682366630235198769623638849768640127905351623081083761368510925;
            6'd31: xpb[108] = 1024'd63279242217729413822648256111618402198896839519004017802365493415732039633595428776684524937897410491995804797091406149392712694711090782616459548563270817517196782838363211852593833155759620239683314574772011224142763645636897977872772684587951779989987893607748120765162515607120274366196965424324346542011;
            6'd32: xpb[108] = 1024'd85331265464127901590927059115995517228651322588284096461817905310590636934245142432386456583419532493260693565942337546885875014031000216661371167067945850490927433021789640837779156675544963750852163046278727690464201319725329650217858669523567877613345552016726617891475262574112643380770849764887324573097;
            6'd33: xpb[108] = 1024'd107383288710526389359205862120372632258405805657564175121270317205449234234894856088088388228941654494525582334793268944379037333350909650706282785572620883464658083205216069822964480195330307262021011517785444156785638993813761322562944654459183975236703210425705115017788009541105012395344734105450302604183;
            6'd34: xpb[108] = 1024'd5368616272800135728685737719935314543461861601108569652590874035330936198235430833775248659806102186347321696186706907293135811829598750196034279060964875504698058819071281470519564523598445051879662380904920776742715817681296221943052069711570623593240965420566554113994228434168748392799928619387686150938;
            6'd35: xpb[108] = 1024'd27420639519198623496964540724312429573216344670388648312043285930189533498885144489477180305328224187612210465037638304786298131149508184240945897565639908478428709002497710455704888043383788563048510852411637243064153491769727894288138054647186721216598623829545051240306975401161117407373812959950664182024;
            6'd36: xpb[108] = 1024'd49472662765597111265243343728689544602970827739668726971495697825048130799534858145179111950850346188877099233888569702279460450469417618285857516070314941452159359185924139440890211563169132074217359323918353709385591165858159566633224039582802818839956282238523548366619722368153486421947697300513642213110;
            6'd37: xpb[108] = 1024'd71524686011995599033522146733066659632725310808948805630948109719906728100184571800881043596372468190141988002739501099772622769789327052330769134574989974425890009369350568426075535082954475585386207795425070175707028839946591238978310024518418916463313940647502045492932469335145855436521581641076620244196;
            6'd38: xpb[108] = 1024'd93576709258394086801800949737443774662479793878228884290400521614765325400834285456582975241894590191406876771590432497265785089109236486375680753079665007399620659552776997411260858602739819096555056266931786642028466514035022911323396009454035014086671599056480542619245216302138224451095465981639598275282;
            6'd39: xpb[108] = 1024'd115628732504792574570079752741820889692234276947508962949852933509623922701483999112284906887416712192671765540441363894758947408429145920420592371584340040373351309736203426396446182122525162607723904738438503108349904188123454583668481994389651111710029257465459039745557963269130593465669350322202576306368;
            6'd40: xpb[108] = 1024'd13614060067066320939559628341383571977290332891053357481173490339505624664824573857971767318281159884493504901834801857673045886907835019910343865072684032413391285350058638044001266450793300397582555601557979728306981011990989483048589409642037760066567012460320478841764182162194329463124544836139959853123;
            6'd41: xpb[108] = 1024'd35666083313464808707838431345760687007044815960333436140625902234364221965474287513673698963803281885758393670685733255166208206227744453955255483577359065387121935533485067029186589970578643908751404073064696194628418686079421155393675394577653857689924670869298975968076929129186698477698429176702937884209;
            6'd42: xpb[108] = 1024'd57718106559863296476117234350137802036799299029613514800078314129222819266124001169375630609325403887023282439536664652659370525547653888000167102082034098360852585716911496014371913490363987419920252544571412660949856360167852827738761379513269955313282329278277473094389676096179067492272313517265915915295;
            6'd43: xpb[108] = 1024'd79770129806261784244396037354514917066553782098893593459530726024081416566773714825077562254847525888288171208387596050152532844867563322045078720586709131334583235900337924999557237010149330931089101016078129127271294034256284500083847364448886052936639987687255970220702423063171436506846197857828893946381;
            6'd44: xpb[108] = 1024'd101822153052660272012674840358892032096308265168173672118983137918940013867423428480779493900369647889553059977238527447645695164187472756089990339091384164308313886083764353984742560529934674442257949487584845593592731708344716172428933349384502150559997646096234467347015170030163805521420082198391871977467;
            6'd45: xpb[108] = 1024'd123874176299058759780953643363269147126062748237453750778435549813798611168073142136481425545891769890817948746089458845138857483507382190134901957596059197282044536267190782969927884049720017953426797959091562059914169382433147844774019334320118248183355304505212964473327916997156174535993966538954850008553;
            6'd46: xpb[108] = 1024'd21859503861332506150433518962831829411118804180998145309756106643680313131413716882168285976756217582639688107482896808052955961986071289624653451084403189322084511881045994617482968377988155743285448822211038679871246206300682744154126749572504896539893059500074403569534135890219910533449161052892233555308;
            6'd47: xpb[108] = 1024'd43911527107730993918712321967208944440873287250278223969208518538538910432063430537870217622278339583904576876333828205546118281305980723669565069589078222295815162064472423602668291897773499254454297293717755146192683880389114416499212734508120994163250717909052900695846882857212279548023045393455211586394;
            6'd48: xpb[108] = 1024'd65963550354129481686991124971586059470627770319558302628660930433397507732713144193572149267800461585169465645184759603039280600625890157714476688093753255269545812247898852587853615417558842765623145765224471612514121554477546088844298719443737091786608376318031397822159629824204648562596929734018189617480;
            6'd49: xpb[108] = 1024'd88015573600527969455269927975963174500382253388838381288113342328256105033362857849274080913322583586434354414035691000532442919945799591759388306598428288243276462431325281573038938937344186276791994236731188078835559228565977761189384704379353189409966034727009894948472376791197017577170814074581167648566;
            6'd50: xpb[108] = 1024'd110067596846926457223548730980340289530136736458118459947565754223114702334012571504976012558844705587699243182886622398025605239265709025804299925103103321217007112614751710558224262457129529787960842708237904545156996902654409433534470689314969287033323693135988392074785123758189386591744698415144145679652;
            6'd51: xpb[108] = 1024'd8052924409200203593028606579902971815192792401662854478886311052996404297353146250662872989709153279520982544280060360939703717744398125294051418591447313257047088228606922205779346785397667577819493571357381165114073726521944332914578104567355935389861448130849831170991342651253122589199892929081529226407;
            6'd52: xpb[108] = 1024'd30104947655598691361307409584280086844947275470942933138338722947855001598002859906364804635231275280785871313130991758432866037064307559338963037096122346230777738412033351190964670305183011088988342042864097631435511400610376005259664089502972033013219106539828328297304089618245491603773777269644507257493;
            6'd53: xpb[108] = 1024'd52156970901997179129586212588657201874701758540223011797791134842713598898652573562066736280753397282050760081981923155926028356384216993383874655600797379204508388595459780176149993824968354600157190514370814097756949074698807677604750074438588130636576764948806825423616836585237860618347661610207485288579;
            6'd54: xpb[108] = 1024'd74208994148395666897865015593034316904456241609503090457243546737572196199302287217768667926275519283315648850832854553419190675704126427428786274105472412178239038778886209161335317344753698111326038985877530564078386748787239349949836059374204228259934423357785322549929583552230229632921545950770463319665;
            6'd55: xpb[108] = 1024'd96261017394794154666143818597411431934210724678783169116695958632430793499952000873470599571797641284580537619683785950912352995024035861473697892610147445151969688962312638146520640864539041622494887457384247030399824422875671022294922044309820325883292081766763819676242330519222598647495430291333441350751;
            6'd56: xpb[108] = 1024'd118313040641192642434422621601788546963965207748063247776148370527289390800601714529172531217319763285845426388534717348405515314343945295518609511114822478125700339145739067131705964384324385133663735928890963496721262096964102694640008029245436423506649740175742316802555077486214967662069314631896419381837;
            6'd57: xpb[108] = 1024'd16298368203466388803902497201351229249021263691607642307468927357171092763942289274859391648184210977667165749928155311319613792822634395008361004603166470165740314759594278779261048712592522923522386792010440116678338920831637594020115444497823071863187495170603755898761296379278703659524509145833802928592;
            6'd58: xpb[108] = 1024'd38350391449864876572181300205728344278775746760887720966921339252029690064592002930561323293706332978932054518779086708812776112142543829053272623107841503139470964943020707764446372232377866434691235263517156582999776594920069266365201429433439169486545153579582253025074043346271072674098393486396780959678;
            6'd59: xpb[108] = 1024'd60402414696263364340460103210105459308530229830167799626373751146888287365241716586263254939228454980196943287630018106305938431462453263098184241612516536113201615126447136749631695752163209945860083735023873049321214269008500938710287414369055267109902811988560750151386790313263441688672277826959758990764;
            6'd60: xpb[108] = 1024'd82454437942661852108738906214482574338284712899447878285826163041746884665891430241965186584750576981461832056480949503799100750782362697143095860117191569086932265309873565734817019271948553457028932206530589515642651943096932611055373399304671364733260470397539247277699537280255810703246162167522737021850;
            6'd61: xpb[108] = 1024'd104506461189060339877017709218859689368039195968727956945278574936605481966541143897667118230272698982726720825331880901292263070102272131188007478621866602060662915493299994720002342791733896968197780678037305981964089617185364283400459384240287462356618128806517744404012284247248179717820046508085715052936;
            6'd62: xpb[108] = 1024'd2491788751334086246497584818422371653095251912272351476599131766487183929881718643353978661137146674548460186725318864206361548580961230677758972110210594100702891107155206367557427120002034758056431541156782601921166441052899182780566799492674110713155883801379183500218503140311915715275241022023098599691;
            6'd63: xpb[108] = 1024'd24543811997732574014776387822799486682849734981552430136051543661345781230531432299055910306659268675813348955576250261699523867900870664722670590614885627074433541290581635352742750639787378269225280012663499068242604115141330855125652784428290208336513542210357680626531250107304284729849125362586076630777;
        endcase
    end

    always_comb begin
        case(flag[36][11:6])
            6'd0: xpb[109] = 1024'd0;
            6'd1: xpb[109] = 1024'd46595835244131061783055190827176601712604218050832508795503955556204378531181145954757841952181390677078237724427181659192686187220780098767582209119560660048164191474008064337928074159572721780394128484170215534564041789229762527470738769363906305959871200619336177752843997074296653744423009703149054661863;
            6'd2: xpb[109] = 1024'd93191670488262123566110381654353203425208436101665017591007911112408757062362291909515683904362781354156475448854363318385372374441560197535164418239121320096328382948016128675856148319145443560788256968340431069128083578459525054941477538727812611919742401238672355505687994148593307488846019406298109323726;
            6'd3: xpb[109] = 1024'd15720810048268443950366645076715372393114227026761842258380011603636240256234298954258454641886497721791563765824051542998994720821119961747586502342350939210801899852452975676153983287200959619872187844123406757327764517468390809447237738408489468612793698443891475228425463148961328216150339282821569501258;
            6'd4: xpb[109] = 1024'd62316645292399505733421835903891974105718445077594351053883967159840618787415444909016296594067888398869801490251233202191680908041900060515168711461911599258966091326461040014082057446773681400266316328293622291891806306698153336917976507772395774572664899063227652981269460223257981960573348985970624163121;
            6'd5: xpb[109] = 1024'd108912480536530567516477026731068575818322663128426859849387922716044997318596590863774138546249279075948039214678414861384367095262680159282750920581472259307130282800469104352010131606346403180660444812463837826455848095927915864388715277136302080532536099682563830734113457297554635704996358689119678824984;
            6'd6: xpb[109] = 1024'd31441620096536887900733290153430744786228454053523684516760023207272480512468597908516909283772995443583127531648103085997989441642239923495173004684701878421603799704905951352307966574401919239744375688246813514655529034936781618894475476816978937225587396887782950456850926297922656432300678565643139002516;
            6'd7: xpb[109] = 1024'd78037455340667949683788480980607346498832672104356193312263978763476859043649743863274751235954386120661365256075284745190675628863020022262755213804262538469767991178914015690236040733974641020138504172417029049219570824166544146365214246180885243185458597507119128209694923372219310176723688268792193664379;
            6'd8: xpb[109] = 1024'd566594900674270068044744402969515466738463029453017979636079254704342237521750908017521973478102488296453573044972969804297975242579786475177297907492157584241508083350862690533875702030157079222435048200004737419251763175409900870974445861562099878509894712338247932432392372587330904028008145315653841911;
            6'd9: xpb[109] = 1024'd47162430144805331851099935230146117179342681080285526775140034810908720768702896862775363925659493165374691297472154628996984162463359885242759507027052817632405699557358927028461949861602878859616563532370220271983293552405172428341713215225468405838381095331674425685276389446883984648451017848464708503774;
            6'd10: xpb[109] = 1024'd93758265388936393634155126057322718891946899131118035570643990367113099299884042817533205877840883842452929021899336288189670349684139984010341716146613477680569891031366991366390024021175600640010692016540435806547335341634934955812451984589374711798252295951010603438120386521180638392874027551613763165637;
            6'd11: xpb[109] = 1024'd16287404948942714018411389479684887859852690056214860238016090858340582493756049862275976615364600210088017338869024512803292696063699748222763800249843096795043407935803838366687858989231116699094622892323411494747016280643800710318212184270051568491303593156229723160857855521548659120178347428137223343169;
            6'd12: xpb[109] = 1024'd62883240193073775801466580306861489572456908107047369033520046414544961024937195817033818567545990887166255063296206171995978883284479846990346009369403756843207599409811902704615933148803838479488751376493627029311058069873563237788950953633957874451174793775565900913701852595845312864601357131286278005032;
            6'd13: xpb[109] = 1024'd109479075437204837584521771134038091285061126157879877829024001970749339556118341771791660519727381564244492787723387831188665070505259945757928218488964416891371790883819967042544007308376560259882879860663842563875099859103325765259689722997864180411045994394902078666545849670141966609024366834435332666895;
            6'd14: xpb[109] = 1024'd32008214997211157968778034556400260252966917082976702496396102461976822749990348816534431257251097931879581104693076055802287416884819709970350302592194036005845307788256814042841842276432076318966810736446818252074780798112191519765449922678541037104097291600121198389283318670509987336328686710958792844427;
            6'd15: xpb[109] = 1024'd78604050241342219751833225383576861965571135133809211291900058018181201281171494771292273209432488608957818829120257714994973604105599808737932511711754696054009499262264878380769916436004798099360939220617033786638822587341954047236188692042447343063968492219457376142127315744806641080751696414107847506290;
            6'd16: xpb[109] = 1024'd1133189801348540136089488805939030933476926058906035959272158509408684475043501816035043946956204976592907146089945939608595950485159572950354595814984315168483016166701725381067751404060314158444870096400009474838503526350819801741948891723124199757019789424676495864864784745174661808056016290631307683822;
            6'd17: xpb[109] = 1024'd47729025045479601919144679633115632646081144109738544754776114065613063006224647770792885899137595653671144870517127598801282137705939671717936804934544975216647207640709789718995825563633035938838998580570225009402545315580582329212687661087030505716890990044012673617708781819471315552479025993780362345685;
            6'd18: xpb[109] = 1024'd94324860289610663702199870460292234358685362160571053550280069621817441537405793725550727851318986330749382594944309257993968324926719770485519014054105635264811399114717854056923899723205757719233127064740440543966587104810344856683426430450936811676762190663348851370552778893767969296902035696929417007548;
            6'd19: xpb[109] = 1024'd16853999849616984086456133882654403326591153085667878217652170113044924731277800770293498588842702698384470911913997482607590671306279534697941098157335254379284916019154701057221734691261273778317057940523416232166268043819210611189186630131613668369813487868567971093290247894135990024206355573452877185080;
            6'd20: xpb[109] = 1024'd63449835093748045869511324709831005039195371136500387013156125669249303262458946725051340541024093375462708636341179141800276858527059633465523307276895914427449107493162765395149808850833995558711186424693631766730309833048973138659925399495519974329684688487904148846134244968432643768629365276601931846943;
            6'd21: xpb[109] = 1024'd110045670337879107652566515537007606751799589187332895808660081225453681793640092679809182493205484052540946360768360800992963045747839732233105516396456574475613298967170829733077883010406717339105314908863847301294351622278735666130664168859426280289555889107240326598978242042729297513052374979750986508806;
            6'd22: xpb[109] = 1024'd32574809897885428036822778959369775719705380112429720476032181716681164987512099724551953230729200420176034677738049025606585392127399496445527600499686193590086815871607676733375717978462233398189245784646822989494032561287601420636424368540103136982607186312459446321715711043097318240356694856274446686338;
            6'd23: xpb[109] = 1024'd79170645142016489819877969786546377432309598163262229271536137272885543518693245679309795182910591097254272402165230684799271579348179595213109809619246853638251007345615741071303792138034955178583374268817038524058074350517363948107163137904009442942478386931795624074559708117393971984779704559423501348201;
            6'd24: xpb[109] = 1024'd1699784702022810204134233208908546400215389088359053938908237764113026712565252724052565920434307464889360719134918909412893925727739359425531893722476472752724524250052588071601627106090471237667305144600014212257755289526229702612923337584686299635529684137014743797297177117761992712084024435946961525733;
            6'd25: xpb[109] = 1024'd48295619946153871987189424036085148112819607139191562734412193320317405243746398678810407872615698141967598443562100568605580112948519458193114102842037132800888715724060652409529701265663193018061433628770229746821797078755992230083662106948592605595400884756350921550141174192058646456507034139096016187596;
            6'd26: xpb[109] = 1024'd94891455190284933770244614863261749825423825190024071529916148876521783774927544633568249824797088819045836167989282227798266300169299556960696311961597792849052907198068716747457775425235914798455562112940445281385838867985754757554400876312498911555272085375687099302985171266355300200930043842245070849459;
            6'd27: xpb[109] = 1024'd17420594750291254154500878285623918793329616115120896197288249367749266968799551678311020562320805186680924484958970452411888646548859321173118396064827411963526424102505563747755610393291430857539492988723420969585519806994620512060161075993175768248323382580906219025722640266723320928234363718768531026991;
            6'd28: xpb[109] = 1024'd64016429994422315937556069112800520505933834165953404992792204923953645499980697633068862514502195863759162209386152111604574833769639419940700605184388072011690615576513628085683684552864152637933621472893636504149561596224383039530899845357082074208194583200242396778566637341019974672657373421917585688854;
            6'd29: xpb[109] = 1024'd110612265238553377720611259939977122218538052216785913788296160480158024031161843587826704466683586540837399933813333770797261020990419518708282814303948732059854807050521692423611758712436874418327749957063852038713603385454145567001638614720988380168065783819578574531410634415316628417080383125066640350717;
            6'd30: xpb[109] = 1024'd33141404798559698104867523362339291186443843141882738455668260971385507225033850632569475204207302908472488250783021995410883367369979282920704898407178351174328323954958539423909593680492390477411680832846827726913284324463011321507398814401665236861117081024797694254148103415684649144384703001590100528249;
            6'd31: xpb[109] = 1024'd79737240042690759887922714189515892899048061192715247251172216527589885756214996587327317156388693585550725975210203654603569554590759381688287107526739011222492515428966603761837667840065112257805809317017043261477326113692773848978137583765571542820988281644133872006992100489981302888807712704739155190112;
            6'd32: xpb[109] = 1024'd2266379602697080272178977611878061866953852117812071918544317018817368950087003632070087893912409953185814292179891879217191900970319145900709191629968630336966032333403450762135502808120628316889740192800018949677007052701639603483897783446248399514039578849352991729729569490349323616112032581262615367644;
            6'd33: xpb[109] = 1024'd48862214846828142055234168439054663579558070168644580714048272575021747481268149586827929846093800630264052016607073538409878088191099244668291400749529290385130223807411515100063576967693350097283868676970234484241048841931402130954636552810154705473910779468689169482573566564645977360535042284411670029507;
            6'd34: xpb[109] = 1024'd95458050090959203838289359266231265292162288219477089509552228131226126012449295541585771798275191307342289741034255197602564275411879343435873609869089950433294415281419579437991651127266071877677997161140450018805090631161164658425375322174061011433781980088025347235417563638942631104958051987560724691370;
            6'd35: xpb[109] = 1024'd17987189650965524222545622688593434260068079144573914176924328622453609206321302586328542535798907674977378058003943422216186621791439107648295693972319569547767932185856426438289486095321587936761928036923425707004771570170030412931135521854737868126833277293244466958155032639310651832262371864084184868902;
            6'd36: xpb[109] = 1024'd64583024895096586005600813515770035972672297195406422972428284178657987737502448541086384487980298352055615782431125081408872809012219206415877903091880229595932123659864490776217560254894309717156056521093641241568813359399792940401874291218644174086704477912580644710999029713607305576685381567233239530765;
            6'd37: xpb[109] = 1024'd111178860139227647788656004342946637685276515246238931767932239734862366268683594495844226440161689029133853506858306740601558996232999305183460112211440889644096315133872555114145634414467031497550185005263856776132855148629555467872613060582550480046575678531916822463843026787903959321108391270382294192628;
            6'd38: xpb[109] = 1024'd33707999699233968172912267765308806653182306171335756435304340226089849462555601540586997177685405396768941823827994965215181342612559069395882196314670508758569832038309402114443469382522547556634115881046832464332536087638421222378373260263227336739626975737135942186580495788271980048412711146905754370160;
            6'd39: xpb[109] = 1024'd80303834943365029955967458592485408365786524222168265230808295782294227993736747495344839129866796073847179548255176624407867529833339168163464405434231168806734023512317466452371543542095269337028244365217047998896577876868183749849112029627133642699498176356472119939424492862568633792835720850054809032023;
            6'd40: xpb[109] = 1024'd2832974503371350340223722014847577333692315147265089898180396273521711187608754540087609867390512441482267865224864849021489876212898932375886489537460787921207540416754313452669378510150785396112175241000023687096258815877049504354872229307810499392549473561691239662161961862936654520140040726578269209555;
            6'd41: xpb[109] = 1024'd49428809747502412123278912842024179046296533198097598693684351829726089718789900494845451819571903118560505589652046508214176063433679031143468698657021447969371731890762377790597452669723507176506303725170239221660300605106812031825610998671716805352420674181027417415005958937233308264563050429727323871418;
            6'd42: xpb[109] = 1024'd96024644991633473906334103669200780758900751248930107489188307385930468249971046449603293771753293795638743314079228167406862250654459129911050907776582108017535923364770442128525526829296228956900432209340454756224342394336574559296349768035623111312291874800363595167849956011529962008986060132876378533281;
            6'd43: xpb[109] = 1024'd18553784551639794290590367091562949726806542174026932156560407877157951443843053494346064509277010163273831631048916392020484597034018894123472991879811727132009440269207289128823361797351745015984363085123430444424023333345440313802109967716299968005343172005582714890587425011897982736290380009399838710813;
            6'd44: xpb[109] = 1024'd65149619795770856073645557918739551439410760224859440952064363433362329975024199449103906461458400840352069355476098051213170784254798992891055200999372387180173631743215353466751435956924466796378491569293645978988065122575202841272848737080206273965214372624918892643431422086194636480713389712548893372676;
            6'd45: xpb[109] = 1024'd111745455039901917856700748745916153152014978275691949747568318989566708506205345403861748413639791517430307079903279710405856971475579091658637410118933047228337823217223417804679510116497188576772620053463861513552106911804965368743587506444112579925085573244255070396275419160491290225136399415697948034539;
            6'd46: xpb[109] = 1024'd34274594599908238240957012168278322119920769200788774414940419480794191700077352448604519151163507885065395396872967935019479317855138855871059494222162666342811340121660264804977345084552704635856550929246837201751787850813831123249347706124789436618136870449474190119012888160859310952440719292221408212071;
            6'd47: xpb[109] = 1024'd80870429844039300024012202995454923832524987251621283210444375036998570231258498403362361103344898562143633121300149594212165505075918954638641703341723326390975531595668329142905419244125426416250679413417052736315829640043593650720086475488695742578008071068810367871856885235155964696863728995370462873934;
            6'd48: xpb[109] = 1024'd3399569404045620408268466417817092800430778176718107877816475528226053425130505448105131840868614929778721438269837818825787851455478718851063787444952945505449048500105176143203254212180942475334610289200028424515510579052459405225846675169372599271059368274029487594594354235523985424168048871893923051466;
            6'd49: xpb[109] = 1024'd49995404648176682191323657244993694513034996227550616673320431084430431956311651402862973793050005606856959162697019478018474038676258817618645996564513605553613239974113240481131328371753664255728738773370243959079552368282221932696585444533278905230930568893365665347438351309820639168591058575042977713329;
            6'd50: xpb[109] = 1024'd96591239892307743974378848072170296225639214278383125468824386640634810487492797357620815745231396283935196887124201137211160225897038916386228205684074265601777431448121304819059402531326386036122867257540459493643594157511984460167324213897185211190801769512701843100282348384117292913014068278192032375192;
            6'd51: xpb[109] = 1024'd19120379452314064358635111494532465193545005203479950136196487131862293681364804402363586482755112651570285204093889361824782572276598680598650289787303884716250948352558151819357237499381902095206798133323435181843275096520850214673084413577862067883853066717920962823019817384485313640318388154715492552724;
            6'd52: xpb[109] = 1024'd65716214696445126141690302321709066906149223254312458931700442688066672212545950357121428434936503328648522928521071021017468759497378779366232498906864544764415139826566216157285311658954623875600926617493650716407316885750612742143823182941768373843724267337257140575863814458781967384741397857864547214587;
            6'd53: xpb[109] = 1024'd112312049940576187924745493148885668618753441305144967727204398244271050743727096311879270387117894005726760652948252680210154946718158878133814708026425204812579331300574280495213385818527345655995055101663866250971358674980375269614561952305674679803595467956593318328707811533078621129164407561013601876450;
            6'd54: xpb[109] = 1024'd34841189500582508309001756571247837586659232230241792394576498735498533937599103356622041124641610373361848969917940904823777293097718642346236792129654823927052848205011127495511220786582861715078985977446841939171039613989241024120322151986351536496646765161812438051445280533446641856468727437537062053982;
            6'd55: xpb[109] = 1024'd81437024744713570092056947398424439299263450281074301190080454291702912468780249311379883076823001050440086694345122564016463480318498741113819001249215483975217039679019191833439294946155583495473114461617057473735081403219003551591060921350257842456517965781148615804289277607743295600891737140686116715845;
            6'd56: xpb[109] = 1024'd3966164304719890476313210820786608267169241206171125857452554782930395662652256356122653814346717418075175011314810788630085826698058505326241085352445103089690556583456038833737129914211099554557045337400033161934762342227869306096821121030934699149569262986367735527026746608111316328196057017209576893377;
            6'd57: xpb[109] = 1024'd50561999548850952259368401647963209979773459257003634652956510339134774193833402310880495766528108095153412735741992447822772013918838604093823294472005763137854748057464103171665204073783821334951173821570248696498804131457631833567559890394841005109440463605703913279870743682407970072619066720358631555240;
            6'd58: xpb[109] = 1024'd97157834792982014042423592475139811692377677307836143448460465895339152725014548265638337718709498772231650460169174107015458201139618702861405503591566423186018939531472167509593278233356543115345302305740464231062845920687394361038298659758747311069311664225040091032714740756704623817042076423507686217103;
            6'd59: xpb[109] = 1024'd19686974352988334426679855897501980660283468232932968115832566386566635918886555310381108456233215139866738777138862331629080547519178467073827587694796042300492456435909014509891113201412059174429233181523439919262526859696260115544058859439424167762362961430259210755452209757072644544346396300031146394635;
            6'd60: xpb[109] = 1024'd66282809597119396209735046724678582372887686283765476911336521942771014450067701265138950408414605816944976501566043990821766734739958565841409796814356702348656647909917078847819187360984780954823361665693655453826568648926022643014797628803330473722234162049595388508296206831369298288769406003180201056498;
            6'd61: xpb[109] = 1024'd112878644841250457992790237551855184085491904334597985706840477498975392981248847219896792360595996494023214225993225650014452921960738664608992005933917362396820839383925143185747261520557502735217490149863870988390610438155785170485536398167236779682105362668931566261140203905665952033192415706329255718361;
            6'd62: xpb[109] = 1024'd35407784401256778377046500974217353053397695259694810374212577990202876175120854264639563098119712861658302542962913874628075268340298428821414090037146981511294356288361990186045096488613018794301421025646846676590291377164650924991296597847913636375156659874150685983877672906033972760496735582852715895893;
            6'd63: xpb[109] = 1024'd82003619645387840160101691801393954766001913310527319169716533546407254706302000219397405050301103538736540267390095533820761455561078527588996299156707641559458547762370054523973170648185740574695549509817062211154333166394413452462035367211819942335027860493486863736721669980330626504919745286001770557756;
        endcase
    end

    always_comb begin
        case(flag[36][16:12])
            5'd0: xpb[110] = 1024'd0;
            5'd1: xpb[110] = 1024'd4532759205394160544357955223756123733907704235624143837088634037634737900174007264140175787824819906371628584359783758434383801940638291801418383259937260673932064666806901524271005616241256633779480385600037899354014105403279206967795566892496799028079157698705983459459138980698647232224065162525230735288;
            5'd2: xpb[110] = 1024'd9065518410788321088715910447512247467815408471248287674177268075269475800348014528280351575649639812743257168719567516868767603881276583602836766519874521347864129333613803048542011232482513267558960771200075798708028210806558413935591133784993598056158315397411966918918277961397294464448130325050461470576;
            5'd3: xpb[110] = 1024'd13598277616182481633073865671268371201723112706872431511265902112904213700522021792420527363474459719114885753079351275303151405821914875404255149779811782021796194000420704572813016848723769901338441156800113698062042316209837620903386700677490397084237473096117950378377416942095941696672195487575692205864;
            5'd4: xpb[110] = 1024'd18131036821576642177431820895024494935630816942496575348354536150538951600696029056560703151299279625486514337439135033737535207762553167205673533039749042695728258667227606097084022464965026535117921542400151597416056421613116827871182267569987196112316630794823933837836555922794588928896260650100922941152;
            5'd5: xpb[110] = 1024'd22663796026970802721789776118780618669538521178120719185443170188173689500870036320700878939124099531858142921798918792171919009703191459007091916299686303369660323334034507621355028081206283168897401928000189496770070527016396034838977834462483995140395788493529917297295694903493236161120325812626153676440;
            5'd6: xpb[110] = 1024'd27196555232364963266147731342536742403446225413744863022531804225808427401044043584841054726948919438229771506158702550606302811643829750808510299559623564043592388000841409145626033697447539802676882313600227396124084632419675241806773401354980794168474946192235900756754833884191883393344390975151384411728;
            5'd7: xpb[110] = 1024'd31729314437759123810505686566292866137353929649369006859620438263443165301218050848981230514773739344601400090518486309040686613584468042609928682819560824717524452667648310669897039313688796436456362699200265295478098737822954448774568968247477593196554103890941884216213972864890530625568456137676615147016;
            5'd8: xpb[110] = 1024'd36262073643153284354863641790048989871261633884993150696709072301077903201392058113121406302598559250973028674878270067475070415525106334411347066079498085391456517334455212194168044929930053070235843084800303194832112843226233655742364535139974392224633261589647867675673111845589177857792521300201845882304;
            5'd9: xpb[110] = 1024'd40794832848547444899221597013805113605169338120617294533797706338712641101566065377261582090423379157344657259238053825909454217465744626212765449339435346065388582001262113718439050546171309704015323470400341094186126948629512862710160102032471191252712419288353851135132250826287825090016586462727076617592;
            5'd10: xpb[110] = 1024'd45327592053941605443579552237561237339077042356241438370886340376347379001740072641401757878248199063716285843597837584343838019406382918014183832599372606739320646668069015242710056162412566337794803856000378993540141054032792069677955668924967990280791576987059834594591389806986472322240651625252307352880;
            5'd11: xpb[110] = 1024'd49860351259335765987937507461317361072984746591865582207974974413982116901914079905541933666073018970087914427957621342778221821347021209815602215859309867413252711334875916766981061778653822971574284241600416892894155159436071276645751235817464789308870734685765818054050528787685119554464716787777538088168;
            5'd12: xpb[110] = 1024'd54393110464729926532295462685073484806892450827489726045063608451616854802088087169682109453897838876459543012317405101212605623287659501617020599119247128087184776001682818291252067394895079605353764627200454792248169264839350483613546802709961588336949892384471801513509667768383766786688781950302768823456;
            5'd13: xpb[110] = 1024'd58925869670124087076653417908829608540800155063113869882152242489251592702262094433822285241722658782831171596677188859646989425228297793418438982379184388761116840668489719815523073011136336239133245012800492691602183370242629690581342369602458387365029050083177784972968806749082414018912847112827999558744;
            5'd14: xpb[110] = 1024'd63458628875518247621011373132585732274707859298738013719240876526886330602436101697962461029547478689202800181036972618081373227168936085219857365639121649435048905335296621339794078627377592872912725398400530590956197475645908897549137936494955186393108207781883768432427945729781061251136912275353230294032;
            5'd15: xpb[110] = 1024'd67991388080912408165369328356341856008615563534362157556329510564521068502610108962102636817372298595574428765396756376515757029109574377021275748899058910108980970002103522864065084243618849506692205784000568490310211581049188104516933503387451985421187365480589751891887084710479708483360977437878461029320;
            5'd16: xpb[110] = 1024'd72524147286306568709727283580097979742523267769986301393418144602155806402784116226242812605197118501946057349756540134950140831050212668822694132158996170782913034668910424388336089859860106140471686169600606389664225686452467311484729070279948784449266523179295735351346223691178355715585042600403691764608;
            5'd17: xpb[110] = 1024'd77056906491700729254085238803854103476430972005610445230506778639790544302958123490382988393021938408317685934116323893384524632990850960624112515418933431456845099335717325912607095476101362774251166555200644289018239791855746518452524637172445583477345680878001718810805362671877002947809107762928922499896;
            5'd18: xpb[110] = 1024'd81589665697094889798443194027610227210338676241234589067595412677425282203132130754523164180846758314689314518476107651818908434931489252425530898678870692130777164002524227436878101092342619408030646940800682188372253897259025725420320204064942382505424838576707702270264501652575650180033172925454153235184;
            5'd19: xpb[110] = 1024'd86122424902489050342801149251366350944246380476858732904684046715060020103306138018663339968671578221060943102835891410253292236872127544226949281938807952804709228669331128961149106708583876041810127326400720087726268002662304932388115770957439181533503996275413685729723640633274297412257238087979383970472;
            5'd20: xpb[110] = 1024'd90655184107883210887159104475122474678154084712482876741772680752694758003480145282803515756496398127432571687195675168687676038812765836028367665198745213478641293336138030485420112324825132675589607712000757987080282108065584139355911337849935980561583153974119669189182779613972944644481303250504614705760;
            5'd21: xpb[110] = 1024'd95187943313277371431517059698878598412061788948107020578861314790329495903654152546943691544321218033804200271555458927122059840753404127829786048458682474152573358002944932009691117941066389309369088097600795886434296213468863346323706904742432779589662311672825652648641918594671591876705368413029845441048;
            5'd22: xpb[110] = 1024'd99720702518671531975875014922634722145969493183731164415949948827964233803828159811083867332146037940175828855915242685556443642694042419631204431718619734826505422669751833533962123557307645943148568483200833785788310318872142553291502471634929578617741469371531636108101057575370239108929433575555076176336;
            5'd23: xpb[110] = 1024'd104253461724065692520232970146390845879877197419355308253038582865598971704002167075224043119970857846547457440275026443990827444634680711432622814978556995500437487336558735058233129173548902576928048868800871685142324424275421760259298038527426377645820627070237619567560196556068886341153498738080306911624;
            5'd24: xpb[110] = 1024'd108786220929459853064590925370146969613784901654979452090127216903233709604176174339364218907795677752919086024634810202425211246575319003234041198238494256174369552003365636582504134789790159210707529254400909584496338529678700967227093605419923176673899784768943603027019335536767533573377563900605537646912;
            5'd25: xpb[110] = 1024'd113318980134854013608948880593903093347692605890603595927215850940868447504350181603504394695620497659290714608994593960859595048515957295035459581498431516848301616670172538106775140406031415844487009640000947483850352635081980174194889172312419975701978942467649586486478474517466180805601629063130768382200;
            5'd26: xpb[110] = 1024'd117851739340248174153306835817659217081600310126227739764304484978503185404524188867644570483445317565662343193354377719293978850456595586836877964758368777522233681336979439631046146022272672478266490025600985383204366740485259381162684739204916774730058100166355569945937613498164828037825694225655999117488;
            5'd27: xpb[110] = 1024'd122384498545642334697664791041415340815508014361851883601393119016137923304698196131784746271270137472033971777714161477728362652397233878638296348018306038196165746003786341155317151638513929112045970411201023282558380845888538588130480306097413573758137257865061553405396752478863475270049759388181229852776;
            5'd28: xpb[110] = 1024'd2850562066911753843223818860357031804717291471740343310349897988795765867563064485909850844437283068962450954616451801583682613496651835884554606261912257936407136101022025341957918063237980024515253188413821335548034101070921022133297303306680923519396512149650478834749363385633489485155134724080866103733;
            5'd29: xpb[110] = 1024'd7383321272305914387581774084113155538624995707364487147438532026430503767737071750050026632262102975334079538976235560018066415437290127685972989521849518610339200767828926866228923679479236658294733574013859234902048206474200229101092870199177722547475669848356462294208502366332136717379199886606096839021;
            5'd30: xpb[110] = 1024'd11916080477700074931939729307869279272532699942988630984527166064065241667911079014190202420086922881705708123336019318452450217377928419487391372781786779284271265434635828390499929295720493292074213959613897134256062311877479436068888437091674521575554827547062445753667641347030783949603265049131327574309;
            5'd31: xpb[110] = 1024'd16448839683094235476297684531625403006440404178612774821615800101699979568085086278330378207911742788077336707695803076886834019318566711288809756041724039958203330101442729914770934911961749925853694345213935033610076417280758643036684003984171320603633985245768429213126780327729431181827330211656558309597;
        endcase
    end

    always_comb begin
        case(flag[37][5:0])
            6'd0: xpb[111] = 1024'd0;
            6'd1: xpb[111] = 1024'd72524147286306568709727283580097979742523267769986301393418144602155806402784116226242812605197118501946057349756540134950140831050212668822694132158996170782913034668910424388336089859860106140471686169600606389664225686452467311484729070279948784449266523179295735351346223691178355715585042600403691764608;
            6'd2: xpb[111] = 1024'd20981598888488396020655639755381526740348108414236918658704434139334717468259093542470553995736562694448965292055586835321217821259205003090228139301661300632135394768249631439041940528203006559633174730813972932964090522684037850004479570876668119631713142944474412672585919308428078414051395374181789044885;
            6'd3: xpb[111] = 1024'd93505746174794964730382923335479506482871376184223220052122578741490523871043209768713366600933681196395022641812126970271358652309417671912922271460657471415048429437160055827378030388063112700104860900414579322628316209136505161489208641156616904080979666123770148023932142999606434129636437974585480809493;
            6'd4: xpb[111] = 1024'd41963197776976792041311279510763053480696216828473837317408868278669434936518187084941107991473125388897930584111173670642435642518410006180456278603322601264270789536499262878083881056406013119266349461627945865928181045368075700008959141753336239263426285888948825345171838616856156828102790748363578089770;
            6'd5: xpb[111] = 1024'd114487345063283360751038563090861033223219484598460138710827012880825241339302303311183920596670243890843987933867713805592576473568622675003150410762318772047183824205409687266419970916266119259738035631228552255592406731820543011493688212033285023712692809068244560696518062308034512543687833348767269854378;
            6'd6: xpb[111] = 1024'd62944796665465188061966919266144580221044325242710755976113302418004152404777280627411661987209688083346895876166760505963653463777615009270684417904983901896406184304748894317125821584609019678899524192441918798892271568052113550013438712630004358895139428833423238017757757925284235242154186122545367134655;
            6'd7: xpb[111] = 1024'd11402248267647015372895275441428127218869165886961373241399591955183063470252257943639403377749132275849803818465807206334730453986607343538218425047649031745628544404088101367831672252951920098061012753655285342192136404283684088533189213226723694077586048598601915338997453542533957940620538896323464414932;
            6'd8: xpb[111] = 1024'd83926395553953584082622559021526106961392433656947674634817736557338869873036374169882215982946250777795861168222347341284871285036820012360912557206645202528541579072998525756167762112812026238532698923255891731856362090736151400017918283506672478526852571777897650690343677233712313656205581496727156179540;
            6'd9: xpb[111] = 1024'd32383847156135411393550915196809653959217274301198291900104026094517780938511351486109957373485694970298769110521394041655948275245812346628446564349310332377763939172337732806873612781154926657694187484469258275156226926967721938537668784103391813709299191543076328011583372850962036354671934270505253459817;
            6'd10: xpb[111] = 1024'd104907994442441980103278198776907633701740542071184593293522170696673587341295467712352769978682813472244826460277934176606089106296025015451140696508306503160676973841248157195209702641015032798165873654069864664820452613420189250022397854383340598158565714722372063362929596542140392070256976870908945224425;
            6'd11: xpb[111] = 1024'd53365446044623807414206554952191180699565382715435210558808460233852498406770445028580511369222257664747734402576980876977166096505017349718674703650971633009899333940587364245915553309357933217327362215283231208120317449651759788542148354980059933341012334487550740684169292159390114768723329644687042504702;
            6'd12: xpb[111] = 1024'd1822897646805634725134911127474727697390223359685827824094749771031409472245422344808252759761701857250642344876027577348243086714009683986208710793636762859121694039926571296621403977700833636488850776496597751420182285883330327061898855576779268523458954252729418005408987776639837467189682418465139784979;
            6'd13: xpb[111] = 1024'd74347044933112203434862194707572707439913491129672129217512894373187215875029538571051065364958820359196699694632567712298383917764222352808902842952632933642034728708836995684957493837560939776960536946097204141084407972335797638546627925856728052972725477432025153356755211467818193182774725018868831549587;
            6'd14: xpb[111] = 1024'd22804496535294030745790550882856254437738331773922746482799183910366126940504515887278806755498264551699607636931614412669460907973214687076436850095298063491257088808176202735663344505903840196122025507310570684384272808567368177066378426453447388155172097197203830677994907085067915881241077792646928829864;
            6'd15: xpb[111] = 1024'd95328643821600599455517834462954234180261599543909047876217328512521933343288632113521619360695383053645664986688154547619601739023427355899130982254294234274170123477086627123999434365763946336593711676911177074048498495019835488551107496733396172604438620376499566029341130776246271596826120393050620594472;
            6'd16: xpb[111] = 1024'd43786095423782426766446190638237781178086440188159665141503618049700844408763609429749360751234827246148572928987201247990678729232419690166664989396959364123392483576425834174705285034106846755755200238124543617348363331251406027070857997330115507786885240141678243350580826393495994295292473166828717874749;
            6'd17: xpb[111] = 1024'd116310242710088995476173474218335760920609707958145966534921762651856650811547725655992173356431945748094630278743741382940819560282632358989359121555955534906305518245336258563041374893966952896226886407725150007012589017703873338555587067610064292236151763320973978701927050084674350010877515767232409639357;
            6'd18: xpb[111] = 1024'd64767694312270822787101830393619307918434548602396583800208052189035561877022702972219914746971389940597538221042788083311896550491624693256893128698620664755527878344675465613747225562309853315388374968938516550312453853935443877075337568206783627418598383086152656023166745701924072709343868541010506919634;
            6'd19: xpb[111] = 1024'd13225145914452650098030186568902854916259389246647201065494341726214472942497680288447656137510834133100446163341834783682973540700617027524427135841285794604750238444014672664453076230652753734549863530151883093612318690167014415595088068803502962601045002851331333344406441319173795407810221314788604199911;
            6'd20: xpb[111] = 1024'd85749293200759218807757470149000834658782657016633502458912486328370279345281796514690468742707952635046503513098374918633114371750829696347121268000281965387663273112925097052789166090512859875021549699752489483276544376619481727079817139083451747050311526030627068695752665010352151123395263915192295964519;
            6'd21: xpb[111] = 1024'd34206744802941046118685826324284381656607497660884119724198775865549190410756773830918210133247396827549411455397421619004191361959822030614655275142947095236885633212264304103495016758855760294183038260965856026576409212851052265599567639680171082232758145795805746016992360627601873821861616688970393244796;
            6'd22: xpb[111] = 1024'd106730892089247614828413109904382361399130765430870421117616920467704996813540890057161022738444515329495468805153961753954332193010034699437349407301943266019798667881174728491831106618715866434654724430566462416240634899303519577084296709960119866682024668975101481368338584318780229537446659289374085009404;
            6'd23: xpb[111] = 1024'd55188343691429442139341466079665908396955606075121038382903210004883907879015867373388764128983959521998376747453008454325409183219027033704883414444608395869021027980513935542536957287058766853816212991779828959540499735535090115604047210556839201864471288740280158689578279936029952235913012063152182289681;
            6'd24: xpb[111] = 1024'd3645795293611269450269822254949455394780446719371655648189499542062818944490844689616505519523403714501284689752055154696486173428019367972417421587273525718243388079853142593242807955401667272977701552993195502840364571766660654123797711153558537046917908505458836010817975553279674934379364836930279569958;
            6'd25: xpb[111] = 1024'd76169942579917838159997105835047435137303714489357957041607644144218625347274960915859318124720522216447342039508595289646627004478232036795111553746269696501156422748763566981578897815261773413449387722593801892504590258219127965608526781433507321496184431684754571362164199244458030649964407437333971334566;
            6'd26: xpb[111] = 1024'd24627394182099665470925462010330982135128555133608574306893933681397536412749938232087059515259966408950249981807641990017703994687224371062645560888934826350378782848102774032284748483604673832610876283807168435804455094450698504128277282030226656678631051449933248683403894861707753348430760211112068614843;
            6'd27: xpb[111] = 1024'd97151541468406234180652745590428961877651822903594875700312078283553342815534054458329872120457084910896307331564182124967844825737437039885339693047930997133291817517013198420620838343464779973082562453407774825468680780903165815613006352310175441127897574629228984034750118552886109064015802811515760379451;
            6'd28: xpb[111] = 1024'd45608993070588061491581101765712508875476663547845492965598367820732253881009031774557613510996529103399215273863228825338921815946429374152873700190596126982514177616352405471326689011807680392244051014621141368768545617134736354132756852906894776310344194394407661355989814170135831762482155585293857659728;
            6'd29: xpb[111] = 1024'd118133140356894630201308385345810488617999931317831794359016512422888060283793148000800426116193647605345272623619768960289062646996642042975567832349592297765427212285262829859662778871667786532715737184221747758432771303587203665617485923186843560759610717573703396707336037861314187478067198185697549424336;
            6'd30: xpb[111] = 1024'd66590591959076457512236741521094035615824771962082411624302801960066971349268125317028167506733091797848180565918815660660139637205634377243101839492257427614649572384602036910368629540010686951877225745435114301732636139818774204137236423783562895942057337338882074028575733478563910176533550959475646704613;
            6'd31: xpb[111] = 1024'd15048043561258284823165097696377582613649612606333028889589091497245882414743102633255908897272535990351088508217862361031216627414626711510635846634922557463871932483941243961074480208353587371038714306648480845032500976050344742656986924380282231124503957104060751349815429095813632874999903733253743984890;
            6'd32: xpb[111] = 1024'd87572190847564853532892381276475562356172880376319330283007236099401688817527218859498721502469654492297145857974402495981357458464839380333329978793918728246784967152851668349410570068213693511510400476249087234696726662502812054141715994660231015573770480283356486701161652786991988590584946333657435749498;
            6'd33: xpb[111] = 1024'd36029642449746680843820737451759109353997721020569947548293525636580599883002196175726462893009098684800053800273449196352434448673831714600863985936583858096007327252190875400116420736556593930671889037462453777996591498734382592661466495256950350756217100048535164022401348404241711289051299107435533029775;
            6'd34: xpb[111] = 1024'd108553789736053249553548021031857089096520988790556248941711670238736406285786312401969275498206217186746111150029989331302575279724044383423558118095580028878920361921101299788452510596416700071143575207063060167660817185186849904146195565536899135205483623227830899373747572095420067004636341707839224794383;
            6'd35: xpb[111] = 1024'd57011241338235076864476377207140636094345829434806866206997959775915317351261289718197016888745661379249019092329036031673652269933036717691092125238245158728142722020440506839158361264759600490305063768276426710960682021418420442665946066133618470387930242993009576694987267712669789703102694481617322074660;
            6'd36: xpb[111] = 1024'd5468692940416904175404733382424183092170670079057483472284249313094228416736267034424758279285105571751927034628082732044729260142029051958626132380910288577365082119779713889864211933102500909466552329489793254260546857649990981185696566730337805570376862758188254016226963329919512401569047255395419354937;
            6'd37: xpb[111] = 1024'd77992840226723472885132016962522162834693937849043784865702393915250034819520383260667570884482224073697984384384622866994870091192241720781320264539906459360278116788690138278200301792962607049938238499090399643924772544102458292670425637010286590019643385937483989367573187021097868117154089855799111119545;
            6'd38: xpb[111] = 1024'd26450291828905300196060373137805709832518778493294402130988683452428945884995360576895312275021668266200892326683669567365947081401234055048854271682571589209500476888029345328906152461305507469099727060303766187224637380334028831190176137607005925202090005702662666688812882638347590815620442629577208399822;
            6'd39: xpb[111] = 1024'd98974439115211868905787656717903689575042046263280703524406828054584752287779476803138124880218786768146949676440209702316087912451446723871548403841567759992413511556939769717242242321165613609571413229904372576888863066786496142674905207886954709651356528881958402040159106329525946531205485229980900164430;
            6'd40: xpb[111] = 1024'd47431890717393696216716012893187236572866886907531320789693117591763663353254454119365866270758230960649857618739256402687164902660439058139082410984232889841635871656278976767948092989508514028732901791117739120188727903018066681194655708483674044833803148647137079361398801946775669229671838003758997444707;
            6'd41: xpb[111] = 1024'd119956038003700264926443296473285216315390154677517622183111262193919469756038570345608678875955349462595914968495796537637305733710651726961776543143229060624548906325189401156284182849368620169204587960718345509852953589470533992679384778763622829283069671826432814712745025637954024945256880604162689209315;
            6'd42: xpb[111] = 1024'd68413489605882092237371652648568763313214995321768239448397551731098380821513547661836420266494793655098822910794843238008382723919644061229310550285894190473771266424528608206990033517711520588366076521931712053152818425702104531199135279360342164465516291591611492033984721255203747643723233377940786489592;
            6'd43: xpb[111] = 1024'd16870941208063919548300008823852310311039835966018856713683841268277291886988524978064161657034237847601730853093889938379459714128636395496844557428559320322993626523867815257695884186054421007527565083145078596452683261933675069718885779957061499647962911356790169355224416872453470342189586151718883769869;
            6'd44: xpb[111] = 1024'd89395088494370488258027292403950290053563103736005158107101985870433098289772641204306974262231356349547788202850430073329600545178849064319538689587555491105906661192778239646031974045914527147999251252745684986116908948386142381203614850237010284097229434536085904706570640563631826057774628752122575534477;
            6'd45: xpb[111] = 1024'd37852540096552315568955648579233837051387944380255775372388275407612009355247618520534715652770800542050696145149476773700677535387841398587072696730220620955129021292117446696737824714257427567160739813959051529416773784617712919723365350833729619279676054301264582027810336180881548756240981525900672814754;
            6'd46: xpb[111] = 1024'd110376687382858884278682932159331816793911212150242076765806420009767815758031734746777528257967919043996753494906016908650818366438054067409766828889216791738042055961027871085073914574117533707632425983559657919080999471070180231208094421113678403728942577480560317379156559872059904471826024126304364579362;
            6'd47: xpb[111] = 1024'd58834138985040711589611288334615363791736052794492694031092709546946726823506712063005269648507363236499661437205063609021895356647046401677300836031881921587264416060367078135779765242460434126793914544773024462380864307301750769727844921710397738911389197245738994700396255489309627170292376900082461859639;
            6'd48: xpb[111] = 1024'd7291590587222538900539644509898910789560893438743311296378999084125637888981689379233011039046807429002569379504110309392972346856038735944834843174547051436486776159706285186485615910803334545955403105986391005680729143533321308247595422307117074093835817010917672021635951106559349868758729673860559139916;
            6'd49: xpb[111] = 1024'd79815737873529107610266928089996890532084161208729612689797143686281444291765805605475823644243925930948626729260650444343113177906251404767528975333543222219399810828616709574821705770663440686427089275586997395344954829985788619732324492587065858543102340190213407372982174797737705584343772274264250904524;
            6'd50: xpb[111] = 1024'd28273189475710934921195284265280437529909001852980229955083433223460355357240782921703565034783370123451534671559697144714190168115243739035062982476208352068622170927955916625527556439006341105588577836800363938644819666217359158252074993183785193725548959955392084694221870414987428282810125048042348184801;
            6'd51: xpb[111] = 1024'd100797336762017503630922567845378417272432269622966531348501577825616161760024899147946377639980488625397592021316237279664330999165456407857757114635204522851535205596866341013863646298866447246060264006400970328309045352669826469736804063463733978174815483134687820045568094106165783998395167648446039949409;
            6'd52: xpb[111] = 1024'd49254788364199330941850924020661964270257110267217148613787867362795072825499876464174119030519932817900499963615283980035407989374448742125291121777869652700757565696205548064569496967209347665221752567614336871608910188901397008256554564060453313357262102899866497366807789723415506696861520422224137229686;
            6'd53: xpb[111] = 1024'd121778935650505899651578207600759944012780378037203450007206011964950879228283992690416931635717051319846557313371824114985548820424661410947985253936865823483670600365115972452905586827069453805693438737214943261273135875353864319741283634340402097806528626079162232718154013414593862412446563022627828994294;
            6'd54: xpb[111] = 1024'd70236387252687726962506563776043491010605218681454067272492301502129790293758970006644673026256495512349465255670870815356625810633653745215519261079530953332892960464455179503611437495412354224854927298428309804573000711585434858261034134937121432988975245844340910039393709031843585110912915796405926274571;
            6'd55: xpb[111] = 1024'd18693838854869554273434919951327038008430059325704684537778591039308701359233947322872414416795939704852373197969917515727702800842646079483053268222196083182115320563794386554317288163755254644016415859641676347872865547817005396780784635533840768171421865609519587360633404649093307809379268570184023554848;
            6'd56: xpb[111] = 1024'd91217986141176122983162203531425017750953327095690985931196735641464507762018063549115227021993058206798430547726457650677843631892858748305747400381192253965028355232704810942653378023615360784488102029242282737537091234269472708265513705813789552620688388788815322711979628340271663524964311170587715319456;
            6'd57: xpb[111] = 1024'd39675437743357950294090559706708564748778167739941603196483025178643418827493040865342968412532502399301338490025504351048920622101851082573281407523857383814250715332044017993359228691958261203649590590455649280836956070501043246785264206410508887803135008553994000033219323957521386223430663944365812599733;
            6'd58: xpb[111] = 1024'd112199585029664519003817843286806544491301435509927904589901169780799225230277157091585781017729620901247395839782044485999061453152063751395975539682853554597163750000954442381695318551818367344121276760056255670501181756953510558269993276690457672252401531733289735384565547648699741939015706544769504364341;
            6'd59: xpb[111] = 1024'd60657036631846346314746199462090091489126276154178521855187459317978136295752134407813522408269065093750303782081091186370138443361056085663509546825518684446386110100293649432401169220161267763282765321269622213801046593185081096789743777287177007434848151498468412705805243265949464637482059318547601644618;
            6'd60: xpb[111] = 1024'd9114488234028173625674555637373638486951116798429139120473748855157047361227111724041263798808509286253211724380137886741215433570048419931043553968183814295608470199632856483107019888504168182444253882482988757100911429416651635309494277883896342617294771263647090027044938883199187335948412092325698924895;
            6'd61: xpb[111] = 1024'd81638635520334742335401839217471618229474384568415440513891893457312853764011227950284076404005627788199269074136678021691356264620261088753737686127179985078521504868543280871443109748364274322915940052083595146765137115869118946794223348163845127066561294442942825378391162574377543051533454692729390689503;
            6'd62: xpb[111] = 1024'd30096087122516569646330195392755165227299225212666057779178182994491764829486205266511817794545071980702177016435724722062433254829253423021271693269845114927743864967882487922148960416707174742077428613296961690065001952100689485313973848760564462249007914208121502699630858191627265749999807466507487969780;
            6'd63: xpb[111] = 1024'd102620234408823138356057478972853144969822492982652359172596327596647571232270321492754630399742190482648234366192264857012574085879466091843965825428841285710656899636792912310485050276567280882549114782897568079729227638553156796798702919040513246698274437387417238050977081882805621465584850066911179734388;
        endcase
    end

    always_comb begin
        case(flag[37][11:6])
            6'd0: xpb[112] = 1024'd0;
            6'd1: xpb[112] = 1024'd51077686011004965666985835148136691967647333626902976437882617133826482297745298808982371790281634675151142308491311557383651076088458426111499832571506415559879259736132119361190900944910181301710603344110934623029092474784727335318453419637232581880721057152595915372216777500055344164051202840689277014665;
            6'd2: xpb[112] = 1024'd102155372022009931333971670296273383935294667253805952875765234267652964595490597617964743580563269350302284616982623114767302152176916852222999665143012831119758519472264238722381801889820362603421206688221869246058184949569454670636906839274465163761442114305191830744433555000110688328102405681378554029330;
            6'd3: xpb[112] = 1024'd29166362348890155602158578039595643158243573754973245185515996336502551555926757516932044156187229716010277518016441237571889387424154943779339372698188205745947104638825140745942463643213338183821612423945564022722916574133285232990381689228468296375343268043670688086543804426237399475034918695442236559664;
            6'd4: xpb[112] = 1024'd80244048359895121269144413187732335125890907381876221623398613470329033853672056325914415946468864391161419826507752794955540463512613369890839205269694621305826364374957260107133364588123519485532215768056498645752009048918012568308835108865700878256064325196266603458760581926292743639086121536131513574329;
            6'd5: xpb[112] = 1024'd7255038686775345537331320931054594348839813883043513933149375539178620814108216224881716522092824756869412727541570917760127698759851461447178912824869995932014949541518162130694026341516495065932621503780193422416740673481843130662309958819704010869965478934745460800870831352419454786018634550195196104663;
            6'd6: xpb[112] = 1024'd58332724697780311204317156079191286316487147509946490371031992673005103111853515033864088312374459432020555036032882475143778774848309887558678745396376411491894209277650281491884927286426676367643224847891128045445833148266570465980763378456936592750686536087341376173087608852474798950069837390884473119328;
            6'd7: xpb[112] = 1024'd109410410708785276871302991227327978284134481136849466808914609806831585409598813842846460102656094107171697344524194032527429850936768313670178577967882827051773469013782400853075828231336857669353828192002062668474925623051297801299216798094169174631407593239937291545304386352530143114121040231573750133993;
            6'd8: xpb[112] = 1024'd36421401035665501139489898970650237507083387638016759118665371875681172370034973741813760678280054472879690245558012155332017086184006405226518285523058201677962054180343302876636489984729833249754233927725757445139657247615128363652691648048172307245308746978416148887414635778656854261053553245637432664327;
            6'd9: xpb[112] = 1024'd87499087046670466806475734118786929474730721264919735556547989009507654667780272550796132468561689148030832554049323712715668162272464831338018118094564617237841313916475422237827390929640014551464837271836692068168749722399855698971145067685404889126029804131012064259631413278712198425104756086326709678992;
            6'd10: xpb[112] = 1024'd14510077373550691074662641862109188697679627766087027866298751078357241628216432449763433044185649513738825455083141835520255397519702922894357825649739991864029899083036324261388052683032990131865243007560386844833481346963686261324619917639408021739930957869490921601741662704838909572037269100390392209326;
            6'd11: xpb[112] = 1024'd65587763384555656741648477010245880665326961392990004304181368212183723925961731258745804834467284188889967763574453392903906473608161349005857658221246407423909158819168443622578953627943171433575846351671321467862573821748413596643073337276640603620652015022086836973958440204894253736088471941079669223991;
            6'd12: xpb[112] = 1024'd116665449395560622408634312158382572632974295019892980742063985346010206223707030067728176624748918864041110072065764950287557549696619775117357490792752822983788418555300562983769854572853352735286449695782256090891666296533140931961526756913873185501373072174682752346175217704949597900139674781768946238656;
            6'd13: xpb[112] = 1024'd43676439722440846676821219901704831855923201521060273051814747414859793184143189966695477200372879229749102973099583073092144784943857866673697198347928197609977003721861465007330516326246328315686855431505950867556397921096971494315001606867876318115274225913161609688285467131076309047072187795832628768990;
            6'd14: xpb[112] = 1024'd94754125733445812343807055049841523823570535147963249489697364548686275481888488775677848990654513904900245281590894630475795861032316292785197030919434613169856263457993584368521417271156509617397458775616885490585490395881698829633455026505108899995995283065757525060502244631131653211123390636521905783655;
            6'd15: xpb[112] = 1024'd21765116060326036611993962793163783046519441649130541799448126617535862442324648674645149566278474270608238182624712753280383096279554384341536738474609987796044848624554486392082079024549485197797864511340580267250222020445529391986929876459112032609896436804236382402612494057258364358055903650585588313989;
            6'd16: xpb[112] = 1024'd72842802071331002278979797941300475014166775276033518237330743751362344740069947483627521356560108945759380491116024310664034172368012810453036571046116403355924108360686605753272979969459666499508467855451514890279314495230256727305383296096344614490617493956832297774829271557313708522107106491274865328654;
            6'd17: xpb[112] = 1024'd123920488082335967945965633089437166981814108902936494675213360885188827037815246292609893146841743620910522799607335868047685248456471236564536403617622818915803368096818725114463880914369847801219071199562449513308406970014984062623836715733577196371338551109428213147046049057369052686158309331964142343319;
            6'd18: xpb[112] = 1024'd50931478409216192214152540832759426204763015404103786984964122954038413998251406191577193722465703986618515700641153990852272483703709328120876111172798193541991953263379627138024542667762823381619476935286144289973138594578814624977311565687580328985239704847907070489156298483495763833090822346027824873653;
            6'd19: xpb[112] = 1024'd102009164420221157881138375980896118172410349031006763422846740087864896295996705000559565512747338661769658009132465548235923559792167754232375943744304609101871212999511746499215443612673004683330080279397078913002231069363541960295764985324812910865960762000502985861373075983551107997142025186717101888318;
            6'd20: xpb[112] = 1024'd29020154747101382149325283724218377395359255532174055732597502156714483256432864899526866088371299027477650910166283671040510795039405845788715651299479983728059798166072648522776105366065980263730486015120773689666962693927372522649239835278816043479861915738981843203483325409677819144074538200780784418652;
            6'd21: xpb[112] = 1024'd80097840758106347816311118872355069363006589159077032170480119290540965554178163708509237878652933702628793218657595228424161871127864271900215483870986399287939057902204767883967006310976161565441089359231708312696055168712099857967693254916048625360582972891577758575700102909733163308125741041470061433317;
            6'd22: xpb[112] = 1024'd7108831084986572084498026615677328585955495660244324480230881359390552514614323607476538454276894068336786119691413351228749106375102363456555191426161773914127643068765669907527668064369137145841495094955403089360786793275930420321168104870051757974484126630056615917810352335859874455058254055533743963651;
            6'd23: xpb[112] = 1024'd58186517095991537751483861763814020553602829287147300918113498493217034812359622416458910244558528743487928428182724908612400182463560789568055023997668189474006902804897789268718569009279318447552098439066337712389879268060657755639621524507284339855205183782652531290027129835915218619109456896223020978316;
            6'd24: xpb[112] = 1024'd109264203106996503418469696911950712521250162914050277355996115627043517110104921225441282034840163418639070736674036465996051258552019215679554856569174605033886162541029908629909469954189499749262701783177272335418971742845385090958074944144516921735926240935248446662243907335970562783160659736912297992981;
            6'd25: xpb[112] = 1024'd36275193433876727686656604655272971744199069415217569665746877695893104070541081124408582610464123784347063637707854588800638493799257307235894564124349979660074747707590810653470131707582475329663107518900967112083703367409215653311549794098520054349827394673727304004354156762097273930093172750975980523315;
            6'd26: xpb[112] = 1024'd87352879444881693353642439803409663711846403042120546103629494829719586368286379933390954400745758459498205946199166146184289569887715733347394396695856395219954007443722930014661032652492656631373710863011901735112795842193942988630003213735752636230548451826323219376570934262152618094144375591665257537980;
            6'd27: xpb[112] = 1024'd14363869771761917621829347546731922934795309543287838413380256898569173328722539832358254976369718825206198847232984268988876805134953824903734104251031769846142592610283832038221694405885632211774116598735596511777527466757773550983478063689755768844449605564802076718681183688279329241076888605728940068314;
            6'd28: xpb[112] = 1024'd65441555782766883288815182694868614902442643170190814851262874032395655626467838641340626766651353500357341155724295826372527881223412251015233936822538185406021852346415951399412595350795813513484719942846531134806619941542500886301931483326988350725170662717397992090897961188334673405128091446418217082979;
            6'd29: xpb[112] = 1024'd116519241793771848955801017843005306870089976797093791289145491166222137924213137450322998556932988175508483464215607383756178957311870677126733769394044600965901112082548070760603496295705994815195323286957465757835712416327228221620384902964220932605891719869993907463114738688390017569179294287107494097644;
            6'd30: xpb[112] = 1024'd43530232120652073223987925586327566093038883298261083598896253235071724884649297349290299132556948541216476365249425506560766192559108768683073476949219975592089697249108972784164158049098970395595729022681160534500444040891058783973859752918224065219792873608472764805224988114516728716111807301171176627978;
            6'd31: xpb[112] = 1024'd94607918131657038890973760734464258060686216925164060036778870368898207182394596158272670922838583216367618673740737063944417268647567194794573309520726391151968956985241092145355058994009151697306332366792095157529536515675786119292313172555456647100513930761068680177441765614572072880163010141860453642643;
            6'd32: xpb[112] = 1024'd21618908458537263159160668477786517283635123426331352346529632437747794142830756057239971498462543582075611574774555186749004503894805286350913017075901765778157542151801994168915720747402127277706738102515789934194268140239616681645788022509459779714415084499547537519552015040698784027095523155924136172977;
            6'd33: xpb[112] = 1024'd72696594469542228826146503625923209251282457053234328784412249571574276440576054866222343288744178257226753883265866744132655579983263712462412849647408181338036801887934113530106621692312308579417341446626724557223360615024344016964241442146692361595136141652143452891768792540754128191146725996613413187642;
            6'd34: xpb[112] = 1024'd123774280480547194493132338774059901218929790680137305222294866705400758738321353675204715079025812932377896191757178301516306656071722138573912682218914596897916061624066232891297522637222489881127944790737659180252453089809071352282694861783924943475857198804739368263985570040809472355197928837302690202307;
            6'd35: xpb[112] = 1024'd50785270807427418761319246517382160441878697181304597532045628774250345698757513574172015654649773298085889092790996424320893891318960230130252389774089971524104646790627134914858184390615465461528350526461353956917184714372901914636169711737928076089758352543218225606095819466936183502130441851366372732641;
            6'd36: xpb[112] = 1024'd101862956818432384428305081665518852409526030808207573969928245908076827996502812383154387444931407973237031401282307981704544967407418656241752222345596387083983906526759254276049085335525646763238953870572288579946277189157629249954623131375160657970479409695814140978312596966991527666181644692055649747306;
            6'd37: xpb[112] = 1024'd28873947145312608696491989408841111632474937309374866279679007976926414956938972282121688020555368338945024302316126104509132202654656747798091929900771761710172491693320156299609747088918622343639359606295983356611008813721459812308097981329163790584380563434292998320422846393118238813114157706119332277640;
            6'd38: xpb[112] = 1024'd79951633156317574363477824556977803600122270936277842717561625110752897254684271091104059810837003014096166610807437661892783278743115173909591762472278177270051751429452275660800648033828803645349962950406917979640101288506187147626551400966396372465101620586888913692639623893173582977165360546808609292305;
            6'd39: xpb[112] = 1024'd6962623483197798631664732300300062823071177437445135027312387179602484215120430990071360386460963379804159511841255784697370513990353265465931470027453551896240336596013177684361309787221779225750368686130612756304832913070017709980026250920399505079002774325367771034749873319300294124097873560872291822639;
            6'd40: xpb[112] = 1024'd58040309494202764298650567448436754790718511064348111465195004313428966512865729799053732176742598054955301820332567342081021590078811691577431302598959967456119596332145297045552210732131960527460972030241547379333925387854745045298479670557632086959723831477963686406966650819355638288149076401561568837304;
            6'd41: xpb[112] = 1024'd109117995505207729965636402596573446758365844691251087903077621447255448810611028608036103967024232730106444128823878899464672666167270117688931135170466383015998856068277416406743111677042141829171575374352482002363017862639472380616933090194864668840444888630559601779183428319410982452200279242250845851969;
            6'd42: xpb[112] = 1024'd36128985832087954233823310339895705981314751192418380212828383516105035771047188507003404542648193095814437029857697022269259901414508209245270842725641757642187441234838318430303773430435117409571981110076176779027749487203302942970407940148867801454346042369038459121293677745537693599132792256314528382303;
            6'd43: xpb[112] = 1024'd87206671843092919900809145488032397948962084819321356650711000649931518068792487315985776332929827770965579338349008579652910977502966635356770675297148173202066700970970437791494674375345298711282584454187111402056841961988030278288861359786100383335067099521634374493510455245593037763183995097003805396968;
            6'd44: xpb[112] = 1024'd14217662169973144168996053231354657171910991320488648960461762718781105029228647214953076908553788136673572239382826702457498212750204726913110382852323547828255286137531339815055336128738274291682990189910806178721573586551860840642336209740103515948968253260113231835620704671719748910116508111067487927302;
            6'd45: xpb[112] = 1024'd65295348180978109835981888379491349139558324947391625398344379852607587326973946023935448698835422811824714547874138259841149288838663153024610215423829963388134545873663459176246237073648455593393593534021740801750666061336588175960789629377336097829689310412709147207837482171775093074167710951756764941967;
            6'd46: xpb[112] = 1024'd116373034191983075502967723527628041107205658574294601836226996986434069624719244832917820489117057486975856856365449817224800364927121579136110047995336378948013805609795578537437138018558636895104196878132675424779758536121315511279243049014568679710410367565305062580054259671830437238218913792446041956632;
            6'd47: xpb[112] = 1024'd43384024518863299771154631270950300330154565075461894145977759055283656585155404731885121064741017852683849757399267940029387600174359670692449755550511753574202390776356480560997799771951612475504602613856370201444490160685146073632717898968571812324311521303783919922164509097957148385151426806509724486966;
            6'd48: xpb[112] = 1024'd94461710529868265438140466419086992297801898702364870583860376189110138882900703540867492855022652527834992065890579497413038676262818096803949588122018169134081650512488599922188700716861793777215205957967304824473582635469873408951171318605804394205032578456379835294381286598012492549202629647199001501631;
            6'd49: xpb[112] = 1024'd21472700856748489706327374162409251520750805203532162893611138257959725843336863439834793430646612893542984966924397620217625911510056188360289295677193543760270235679049501945749362470254769357615611693690999601138314260033703971304646168559807526818933732194858692636491536024139203696135142661262684031965;
            6'd50: xpb[112] = 1024'd72550386867753455373313209310545943488398138830435139331493755391786208141082162248817165220928247568694127275415709177601276987598514614471789128248699959320149495415181621306940263415164950659326215037801934224167406734818431306623099588197040108699654789347454608008708313524194547860186345501951961046630;
            6'd51: xpb[112] = 1024'd123628072878758421040299044458682635456045472457338115769376372525612690438827461057799537011209882243845269583907020734984928063686973040583288960820206374880028755151313740668131164360075131961036818381912868847196499209603158641941553007834272690580375846500050523380925091024249892024237548342641238061295;
            6'd52: xpb[112] = 1024'd50639063205638645308485952202004894678994378958505408079127134594462277399263620956766837586833842609553262484940838857789515298934211132139628668375381749506217340317874642691691826113468107541437224117636563623861230834166989204295027857788275823194277000238529380723035340450376603171170061356704920591629;
            6'd53: xpb[112] = 1024'd101716749216643610975471787350141586646641712585408384517009751728288759697008919765749209377115477284704404793432150415173166375022669558251128500946888165066096600054006762052882727058378288843147827461747498246890323308951716539613481277425508405074998057391125296095252117950431947335221264197394197606294;
            6'd54: xpb[112] = 1024'd28727739543523835243658695093463845869590619086575676826760513797138346657445079664716509952739437650412397694465968537977753610269907649807468208502063539692285185220567664076443388811771264423548233197471193023555054933515547101966956127379511537688899211129604153437362367376558658482153777211457880136628;
            6'd55: xpb[112] = 1024'd79805425554528800910644530241600537837237952713478653264643130930964828955190378473698881743021072325563540002957280095361404686358366075918968041073569955252164444956699783437634289756681445725258836541582127646584147408300274437285409547016744119569620268282200068809579144876614002646204980052147157151293;
            6'd56: xpb[112] = 1024'd6816415881409025178831437984922797060186859214645945574393892999814415915626538372666182318645032691271532903991098218165991921605604167475307748628745329878353030123260685461194951510074421305659242277305822423248879032864104999638884396970747252183521422020678926151689394302740713793137493066210839681627;
            6'd57: xpb[112] = 1024'd57894101892413990845817273133059489027834192841548922012276510133640898213371837181648554108926667366422675212482409775549642997694062593586807581200251745438232289859392804822385852454984602607369845621416757046277971507648832334957337816607979834064242479173274841523906171802796057957188695906900116696292;
            6'd58: xpb[112] = 1024'd108971787903418956512803108281196180995481526468451898450159127267467380511117135990630925899208302041573817520973721332933294073782521019698307413771758160998111549595524924183576753399894783909080448965527691669307063982433559670275791236245212415944963536325870756896122949302851402121239898747589393710957;
            6'd59: xpb[112] = 1024'd35982778230299180780990016024518440218430432969619190759909889336316967471553295889598226474832262407281810422007539455737881309029759111254647121326933535624300134762085826207137415153287759489480854701251386445971795606997390232629266086199215548558864690064349614238233198728978113268172411761653076241291;
            6'd60: xpb[112] = 1024'd87060464241304146447975851172655132186077766596522167197792506470143449769298594698580598265113897082432952730498851013121532385118217537366146953898439951184179394498217945568328316098197940791191458045362321069000888081782117567947719505836448130439585747216945529610449976229033457432223614602342353255956;
            6'd61: xpb[112] = 1024'd14071454568184370716162758915977391409026673097689459507543268538993036729734754597547898840737857448140945631532669135926119620365455628922486661453615325810367979664778847591888977851590916371591863781086015845665619706345948130301194355790451263053486900955424386952560225655160168579156127616406035786290;
            6'd62: xpb[112] = 1024'd65149140579189336383148594064114083376674006724592435945425885672819519027480053406530270631019492123292087940023980693309770696453914055033986494025121741370247239400910966953079878796501097673302467125196950468694712181130675465619647775427683844934207958108020302324777003155215512743207330457095312800955;
            6'd63: xpb[112] = 1024'd116226826590194302050134429212250775344321340351495412383308502806646001325225352215512642421301126798443230248515292250693421772542372481145486326596628156930126499137043086314270779741411278975013070469307885091723804655915402800938101195064916426814929015260616217696993780655270856907258533297784589815620;
        endcase
    end

    always_comb begin
        case(flag[37][16:12])
            5'd0: xpb[113] = 1024'd0;
            5'd1: xpb[113] = 1024'd43237816917074526318321336955573034567270246852662704693059264875495588285661512114479942996925087164151223149549110373498009007789610572701826034151803531556315084303603988337831441494804254555413476205031579868388536280479233363291576045018919559428830168999095075039104030081397568054191046311848272345954;
            5'd2: xpb[113] = 1024'd86475633834149052636642673911146069134540493705325409386118529750991176571323024228959885993850174328302446299098220746996018015579221145403652068303607063112630168607207976675662882989608509110826952410063159736777072560958466726583152090037839118857660337998190150078208060162795136108382092623696544691908;
            5'd3: xpb[113] = 1024'd5646755067098837556165083461904670957112313432252429951045939561509869519675397433424757776117587183010520041189837685914963182527611383550317977439079553735254578341240747675864085292895557944930231006707499758801247991216803316909749565373529229019670603583168167087205562170264071145454449108919222553531;
            5'd4: xpb[113] = 1024'd48884571984173363874486420417477705524382560284915134644105204437005457805336909547904700773042674347161743190738948059412972190317221956252144011590883085291569662644844736013695526787699812500343707211739079627189784271696036680201325610392448788448500772582263242126309592251661639199645495420767494899485;
            5'd5: xpb[113] = 1024'd92122388901247890192807757373050740091652807137577839337164469312501046090998421662384643769967761511312966340288058432910981198106832528953970045742686616847884746948448724351526968282504067055757183416770659495578320552175270043492901655411368347877330941581358317165413622333059207253836541732615767245439;
            5'd6: xpb[113] = 1024'd11293510134197675112330166923809341914224626864504859902091879123019739039350794866849515552235174366021040082379675371829926365055222767100635954878159107470509156682481495351728170585791115889860462013414999517602495982433606633819499130747058458039341207166336334174411124340528142290908898217838445107062;
            5'd7: xpb[113] = 1024'd54531327051272201430651503879382376481494873717167564595151143998515327325012306981329458549160261530172263231928785745327935372844833339802461989029962639026824240986085483689559612080595370445273938218446579385991032262912839997111075175765978017468171376165431409213515154421925710345099944529686717453016;
            5'd8: xpb[113] = 1024'd97769143968346727748972840834955411048765120569830269288210408874010915610673819095809401546085348694323486381477896118825944380634443912504288023181766170583139325289689472027391053575399625000687414423478159254379568543392073360402651220784897576897001545164526484252619184503323278399290990841534989798970;
            5'd9: xpb[113] = 1024'd16940265201296512668495250385714012871336940296757289853137818684529608559026192300274273328352761549031560123569513057744889547582834150650953932317238661205763735023722243027592255878686673834790693020122499276403743973650409950729248696120587687059011810749504501261616686510792213436363347326757667660593;
            5'd10: xpb[113] = 1024'd60178082118371038986816587341287047438607187149419994546197083560025196844687704414754216325277848713182783273118623431242898555372444723352779966469042192762078819327326231365423697373490928390204169225154079144792280254129643314020824741139507246487841979748599576300720716592189781490554393638605940006547;
            5'd11: xpb[113] = 1024'd103415899035445565305137924296860082005877434002082699239256348435520785130349216529234159322202935877334006422667733804740907563162055296054606000620845724318393903630930219703255138868295182945617645430185659013180816534608876677312400786158426805916672148747694651339824746673587349544745439950454212352501;
            5'd12: xpb[113] = 1024'd22587020268395350224660333847618683828449253729009719804183758246039478078701589733699031104470348732042080164759350743659852730110445534201271909756318214941018313364962990703456341171582231779720924026829999035204991964867213267638998261494116916078682414332672668348822248681056284581817796435676890214124;
            5'd13: xpb[113] = 1024'd65824837185469876542981670803191718395719500581672424497243023121535066364363101848178974101395435896193303314308461117157861737900056106903097943908121746497333397668566979041287782666386486335134400231861578903593528245346446630930574306513036475507512583331767743387926278762453852636008842747525162560078;
            5'd14: xpb[113] = 1024'd109062654102544402861303007758764752962989747434335129190302287997030654650024613962658917098320523060344526463857571490655870745689666679604923978059925278053648481972170967379119224161190740890547876436893158771982064525825679994222150351531956034936342752330862818427030308843851420690199889059373434906032;
            5'd15: xpb[113] = 1024'd28233775335494187780825417309523354785561567161262149755229697807549347598376987167123788880587935915052600205949188429574815912638056917751589887195397768676272891706203738379320426464477789724651155033537498794006239956084016584548747826867646145098353017915840835436027810851320355727272245544596112767655;
            5'd16: xpb[113] = 1024'd71471592252568714099146754265096389352831814013924854448288962683044935884038499281603731877513023079203823355498298803072824920427667490453415921347201300232587976009807726717151867959282044280064631238569078662394776236563249947840323871886565704527183186914935910475131840932717923781463291856444385113609;
            5'd17: xpb[113] = 1024'd114709409169643240417468091220669423920102060866587559141348227558540524169700011396083674874438110243355046505047409176570833928217278063155241955499004831788903060313411715054983309454086298835478107443600658530783312517042483311131899916905485263956013355914030985514235871014115491835654338168292657459563;
            5'd18: xpb[113] = 1024'd33880530402593025336990500771428025742673880593514579706275637369059217118052384600548546656705523098063120247139026115489779095165668301301907864634477322411527470047444486055184511757373347669581386040244998552807487947300819901458497392241175374118023621499009002523233373021584426872726694653515335321186;
            5'd19: xpb[113] = 1024'd77118347319667551655311837727001060309944127446177284399334902244554805403713896715028489653630610262214343396688136488987788102955278874003733898786280853967842554351048474393015953252177602224994862245276578421196024227780053264750073437260094933546853790498104077562337403102981994926917740965363607667140;
            5'd20: xpb[113] = 1024'd120356164236742077973633174682574094877214374298839989092394167120050393689375408829508432650555697426365566546237246862485797110744889446705559932938084385524157638654652462730847394746981856780408338450308158289584560508259286628041649482279014492975683959497199152601441433184379562981108787277211880013094;
            5'd21: xpb[113] = 1024'd39527285469691862893155584233332696699786194025767009657321576930569086637727782033973304432823110281073640288328863801404742277693279684852225842073556876146782048388685233731048597050268905614511617046952498311608735938517623218368246957614704603137694225082177169610438935191848498018181143762434557874717;
            5'd22: xpb[113] = 1024'd82765102386766389211476921188905731267056440878429714350380841806064674923389294148453247429748197445224863437877974174902751285482890257554051876225360407703097132692289222068880038545073160169925093251984078179997272218996856581659823002633624162566524394081272244649542965273246066072372190074282830220671;
            5'd23: xpb[113] = 1024'd1936223619716174130999330739664333089628260605356734915308251616583367871741667352918119212015610299932937179969591113821696452431280495700717785360832898325721542426321993069081240848360209004028371848628418202021447649255193171986420477969314272728534659666250261658540467280715001109444546559505508082294;
            5'd24: xpb[113] = 1024'd45174040536790700449320667695237367656898507458019439608367516492078956157403179467398062208940697464084160329518701487319705460220891068402543819512636429882036626729925981406912682343164463559441848053659998070409983929734426535277996522988233832157364828665345336697644497362112569163635592871353780428248;
            5'd25: xpb[113] = 1024'd88411857453865226767642004650810402224168754310682144301426781367574544443064691581878005205865784628235383479067811860817714468010501641104369853664439961438351711033529969744744123837968718114855324258691577938798520210213659898569572568007153391586194997664440411736748527443510137217826639183202052774202;
            5'd26: xpb[113] = 1024'd7582978686815011687164414201569004046740574037609164866354191178093237391417064786342876988133197482943457221159428799736659634958891879251035762799912452060976120767562740744945326141255766948958602855335917960822695640471996488896170043342843501748205263249418428745746029450979072254898995668424730635825;
            5'd27: xpb[113] = 1024'd50820795603889538005485751157142038614010820890271869559413456053588825677078576900822819985058284647094680370708539173234668642748502451952861796951715983617291205071166729082776767636060021504372079060367497829211231920951229852187746088361763061177035432248513503784850059532376640309090041980273002981779;
            5'd28: xpb[113] = 1024'd94058612520964064323807088112715073181281067742934574252472720929084413962740089015302762981983371811245903520257649546732677650538113024654687831103519515173606289374770717420608209130864276059785555265399077697599768201430463215479322133380682620605865601247608578823954089613774208363281088292121275327733;
            5'd29: xpb[113] = 1024'd13229733753913849243329497663473675003852887469861594817400130739603106911092462219767634764250784665953977262349266485651622817486503262801353740238992005796230699108803488420809411434151324893888833862043417719623943631688799805805919608716372730767875866832586595832951591621243143400353444777343953189356;
            5'd30: xpb[113] = 1024'd56467550670988375561650834619046709571123134322524299510459395615098695196753974334247577761175871830105200411898376859149631825276113835503179774390795537352545783412407476758640852928955579449302310067074997588012479912168033169097495653735292290196706035831681670872055621702640711454544491089192225535310;
            5'd31: xpb[113] = 1024'd99705367588062901879972171574619744138393381175187004203518660490594283482415486448727520758100958994256423561447487232647640833065724408205005808542599068908860867716011465096472294423759834004715786272106577456401016192647266532389071698754211849625536204830776745911159651784038279508735537401040497881264;
        endcase
    end

    always_comb begin
        case(flag[38][5:0])
            6'd0: xpb[114] = 1024'd0;
            6'd1: xpb[114] = 1024'd71471592252568714099146754265096389352831814013924854448288962683044935884038499281603731877513023079203823355498298803072824920427667490453415921347201300232587976009807726717151867959282044280064631238569078662394776236563249947840323871886565704527183186914935910475131840932717923781463291856444385113609;
            6'd2: xpb[114] = 1024'd18876488821012686799494581125378345960965200902114024768446070301112976430767859653192392540368371848964497303539104171566586000014114646351671717678071559531485277450044236096673496727046882838819064868750917478425191622905603122715669174089901959787546470415754762920157153791507214545807893886263175742887;
            6'd3: xpb[114] = 1024'd90348081073581400898641335390474735313797014916038879216735032984157912314806358934796124417881394928168320659037402974639410920441782136805087639025272859764073253459851962813825364686328927118883696107319996140819967859468853070555993045976467664314729657330690673395288994724225138327271185742707560856496;
            6'd4: xpb[114] = 1024'd37752977642025373598989162250756691921930401804228049536892140602225952861535719306384785080736743697928994607078208343133172000028229292703343435356143119062970554900088472193346993454093765677638129737501834956850383245811206245431338348179803919575092940831509525840314307583014429091615787772526351485774;
            6'd5: xpb[114] = 1024'd109224569894594087698135916515853081274762215818152903985181103285270888745574218587988516958249766777132817962576507146205996920455896783156759356703344419295558530909896198910498861413375809957702760976070913619245159482374456193271662220066369624102276127746445436315446148515732352873079079628970736599383;
            6'd6: xpb[114] = 1024'd56629466463038060398483743376135037882895602706342074305338210903338929292303578959577177621105115546893491910617312514699758000042343939055015153034214678594455832350132708290020490181140648516457194606252752435275574868716809368147007522269705879362639411247264288760471461374521643637423681658789527228661;
            6'd7: xpb[114] = 1024'd4034363031482033098831570236416994491028989594531244625495318521406969839032939331165838283960464316654165858658117883193519079628791094953270949365084937893353133790369217669542118948905487075211628236434591251305990255059162543022352824473042134623002694748083141205496774233310934401768283688608317857939;
            6'd8: xpb[114] = 1024'd75505955284050747197978324501513383843860803608456099073784281204451905723071438612769570161473487395857989214156416686266344000056458585406686870712286238125941109800176944386693986908187531355276259475003669913700766491622412490862676696359607839150185881663019051680628615166028858183231575545052702971548;
            6'd9: xpb[114] = 1024'd22910851852494719898326151361795340451994190496645269393941388822519946269800798984358230824328836165618663162197222054760105079642905741304942667043156497424838411240413453766215615675952369914030693105185508729731181877964765665738021998562944094410549165163837904125653928024818148947576177574871493600826;
            6'd10: xpb[114] = 1024'd94382444105063433997472905626891729804826004510570123842230351505564882153839298265961962701841859244822486517695520857832930000070573231758358588390357797657426387250221180483367483635234414194095324343754587392125958114528015613578345870449509798937732352078773814600785768957536072729039469431315878714435;
            6'd11: xpb[114] = 1024'd41787340673507406697820732487173686412959391398759294162387459123632922700568658637550623364697208014583160465736326226326691079657020387656614384721228056956323688690457689862889112402999252752849757973936426208156373500870368788453691172652846054198095635579592667045811081816325363493384071461134669343713;
            6'd12: xpb[114] = 1024'd113258932926076120796967486752270075765791205412684148610676421806677858584607157919154355242210231093786983821234625029399516000084687878110030306068429357188911664700265416580040980362281297032914389212505504870551149737433618736294015044539411758725278822494528577520942922749043287274847363317579054457322;
            6'd13: xpb[114] = 1024'd60663829494520093497315313612552032373924592300873318930833529424745899131336518290743015905065579863547657769275430397893277079671135034008286102399299616487808966140501925959562609130046135591668822842687343686581565123775971911169360346742748013985642105995347429965968235607832578039191965347397845086600;
            6'd14: xpb[114] = 1024'd8068726062964066197663140472833988982057979189062489250990637042813939678065878662331676567920928633308331717316235766387038159257582189906541898730169875786706267580738435339084237897810974150423256472869182502611980510118325086044705648946084269246005389496166282410993548466621868803536567377216635715878;
            6'd15: xpb[114] = 1024'd79540318315532780296809894737930378334889793202987343699279599725858875562104377943935408445433951712512155072814534569459863079685249680359957820077371176019294243590546162056236105857093018430487887711438261165006756746681575033885029520832649973773188576411102192886125389399339792584999859233661020829487;
            6'd16: xpb[114] = 1024'd26945214883976752997157721598212334943023180091176514019436707343926916108833738315524069108289300482272829020855339937953624159271696836258213616408241435318191545030782671435757734624857856989242321341620099981037172133023928208760374823035986229033551859911921045331150702258129083349344461263479811458765;
            6'd17: xpb[114] = 1024'd98416807136545467096304475863308724295854994105101368467725670026971851992872237597127800985802323561476652376353638741026449079699364326711629537755442735550779521040590398152909602584139901269306952580189178643431948369587178156600698694922551933560735046826856955806282543190847007130807753119924196572374;
            6'd18: xpb[114] = 1024'd45821703704989439796652302723590680903988380993290538787882777645039892539601597968716461648657672331237326324394444109520210159285811482609885334086312994849676822480826907532431231351904739828061386210371017459462363755929531331476043997125888188821098330327675808251307856049636297895152355149742987201652;
            6'd19: xpb[114] = 1024'd117293295957558153895799056988687070256820195007215393236171740328084828423640097250320193526170695410441149679892742912593035079713478973063301255433514295082264798490634634249583099311186784108126017448940096121857139992492781279316367869012453893348281517242611718726439696982354221676615647006187372315261;
            6'd20: xpb[114] = 1024'd64698192526002126596146883848969026864953581895404563556328847946152868970369457621908854189026044180201823627933548281086796159299926128961557051764384554381162099930871143629104728078951622666880451079121934937887555378835134454191713171215790148608644800743430571171465009841143512440960249036006162944539;
            6'd21: xpb[114] = 1024'd12103089094446099296494710709250983473086968783593733876485955564220909517098817993497514851881392949962497575974353649580557238886373284859812848095254813680059401371107653008626356846716461225634884709303773753917970765177487629067058473419126403869008084244249423616490322699932803205304851065824953573817;
            6'd22: xpb[114] = 1024'd83574681347014813395641464974347372825918782797518588324774918247265845401137317275101246729394416029166320931472652452653382159314040775313228769442456113912647377380915379725778224805998505505699515947872852416312747001740737576907382345305692108396191271159185334091622163632650726986768142922269338687426;
            6'd23: xpb[114] = 1024'd30979577915458786095989291834629329434052169685707758644932025865333885947866677646689907392249764798926994879513457821147143238900487931211484565773326373211544678821151889105299853573763344064453949578054691232343162388083090751782727647509028363656554554660004186536647476491440017751112744952088129316704;
            6'd24: xpb[114] = 1024'd102451170168027500195136046099725718786883983699632613093220988548378821831905176928293639269762787878130818235011756624219968159328155421664900487120527673444132654830959615822451721533045388344518580816623769894737938624646340699623051519395594068183737741574940097011779317424157941532576036808532514430313;
            6'd25: xpb[114] = 1024'd49856066736471472895483872960007675395017370587821783413378096166446862378634537299882299932618136647891492183052561992713729238914602577563156283451397932743029956271196125201973350300810226903273014446805608710768354010988693874498396821598930323444101025075758949456804630282947232296920638838351305059591;
            6'd26: xpb[114] = 1024'd121327658989040186994630627225104064747849184601746637861667058849491798262673036581486031810131159727095315538550860795786554159342270068016572204798599232975617932281003851919125218260092271183337645685374687373163130247551943822338720693485496027971284211990694859931936471215665156078383930694795690173200;
            6'd27: xpb[114] = 1024'd68732555557484159694978454085386021355982571489935808181824166467559838809402396953074692472986508496855989486591666164280315238928717223914828001129469492274515233721240361298646847027857109742092079315556526189193545633894296997214065995688832283231647495491513712376961784074454446842728532724614480802478;
            6'd28: xpb[114] = 1024'd16137452125928132395326280945667977964115958378124978501981274085627879356131757324663353135841857266616663434632471532774076318515164379813083797460339751573412535161476870678168475795621948300846512945738365005223961020236650172089411297892168538492010778992332564821987096933243737607073134754433271431756;
            6'd29: xpb[114] = 1024'd87609044378496846494473035210764367316947772392049832950270236768672815240170256606267085013354880345820486790130770335846901238942831870266499718807541051806000511171284597395320343754903992580911144184307443667618737256799900119929735169778734243019193965907268475297118937865961661388536426610877656545365;
            6'd30: xpb[114] = 1024'd35013940946940819194820862071046323925081159280239003270427344386740855786899616977855745676210229115581160738171575704340662318529279026164755515138411311104897812611521106774841972522668831139665577814489282483649152643142253294805080471982070498279557249408087327742144250724750952152881028640696447174643;
            6'd31: xpb[114] = 1024'd106485533199509533293967616336142713277912973294163857718716307069785791670938116259459477553723252194784984093669874507413487238956946516618171436485612611337485788621328833491993840481950875419730209053058361146043928879705503242645404343868636202806740436323023238217276091657468875934344320497140832288252;
            6'd32: xpb[114] = 1024'd53890429767953505994315443196424669886046360182353028038873414687853832217667476631048138216578600964545658041710679875907248318543393672516427232816482870636383090061565342871515469249715713978484642683240199962074344266047856417520749646071972458067103719823842090662301404516258166698688922526959622917530;
            6'd33: xpb[114] = 1024'd1295326336397478694663270056706626494179747070542198359030522305921872764396837002636798879433949734306331989751485244401009398129840828414683029147353129935280391501801852251037098017480552537239076313422038778104759652390209592396094948275308713327467003324660943107326717375047457463033524556778413546808;
            6'd34: xpb[114] = 1024'd72766918588966192793810024321803015847011561084467052807319484988966808648435336284240530756946972813510155345249784047473834318557508318868098950494554430167868367511609578968188965976762596817303707551991117440499535888953459540236418820161874417854650190239596853582458558307765381244496816413222798660417;
            6'd35: xpb[114] = 1024'd20171815157410165494157851182084972455144947972656223127476592607034849195164696655829191419802321583270829293290589415967595398143955474766354746825424689466765668951846088347710594744527435376058141182172956256529951275295812715111764122365210673115013473740415706027483871166554672008841418443041589289695;
            6'd36: xpb[114] = 1024'd91643407409978879593304605447181361807976761986581077575765555290079785079203195937432923297315344662474652648788888219040420318571622965219770668172625989699353644961653815064862462703809479656122772420742034918924727511859062662952087994251776377642196660655351616502615712099272595790304710299485974403304;
            6'd37: xpb[114] = 1024'd39048303978422852293652432307463318416110148874770247895922662908147825625932556309021583960170693432235326596829693587534181398158070121118026464503496248998250946401890324444384091471574318214877206050923873734955142898201415837827433296455112632902559944156170468947641024958061886554649312329304765032582;
            6'd38: xpb[114] = 1024'd110519896230991566392799186572559707768941962888695102344211625591192761509971055590625315837683716511439149952327992390607006318585737611571442385850697549230838922411698051161535959430856362494941837289492952397349919134764665785667757168341678337429743131071106379422772865890779810336112604185749150146191;
            6'd39: xpb[114] = 1024'd57924792799435539093147013432841664377075349776884272664368733209260802056700415962213976500539065281199823900368797759100767398172184767469698182181567808529736223851934560541057588198621201053696270919674791213380334521107018960543102470545014592690106414571925231867798178749569101100457206215567940775469;
            6'd40: xpb[114] = 1024'd5329689367879511793494840293123620985208736665073442984525840827328842603429776333802637163394414050960497848409603127594528477758631923367953978512438067828633525292171069920579216966386039612450704549856630029410749907449372135418447772748350847950469698072744084312823491608358391864801808245386731404747;
            6'd41: xpb[114] = 1024'd76801281620448225892641594558220010338040550678998297432814803510373778487468275615406369040907437130164321203907901930667353398186299413821369899859639368061221501301978796637731084925668083892515335788425708691805526144012622083258771644634916552477652884987679994787955332541076315646265100101831116518356;
            6'd42: xpb[114] = 1024'd24206178188892198592989421418501966946173937567187467752971911128441819034197635986995029703762785899924995151948707299161114477772746569719625696190509627360118802742215306017252713693432922451269769418607547507835941530354975258134116946838252807738016168488498847232980645399865606410609702131649907147634;
            6'd43: xpb[114] = 1024'd95677770441460912692136175683598356299005751581112322201260873811486754918236135268598761581275808979128818507447006102233939398200414060173041617537710927592706778752023032734404581652714966731334400657176626170230717766918225205974440818724818512265199355403434757708112486332583530192072993988094292261243;
            6'd44: xpb[114] = 1024'd43082667009904885392484002543880312907139138469301492521417981429554795464965495640187422244131157748889492455487811470727700477786861216071297413868581186891604080192259542113926210420479805290088834287358464986261133153260578380849786120928154767525562638904253610153137799191372820956417596017913082890521;
            6'd45: xpb[114] = 1024'd114554259262473599491630756808976702259970952483226346969706944112599731349003994921791154121644180828093315810986110273800525398214528706524713335215782487124192056202067268831078078379761849570153465525927543648655909389823828328690109992814720472052745825819189520628269640124090744737880887874357468004130;
            6'd46: xpb[114] = 1024'd61959155830917572191978583669258658868104339371415517289864051730667771895733355293379814784499529597853989759026915642294286477800975862422969131546652746423089357642303778210599707147526688128907899156109382464686324776166181503565455295018056727313109109320008373073294952982880035502225489904176258633408;
            6'd47: xpb[114] = 1024'd9364052399361544892326410529540615476237726259604687610021159348735812442462715664968475447354878367614663707067721010788047557387423018321224927877523005721986659082540287590121335915291526687662332786291221280716740162508534678440800597221392982573472392820827225518320265841669326266570091933995049262686;
            6'd48: xpb[114] = 1024'd80835644651930258991473164794637004829069540273529542058310122031780748326501214946572207324867901446818487062566019813860872477815090508774640849224724305954574635092348014307273203874573570967726964024860299943111516399071784626281124469107958687100655579735763135993452106774387250048033383790439434376295;
            6'd49: xpb[114] = 1024'd28240541220374231691820991654918961437202927161718712378467229649848788873230575318160867987723250216579161010606825182354633557401537664672896645555594565253471936532584523686794832642338409526481397655042138759141931785414137801156469771311294942361018863236581988438477419633176540812377985820258225005573;
            6'd50: xpb[114] = 1024'd99712133472942945790967745920015350790034741175643566826756192332893724757269074599764599865236273295782984366105123985427458477829205155126312566902795865486059912542392250403946700601620453806546028893611217421536708021977387748996793643197860646888202050151517898913609260565894464593841277676702610119182;
            6'd51: xpb[114] = 1024'd47117030041386918491315572780297307398168128063832737146913299950961765303998434971353260528091622065543658314145929353921219557415652311024568363233666124784957213982628759783468329369385292365300462523793056237567123408319740923872138945401196902148565333652336751358634573424683755358185879706521400748460;
            6'd52: xpb[114] = 1024'd118588622293955632590462327045393696750999942077757591595202262634006701188036934252956992405604645144747481669644228156994044477843319801477984284580867425017545189992436486500620197328667336645365093762362134899961899644882990871712462817287762606675748520567272661833766414357401679139649171562965785862069;
            6'd53: xpb[114] = 1024'd65993518862399605290810153905675653359133328965946761915359370252074741734766294624545653068459993914508155617685033525487805557429766957376240080911737684316442491432672995880141826096432175204119527392543973715992315031225344046587808119491098861936111804068091514278791727216190969903993773592784576491347;
            6'd54: xpb[114] = 1024'd13398415430843577991157980765957609967266715854135932235516477870142782281495654996134313731315342684268829565725838893981566637016214113274495877242607943615339792872909505259663454864197013762873961022725812532022730417567697221463153421694435117196475087568910366723817040074980260668338375622603367120625;
            6'd55: xpb[114] = 1024'd84870007683412292090304735031053999320098529868060786683805440553187718165534154277738045608828365763472652921224137697054391557443881603727911798589809243847927768882717231976815322823479058042938592261294891194417506654130947169303477293581000821723658274483846277198948881007698184449801667479047752234234;
            6'd56: xpb[114] = 1024'd32274904251856264790652561891335955928231916756249957003962548171255758712263514649326706271683714533233326869264943065548152637030328759626167594920679503146825070322953741356336951591243896601693025891476730010447922040473300344178822595784337076984021557984665129643974193866487475214146269508866542863512;
            6'd57: xpb[114] = 1024'd103746496504424978889799316156432345281063730770174811452251510854300694596302013930930438149196737612437150224763241868620977557457996250079583516267880803379413046332761468073488819550525940881757657130045808672842698277036550292019146467670902781511204744899601040119106034799205398995609561365310927977121;
            6'd58: xpb[114] = 1024'd51151393072868951590147143016714301889197117658363981772408618472368735143031374302519098812052086382197824172804047237114738637044443405977839312598751062678310347772997977453010448318290779440512090760227647488873113663378903466894491769874239036771568028400419892564131347657994689759954163395129718606399;
            6'd59: xpb[114] = 1024'd122622985325437665689293897281810691242028931672288836220697581155413671027069873584122830689565109461401647528302346040187563557472110896431255233945952362910898323782805704170162316277572823720576721998796726151267889899942153414734815641760804741298751215315355803039263188590712613541417455251574103720008;
            6'd60: xpb[114] = 1024'd70027881893881638389641724142092647850162318560478006540854688773481711573799233955711491352420458231162321476343151408681324637058558052329511030276822622209795625223042213549683945045337662279331155628978564967298305286284506589610160943964140996559114498816174655484288501449501904305762057281392894349286;
            6'd61: xpb[114] = 1024'd17432778462325611089989551002374604458295705448667176861011796391549752120528594327300152015275807000922995424383956777175085716645005208227766826607692881508692926663278722929205573813102500838085589259160403783328720672626859764485506246167477251819477782316993507929313814308291195070106659311211684978564;
            6'd62: xpb[114] = 1024'd88904370714894325189136305267470993811127519462592031309300759074594688004567093608903883892788830080126818779882255580247910637072672698681182747954894181741280902673086449646357441772384545118150220497729482445723496909190109712325830118054042956346660969231929418404445655241009118851569951167656070092173;
            6'd63: xpb[114] = 1024'd36309267283338297889484132127752950419260906350781201629457866692662728551296453980492544555644178849887492727923060948741671716659119854579438544285764441040178204113322959025879070540149383676904654127911321261753912295532462887201175420257379211607024252732748270849470968099798409615914553197474860721451;
        endcase
    end

    always_comb begin
        case(flag[38][11:6])
            6'd0: xpb[115] = 1024'd0;
            6'd1: xpb[115] = 1024'd107780859535907011988630886392849339772092720364706056077746829375707664435334953262096276433157201929091316083421359751814496637086787345032854465632965741272766180123130685743030938499431427956969285366480399924148688532095712835041499292143944916134207439647684181324602809032516333397377845053919245835060;
            6'd2: xpb[115] = 1024'd91495023387689282578462845380884246799487013603676428027361803686438433533360767614177481651656729548739482759385226069049929433332354355510548806249600441611841685676690154148431637807345650192628373124573560001933016213970528897118020014604660383001594975881251304619099089991104033777637000281212897185789;
            6'd3: xpb[115] = 1024'd75209187239471553168294804368919153826881306842646799976976777997169202631386581966258686870156257168387649435349092386285362229577921365988243146866235141950917191230249622553832337115259872428287460882666720079717343895845344959194540737065375849868982512114818427913595370949691734157896155508506548536518;
            6'd4: xpb[115] = 1024'd58923351091253823758126763356954060854275600081617171926591752307899971729412396318339892088655784788035816111312958703520795025823488376465937487482869842289992696783809090959233036423174094663946548640759880157501671577720161021271061459526091316736370048348385551208091651908279434538155310735800199887247;
            6'd5: xpb[115] = 1024'd42637514943036094347958722344988967881669893320587543876206726618630740827438210670421097307155312407683982787276825020756227822069055386943631828099504542629068202337368559364633735731088316899605636398853040235285999259594977083347582181986806783603757584581952674502587932866867134918414465963093851237976;
            6'd6: xpb[115] = 1024'd26351678794818364937790681333023874909064186559557915825821700929361509925464025022502302525654840027332149463240691337991660618314622397421326168716139242968143707890928027770034435039002539135264724156946200313070326941469793145424102904447522250471145120815519797797084213825454835298673621190387502588705;
            6'd7: xpb[115] = 1024'd10065842646600635527622640321058781936458479798528287775436675240092279023489839374583507744154367646980316139204557655227093414560189407899020509332773943307219213444487496175435134346916761370923811915039360390854654623344609207500623626908237717338532657049086921091580494784042535678932776417681153939434;
            6'd8: xpb[115] = 1024'd117846702182507647516253526713908121708551200163234343853183504615799943458824792636679784177311569576071632222625917407041590051646976752931874974965739684579985393567618181918466072846348189327893097281519760315003343155440322042542122919052182633472740096696771102416183303816558869076310621471600399774494;
            6'd9: xpb[115] = 1024'd101560866034289918106085485701943028735945493402204715802798478926530712556850606988760989395811097195719798898589783724277022847892543763409569315582374384919060899121177650323866772154262411563552185039612920392787670837315138104618643641512898100340127632930338225710679584775146569456569776698894051125223;
            6'd10: xpb[115] = 1024'd85275029886072188695917444689977935763339786641175087752413453237261481654876421340842194614310624815367965574553650041512455644138110773887263656199009085258136404674737118729267471462176633799211272797706080470571998519189954166695164363973613567207515169163905349005175865733734269836828931926187702475952;
            6'd11: xpb[115] = 1024'd68989193737854459285749403678012842790734079880145459702028427547992250752902235692923399832810152435016132250517516358747888440383677784364957996815643785597211910228296587134668170770090856034870360555799240548356326201064770228771685086434329034074902705397472472299672146692321970217088087153481353826681;
            6'd12: xpb[115] = 1024'd52703357589636729875581362666047749818128373119115831651643401858723019850928050045004605051309680054664298926481382675983321236629244794842652337432278485936287415781856055540068870078005078270529448313892400626140653882939586290848205808895044500942290241631039595594168427650909670597347242380775005177410;
            6'd13: xpb[115] = 1024'd36417521441419000465413321654082656845522666358086203601258376169453788948953864397085810269809207674312465602445248993218754032874811805320346678048913186275362921335415523945469569385919300506188536071985560703924981564814402352924726531355759967809677777864606718888664708609497370977606397608068656528139;
            6'd14: xpb[115] = 1024'd20131685293201271055245280642117563872916959597056575550873350480184558046979678749167015488308735293960632278409115310454186829120378815798041018665547886614438426888974992350870268693833522741847623830078720781709309246689218415001247253816475434677065314098173842183160989568085071357865552835362307878868;
            6'd15: xpb[115] = 1024'd3845849144983541645077239630152470900311252836026947500488324790915327145005493101248220706808262913608798954372981627689619625365945826275735359282182586953513932442534460756270968001747744977506711588171880859493636928564034477077767976277190901544452850331740965477657270526672771738124708062655959229597;
            6'd16: xpb[115] = 1024'd111626708680890553633708126023001810672403973200733003578235154166622991580340446363344497139965464842700115037794341379504116262452733171308589824915148328226280112565665146499301906501179172934475996954652280783642325460659747312119267268421135817678660289979425146802260079559189105135502553116575205064657;
            6'd17: xpb[115] = 1024'd95340872532672824223540085011036717699798266439703375527850128477353760678366260715425702358464992462348281713758207696739549058698300181786284165531783028565355618119224614904702605809093395170135084712745440861426653142534563374195787990881851284546047826212992270096756360517776805515761708343868856415386;
            6'd18: xpb[115] = 1024'd79055036384455094813372043999071624727192559678673747477465102788084529776392075067506907576964520081996448389722074013974981854943867192263978506148417728904431123672784083310103305117007617405794172470838600939210980824409379436272308713342566751413435362446559393391252641476364505896020863571162507766115;
            6'd19: xpb[115] = 1024'd62769200236237365403204002987106531754586852917644119427080077098815298874417889419588112795464047701644615065685940331210414651189434202741672846765052429243506629226343551715504004424921839641453260228931761016995308506284195498348829435803282218280822898680126516685748922434952206276280018798456159116844;
            6'd20: xpb[115] = 1024'd46483364088019635993035961975141438781981146156614491376695051409546067972443703771669318013963575321292781741649806648445847447435001213219367187381687129582582134779903020120904703732836061877112347987024921094779636188159011560425350158263997685148210434913693639980245203393539906656539174025749810467573;
            6'd21: xpb[115] = 1024'd30197527939801906582867920963176345809375439395584863326310025720276837070469518123750523232463102940940948417613672965681280243680568223697061527998321829921657640333462488526305403040750284112771435745118081172563963870033827622501870880724713152015597971147260763274741484352127607036798329253043461818302;
            6'd22: xpb[115] = 1024'd13911691791584177172699879951211252836769732634555235275925000031007606168495332475831728450962630560589115093577539282916713039926135234174755868614956530260733145887021956931706102348664506348430523503211241250348291551908643684578391603185428618882985507380827886569237765310715307417057484480337113169031;
            6'd23: xpb[115] = 1024'd121692551327491189161330766344060592608862452999261291353671829406715270603830285737928004884119832489680431176998899034731209677012922579207610334247922271533499326010152642674737040848095934305399808869691641174496980084004356519619890895329373535017192947028512067893840574343231640814435329534256359004091;
            6'd24: xpb[115] = 1024'd105406715179273459751162725332095499636256746238231663303286803717446039701856100090009210102619360109328597852962765351966642473258489589685304674864556971872574831563712111080137740156010156541058896627784801252281307765879172581696411617790089001884580483262079191188336855301819341194694484761550010354820;
            6'd25: xpb[115] = 1024'd89120879031055730340994684320130406663651039477202035252901778028176808799881914442090415321118887728976764528926631669202075269504056600162999015481191672211650337117271579485538439463924378776717984385877961330065635447753988643772932340250804468751968019495646314482833136260407041574953639988843661705549;
            6'd26: xpb[115] = 1024'd72835042882838000930826643308165313691045332716172407202516752338907577897907728794171620539618415348624931204890497986437508065749623610640693356097826372550725842670831047890939138771838601012377072143971121407849963129628804705849453062711519935619355555729213437777329417218994741955212795216137313056278;
            6'd27: xpb[115] = 1024'd56549206734620271520658602296200220718439625955142779152131726649638346995933543146252825758117942968273097880854364303672940861995190621118387696714461072889801348224390516296339838079752823248036159902064281485634290811503620767925973785172235402486743091962780561071825698177582442335471950443430964407007;
            6'd28: xpb[115] = 1024'd40263370586402542110490561284235127745833919194113151101746700960369116093959357498334030976617470587921264556818230620908373658240757631596082037331095773228876853777949984701740537387667045483695247660157441563418618493378436830002494507632950869354130628196347684366321979136170142715731105670724615757736;
            6'd29: xpb[115] = 1024'd23977534438184812700322520272270034773228212433083523051361675271099885191985171850415236195116998207569431232782096938143806454486324642073776377947730473567952359331509453107141236695581267719354335418250601641202946175253252892079015230093666336221518164429914807660818260094757843095990260898018267108465;
            6'd30: xpb[115] = 1024'd7691698289967083290154479260304941800622505672053895000976649581830654290010986202496441413616525827217597908745963255379239250731891652551470718564365173907027864885068921512541936003495489955013423176343761718987273857128068954155535952554381803088905700663481930955314541053345543476249416125311918459194;
            6'd31: xpb[115] = 1024'd115472557825874095278785365653154281572715226036759951078723478957538318725345939464592717846773727756308913992167323007193735887818678997584325184197330915179794045008199607255572874502926917911982708542824161643135962389223781789197035244698326719223113140311166112279917350085861876873627261179231164294254;
            6'd32: xpb[115] = 1024'd99186721677656365868617324641189188600109519275730323028338453268269087823371753816673923065273255375957080668131189324429168684064246008062019524813965615518869550561759075660973573810841140147641796300917321720920290071098597851273555967159042186090500676544733235574413631044449577253886416406524815644983;
            6'd33: xpb[115] = 1024'd82900885529438636458449283629224095627503812514700694977953427578999856921397568168755128283772782995605247344095055641664601480309813018539713865430600315857945056115318544066374273118755362383300884059010481798704617752973413913350076689619757652957888212778300358868909912003037277634145571633818466995712;
            6'd34: xpb[115] = 1024'd66615049381220907048281242617259002654898105753671066927568401889730626019423382520836333502272310615253414020058921958900034276555380029017408206047235016197020561668878012471774972426669584618959971817103641876488945434848229975426597412080473119825275749011867482163406192961624978014404726861112118346441;
            6'd35: xpb[115] = 1024'd50329213233003177638113201605293909682292398992641438877183376200461395117449196872917538720771838234901580696022788276135467072800947039495102546663869716536096067222437480877175671734583806854619059575196801954273273116723046037503118134541188586692663285245434605457902473920212678394663882088405769697170;
            6'd36: xpb[115] = 1024'd34043377084785448227945160593328816709686692231611810826798350511192164215475011224998743939271365854549747371986654593370899869046514049972796887280504416875171572775996949282576371042498029090278147333289962032057600798597862099579638857001904053560050821479001728752398754878800378774923037315699421047899;
            6'd37: xpb[115] = 1024'd17757540936567718817777119581363723737080985470582182776413324821922933313500825577079949157770893474197914047950520910606332665292081060450491227897139117214247078329556417687977070350412251325937235091383122109841928480472678161656159579462619520427438357712568852046895035837388079155182192542993072398628;
            6'd38: xpb[115] = 1024'd1471704788349989407609078569398630764475278709552554726028299132653702411526639929161154376270421093846080723914387227841765461537648070928185568513773817553322583883115886093377769658326473561596322849476282187626256162347494223732680301923334987294825893946135975341391316795975779535441347770286723749357;
            6'd39: xpb[115] = 1024'd109252564324257001396239964962247970536567999074258610803775128508361366846861593191257430809427623022937396807335746979656262098624435415961040034146739558826088764006246571836408708157757901518565608215956682111774944694443207058774179594067279903429033333593820156665994125828492112932819192824205969584417;
            6'd40: xpb[115] = 1024'd92966728176039271986071923950282877563962292313228982753390102819092135944887407543338636027927150642585563483299613296891694894870002426438734374763374259165164269559806040241809407465672123754224695974049842189559272376318023120850700316527995370296420869827387279960490406787079813313078348051499620935146;
            6'd41: xpb[115] = 1024'd76680892027821542575903882938317784591356585552199354703005077129822905042913221895419841246426678262233730159263479614127127691115569436916428715380008959504239775113365508647210106773586345989883783732143002267343600058192839182927221038988710837163808406060954403254986687745667513693337503278793272285875;
            6'd42: xpb[115] = 1024'd60395055879603813165735841926352691618750878791169726652620051440553674140939036247501046464926205881881896835227345931362560487361136447394123055996643659843315280666924977052610806081500568225542871490236162345127927740067655245003741761449426304031195942294521526549482968704255214073596658506086923636604;
            6'd43: xpb[115] = 1024'd44109219731386083755567800914387598646145172030140098602235025751284443238964850599582251683425733501530063511191212248597993283606703457871817396613278360182390786220484445458011505389414790461201959248329322422912255421942471307080262483910141770898583478528088649843979249662842914453855813733380574987333;
            6'd44: xpb[115] = 1024'd27823383583168354345399759902422505673539465269110470551850000062015212336990664951663456901925261121178230187155078565833426079852270468349511737229913060521466291774043913863412204697329012696861047006422482500696583103817287369156783206370857237765971014761655773138475530621430614834114968960674226338062;
            6'd45: xpb[115] = 1024'd11537547434950624935231718890457412700933758508080842501464974372745981435016479303744662120424788740826396863118944883068858876097837478827206077846547760860541797327603382268812904005243234932520134764515642578480910785692103431233303928831572704633358550995222896432971811580018315214374124187967877688791;
            6'd46: xpb[115] = 1024'd119318406970857636923862605283306752473026478872786898579211803748453645870351432565840938553581990669917712946540304634883355513184624823860060543479513502133307977450734068011843842504674662889489420130996042502629599317787816266274803220975517620767565990642907077757574620612534648611751969241887123523851;
            6'd47: xpb[115] = 1024'd103032570822639907513694564271341659500420772111757270528826778059184414968377246917922143772081518289565879622504170952118788309430191834337754884096148202472383483004293536417244541812588885125148507889089202580413926999662632328351323943436233087634953526876474201052070901571122348992011124469180774874580;
            6'd48: xpb[115] = 1024'd86746734674422178103526523259376566527815065350727642478441752369915184066403061270003348990581045909214046298468037269354221105675758844815449224712782902811458988557853004822645241120503107360807595647182362658198254681537448390427844665896948554502341063110041324346567182529710049372270279696474426225309;
            6'd49: xpb[115] = 1024'd70460898526204448693358482247411473555209358589698014428056726680645953164428875622084554209080573528862212974431903586589653901921325855293143565329417603150534494111412473228045940428417329596466683405275522735982582363412264452504365388357664021369728599343608447641063463488297749752529434923768077576038;
            6'd50: xpb[115] = 1024'd54175062377986719283190441235446380582603651828668386377671700991376722262454689974165759427580101148510379650395769903825086698166892865770837905946052303489609999664971941633446639736331551832125771163368682813766910045287080514580886110818379488237116135577175570935559744446885450132788590151061728926767;
            6'd51: xpb[115] = 1024'd37889226229768989873022400223481287609997945067638758327286675302107491360480504326246964646079628768158546326359636221060519494412459876248532246562687003828685505218531410038847339044245774067784858921461842891551237727161896576657406833279094955104503671810742694230056025405473150513047745378355380277496;
            6'd52: xpb[115] = 1024'd21603390081551260462854359211516194637392238306609130276901649612838260458506318678328169864579156387806713002323502538295952290658026886726226587179321704167761010772090878444248038352159996303443946679555002969335565409036712638733927555739810421971891208044309817524552306364060850893306900605649031628225;
            6'd53: xpb[115] = 1024'd5317553933333531052686318199551101664786531545579502226516623923569029556532133030409375083078684007454879678287368855531385086903593897203920927795956404506836516325650346849648737660074218539103034437648163047119893090911528700810448278200525888839278744277876940819048587322648551273566055832942682978954;
            6'd54: xpb[115] = 1024'd113098413469240543041317204592400441436879251910285558304263453299276693991867086292505651516235885936546195761708728607345881723990381242236775393428922145779602696448781032592679676159505646496072319804128562971268581623007241535851947570344470804973486183925561122143651396355164884670943900886861928814014;
            6'd55: xpb[115] = 1024'd96812577321022813631149163580435348464273545149255930253878427610007463089892900644586856734735413556194362437672594924581314520235948252714469734045556846118678202002340500998080375467419868731731407562221723049052909304882057597928468292805186271840873720159128245438147677313752585051203056114155580164743;
            6'd56: xpb[115] = 1024'd80526741172805084220981122568470255491667838388226302203493401920738232187918714996668061953234941175842529113636461241816747316481515263192164074662191546457753707555899969403481074775334090967390495320314883126837236986756873660004989015265901738708261256392695368732643958272340285431462211341449231515472;
            6'd57: xpb[115] = 1024'd64240905024587354810813081556505162519062131627196674153108376231469001285944529348749267171734468795490695789600327559052180112727082273669858415278826246796829213109459437808881774083248313203049583078408043204621564668631689722081509737726617205575648792626262492027140239230927985811721366568742882866201;
            6'd58: xpb[115] = 1024'd47955068876369625400645040544540069546456424866167046102723350542199770383970343700830472390233996415138862465564193876287612908972649284147552755895460947135904718663018906214282473391162535438708670836501203282405892350506505784158030460187332672443036328859829615321636520189515686191980521796036534216930;
            6'd59: xpb[115] = 1024'd31669232728151895990476999532574976573850718105137418052338324852930539481996158052911677608733524034787029141528060193523045705218216294625247096512095647474980224216578374619683172699076757674367758594594363360190220032381321846234551182648048139310423865093396738616132801148103386572239677023330185567659;
            6'd60: xpb[115] = 1024'd15383396579934166580308958520609883601245011344107790001953299163661308580021972404992882827233051654435195817491926510758478501463783305102941437128730347814055729770137843025083872006990979910026846352687523437974547714256137908311071905108763606177811401326963861910629082106691086952498832250623836918388;
            6'd61: xpb[115] = 1024'd123164256115841178568939844913459223373337731708813846079700128539368973015356925667089159260390253583526511900913286262572975138550570650135795902761696089086821909893268528768114810506422407866996131719167923362123236246351850743352571197252708522312018840974648043235231891139207420349876677304543082753448;
            6'd62: xpb[115] = 1024'd106878419967623449158771803901494130400732024947784218029315102850099742113382740019170364478889781203174678576877152579808407934796137660613490243378330789425897415446827997173515509814336630102655219477261083439907563928226666805429091919713423989179406377208215166529728172097795120730135832531836734104177;
            6'd63: xpb[115] = 1024'd90592583819405719748603762889529037428126318186754589978930077160830511211408554371251569697389308822822845252841018897043840731041704671091184583994965489764972921000387465578916209122250852338314307235354243517691891610101482867505612642174139456046793913441782289824224453056382821110394987759130385454906;
        endcase
    end

    always_comb begin
        case(flag[38][16:12])
            5'd0: xpb[116] = 1024'd0;
            5'd1: xpb[116] = 1024'd74306747671187990338435721877563944455520611425724961928545051471561280309434368723332774915888836442471011928804885214279273527287271681568878924611600190104048426553946933984316908430165074573973394993447403595476219291976298929582133364634854922914181449675349413118720734014970521490654142986424036805635;
            5'd2: xpb[116] = 1024'd24546799658251239278072516350313456166342795725714239728958247878145665281559598536650478617119998575498874450152276993979483213733323028582597724206869339274406178538322650631003577668812943426636592378507567344588077733731701086199288159586480396561542995936581768207334939956012409964189596146222479126939;
            5'd3: xpb[116] = 1024'd98853547329439229616508238227877400621863407151439201657503299349706945590993967259983253533008835017969886378957162208258756741020594710151476648818469529378454605092269584615320486098978018000609987371954970940064297025708000015781421524221335319475724445611931181326055673970982931454843739132646515932574;
            5'd4: xpb[116] = 1024'd49093599316502478556145032700626912332685591451428479457916495756291330563119197073300957234239997150997748900304553987958966427466646057165195448413738678548812357076645301262007155337625886853273184757015134689176155467463402172398576319172960793123085991873163536414669879912024819928379192292444958253878;
            5'd5: xpb[116] = 1024'd123400346987690468894580754578190856788206202877153441386461547227852610872553565796633732150128833593468760829109439202238239954753917738734074373025338868652860783630592235246324063767790961427246579750462538284652374759439701101980709683807815716037267441548512949533390613926995341419033335278868995059513;
            5'd6: xpb[116] = 1024'd73640398974753717834217549050940368499028387177142719186874743634436995844678795609951435851359995726496623350456830981938449641199969085747793172620608017823218535614967951893010733006438830279909777135522702033764233201195103258597864478759441189684628987809745304622004819868037229892568788438667437380817;
            5'd7: xpb[116] = 1024'd23880450961816966773854343523689880209850571477131996987287940041021380816804025423269139552591157859524485871804222761638659327646020432761511972215877166993576287599343668539697402245086699132572974520582865782876091642950505415215019273711066663331990534070977659710619025809079118366104241598465879702121;
            5'd8: xpb[116] = 1024'd98187198633004957112290065401253824665371182902856958915832991512582661126238394146601914468479994301995497800609107975917932854933292114330390896827477357097624714153290602524014310675251773706546369514030269378352310934926804344797152638345921586246171983746327072829339759824049639856758384584889916507756;
            5'd9: xpb[116] = 1024'd48427250620068206051926859874003336376193367202846236716246187919167046098363623959919618169711156435023360321956499755618142541379343461344109696422746506267982466137666319170700979913899642559209566899090433127464169376682206501414307433297547059893533530007559427917953965765091528330293837744688358829060;
            5'd10: xpb[116] = 1024'd122733998291256196390362581751567280831713978628571198644791239390728326407797992683252393085599992877494372250761384969897416068666615142912988621034346696372030892691613253155017888344064717133182961892537836722940388668658505430996440797932401982807714979682908841036674699780062049820947980731112395634695;
            5'd11: xpb[116] = 1024'd72974050278319445329999376224316792542536162928560476445204435797312711379923222496570096786831155010522234772108776749597625755112666489926707420629615845542388644675988969801704557582712585985846159277598000472052247110413907587613595592884027456455076525944141196125288905721103938294483433890910837955999;
            5'd12: xpb[116] = 1024'd23214102265382694269636170697066304253358347228549754245617632203897096352048452309887800488062317143550097293456168529297835441558717836940426220224884994712746396660364686448391226821360454838509356662658164221164105552169309744230750387835652930102438072205373551213903111662145826768018887050709280277303;
            5'd13: xpb[116] = 1024'd97520849936570684608071892574630248708878958654274716174162683675458376661482821033220575403951153586021109222261053743577108968845989518509305144836485184816794823214311620432708135251525529412482751656105567816640324844145608673812883752470507853016619521880722964332623845677116348258673030037133317082938;
            5'd14: xpb[116] = 1024'd47760901923633933547708687047379760419701142954263993974575880082042761633608050846538279105182315719048971743608445523277318655292040865523023944431754333987152575198687337079394804490173398265145949041165731565752183285901010830430038547422133326663981068141955319421238051618158236732208483196931759404242;
            5'd15: xpb[116] = 1024'd122067649594821923886144408924943704875221754379988955903120931553604041943042419569871054021071152161519983672413330737556592182579312547091902869043354524091201001752634271063711712920338472839119344034613135161228402577877309760012171912056988249578162517817304732539958785633128758222862626183355796209877;
            5'd16: xpb[116] = 1024'd72307701581885172825781203397693216586043938679978233703534127960188426915167649383188757722302314294547846193760722517256801869025363894105621668638623673261558753737009987710398382158986341691782541419673298910340261019632711916629326707008613723225524064078537087628572991574170646696398079343154238531181;
            5'd17: xpb[116] = 1024'd22547753568948421765417997870442728296866122979967511503947324366772811887292879196506461423533476427575708715108114296957011555471415241119340468233892822431916505721385704357085051397634210544445738804733462659452119461388114073246481501960239196872885610339769442717187197515212535169933532502952680852485;
            5'd18: xpb[116] = 1024'd96854501240136412103853719748006672752386734405692473432492375838334092196727247919839236339422312870046720643912999511236285082758686922688219392845493012535964932275332638341401959827799285118419133798180866254928338753364413002828614866595094119787067060015118855835907931530183056660587675489376717658120;
            5'd19: xpb[116] = 1024'd47094553227199661043490514220756184463208918705681751232905572244918477168852477733156940040653475003074583165260391290936494769204738269701938192440762161706322684259708354988088629066447153971082331183241030004040197195119815159445769661546719593434428606276351210924522137471224945134123128649175159979424;
            5'd20: xpb[116] = 1024'd121401300898387651381926236098320128918729530131406713161450623716479757478286846456489714956542311445545595094065276505215768296492009951270817117052362351810371110813655288972405537496612228545055726176688433599516416487096114089027903026181574516348610055951700624043242871486195466624777271635599196785059;
            5'd21: xpb[116] = 1024'd71641352885450900321563030571069640629551714431395990961863820123064142450412076269807418657773473578573457615412668284915977982938061298284535916647631500980728862798031005619092206735260097397718923561748597348628274928851516245645057821133199989995971602212932979131857077427237355098312724795397639106363;
            5'd22: xpb[116] = 1024'd21881404872514149261199825043819152340373898731385268762277016529648527422537306083125122359004635711601320136760060064616187669384112645298254716242900650151086614782406722265778875973907966250382120946808761097740133370606918402262212616084825463643333148474165334220471283368279243571848177955196081427667;
            5'd23: xpb[116] = 1024'd96188152543702139599635546921383096795894510157110230690822068001209807731971674806457897274893472154072332065564945278895461196671384326867133640854500840255135041336353656250095784404073040824355515940256164693216352662583217331844345980719680386557514598149514747339192017383249765062502320941620118233302;
            5'd24: xpb[116] = 1024'd46428204530765388539272341394132608506716694457099508491235264407794192704096904619775600976124634287100194586912337058595670883117435673880852440449769989425492793320729372896782453642720909677018713325316328442328211104338619488461500775671305860204876144410747102427806223324291653536037774101418560554606;
            5'd25: xpb[116] = 1024'd120734952201953378877708063271696552962237305882824470419780315879355473013531273343108375892013470729571206515717222272874944410404707355449731365061370179529541219874676306881099362072885984250992108318763732037804430396314918418043634140306160783119057594086096515546526957339262175026691917087842597360241;
            5'd26: xpb[116] = 1024'd70975004189016627817344857744446064673059490182813748220193512285939857985656503156426079593244632862599069037064614052575154096850758702463450164656639328699898971859052023527786031311533853103655305703823895786916288838070320574660788935257786256766419140347328870635141163280304063500227370247641039681545;
            5'd27: xpb[116] = 1024'd21215056176079876756981652217195576383881674482803026020606708692524242957781732969743783294475794995626931558412005832275363783296810049477168964251908477870256723843427740174472700550181721956318503088884059536028147279825722731277943730209411730413780686608561225723755369221345951973762823407439482002849;
            5'd28: xpb[116] = 1024'd95521803847267867095417374094759520839402285908527987949151760164085523267216101693076558210364631438097943487216891046554637310584081731046047888863508667974305150397374674158789608980346796530291898082331463131504366571802021660860077094844266653327962136283910638842476103236316473464416966393863518808484;
            5'd29: xpb[116] = 1024'd45761855834331116035054168567509032550224470208517265749564956570669908239341331506394261911595793571125806008564282826254846997030133078059766688458777817144662902381750390805476278218994665382955095467391626880616225013557423817477231889795892126975323682545142993931090309177358361937952419553661961129788;
            5'd30: xpb[116] = 1024'd120068603505519106373489890445072977005745081634242227678110008042231188548775700229727036827484630013596817937369168040534120524317404759628645613070378007248711328935697324789793186649159739956928490460839030476092444305533722747059365254430747049889505132220492407049811043192328883428606562540085997935423;
            5'd31: xpb[116] = 1024'd70308655492582355313126684917822488716567265934231505478523204448815573520900930043044740528715792146624680458716559820234330210763456106642364412665647156419069080920073041436479855887807608809591687845899194225204302747289124903676520049382372523536866678481724762138425249133370771902142015699884440256727;
        endcase
    end

    always_comb begin
        case(flag[39][5:0])
            6'd0: xpb[117] = 1024'd0;
            6'd1: xpb[117] = 1024'd72307701581885172825781203397693216586043938679978233703534127960188426915167649383188757722302314294547846193760722517256801869025363894105621668638623673261558753737009987710398382158986341691782541419673298910340261019632711916629326707008613723225524064078537087628572991574170646696398079343154238531181;
            6'd2: xpb[117] = 1024'd20548707479645604252763479390572000427389450234220783278936400855399958493026159856362444229946954279652542980063951599934539897209507453656083212260916305589426832904448758083166525126455477662254885230959357974316161189044527060293674844333997997184228224742957117227039455074412660375677468859682882578031;
            6'd3: xpb[117] = 1024'd92856409061530777078544682788265217013433388914199016982470528815588385408193809239551201952249268574200389173824674117191341766234871347761704880899539978850985586641458745793564907285441819354037426650632656884656422208677238976923001551342611720409752288821494204855612446648583307072075548202837121109212;
            6'd4: xpb[117] = 1024'd41097414959291208505526958781144000854778900468441566557872801710799916986052319712724888459893908559305085960127903199869079794419014907312166424521832611178853665808897516166333050252910955324509770461918715948632322378089054120587349688667995994368456449485914234454078910148825320751354937719365765156062;
            6'd5: xpb[117] = 1024'd113405116541176381331308162178837217440822839148419800261406929670988343901219969095913646182196222853852932153888625717125881663444378801417788093160456284440412419545907503876731432411897297016292311881592014858972583397721766037216676395676609717593980513564451322082651901722995967447753017062520003687243;
            6'd6: xpb[117] = 1024'd61646122438936812758290438171716001282168350702662349836809202566199875479078479569087332689840862838957628940191854799803619691628522360968249636782748916768280498713346274249499575379366432986764655692878073922948483567133581180881024533001993991552684674228871351681118365223237981127032406579048647734093;
            6'd7: xpb[117] = 1024'd9887128336697244185272714164594785123513862256904899412211475461411407056936990042261019197485502824062325726495083882481357719812665920518711180405041549096148577880785044622267718346835568957236999504164132986924383736545396324545372670327378265511388834893291381279584828723479994806311796095577291780943;
            6'd8: xpb[117] = 1024'd82194829918582417011053917562288001709557800936883133115745603421599833972104639425449776919787817118610171920255806399738159588838029814624332849043665222357707331617795032332666100505821910649019540923837431897264644756178108241174699377335991988736912898971828468908157820297650641502709875438731530312124;
            6'd9: xpb[117] = 1024'd30435835816342848438036193555166785550903312491125682691147876316811365549963149898623463427432457103714868706559035482415897617022173374174794392665957854685575410785233802705434243473291046619491884735123490961240544925589923384839047514661376262695617059636248498506624283797892655181989264955260174358974;
            6'd10: xpb[117] = 1024'd102743537398228021263817396952860002136947251171103916394682004276999792465130799281812221149734771398262714900319757999672699486047537268280416061304581527947134164522243790415832625632277388311274426154796789871580805945222635301468374221669989985921141123714785586135197275372063301878387344298414412890155;
            6'd11: xpb[117] = 1024'd50984543295988452690799672945738785978292762725346465970084277172211324042989309754985907657379411383367411686622987082350437514231680827830877604926874160275002243689682560788600768599746524281746769966082848935556706114634450445132722358995374259879845284379205615733663738872305315557666733814943056937005;
            6'd12: xpb[117] = 1024'd123292244877873625516580876343432002564336701405324699673618405132399750958156959138174665379681725677915257880383709599607239383257044721936499273565497833536560997426692548498999150758732865973529311385756147845896967134267162361762049066003987983105369348457742703362236730446475962254064813158097295468186;
            6'd13: xpb[117] = 1024'd71533250775634056943563152336310786405682212959567249249020678027611282536015469611348351887326365663019954666686938682284977411441188281486960817187790465864429076594131318871767293726202001944001655197042206909872867303678977505426397203329372257064073509122162732960703193946717975933344202674625939515036;
            6'd14: xpb[117] = 1024'd19774256673394488370545428329189570247027724513809798824422950922822814113873980084522038394971005648124651452990167764962715439625331841037422360810083098192297155761570089244535436693671137914473999008328265973848767473090792649090745340654756531022777669786582762559169657446959989612623592191154583561886;
            6'd15: xpb[117] = 1024'd92081958255279661196326631726882786833071663193788032527957078883011241029041629467710796117273319942672497646750890282219517308650695735143044029448706771453855909498580076954933818852657479606256540428001564884189028492723504565720072047663370254248301733865119850187742649021130636309021671534308822093067;
            6'd16: xpb[117] = 1024'd40322964153040092623308907719761570674417174748030582103359351778222772606900139940884482624917959927777194433054119364897255336834839294693505573070999403781723988666018847327701961820126615576728884239287623948164928662135319709384420184988754528207005894529539879786209112521372649988301061050837466139917;
            6'd17: xpb[117] = 1024'd112630665734925265449090111117454787260461113428008815806893479738411199522067789324073240347220274222325040626814841882154057205860203188799127241709623077043282742403028835038100343979112957268511425658960922858505189681768031626013746891997368251432529958608076967414782104095543296684699140393991704671098;
            6'd18: xpb[117] = 1024'd60871671632685696876072387110333571101806624982251365382295752633622731099926299797246926854864914207429737413118070964831795234044346748349588785331915709371150821570467605410868486946582093238983769470246981922481089851179846769678095029322752525391234119272496997013248567595785310363978529910520348717948;
            6'd19: xpb[117] = 1024'd9112677530446128303054663103212354943152136536493914957698025528834262677784810270420613362509554192534434199421300047509533262228490307900050328954208341699018900737906375783636629914051229209456113281533040986456990020591661913342443166648136799349938279936917026611715031096027324043257919427048992764798;
            6'd20: xpb[117] = 1024'd81420379112331301128835866500905571529196075216472148661232153489022689592952459653609371084811868487082280393182022564766335131253854202005671997592832014960577654474916363494035012073037570901238654701206339896797251040224373829971769873656750522575462344015454114240288022670197970739655998770203231295979;
            6'd21: xpb[117] = 1024'd29661385010091732555818142493784355370541586770714698236634426384234221170810970126783057592456508472186977179485251647444073159437997761556133541215124647288445733642355133866803155040506706871710998512492398960773151209636188973636118010982134796534166504679874143838754486170439984418935388286731875342829;
            6'd22: xpb[117] = 1024'd101969086591976905381599345891477571956585525450692931940168554344422648085978619509971815314758822766734823373245974164700875028463361655661755209853748320550004487379365121577201537199493048563493539932165697871113412229268900890265444717990748519759690568758411231467327477744610631115333467629886113874010;
            6'd23: xpb[117] = 1024'd50210092489737336808581621884356355797931037004935481515570827239634179663837129983145501822403462751839520159549203247378613056647505215212216753476040952877872566546803891949969680166962184533965883743451756935089312398680716033929792855316132793718394729422831261065793941244852644794612857146414757920860;
            6'd24: xpb[117] = 1024'd122517794071622509634362825282049572383974975684913715219104955199822606579004779366334259544705777046387366353309925764635414925672869109317838422114664626139431320283813879660368062325948526225748425163125055845429573418313427950559119562324746516943918793501368348694366932819023291491010936489568996452041;
            6'd25: xpb[117] = 1024'd70758799969382941061345101274928356225320487239156264794507228095034138156863289839507946052350417031492063139613154847313152953857012668868299965736957258467299399451252650033136205293417662196220768974411114909405473587725243094223467699650130790902622954165788378292833396319265305170290326006097640498891;
            6'd26: xpb[117] = 1024'd18999805867143372488327377267807140066665998793398814369909500990245669734721800312681632559995057016596759925916383929990890982041156228418761509359249890795167478618691420405904348260886798166693112785697173973381373757137058237887815836975515064861327114830208407891299859819507318849569715522626284545741;
            6'd27: xpb[117] = 1024'd91307507449028545314108580665500356652709937473377048073443628950434096649889449695870390282297371311144606119677106447247692851066520122524383177997873564056726232355701408116302730419873139858475654205370472883721634776769770154517142543984128788086851178908745495519872851393677965545967794865780523076922;
            6'd28: xpb[117] = 1024'd39548513346788976741090856658379140494055449027619597648845901845645628227747960169044076789942011296249302905980335529925430879250663682074844721620166196384594311523140178489070873387342275828947998016656531947697534946181585298181490681309513062045555339573165525118339314893919979225247184382309167123772;
            6'd29: xpb[117] = 1024'd111856214928674149566872060056072357080099387707597831352380029805834055142915609552232834512244325590797149099741058047182232748276027576180466390258789869646153065260150166199469255546328617520730539436329830858037795965814297214810817388318126785271079403651702612746912306468090625921645263725463405654953;
            6'd30: xpb[117] = 1024'd60097220826434580993854336048951140921444899261840380927782302701045586720774120025406521019888965575901845886044287129859970776460171135730927933881082501974021144427588936572237398513797753491202883247615889922013696135226112358475165525643511059229783564316122642345378769968332639600924653241992049701803;
            6'd31: xpb[117] = 1024'd8338226724195012420836612041829924762790410816082930503184575596257118298632630498580207527533605561006542672347516212537708804644314695281389477503375134301889223595027706945005541481266889461675227058901948985989596304637927502139513662968895333188487724980542671943845233468574653280204042758520693748653;
            6'd32: xpb[117] = 1024'd80645928306080185246617815439523141348834349496061164206718703556445545213800279881768965249835919855554388866108238729794510673669678589387011146141998807563447977332037694655403923640253231153457768478575247896329857324270639418768840369977509056414011789059079759572418225042745299976602122101674932279834;
            6'd33: xpb[117] = 1024'd28886934203840616673600091432401925190179861050303713782120976451657076791658790354942651757480559840659085652411467812472248701853822148937472689764291439891316056499476465028172066607722367123930112289861306960305757493682454562433188507302893330372715949723499789170884688542987313655881511618203576326684;
            6'd34: xpb[117] = 1024'd101194635785725789499381294830095141776223799730281947485655104411845503706826439738131409479782874135206931846172190329729050570879186043043094358402915113152874810236486452738570448766708708815712653709534605870646018513315166479062515214311507053598240013802036876799457680117157960352279590961357814857865;
            6'd35: xpb[117] = 1024'd49435641683486220926363570822973925617569311284524497061057377307057035284684950211305095987427514120311628632475419412406788599063329602593555902025207745480742889403925223111338591734177844786184997520820664934621918682726981622726863351636891327556944174466456906397924143617399974031558980477886458904715;
            6'd36: xpb[117] = 1024'd121743343265371393752144774220667142203613249964502730764591505267245462199852599594493853709729828414859474826236141929663590468088693496699177570663831418742301643140935210821736973893164186477967538940493963844962179702359693539356190058645505050782468238544993994026497135191570620727957059821040697435896;
            6'd37: xpb[117] = 1024'd69984349163131825179127050213545926044958761518745280339993778162456993777711110067667540217374468399964171612539371012341328496272837056249639114286124051070169722308373981194505116860633322448439882751780022908938079871771508683020538195970889324741172399209414023624963598691812634407236449337569341482746;
            6'd38: xpb[117] = 1024'd18225355060892256606109326206424709886304273072987829915396051057668525355569620540841226725019108385068868398842600095019066524456980615800100657908416683398037801475812751567273259828102458418912226563066081972913980041183323826684886333296273598699876559873834053223430062192054648086515838854097985529596;
            6'd39: xpb[117] = 1024'd90533056642777429431890529604117926472348211752966063618930179017856952270737269924029984447321422679616714592603322612275868393482344509905722326547040356659596555212822739277671641987088800110694767982739380883254241060816035743314213040304887321925400623952371140852003053766225294782913918197252224060777;
            6'd40: xpb[117] = 1024'd38774062540537860858872805596996710313693723307208613194332451913068483848595780397203670954966062664721411378906551694953606421666488069456183870169332988987464634380261509650439784954557936081167111794025439947230141230227850886978561177630271595884104784616791170450469517266467308462193307713780868107627;
            6'd41: xpb[117] = 1024'd111081764122423033684654008994689926899737661987186846897866579873256910763763429780392428677268376959269257572667274212210408290691851963561805538807956662249023388117271497360838167113544277772949653213698738857570402249860562803607887884638885319109628848695328258079042508840637955158591387056935106638808;
            6'd42: xpb[117] = 1024'd59322770020183465111636284987568710741083173541429396473268852768468442341621940253566115184913016944373954358970503294888146318875995523112267082430249294576891467284710267733606310081013413743421997024984797921546302419272377947272236021964269593068333009359748287677508972340879968837870776573463750685658;
            6'd43: xpb[117] = 1024'd7563775917943896538618560980447494582428685095671946048671125663679973919480450726739801692557656929478651145273732377565884347060139082662728626052541926904759546452149038106374453048482549713894340836270856985522202588684193090936584159289653867027037170024168317275975435841121982517150166089992394732508;
            6'd44: xpb[117] = 1024'd79871477499829069364399764378140711168472623775650179752205253623868400834648100109928559414859971224026497339034454894822686216085502976768350294691165600166318300189159025816772835207468891405676882255944155895862463608316905007565910866298267590252561234102705404904548427415292629213548245433146633263689;
            6'd45: xpb[117] = 1024'd28112483397589500791382040371019495009818135329892729327607526519079932412506610583102245922504611209131194125337683977500424244269646536318811838313458232494186379356597796189540978174938027376149226067230214959838363777728720151230259003623651864211265394767125434503014890915534642892827634949675277310539;
            6'd46: xpb[117] = 1024'd100420184979474673617163243768712711595862074009870963031141654479268359327674259966291003644806925503679040319098406494757226113295010430424433506952081905755745133093607783899939360333924369067931767486903513870178624797361432067859585710632265587436789458845662522131587882489705289589225714292829515841720;
            6'd47: xpb[117] = 1024'd48661190877235105044145519761591495437207585564113512606543927374479890905532770439464690152451565488783737105401635577434964141479153989974895050574374538083613212261046554272707503301393505038404111298189572934154524966773247211523933847957649861395493619510082551730054345989947303268505103809358159888570;
            6'd48: xpb[117] = 1024'd120968892459120277869926723159284712023251524244091746310078055334668317820700419822653447874753879783331583299162358094691766010504517884080516719212998211345171965998056541983105885460379846730186652717862871844494785986405959128153260554966263584621017683588619639358627337564117949964903183152512398419751;
            6'd49: xpb[117] = 1024'd69209898356880709296908999152163495864597035798334295885480328229879849398558930295827134382398519768436280085465587177369504038688661443630978262835290843673040045165495312355874028427848982700658996529148930908470686155817774271817608692291647858579721844253039668957093801064359963644182572669041042466601;
            6'd50: xpb[117] = 1024'd17450904254641140723891275145042279705942547352576845460882601125091380976417440769000820890043159753540976871768816260047242066872805003181439806457583476000908124332934082728642171395318118671131340340434989972446586325229589415481956829617032132538426004917459698555560264564601977323461962185569686513451;
            6'd51: xpb[117] = 1024'd89758605836526313549672478542735496291986486032555079164416729085279807891585090152189578612345474048088823065529538777304043935898168897287061475096207149262466878069944070439040553554304460362913881760108288882786847344862301332111283536625645855763950068995996786184133256138772624019860041528723925044632;
            6'd52: xpb[117] = 1024'd37999611734286744976654754535614280133331997586797628739819001980491339469443600625363265119990114033193519851832767859981781964082312456837523018718499781590334957237382840811808696521773596333386225571394347946762747514274116475775631673951030129722654229660416815782599719639014637699139431045252569091482;
            6'd53: xpb[117] = 1024'd110307313316171917802435957933307496719375936266775862443353129940679766384611250008552022842292428327741366045593490377238583833107676350943144687357123454851893710974392828522207078680759938025168766991067646857103008533906828392404958380959643852948178293738953903411172711213185284395537510388406807622663;
            6'd54: xpb[117] = 1024'd58548319213932349229418233926186280560721447821018412018755402835891297962469760481725709349937068312846062831896719459916321861291819910493606230979416087179761790141831598894975221648229073995641110802353705921078908703318643536069306518285028126906882454403373933009639174713427298074816899904935451669513;
            6'd55: xpb[117] = 1024'd6789325111692780656400509919065064402066959375260961594157675731102829540328270954899395857581708297950759618199948542594059889475963470044067774601708719507629869309270369267743364615698209966113454613639764985054808872730458679733654655610412400865586615067793962608105638213669311754096289421464095716363;
            6'd56: xpb[117] = 1024'd79097026693577953482181713316758280988110898055239195297691803691291256455495920338088153579884022592498605811960671059850861758501327364149689443240332392769188623046280356978141746774684551657895996033313063895395069892363170596362981362619026124091110679146331050236678629787839958450494368764618334247544;
            6'd57: xpb[117] = 1024'd27338032591338384909163989309637064829456409609481744873094076586502788033354430811261840087528662577603302598263900142528599786685470923700150986862625025097056702213719127350909889742153687628368339844599122959370970061774985740027329499944410398049814839810751079835145093288081972129773758281146978294394;
            6'd58: xpb[117] = 1024'd99645734173223557734945192707330281415500348289459978576628204546691214948522080194450597809830976872151148792024622659785401655710834817805772655501248698358615455950729115061308271901140029320150881264272421869711231081407697656656656206953024121275338903889288167463718084862252618826171837624301216825575;
            6'd59: xpb[117] = 1024'd47886740070983989161927468700209065256845859843702528152030477441902746526380590667624284317475616857255845578327851742463139683894978377356234199123541330686483535118167885434076414868609165290623225075558480933687131250819512800321004344278408395234043064553708197062184548362494632505451227140829860872425;
            6'd60: xpb[117] = 1024'd120194441652869161987708672097902281842889798523680761855564605402091173441548240050813042039777931151803691772088574259719941552920342271461855867762165003948042288855177873144474797027595506982405766495231779844027392270452224716950331051287022118459567128632245284690757539936665279201849306483984099403606;
            6'd61: xpb[117] = 1024'd68435447550629593414690948090781065684235310077923311430966878297302705019406750523986728547422571136908388558391803342397679581104485831012317411384457636275910368022616643517242939995064642952878110306517838908003292439864039860614679188612406392418271289296665314289224003436907292881128696000512743450456;
            6'd62: xpb[117] = 1024'd16676453448390024841673224083659849525580821632165861006369151192514236597265260997160415055067211122013085344695032425075417609288629390562778955006750268603778447190055413890011082962533778923350454117803897971979192609275855004279027325937790666376975449961085343887690466937149306560408085517041387497306;
            6'd63: xpb[117] = 1024'd88984155030275197667454427481353066111624760312144094709903279152702663512432910380349172777369525416560931538455754942332219478313993284668400623645373941865337200927065401600409465121520120615132995537477196882319453628908566920908354032946404389602499514039622431516263458511319953256806164860195626028487;
        endcase
    end

    always_comb begin
        case(flag[39][11:6])
            6'd0: xpb[118] = 1024'd0;
            6'd1: xpb[118] = 1024'd37225160928035629094436703474231849952970271866386644285305552047914195090291420853522859285014165401665628324758984025009957506498136844218862167267666574193205280094504171973177608088989256585605339348763255946295353798320382064572702170271788663561203674704042461114729922011561966936085554376724270075337;
            6'd2: xpb[118] = 1024'd74450321856071258188873406948463699905940543732773288570611104095828390180582841707045718570028330803331256649517968050019915012996273688437724334535333148386410560189008343946355216177978513171210678697526511892590707596640764129145404340543577327122407349408084922229459844023123933872171108753448540150674;
            6'd3: xpb[118] = 1024'd111675482784106887283310110422695549858910815599159932855916656143742585270874262560568577855042496204996884974276952075029872519494410532656586501802999722579615840283512515919532824266967769756816018046289767838886061394961146193718106510815365990683611024112127383344189766034685900808256663130172810226011;
            6'd4: xpb[118] = 1024'd24833948028017774978947886492112967067182660339810893013090353126679885023856544504076365925398987297219363891578442665460766185151327042320288544054335255839130445808445470555080193164439820621111159786665783938817054343060631485325830111403925204977994795402052786428813159972319234727223527680271485817017;
            6'd5: xpb[118] = 1024'd62059108956053404073384589966344817020152932206197537298395905174594080114147965357599225210413152698884992216337426690470723691649463886539150711322001830032335725902949642528257801253429077206716499135429039885112408141381013549898532281675713868539198470106095247543543081983881201663309082056995755892354;
            6'd6: xpb[118] = 1024'd99284269884089033167821293440576666973123204072584181583701457222508275204439386211122084495427318100550620541096410715480681198147600730758012878589668404225541005997453814501435409342418333792321838484192295831407761939701395614471234451947502532100402144810137708658273003995443168599394636433720025967691;
            6'd7: xpb[118] = 1024'd12442735127999920863459069509994084181395048813235141740875154205445574957421668154629872565783809192773099458397901305911574863804517240421714920841003937485055611522386769136982778239890384656616980224568311931338754887800880906078958052536061746394785916100063111742896397933076502518361500983818701558697;
            6'd8: xpb[118] = 1024'd49667896056035549957895772984225934134365320679621786026180706253359770047713089008152731850797974594438727783156885330921532370302654084640577088108670511678260891616890941110160386328879641242222319573331567877634108686121262970651660222807850409955989590804105572857626319944638469454447055360542971634034;
            6'd9: xpb[118] = 1024'd86893056984071179052332476458457784087335592546008430311486258301273965138004509861675591135812139996104356107915869355931489876800790928859439255376337085871466171711395113083337994417868897827827658922094823823929462484441645035224362393079639073517193265508148033972356241956200436390532609737267241709371;
            6'd10: xpb[118] = 1024'd51522227982066747970252527875201295607437286659390468659955284211264890986791805183379206168631088326835025217359946362383542457707438523141297627672619130980777236328067718885363315340948692122800662470839923860455432541130326832085993668198287811577036798073437056979635893833770309499474287365917300377;
            6'd11: xpb[118] = 1024'd37276683156017695842406956002107051248577709153046034753965507332125459981278212658706238491182796489992463349976343971372341048955844282742003464895339193324186057330832239692062971404330205277728140011234095870155809230861512391404788163939986951372780711502115898171709557905395737245585028664090187375714;
            6'd12: xpb[118] = 1024'd74501844084053324936843659476338901201547981019432679039271059380039655071569633512229097776196961891658091674735327996382298555453981126960865632163005767517391337425336411665240579493319461863333479359997351816451163029181894455977490334211775614933984386206158359286439479916957704181670583040814457451051;
            6'd13: xpb[118] = 1024'd111727005012088954031280362950570751154518252885819323324576611427953850161861054365751957061211127293323719999494312021392256061952117971179727799430672341710596617519840583638418187582308718448938818708760607762746516827502276520550192504483564278495188060910200820401169401928519671117756137417538727526388;
            6'd14: xpb[118] = 1024'd24885470255999841726918139019988168362790097626470283481750308410891149914843336309259745131567618385546198916795802611823149727609034480843429841682007874970111223044773538273965556479780769313233960449136623862677509775601761812157916105072123492789571832200126223485792795866153005036723001967637403117394;
            6'd15: xpb[118] = 1024'd62110631184035470821354842494220018315760369492856927767055860458805345005134757162782604416581783787211827241554786636833107234107171325062292008949674449163316503139277710247143164568770025898839299797899879808972863573922143876730618275343912156350775506904168684600522717877714971972808556344361673192731;
            6'd16: xpb[118] = 1024'd99335792112071099915791545968451868268730641359243572052361412506719540095426178016305463701595949188877455566313770661843064740605308169281154176217341023356521783233781882220320772657759282484444639146663135755268217372242525941303320445615700819911979181608211145715252639889276938908894110721085943268068;
            6'd17: xpb[118] = 1024'd12494257355981987611429322037869285477002486099894532209535109489656839848408459959813251771952440281099934483615261252273958406262224678944856218468676556616036388758714836855868141555231333348739780887039151855199210320342011232911044046204260034206362952898136548799876033826910272827860975271184618859074;
            6'd18: xpb[118] = 1024'd49719418284017616705866025512101135429972757966281176494840661537571034938699880813336111056966605682765562808374245277283915912760361523163718385736343130809241668853219008829045749644220589934345120235802407801494564118662393297483746216476048697767566627602179009914605955838472239763946529647908888934411;
            6'd19: xpb[118] = 1024'd86944579212053245800302728986332985382943029832667820780146213585485230028991301666858970341980771084431191133133229302293873419258498367382580553004009705002446948947723180802223357733209846519950459584565663747789917916982775362056448386747837361328770302306221471029335877850034206700032084024633159009748;
            6'd20: xpb[118] = 1024'd103044455964133495940505055750402591214874573318780937319910568422529781973583610366758412337262176653670050434719892724767084915414877046282595255345238261961554472656135437770726630681897384245601324941679847720910865082260653664171987336396575623154073596146874113959271787667540618998948574731834600754;
            6'd21: xpb[118] = 1024'd37328205383999762590377208529982252544185146439705425222625462616336724872265004463889617697351427578319298375193703917734724591413551721265144762523011812455166834567160307410948334719671153969850940673704935794016264663402642718236874157608185239184357748300189335228689193799229507555084502951456104676091;
            6'd22: xpb[118] = 1024'd74553366312035391684813912004214102497155418306092069507931014664250919962556425317412476982365592979984926699952687942744682097911688565484006929790678386648372114661664479384125942808660410555456280022468191740311618461723024782809576327879973902745561423004231796343419115810791474491170057328180374751428;
            6'd23: xpb[118] = 1024'd111778527240071020779250615478445952450125690172478713793236566712165115052847846170935336267379758381650555024711671967754639604409825409702869097058344960841577394756168651357303550897649667141061619371231447686606972260043406847382278498151762566306765097708274257458149037822353441427255611704904644826765;
            6'd24: xpb[118] = 1024'd24936992483981908474888391547863369658397534913129673950410263695102414805830128114443124337736249473873033942013162558185533270066741919366571139309680494101092000281101605992850919795121718005356761111607463786537965208142892138990002098740321780601148868998199660542772431759986775346222476255003320417771;
            6'd25: xpb[118] = 1024'd62162153412017537569325095022095219611367806779516318235715815743016609896121548967965983622750414875538662266772146583195490776564878763585433306577347068294297280375605777966028527884110974590962100460370719732833319006463274203562704269012110444162352543702242121657502353771548742282308030631727590493108;
            6'd26: xpb[118] = 1024'd99387314340053166663761798496327069564338078645902962521021367790930804986412969821488842907764580277204290591531130608205448283063015607804295473845013642487502560470109949939206135973100231176567439809133975679128672804783656268135406439283899107723556218406284582772232275783110709218393585008451860568445;
            6'd27: xpb[118] = 1024'd12545779583964054359399574565744486772609923386553922678195064773868104739395251764996630978121071369426769508832621198636341948719932117467997516096349175747017165995042904574753504870572282040862581549509991779059665752883141559743130039872458322017939989696209985856855669720744043137360449558550536159451;
            6'd28: xpb[118] = 1024'd49770940511999683453836278039976336725580195252940566963500616821782299829686672618519490263135236771092397833591605223646299455218068961686859683364015749940222446089547076547931112959561538626467920898273247725355019551203523624315832210144246985579143664400252446971585591732306010073446003935274806234788;
            6'd29: xpb[118] = 1024'd86996101440035312548272981514208186678550467119327211248806168869696494919978093472042349548149402172758026158350589248656256961716205805905721850631682324133427726184051248521108721048550795212073260247036503671650373349523905688888534380416035649140347339104294908086315513743867977009531558311999076310125;
            6'd30: xpb[118] = 1024'd154566683946200243910757583625603886822311859978171405979865852633794672960375415550137618505893264980505075652079839087150627373122315569423892883017857392942331708984203156656089946022846076368401987412519771581366297623390980496257981004594863434731110394220311170938907681501310928498422862097751901131;
            6'd31: xpb[118] = 1024'd37379727611981829338347461057857453839792583726364815691285417900547989763251796269072996903520058666646133400411063864097108133871259159788286060150684431586147611803488375129833698035012102661973741336175775717876720095943773045068960151276383526995934785098262772285668829693063277864583977238822021976468;
            6'd32: xpb[118] = 1024'd74604888540017458432784164532089303792762855592751459976590969948462184853543217122595856188534224068311761725170047889107065640369396004007148227418351005779352891897992547103011306124001359247579080684939031664172073894264155109641662321548172190557138459802305233400398751704625244800669531615546292051805;
            6'd33: xpb[118] = 1024'd111830049468053087527220868006321153745733127459138104261896521996376379943834637976118715473548389469977390049929031914117023146867532848226010394686017579972558171992496719076188914212990615833184420033702287610467427692584537174214364491819960854118342134506347694515128673716187211736755085992270562127142;
            6'd34: xpb[118] = 1024'd24988514711963975222858644075738570954004972199789064419070218979313679696816919919626503543904880562199868967230522504547916812524449357889712436937353113232072777517429673711736283110462666697479561774078303710398420640684022465822088092408520068412725905796273097599752067653820545655721950542369237718148;
            6'd35: xpb[118] = 1024'd62213675639999604317295347549970420906975244066175708704375771027227874787108340773149362828919045963865497291989506529557874319022586202108574604205019687425278057611933845684913891199451923283084901122841559656693774439004404530394790262680308731973929580500315558714481989665382512591807504919093507793485;
            6'd36: xpb[118] = 1024'd99438836568035233411732051024202270859945515932562352989681323075142069877399761626672222113933211365531125616748490554567831825520723046327436771472686261618483337706438017658091499288441179868690240471604815602989128237324786594967492432952097395535133255204358019829211911676944479527893059295817777868822;
            6'd37: xpb[118] = 1024'd12597301811946121107369827093619688068217360673213313146855020058079369630382043570180010184289702457753604534049981144998725491177639555991138813724021794877997943231370972293638868185913230732985382211980831702920121185424271886575216033540656609829517026494283422913835305614577813446859923845916453459828;
            6'd38: xpb[118] = 1024'd49822462739981750201806530567851538021187632539599957432160572105993564720673464423702869469303867859419232858808965170008682997675776400210000980991688369071203223325875144266816476274902487318590721560744087649215474983744653951147918203812445273390720701198325884028565227626139780382945478222640723535165;
            6'd39: xpb[118] = 1024'd87047623668017379296243234042083387974157904405986601717466124153907759810964885277225728754318033261084861183567949195018640504173913244428863148259354943264408503420379316239994084363891743904196060909507343595510828782065036015720620374084233936951924375902368345143295149637701747319031032599364993610502;
            6'd40: xpb[118] = 1024'd206088911928266991881010111500805182429749146637561874639821136845059563947167220733516824674524353307340100869439785449534169830829754092565190510690476523923108945312270875541453261363794768491202649883359695441821730164521307328343974672793151246308147192293748227918543575335081237997897149463669201508;
            6'd41: xpb[118] = 1024'd37431249839963896086317713585732655135400021013024206159945373184759254654238588074256376109688689754972968425628423810459491676328966598311427357778357050717128389039816442848719061350353051354096541998646615641737175528484903371901046144944581814807511821896336209342648465586897048174083451526187939276845;
            6'd42: xpb[118] = 1024'd74656410767999525180754417059964505088370292879410850445250925232673449744530008927779235394702855156638596750387407835469449182827103442530289525046023624910333669134320614821896669439342307939701881347409871588032529326805285436473748315216370478368715496600378670457378387598459015110169005902912209352182;
            6'd43: xpb[118] = 1024'd111881571696035154275191120534196355041340564745797494730556477280587644834821429781302094679717020558304225075146391860479406689325240286749151692313690199103538949228824786795074277528331564525307220696173127534327883125125667501046450485488159141929919171304421131572108309610020982046254560279636479427519;
            6'd44: xpb[118] = 1024'd25040036939946041970828896603613772249612409486448454887730174263524944587803711724809882750073511650526703992447882450910300354982156796412853734565025732363053554753757741430621646425803615389602362436549143634258876073225152792654174086076718356224302942594346534656731703547654315965221424829735155018525;
            6'd45: xpb[118] = 1024'd62265197867981671065265600077845622202582681352835099173035726311439139678095132578332742035087677052192332317206866475920257861480293640631715901832692306556258834848261913403799254514792871975207701785312399580554229871545534857226876256348507019785506617298388995771461625559216282901306979206459425093862;
            6'd46: xpb[118] = 1024'd99490358796017300159702303552077472155552953219221743458341278359353334768386553431855601320101842453857960641965850500930215367978430484850578069100358880749464114942766085376976862603782128560813041134075655526849583669865916921799578426620295683346710292002431456886191547570778249837392533583183695169199;
            6'd47: xpb[118] = 1024'd12648824039928187855340079621494889363824797959872703615514975342290634521368835375363389390458333546080439559267341091361109033635346994514280111351694414008978720467699040012524231501254179425108182874451671626780576617965402213407302027208854897641094063292356859970814941508411583756359398133282370760205;
            6'd48: xpb[118] = 1024'd49873984967963816949776783095726739316795069826259347900820527390204829611660256228886248675472498947746067884026325116371066540133483838733142278619360988202184000562203211985701839590243436010713522223214927573075930416285784277980004197480643561202297737996399321085544863519973550692444952510006640835542;
            6'd49: xpb[118] = 1024'd87099145895999446044213486569958589269765341692645992186126079438119024701951677082409107960486664349411696208785309141381024046631620682952004445887027562395389280656707383958879447679232692596318861571978183519371284214606166342552706367752432224763501412700441782200274785531535517628530506886730910910879;
            6'd50: xpb[118] = 1024'd257611139910333739851262639376006478037186433296952343299776421056324454933959025916896030843155441634175126086799731811917712288537192615706488138363095654903886181640338594426816576704743460614003312354199619302277162705651634160429968340991439057885183990367185284898179469168851547497371436829586501885;
            6'd51: xpb[118] = 1024'd37482772067945962834287966113607856431007458299683596628605328468970519545225379879439755315857320843299803450845783756821875218786674036834568655406029669848109166276144510567604424665694000046219342661117455565597630961026033698733132138612780102619088858694409646399628101480730818483582925813553856577222;
            6'd52: xpb[118] = 1024'd74707932995981591928724669587839706383977730166070240913910880516884714635516800732962614600871486244965431775604767781831832725284810881053430822673696244041314446370648682540782032754683256631824682009880711511892984759346415763305834308884568766180292533398452107514358023492292785419668480190278126652559;
            6'd53: xpb[118] = 1024'd111933093924017221023161373062071556336948002032456885199216432564798909725808221586485473885885651646631060100363751806841790231782947725272292989941362818234519726465152854513959640843672513217430021358643967458188338557666797827878536479156357429741496208102494568629087945503854752355754034567002396727896;
            6'd54: xpb[118] = 1024'd25091559167928108718799149131488973545219846773107845356390129547736209478790503529993261956242142738853539017665242397272683897439864234935995032192698351494034331990085809149507009741144564081725163099019983558119331505766283119486260079744916644035879979392419971713711339441488086274720899117101072318902;
            6'd55: xpb[118] = 1024'd62316720095963737813235852605720823498190118639494489641695681595650404569081924383516121241256308140519167342424226422282641403938001079154857199460364925687239612084589981122684617830133820667330502447783239504414685304086665184058962250016705307597083654096462432828441261453050053210806453493825342394239;
            6'd56: xpb[118] = 1024'd99541881023999366907672556079952673451160390505881133927001233643564599659373345237038980526270473542184795667183210447292598910436137923373719366728031499880444892179094153095862225919123077252935841796546495450710039102407047248631664420288493971158287328800504893943171183464612020146892007870549612469576;
            6'd57: xpb[118] = 1024'd12700346267910254603310332149370090659432235246532094084174930626501899412355627180546768596626964634407274584484701037723492576093054433037421408979367033139959497704027107731409594816595128117230983536922511550641032050506532540239388020877053185452671100090430297027794577402245354065858872420648288060582;
            6'd58: xpb[118] = 1024'd49925507195945883697747035623601940612402507112918738369480482674416094502647048034069627881641130036072902909243685062733450082591191277256283576247033607333164777798531279704587202905584384702836322885685767496936385848826914604812090191148841849013874774794472758142524499413807321001944426797372558135919;
            6'd59: xpb[118] = 1024'd87150668123981512792183739097833790565372778979305382654786034722330289592938468887592487166655295437738531234002669087743407589089328121475145743514700181526370057893035451677764810994573641288441662234449023443231739647147296669384792361420630512575078449498515219257254421425369287938029981174096828211256;
            6'd60: xpb[118] = 1024'd309133367892400487821515167251207773644623719956342811959731705267589345920750831100275237011786529961010151304159678174301254746244631138847785766035714785884663417968406313312179892045692152736803974825039543162732595246781960992515962009189726869462220788440622341877815363002621856996845724195503802262;
            6'd61: xpb[118] = 1024'd37534294295928029582258218641483057726614895586342987097265283753181784436212171684623134522025951931626638476063143703184258761244381475357709953033702288979089943512472578286489787981034948738342143323588295489458086393567164025565218132280978390430665895492483083456607737374564588793082400100919773877599;
            6'd62: xpb[118] = 1024'd74759455223963658676694922115714907679585167452729631382570835801095979526503592538145993807040117333292266800822127728194216267742518319576572120301368863172295223606976750259667396070024205323947482672351551435753440191887546090137920302552767053991869570196525544571337659386126555729167954477644043952936;
            6'd63: xpb[118] = 1024'd111984616151999287771131625589946757632555439319116275667876387849010174616795013391668853092054282734957895125581111753204173774240655163795434287569035437365500503701480922232845004159013461909552822021114807382048793990207928154710622472824555717553073244900568005686067581397688522665253508854368314028273;
        endcase
    end

    always_comb begin
        case(flag[39][16:12])
            5'd0: xpb[119] = 1024'd0;
            5'd1: xpb[119] = 1024'd25143081395910175466769401659364174840827284059767235825050084831947474369777295335176641162410773827180374042882602343635067439897571673459136329820370970625015109226413876868392373056485512773847963761490823481979786938307413446318346073413114931847457016190493408770690975335321856584220373404466989619279;
            5'd2: xpb[119] = 1024'd50286162791820350933538803318728349681654568119534471650100169663894948739554590670353282324821547654360748085765204687270134879795143346918272659640741941250030218452827753736784746112971025547695927522981646963959573876614826892636692146826229863694914032380986817541381950670643713168440746808933979238558;
            5'd3: xpb[119] = 1024'd75429244187730526400308204978092524522481852179301707475150254495842423109331886005529923487232321481541122128647807030905202319692715020377408989461112911875045327679241630605177119169456538321543891284472470445939360814922240338955038220239344795542371048571480226312072926005965569752661120213400968857837;
            5'd4: xpb[119] = 1024'd100572325583640701867077606637456699363309136239068943300200339327789897479109181340706564649643095308721496171530409374540269759590286693836545319281483882500060436905655507473569492225942051095391855045963293927919147753229653785273384293652459727389828064761973635082763901341287426336881493617867958477116;
            5'd5: xpb[119] = 1024'd1648711295426135935048080892006441459437993173100494997118569094760476511577337765868134597396194826458720806955518283596273358646638032740521524085523812191384871562498167004331626090910358147929621199066877563534573841316170458626751797382345209970465177538349985823348348602680649903983177195709353612064;
            5'd6: xpb[119] = 1024'd26791792691336311401817482551370616300265277232867730822168653926707950881354633101044775759806968653639094849838120627231340798544209706199657853905894782816399980788912043872723999147395870921777584960557701045514360779623583904945097870795460141817922193728843394594039323938002506488203550600176343231343;
            5'd7: xpb[119] = 1024'd51934874087246486868586884210734791141092561292634966647218738758655425251131928436221416922217742480819468892720722970866408238441781379658794183726265753441415090015325920741116372203881383695625548722048524527494147717930997351263443944208575073665379209919336803364730299273324363072423924004643332850622;
            5'd8: xpb[119] = 1024'd77077955483156662335356285870098965981919845352402202472268823590602899620909223771398058084628516307999842935603325314501475678339353053117930513546636724066430199241739797609508745260366896469473512483539348009473934656238410797581790017621690005512836226109830212135421274608646219656644297409110322469901;
            5'd9: xpb[119] = 1024'd102221036879066837802125687529463140822747129412169438297318908422550373990686519106574699247039290135180216978485927658136543118236924726577066843367007694691445308468153674477901118316852409243321476245030171491453721594545824243900136091034804937360293242300323620906112249943968076240864670813577312089180;
            5'd10: xpb[119] = 1024'd3297422590852271870096161784012882918875986346200989994237138189520953023154675531736269194792389652917441613911036567192546717293276065481043048171047624382769743124996334008663252181820716295859242398133755127069147682632340917253503594764690419940930355076699971646696697205361299807966354391418707224128;
            5'd11: xpb[119] = 1024'd28440503986762447336865563443377057759703270405968225819287223021468427392931970866912910357203163480097815656793638910827614157190847738940179377991418595007784852351410210877055625238306229069707206159624578609048934620939754363571849668177805351788387371267193380417387672540683156392186727795885696843407;
            5'd12: xpb[119] = 1024'd53583585382672622803634965102741232600530554465735461644337307853415901762709266202089551519613937307278189699676241254462681597088419412399315707811789565632799961577824087745447998294791741843555169921115402091028721559247167809890195741590920283635844387457686789188078647876005012976407101200352686462686;
            5'd13: xpb[119] = 1024'd78726666778582798270404366762105407441357838525502697469387392685363376132486561537266192682024711134458563742558843598097749036985991085858452037632160536257815070804237964613840371351277254617403133682606225573008508497554581256208541815004035215483301403648180197958769623211326869560627474604819676081965;
            5'd14: xpb[119] = 1024'd103869748174492973737173768421469582282185122585269933294437477517310850502263856872442833844435484961638937785441445941732816476883562759317588367452531506882830180030651841482232744407762767391251097444097049054988295435861994702526887888417150147330758419838673606729460598546648726144847848009286665701244;
            5'd15: xpb[119] = 1024'd4946133886278407805144242676019324378313979519301484991355707284281429534732013297604403792188584479376162420866554850788820075939914098221564572256571436574154614687494501012994878272731074443788863597200632690603721523948511375880255392147035629911395532615049957470045045808041949711949531587128060836192;
            5'd16: xpb[119] = 1024'd30089215282188583271913644335383499219141263579068720816405792116228903904509308632781044954599358306556536463749157194423887515837485771680700902076942407199169723913908377881387251329216587217636827358691456172583508462255924822198601465560150561758852548805543366240736021143363806296169904991595050455471;
            5'd17: xpb[119] = 1024'd55232296678098758738683045994747674059968547638835956641455876948176378274286603967957686117010132133736910506631759538058954955735057445139837231897313377824184833140322254749779624385702099991484791120182279654563295400563338268516947538973265493606309564996036775011426996478685662880390278396062040074750;
            5'd18: xpb[119] = 1024'd80375378074008934205452447654111848900795831698603192466505961780123852644063899303134327279420905960917284549514361881694022395632629118598973561717684348449199942366736131618171997442187612765332754881673103136543082338870751714835293612386380425453766581186530183782117971814007519464610651800529029694029;
            5'd19: xpb[119] = 1024'd105518459469919109672221849313476023741623115758370428291556046612071327013841194638310968441831679788097658592396964225329089835530200792058109891538055319074215051593150008486564370498673125539180718643163926618522869277178165161153639685799495357301223597377023592552808947149329376048831025204996019313308;
            5'd20: xpb[119] = 1024'd6594845181704543740192323568025765837751972692401979988474276379041906046309351063472538389584779305834883227822073134385093434586552130962086096342095248765539486249992668017326504363641432591718484796267510254138295365264681834507007189529380839881860710153399943293393394410722599615932708782837414448256;
            5'd21: xpb[119] = 1024'd31737926577614719206961725227389940678579256752169215813524361210989380416086646398649179551995553133015257270704675478020160874484123804421222426162466219390554595476406544885718877420126945365566448557758333736118082303572095280825353262942495771729317726343893352064084369746044456200153082187304404067535;
            5'd22: xpb[119] = 1024'd56881007973524894673731126886754115519406540811936451638574446042936854785863941733825820714406326960195631313587277821655228314381695477880358755982837190015569704702820421754111250476612458139414412319249157218097869241879508727143699336355610703576774742534386760834775345081366312784373455591771393686814;
            5'd23: xpb[119] = 1024'd82024089369435070140500528546118290360233824871703687463624530874884329155641237069002461876817100787376005356469880165290295754279267151339495085803208160640584813929234298622503623533097970913262376080739980700077656180186922173462045409768725635424231758724880169605466320416688169368593828996238383306093;
            5'd24: xpb[119] = 1024'd107167170765345245607269930205482465201061108931470923288674615706831803525418532404179103039227874614556379399352482508925363194176838824798631415623579131265599923155648175490895996589583483687110339842230804182057443118494335619780391483181840567271688774915373578376157295752010025952814202400705372925372;
            5'd25: xpb[119] = 1024'd8243556477130679675240404460032207297189965865502474985592845473802382557886688829340672986980974132293604034777591417981366793233190163702607620427619060956924357812490835021658130454551790739648105995334387817672869206580852293133758986911726049852325887691749929116741743013403249519915885978546768060320;
            5'd26: xpb[119] = 1024'd33386637873040855142009806119396382138017249925269710810642930305749856927663984164517314149391747959473978077660193761616434233130761837161743950247990031581939467038904711890050503511037303513496069756825211299652656144888265739452105060324840981699782903882243337887432718348725106104136259383013757679599;
            5'd27: xpb[119] = 1024'd58529719268951030608779207778760556978844533985036946635693015137697331297441279499693955311802521786654352120542796105251501673028333510620880280068361002206954576265318588758442876567522816287344033518316034781632443083195679185770451133737955913547239920072736746658123693684046962688356632787480747298878;
            5'd28: xpb[119] = 1024'd83672800664861206075548609438124731819671818044804182460743099969644805667218574834870596474213295613834726163425398448886569112925905184080016609888731972831969685491732465626835249624008329061191997279806858263612230021503092632088797207151070845394696936263230155428814669019368819272577006191947736918157;
            5'd29: xpb[119] = 1024'd108815882060771381542318011097488906660499102104571418285793184801592280036995870170047237636624069441015100206308000792521636552823476857539152939709102943456984794718146342495227622680493841835039961041297681745592016959810506078407143280564185777242153952453723564199505644354690675856797379596414726537436;
            5'd30: xpb[119] = 1024'd9892267772556815610288485352038648756627959038602969982711414568562859069464026595208807584377168958752324841733109701577640151879828196443129144513142873148309229374989002025989756545462148887577727194401265381207443047897022751760510784294071259822791065230099914940090091616083899423899063174256121672384;
            5'd31: xpb[119] = 1024'd35035349168466991077057887011402823597455243098370205807761499400510333439241321930385448746787942785932698884615712045212707591777399869902265474333513843773324338601402878894382129601947661661425690955892088863187229986204436198078856857707186191670248081420593323710781066951405756008119436578723111291663;
        endcase
    end

    always_comb begin
        case(flag[40][5:0])
            6'd0: xpb[120] = 1024'd0;
            6'd1: xpb[120] = 1024'd30089215282188583271913644335383499219141263579068720816405792116228903904509308632781044954599358306556536463749157194423887515837485771680700902076942407199169723913908377881387251329216587217636827358691456172583508462255924822198601465560150561758852548805543366240736021143363806296169904991595050455471;
            6'd2: xpb[120] = 1024'd60178430564377166543827288670766998438282527158137441632811584232457807809018617265562089909198716613113072927498314388847775031674971543361401804153884814398339447827816755762774502658433174435273654717382912345167016924511849644397202931120301123517705097611086732481472042286727612592339809983190100910942;
            6'd3: xpb[120] = 1024'd90267645846565749815740933006150497657423790737206162449217376348686711713527925898343134863798074919669609391247471583271662547512457315042102706230827221597509171741725133644161753987649761652910482076074368517750525386767774466595804396680451685276557646416630098722208063430091418888509714974785151366413;
            6'd4: xpb[120] = 1024'd120356861128754333087654577341533996876565054316274883265623168464915615618037234531124179818397433226226145854996628777695550063349943086722803608307769628796678895655633511525549005316866348870547309434765824690334033849023699288794405862240602247035410195222173464962944084573455225184679619966380201821884;
            6'd5: xpb[120] = 1024'd26379380726818174960769294272103063351007890769607919953897105516167624185237404253890153558339117223339532911288292537540373738346208523848344385368380995062157944999970672069306017454565730366873939185070041016553181461058727338028028758117523359527442840613599773173573577642890398463730835131349657793024;
            6'd6: xpb[120] = 1024'd56468596009006758232682938607486562570149154348676640770302897632396528089746712886671198512938475529896069375037449731964261254183694295529045287445323402261327668913879049950693268783782317584510766543761497189136689923314652160226630223677673921286295389419143139414309598786254204759900740122944708248495;
            6'd7: xpb[120] = 1024'd86557811291195341504596582942870061789290417927745361586708689748625431994256021519452243467537833836452605838786606926388148770021180067209746189522265809460497392827787427832080520112998904802147593902452953361720198385570576982425231689237824483045147938224686505655045619929618011056070645114539758703966;
            6'd8: xpb[120] = 1024'd116647026573383924776510227278253561008431681506814082403114481864854335898765330152233288422137192143009142302535764120812036285858665838890447091599208216659667116741695805713467771442215492019784421261144409534303706847826501804623833154797975044804000487030229871895781641072981817352240550106134809159437;
            6'd9: xpb[120] = 1024'd22669546171447766649624944208822627482874517960147119091388418916106344465965499874999262162078876140122529358827427880656859960854931276015987868659819582925146166086032966257224783579914873516111051011448625860522854459861529853857456050674896157296033132421656180106411134142416990631291765271104265130577;
            6'd10: xpb[120] = 1024'd52758761453636349921538588544206126702015781539215839907794211032335248370474808507780307116678234446679065822576585075080747476692417047696688770736761990124315889999941344138612034909131460733747878370140082033106362922117454676056057516235046719054885681227199546347147155285780796927461670262699315586048;
            6'd11: xpb[120] = 1024'd82847976735824933193452232879589625921157045118284560724200003148564152274984117140561352071277592753235602286325742269504634992529902819377389672813704397323485613913849722019999286238348047951384705728831538205689871384373379498254658981795197280813738230032742912587883176429144603223631575254294366041519;
            6'd12: xpb[120] = 1024'd112937192018013516465365877214973125140298308697353281540605795264793056179493425773342397025876951059792138750074899463928522508367388591058090574890646804522655337827758099901386537567564635169021533087522994378273379846629304320453260447355347842572590778838286278828619197572508409519801480245889416496990;
            6'd13: xpb[120] = 1024'd18959711616077358338480594145542191614741145150686318228879732316045064746693595496108370765818635056905525806366563223773346183363654028183631351951258170788134387172095260445143549705264016665348162837827210704492527458664332369686883343232268955064623424229712587039248690641943582798852695410858872468130;
            6'd14: xpb[120] = 1024'd49048926898265941610394238480925690833882408729755039045285524432273968651202904128889415720417993363462062270115720418197233699201139799864332254028200577987304111086003638326530801034480603882984990196518666877076035920920257191885484808792419516823475973035255953279984711785307389095022600402453922923601;
            6'd15: xpb[120] = 1024'd79138142180454524882307882816309190053023672308823759861691316548502872555712212761670460675017351670018598733864877612621121215038625571545033156105142985186473834999912016207918052363697191100621817555210123049659544383176182014084086274352570078582328521840799319520720732928671195391192505394048973379072;
            6'd16: xpb[120] = 1024'd109227357462643108154221527151692689272164935887892480678097108664731776460221521394451505629616709976575135197614034807045008730876111343225734058182085392385643558913820394089305303692913778318258644913901579222243052845432106836282687739912720640341181070646342685761456754072035001687362410385644023834543;
            6'd17: xpb[120] = 1024'd15249877060706950027336244082261755746607772341225517366371045715983785027421691117217479369558393973688522253905698566889832405872376780351274835242696758651122608258157554633062315830613159814585274664205795548462200457467134885516310635789641752833213716037768993972086247141470174966413625550613479805683;
            6'd18: xpb[120] = 1024'd45339092342895533299249888417645254965749035920294238182776837832212688931930999749998524324157752280245058717654855761313719921709862552031975737319639165850292332172065932514449567159829747032222102022897251721045708919723059707714912101349792314592066264843312360212822268284833981262583530542208530261154;
            6'd19: xpb[120] = 1024'd75428307625084116571163532753028754184890299499362958999182629948441592836440308382779569278757110586801595181404012955737607437547348323712676639396581573049462056085974310395836818489046334249858929381588707893629217381978984529913513566909942876350918813648855726453558289428197787558753435533803580716625;
            6'd20: xpb[120] = 1024'd105517522907272699843077177088412253404031563078431679815588422064670496740949617015560614233356468893358131645153170150161494953384834095393377541473523980248631779999882688277224069818262921467495756740280164066212725844234909352112115032470093438109771362454399092694294310571561593854923340525398631172096;
            6'd21: xpb[120] = 1024'd11540042505336541716191894018981319878474399531764716503862359115922505308149786738326587973298152890471518701444833910006318628381099532518918318534135346514110829344219848820981081955962302963822386490584380392431873456269937401345737928347014550601804007845825400904923803640996767133974555690368087143236;
            6'd22: xpb[120] = 1024'd41629257787525124988105538354364819097615663110833437320268151232151409212659095371107632927897511197028055165193991104430206144218585304199619220611077753713280553258128226702368333285178890181459213849275836565015381918525862223544339393907165112360656556651368767145659824784360573430144460681963137598707;
            6'd23: xpb[120] = 1024'd71718473069713708260019182689748318316756926689902158136673943348380313117168404003888677882496869503584591628943148298854093660056071075880320122688020160912450277172036604583755584614395477399096041207967292737598890380781787045742940859467315674119509105456912133386395845927724379726314365673558188054178;
            6'd24: xpb[120] = 1024'd101807688351902291531932827025131817535898190268970878953079735464609217021677712636669722837096227810141128092692305493277981175893556847561021024764962568111620001085944982465142835943612064616732868566658748910182398843037711867941542325027466235878361654262455499627131867071088186022484270665153238509649;
            6'd25: xpb[120] = 1024'd7830207949966133405047543955700884010341026722303915641353672515861225588877882359435696577037911807254515148983969253122804850889822284686561801825573934377099050430282143008899848081311446113059498316962965236401546455072739917175165220904387348370394299653881807837761360140523359301535485830122694480789;
            6'd26: xpb[120] = 1024'd37919423232154716676961188291084383229482290301372636457759464632090129493387190992216741531637270113811051612733126447546692366727308056367262703902516341576268774344190520890287099410528033330696325675654421408985054917328664739373766686464537910129246848459425174078497381283887165597705390821717744936260;
            6'd27: xpb[120] = 1024'd68008638514343299948874832626467882448623553880441357274165256748319033397896499624997786486236628420367588076482283641970579882564793828047963605979458748775438498258098898771674350739744620548333153034345877581568563379584589561572368152024688471888099397264968540319233402427250971893875295813312795391731;
            6'd28: xpb[120] = 1024'd98097853796531883220788476961851381667764817459510078090571048864547937302405808257778831440835986726924124540231440836394467398402279599728664508056401155974608222172007276653061602068961207765969980393037333754152071841840514383770969617584839033646951946070511906559969423570614778190045200804907845847202;
            6'd29: xpb[120] = 1024'd4120373394595725093903193892420448142207653912843114778844985915799945869605977980544805180777670724037511596523104596239291073398545036854205285117012522240087271516344437196818614206660589262296610143341550080371219453875542433004592513461760146138984591461938214770598916640049951469096415969877301818342;
            6'd30: xpb[120] = 1024'd34209588676784308365816838227803947361348917491911835595250778032028849774115286613325850135377029030594048060272261790663178589236030808534906187193954929439256995430252815078205865535877176479933437502033006252954727916131467255203193979021910707897837140267481581011334937783413757765266320961472352273813;
            6'd31: xpb[120] = 1024'd64298803958972891637730482563187446580490181070980556411656570148257753678624595246106895089976387337150584524021418985087066105073516580215607089270897336638426719344161192959593116865093763697570264860724462425538236378387392077401795444582061269656689689073024947252070958926777564061436225953067402729284;
            6'd32: xpb[120] = 1024'd94388019241161474909644126898570945799631444650049277228062362264486657583133903878887940044575745643707120987770576179510953620911002351896307991347839743837596443258069570840980368194310350915207092219415918598121744840643316899600396910142211831415542237878568313492806980070141370357606130944662453184755;
            6'd33: xpb[120] = 1024'd410538839225316782758843829140012274074281103382313916336299315738666150334073601653913784517429640820508044062239939355777295907267789021848768408451110103075492602406731384737380332009732411533721969720134924340892452678344948834019806019132943907574883269994621703436473139576543636657346109631909155895;
            6'd34: xpb[120] = 1024'd30499754121413900054672488164523511493215544682451034732742091431967570054843382234434958739116787947377044507811397133779664811744753560702549670485393517302245216516315109266124631661226319629170549328411591096924400914934269771032621271579283505666427432075537987944172494282940349932827251101226959611366;
            6'd35: xpb[120] = 1024'd60588969403602483326586132499907010712356808261519755549147883548196473959352690867216003693716146253933580971560554328203552327582239332383250572562335924501414940430223487147511882990442906846807376687103047269507909377190194593231222737139434067425279980881081354184908515426304156228997156092822010066837;
            6'd36: xpb[120] = 1024'd90678184685791066598499776835290509931498071840588476365553675664425377863861999499997048648315504560490117435309711522627439843419725104063951474639278331700584664344131865028899134319659494064444204045794503442091417839446119415429824202699584629184132529686624720425644536569667962525167061084417060522308;
            6'd37: xpb[120] = 1024'd120767399967979649870413421170674009150639335419657197181959467780654281768371308132778093602914862867046653899058868717051327359257210875744652376716220738899754388258040242910286385648876081282081031404485959614674926301702044237628425668259735190942985078492168086666380557713031768821336966076012110977779;
            6'd38: xpb[120] = 1024'd26789919566043491743528138101243075625082171872990233870233404831906290335571477855544067342856546864160040955350532476896151034253476312870193153776832105165233437602377403454043397786575462778407661154790175940894073913737072286862048564136656303435017723883594394877010050782466942100388181240981566948919;
            6'd39: xpb[120] = 1024'd56879134848232075015441782436626574844223435452058954686639196948135194240080786488325112297455905170716577419099689671320038550090962084550894055853774512364403161516285781335430649115792049996044488513481632113477582375992997109060650029696806865193870272689137761117746071925830748396558086232576617404390;
            6'd40: xpb[120] = 1024'd86968350130420658287355426772010074063364699031127675503044989064364098144590095121106157252055263477273113882848846865743926065928447856231594957930716919563572885430194159216817900445008637213681315872173088286061090838248921931259251495256957426952722821494681127358482093069194554692727991224171667859861;
            6'd41: xpb[120] = 1024'd117057565412609241559269071107393573282505962610196396319450781180593002049099403753887202206654621783829650346598004060167813581765933627912295860007659326762742609344102537098205151774225224431318143230864544458644599300504846753457852960817107988711575370300224493599218114212558360988897896215766718315332;
            6'd42: xpb[120] = 1024'd23080085010673083432383788037962639756948799063529433007724718231845010616299573476653175946596305780943037402889667820012637256762199065037836637068270693028221658688439697641962163911924605927644772981168760784863746912539874802691475856694029101203608015691650801809847607281993534267949111380736174286472;
            6'd43: xpb[120] = 1024'd53169300292861666704297432373346138976090062642598153824130510348073914520808882109434220901195664087499573866638825014436524772599684836718537539145213100227391382602348075523349415241141193145281600339860216957447255374795799624890077322254179662962460564497194168050583628425357340564119016372331224741943;
            6'd44: xpb[120] = 1024'd83258515575050249976211076708729638195231326221666874640536302464302818425318190742215265855795022394056110330387982208860412288437170608399238441222155507426561106516256453404736666570357780362918427698551673130030763837051724447088678787814330224721313113302737534291319649568721146860288921363926275197414;
            6'd45: xpb[120] = 1024'd113347730857238833248124721044113137414372589800735595456942094580531722329827499374996310810394380700612646794137139403284299804274656380079939343299097914625730830430164831286123917899574367580555255057243129302614272299307649269287280253374480786480165662108280900532055670712084953156458826355521325652885;
            6'd46: xpb[120] = 1024'd19370250455302675121239437974682203888815426254068632145216031631783730897027669097762284550336064697726033850428803163129123479270921817205480120359709280891209879774501991829880930037273749076881884807547345628833419911342677318520903149251401898972198307499707208742685163781520126435510041520490781624025;
            6'd47: xpb[120] = 1024'd49459465737491258393153082310065703107956689833137352961621823748012634801536977730543329504935423004282570314177960357553010995108407588886181022436651688090379603688410369711268181366490336294518712166238801801416928373598602140719504614811552460731050856305250574983421184924883932731679946512085832079496;
            6'd48: xpb[120] = 1024'd79548681019679841665066726645449202327097953412206073778027615864241538706046286363324374459534781310839106777927117551976898510945893360566881924513594095289549327602318747592655432695706923512155539524930257974000436835854526962918106080371703022489903405110793941224157206068247739027849851503680882534967;
            6'd49: xpb[120] = 1024'd109637896301868424936980370980832701546239216991274794594433407980470442610555594996105419414134139617395643241676274746400786026783379132247582826590536502488719051516227125474042684024923510729792366883621714146583945298110451785116707545931853584248755953916337307464893227211611545324019756495275932990438;
            6'd50: xpb[120] = 1024'd15660415899932266810095087911401768020682053444607831282707345031722451177755764718871393154075823614509030297967938506245609701779644569373123603651147868754198100860564286017799696162622892226118996633925930472803092910145479834350330441808774696740788599307763615675522720281046718603070971660245388961578;
            6'd51: xpb[120] = 1024'd45749631182120850082008732246785267239823317023676552099113137147951355082265073351652438108675181921065566761717095700669497217617130341053824505728090275953367824774472663899186947491839479443755823992617386645386601372401404656548931907368925258499641148113306981916258741424410524899240876651840439417049;
            6'd52: xpb[120] = 1024'd75838846464309433353922376582168766458964580602745272915518929264180258986774381984433483063274540227622103225466252895093384733454616112734525407805032683152537548688381041780574198821056066661392651351308842817970109834657329478747533372929075820258493696918850348156994762567774331195410781643435489872520;
            6'd53: xpb[120] = 1024'd105928061746498016625836020917552265678105844181813993731924721380409162891283690617214528017873898534178639689215410089517272249292101884415226309881975090351707272602289419661961450150272653879029478710000298990553618296913254300946134838489226382017346245724393714397730783711138137491580686635030540327991;
            6'd54: xpb[120] = 1024'd11950581344561858498950737848121332152548680635147030420198658431661171458483860339980501757815582531292026745507073849362095924288367321540767086942586456617186321946626580205718462287972035375356108460304515316772765908948282350179757734366147494509378891115820022608360276780573310770631901799999996299131;
            6'd55: xpb[120] = 1024'd42039796626750441770864382183504831371689944214215751236604450547890075362993168972761546712414940837848563209256231043785983440125853093221467989019528863816356045860534958087105713617188622592992935818995971489356274371204207172378359199926298056268231439921363388849096297923937117066801806791595046754602;
            6'd56: xpb[120] = 1024'd72129011908939025042778026518888330590831207793284472053010242664118979267502477605542591667014299144405099673005388238209870955963338864902168891096471271015525769774443335968492964946405209810629763177687427661939782833460131994576960665486448618027083988726906755089832319067300923362971711783190097210073;
            6'd57: xpb[120] = 1024'd102218227191127608314691670854271829809972471372353192869416034780347883172011786238323636621613657450961636136754545432633758471800824636582869793173413678214695493688351713849880216275621797028266590536378883834523291295716056816775562131046599179785936537532450121330568340210664729659141616774785147665544;
            6'd58: xpb[120] = 1024'd8240746789191450187806387784840896284415307825686229557689971831599891739211955961089610361555341448075023193046209192478582146797090073708410570234025044480174543032688874393637228413321178524593220286683100160742438907751084866009185026923520292277969182923876429541197833280099902938192831939754603636684;
            6'd59: xpb[120] = 1024'd38329962071380033459720032120224395503556571404754950374095763947828795643721264593870655316154699754631559656795366386902469662634575845389111472310967451679344266946597252275024479742537765742230047645374556333325947370007009688207786492483670854036821731729419795781933854423463709234362736931349654092155;
            6'd60: xpb[120] = 1024'd68419177353568616731633676455607894722697834983823671190501556064057699548230573226651700270754058061188096120544523581326357178472061617069812374387909858878513990860505630156411731071754352959866875004066012505909455832262934510406387958043821415795674280534963162022669875566827515530532641922944704547626;
            6'd61: xpb[120] = 1024'd98508392635757200003547320790991393941839098562892392006907348180286603452739881859432745225353416367744632584293680775750244694309547388750513276464852266077683714774414008037798982400970940177503702362757468678492964294518859332604989423603971977554526829340506528263405896710191321826702546914539755003097;
            6'd62: xpb[120] = 1024'd4530912233821041876662037721560460416281935016225428695181285231538612019940051582198718965295100364858019640585344535595068369305812825876054053525463632343162764118751168581555994538670321673830332113061685004712111906553887381838612319480893090046559474731932836474035389779626495105753762079509210974237;
            6'd63: xpb[120] = 1024'd34620127516009625148575682056943959635423198595294149511587077347767515924449360214979763919894458671414556104334501730018955885143298597556754955602406039542332488032659546462943245867886908891467159471753141177295620368809812204037213785041043651805412023537476202714771410922990301401923667071104261429708;
        endcase
    end

    always_comb begin
        case(flag[40][11:6])
            6'd0: xpb[121] = 1024'd0;
            6'd1: xpb[121] = 1024'd64709342798198208420489326392327458854564462174362870327992869463996419828958668847760808874493816977971092568083658924442843400980784369237455857679348446741502211946567924344330497197103496109103986830444597349879128831065737026235815250601194213564264572343019568955507432066354107698093572062699311885179;
            6'd2: xpb[121] = 1024'd5351989912271675442179725379840484964430497222990056527853883863015944320608198785506546534329959646499035728709824414306622961120348403919751590342365852549313749323564631351030755202689786496897776052501954853393896811910577279506651931519158977861709241271922079880908336058779582379068454298773029286027;
            6'd3: xpb[121] = 1024'd70061332710469883862669051772167943818994959397352926855846753327012364149566867633267355408823776624470128296793483338749466362101132773157207448021714299290815961270132555695361252399793282606001762882946552203273025642976314305742467182120353191425973813614941648836415768125133690077162026361472341171206;
            6'd4: xpb[121] = 1024'd10703979824543350884359450759680969928860994445980113055707767726031888641216397571013093068659919292998071457419648828613245922240696807839503180684731705098627498647129262702061510405379572993795552105003909706787793623821154559013303863038317955723418482543844159761816672117559164758136908597546058572054;
            6'd5: xpb[121] = 1024'd75413322622741559304848777152008428783425456620342983383700637190028308470175066418773901943153736270969164025503307753056089323221481177076959038364080151840129710593697187046392007602483069102899538935448507056666922454886891585249119113639512169287683054886863728717324104183913272456230480660245370457233;
            6'd6: xpb[121] = 1024'd16055969736815026326539176139521454893291491668970169583561651589047832961824596356519639602989878939497107186129473242919868883361045211759254771027097557647941247970693894053092265608069359490693328157505864560181690435731731838519955794557476933585127723815766239642725008176338747137205362896319087858081;
            6'd7: xpb[121] = 1024'd80765312535013234747028502531848913747855953843333039911554521053044252790783265204280448477483695917468199754213132167362712284341829580996710628706446004389443459917261818397422762805172855599797314987950461910060819266797468864755771045158671147149392296158785808598232440242692854835298934959018399743260;
            6'd8: xpb[121] = 1024'd21407959649086701768718901519361939857721988891960226111415535452063777282432795142026186137319838585996142914839297657226491844481393615679006361369463410197254997294258525404123020810759145987591104210007819413575587247642309118026607726076635911446836965087688319523633344235118329516273817195092117144108;
            6'd9: xpb[121] = 1024'd86117302447284910189208227911689398712286451066323096439408404916060197111391463989786995011813655563967235482922956581669335245462177984916462219048811856938757209240826449748453518007862642096695091040452416763454716078708046144262422976677830125011101537430707888479140776301472437214367389257791429029287;
            6'd10: xpb[121] = 1024'd26759949561358377210898626899202424822152486114950282639269419315079721603040993927532732671649798232495178643549122071533114805601742019598757951711829262746568746617823156755153776013448932484488880262509774266969484059552886397533259657595794889308546206359610399404541680293897911895342271493865146430135;
            6'd11: xpb[121] = 1024'd91469292359556585631387953291529883676716948289313152967262288779076141431999662775293541546143615210466271211632780995975958206582526388836213809391177709488070958564391081099484273210552428593592867092954371616848612890618623423769074908196989102872810778702629968360049112360252019593435843556564458315314;
            6'd12: xpb[121] = 1024'd32111939473630052653078352279042909786582983337940339167123303178095665923649192713039279205979757878994214372258946485839737766722090423518509542054195115295882495941387788106184531216138718981386656315011729120363380871463463677039911589114953867170255447631532479285450016352677494274410725792638175716162;
            6'd13: xpb[121] = 1024'd96821282271828261073567678671370368641147445512303209495116172642092085752607861560800088080473574856965306940342605410282581167702874792755965399733543562037384707887955712450515028413242215090490643145456326470242509702529200703275726839716148080734520019974552048240957448419031601972504297855337487601341;
            6'd14: xpb[121] = 1024'd37463929385901728095258077658883394751013480560930395694977187041111610244257391498545825740309717525493250100968770900146360727842438827438261132396560967845196245264952419457215286418828505478284432367513683973757277683374040956546563520634112845031964688903454559166358352411457076653479180091411205002189;
            6'd15: xpb[121] = 1024'd102173272184099936515747404051210853605577942735293266022970056505108030073216060346306634614803534503464342669052429824589204128823223196675716990075909414586698457211520343801545783615932001587388419197958281323636406514439777982782378771235307058596229261246474128121865784477811184351572752154110516887368;
            6'd16: xpb[121] = 1024'd42815919298173403537437803038723879715443977783920452222831070904127554564865590284052372274639677171992285829678595314452983688962787231358012722738926820394509994588517050808246041621518291975182208420015638827151174495284618236053215452153271822893673930175376639047266688470236659032547634390184234288216;
            6'd17: xpb[121] = 1024'd107525262096371611957927129431051338570008439958283322550823940368123974393824259131813181149133494149963378397762254238895827089943571600595468580418275267136012206535084975152576538818621788084286195250460236177030303326350355262289030702754466036457938502518396208002774120536590766730641206452883546173395;
            6'd18: xpb[121] = 1024'd48167909210445078979617528418564364679874475006910508750684954767143498885473789069558918808969636818491321558388419728759606650083135635277764313081292672943823743912081682159276796824208078472079984472517593680545071307195195515559867383672430800755383171447298718928175024529016241411616088688957263574243;
            6'd19: xpb[121] = 1024'd112877252008643287400106854810891823534438937181273379078677824231139918714432457917319727683463453796462414126472078653202450051063920004515220170760641119685325955858649606503607294021311574581183971302962191030424200138260932541795682634273625014319647743790318287883682456595370349109709660751656575459422;
            6'd20: xpb[121] = 1024'd53519899122716754421797253798404849644304972229900565278538838630159443206081987855065465343299596464990357287098244143066229611203484039197515903423658525493137493235646313510307552026897864968977760525019548533938968119105772795066519315191589778617092412719220798809083360587795823790684542987730292860270;
            6'd21: xpb[121] = 1024'd118229241920914962842286580190732308498869434404263435606531708094155863035040656702826274217793413442961449855181903067509073012184268408434971761103006972234639705182214237854638049224001361078081747355464145883818096950171509821302334565792783992181356985062240367764590792654149931488778115050429604745449;
            6'd22: xpb[121] = 1024'd58871889034988429863976979178245334608735469452890621806392722493175387526690186640572011877629556111489393015808068557372852572323832443117267493766024378042451242559210944861338307229587651465875536577521503387332864931016350074573171246710748756478801653991142878689991696646575406169752997286503322146297;
            6'd23: xpb[121] = 1024'd123581231833186638284466305570572793463299931627253492134385591957171807355648855488332820752123373089460485583891727481815695973304616812354723351445372824783953454505778869205668804426691147574979523407966100737211993762082087100808986497311942970043066226334162447645499128712929513867846569349202634031476;
            6'd24: xpb[121] = 1024'd64223878947260105306156704558085819573165966675880678334246606356191331847298385426078558411959515757988428744517892971679475533444180847037019084108390230591764991882775576212369062432277437962773312630023458240726761742926927354079823178229907734340510895263064958570900032705354988548821451585276351432324;
            6'd25: xpb[121] = 1024'd4866526061333572327847103545598845683032001724507864534107620755210856338947915363824296071795658426516371905144058461543255093583744881719314816771407636399576529259772283219069320437863728350567101852080815744241529723771767607350659859147872498637955564191967469496300936697780463229796333821350068833172;
            6'd26: xpb[121] = 1024'd69575868859531780748336429937926304537596463898870734862100490219207276167906584211585104946289475404487464473227717385986098494564529250956770674450756083141078741206340207563399817634967224459671088682525413094120658554837504633586475109749066712202220136534987038451808368764134570927889905884049380718351;
            6'd27: xpb[121] = 1024'd10218515973605247770026828925439330647462498947497921061961504618226800659556114149330842606125618073015407633853882875849878054704093285639066407113773488948890278583336914570100075640553514847464877904582770597635426535682344886857311790667031476499664805463889549377209272756560045608864788120123098119199;
            6'd28: xpb[121] = 1024'd74927858771803456190516155317766789502026961121860791389954374082223220488514782997091651480619435050986500201937541800292721455684877654876522264793121935690392490529904838914430572837657010956568864735027367947514555366748081913093127041268225690063929377806909118332716704822914153306958360182822410004378;
            6'd29: xpb[121] = 1024'd15570505885876923212206554305279815611892996170487977589815388481242744980164312934837389140455577719514443362563707290156501015824441689558817997456139341498204027906901545921130830843243301344362653957084725451029323347592922166363963722186190454361374046735811629258117608815339627987933242418896127405226;
            6'd30: xpb[121] = 1024'd80279848684075131632695880697607274466457458344850847917808257945239164809122981782598198014949394697485535930647366214599344416805226058796273855135487788239706239853469470265461328040346797453466640787529322800908452178658659192599778972787384667925638619078831198213625040881693735686026814481595439290405;
            6'd31: xpb[121] = 1024'd20922495798148598654386279685120300576323493393478034117669272344258689300772511720343935674785537366013479091273531704463123976944790093478569587798505194047517777230466177272161586045933087841260430009586680304423220159503499445870615653705349432223083288007733709139025944874119210367001696717669156691253;
            6'd32: xpb[121] = 1024'd85631838596346807074875606077447759430887955567840904445662141808255109129731180568104744549279354343984571659357190628905967377925574462716025445477853640789019989177034101616492083243036583950364416840031277654302348990569236472106430904306543645787347860350753278094533376940473318065095268780368468576432;
            6'd33: xpb[121] = 1024'd26274485710420274096566005064960785540753990616468090645523156207274633621380710505850482209115497012512514819983356118769746938065138497398321178140871046596831526554030808623192341248622874338158206062088635157817116971414076725377267585224508410084792529279655789019934280932898792746070151016442185977280;
            6'd34: xpb[121] = 1024'd90983828508618482517055331457288244395318452790830960973516025671271053450339379353611291083609313990483607388067015043212590339045922866635777035820219493338333738500598732967522838445726370447262192892533232507696245802479813751613082835825702623649057101622675357975441712999252900444163723079141497862459;
            6'd35: xpb[121] = 1024'd31626475622691949538745730444801270505184487839458147173377040070290577941988909291357028743445456659011550548693180533076369899185486901318072768483236899146145275877595439974223096451312660835055982114590590011211013783324654004883919516743667387946501770551577868900842616991678375125138605315215215263307;
            6'd36: xpb[121] = 1024'd96335818420890157959235056837128729359748950013821017501369909534286997770947578139117837617939273636982643116776839457519213300166271270555528626162585345887647487824163364318553593648416156944159968945035187361090142614390391031119734767344861601510766342894597437856350049058032482823232177377914527148486;
            6'd37: xpb[121] = 1024'd36978465534963624980925455824641755469614985062448203701230923933306522262597108076863575277775416305510586277403004947382992860305835305237824358825602751695459025201160071325253851654002447331953758167092544864604910595235231284390571448262826365808211011823499948781750953050457957504207059613988244549334;
            6'd38: xpb[121] = 1024'd101687808333161833401414782216969214324179447236811074029223793397302942091555776924624384152269233283481678845486663871825836261286619674475280216504951198436961237147727995669584348851105943441057744997537142214484039426300968310626386698864020579372475584166519517737258385116812065202300631676687556434513;
            6'd39: xpb[121] = 1024'd42330455447235300423105181204482240434045482285438260229084807796322466583205306862370121812105375952009622006112829361689615821426183709157575949167968604244772774524724702676284606856692233828851534219594499717998807407145808563897223379781985343669920253095422028662659289109237539883275513912761273835361;
            6'd40: xpb[121] = 1024'd107039798245433508843594507596809699288609944459801130557077677260318886412163975710130930686599192929980714574196488286132459222406968078395031806847317050986274986471292627020615104053795729937955521050039097067877936238211545590133038630383179557234184825438441597618166721175591647581369085975460585720540;
            6'd41: xpb[121] = 1024'd47682445359506975865284906584322725398475979508428316756938691659338410903813505647876668346435335598508657734822653775996238782546532113077327539510334456794086523848289334027315362059382020325749310272096454571392704219056385843403875311301144321531629494367344108543567625168017122262343968211534303121388;
            6'd42: xpb[121] = 1024'd112391788157705184285774232976650184253040441682791187084931561123334830732772174495637477220929152576479750302906312700439082183527316482314783397189682903535588735794857258371645859256485516434853297102541051921271833050122122869639690561902338535095894066710363677499075057234371229960437540274233615006567;
            6'd43: xpb[121] = 1024'd53034435271778651307464631964163210362906476731418373284792575522354355224421704433383214880765295245007693463532478190302861743666880516997079129852700309343400273171853965378346117262071806822647086324598409424786601030966963122910527242820303299393338735639266188424475961226796704641412422510307332407415;
            6'd44: xpb[121] = 1024'd117743778069976859727953958356490669217470938905781243612785444986350775053380373281144023755259112222978786031616137114745705144647664886234534987532048756084902485118421889722676614459175302931751073155043006774665729862032700149146342493421497512957603307982285757379983393293150812339505994573006644292594;
            6'd45: xpb[121] = 1024'd58386425184050326749644357344003695327336973954408429812646459385370299545029903218889761415095254891506729192242302604609484704787228920916830720195066161892714022495418596729376872464761593319544862377100364278180497842877540402417179174339462277255047976911188268305384297285576287020480876809080361693442;
            6'd46: xpb[121] = 1024'd123095767982248535170133683736331154181901436128771300140639328849366719373988572066650570289589071869477821760325961529052328105768013290154286577874414608634216234441986521073707369661865089428648849207544961628059626673943277428652994424940656490819312549254207837260891729351930394718574448871779673578621;
            6'd47: xpb[121] = 1024'd63738415096322002191824082723844180291767471177398486340500343248386243865638102004396307949425214538005764920952127018916107665907577324836582310537432014442027771818983228080407627667451379816442638429602319131574394654788117681923831105858621255116757218183110348186292633344355869399549331107853390979469;
            6'd48: xpb[121] = 1024'd4381062210395469213514481711357206401633506226025672540361357647405768357287631942142045609261357206533708081578292508779887226047141359518878043200449420249839309195979935087107885673037670204236427651659676635089162635632957935194667786776586019414201887112012859111693537336781344080524213343927108380317;
            6'd49: xpb[121] = 1024'd69090405008593677634003808103684665256197968400388542868354227111402188186246300789902854483755174184504800649661951433222730627027925728756333900879797866991341521142547859431438382870141166313340414482104273984968291466698694961430483037377780232978466459455032428067200969403135451778617785406626420265496;
            6'd50: xpb[121] = 1024'd9733052122667144655694207091197691366064003449015729068215241510421712677895830727648592143591316853032743810288116923086510187167489763438629633542815272799153058519544566438138640875727456701134203704161631488483059447543535214701319718295744997275911128383934938992601873395560926459592667642700137666344;
            6'd51: xpb[121] = 1024'd74442394920865353076183533483525150220628465623378599396208110974418132506854499575409401018085133831003836378371775847529353588148274132676085491222163719540655270466112490782469138072830952810238190534606228838362188278609272240937134968896939210840175700726954507948109305461915034157686239705399449551523;
            6'd52: xpb[121] = 1024'd15085042034938820097873932471038176330494500672005785596069125373437656998504029513155138677921276499531779538997941337393133148287838167358381223885181125348466807843109197789169396078417243198031979756663586341876956259454112494207971649814903975137620369655857018873510209454340508838661121941473166952371;
            6'd53: xpb[121] = 1024'd79794384833137028518363258863365635185058962846368655924061994837434076827462698360915947552415093477502872107081600261835976549268622536595837081564529572089969019789677122133499893275520739307135966587108183691756085090519849520443786900416098188701884941998876587829017641520694616536754694004172478837550;
            6'd54: xpb[121] = 1024'd20437031947210495540053657850878661294924997894995842123923009236453601319112228298661685212251236146030815267707765751699756109408186571278132814227546977897780557166673829140200151281107029694929755809165541195270853071364689773714623581334062952999329610927779098754418545513120091217729576240246196238398;
            6'd55: xpb[121] = 1024'd85146374745408703960542984243206120149489460069358712451915878700450021148070897146422494086745053124001907835791424676142599510388970940515588671906895424639282769113241753484530648478210525804033742639610138545149981902430426799950438831935257166563594183270798667709925977579474198915823148302945508123577;
            6'd56: xpb[121] = 1024'd25789021859482170982233383230719146259355495117985898651776893099469545639720427084168231746581195792529850996417590166006379070528534975197884404569912830447094306490238460491230906483796816191827531861667496048664749883275267053221275512853221930861038852199701178635326881571899673596798030539019225524425;
            6'd57: xpb[121] = 1024'd90498364657680379402722709623046605113919957292348768979769762563465965468679095931929040621075012770500943564501249090449222471509319344435340262249261277188596518436806384835561403680900312300931518692112093398543878714341004079457090763454416144425303424542720747590834313638253781294891602601718537409604;
            6'd58: xpb[121] = 1024'd31141011771753846424413108610559631223785992340975955179630776962485489960328625869674778280911155439028886725127414580313002031648883379117635994912278682996408055813803091842261661686486602688725307914169450902058646695185844332727927444372380908722748093471623258516235217630679255975866484837792254810452;
            6'd59: xpb[121] = 1024'd95850354569952054844902435002887090078350454515338825507623646426481909789287294717435587155404972416999979293211073504755845432629667748355091852591627129737910267760371016186592158883590098797829294744614048251937775526251581358963742694973575122287012665814642827471742649697033363673960056900491566695631;
            6'd60: xpb[121] = 1024'd36493001684025521866592833990400116188216489563966011707484660825501434280936824655181324815241115085527922453837238994619624992769231783037387585254644535545721805137367723193292416889176389185623083966671405755452543507096421612234579375891539886584457334743545338397143553689458838354934939136565284096479;
            6'd61: xpb[121] = 1024'd101202344482223730287082160382727575042780951738328882035477530289497854109895493502942133689734932063499015021920897919062468393750016152274843442933992982287224017083935647537622914086279885294727070797116003105331672338162158638470394626492734100148721907086564907352650985755812946053028511199264595981658;
            6'd62: xpb[121] = 1024'd41844991596297197308772559370240601152646986786956068235338544688517378601545023440687871349571074732026958182547063408926247953889580186957139175597010388095035554460932354544323172091866175682520860019173360608846440319006998891741231307410698864446166576015467418278051889748238420734003393435338313382506;
            6'd63: xpb[121] = 1024'd106554334394495405729261885762568060007211448961318938563331414152513798430503692288448680224064891709998050750630722333369091354870364556194595033276358834836537766407500278888653669288969671791624846849617957958725569150072735917977046558011893078010431148358486987233559321814592528432096965498037625267685;
        endcase
    end

    always_comb begin
        case(flag[40][16:12])
            5'd0: xpb[122] = 1024'd0;
            5'd1: xpb[122] = 1024'd47196981508568872750952284750081086117077484009946124763192428551533322922153222226194417883901034378525993911256887823232870915009928590876890765939376240644349303784496985895353927294555962179418636071675315462240337130917576171247883238929857842307875817287389498158960225807018003113071847734111342668533;
            5'd2: xpb[122] = 1024'd94393963017137745501904569500162172234154968019892249526384857103066645844306444452388835767802068757051987822513775646465741830019857181753781531878752481288698607568993971790707854589111924358837272143350630924480674261835152342495766477859715684615751634574778996317920451614036006226143695468222685337066;
            5'd3: xpb[122] = 1024'd17524248841581876854057926845428825606534024904102690161445430589623073429150527768568182437045428826134832326313170035119548904188565438075512172801797680999357236783919740348431542692150680816945710606638706540356650542531831740778671147106344077656807548448051436446774149347125376322096853375708433521268;
            5'd4: xpb[122] = 1024'd64721230350150749605010211595509911723611508914048814924637859141156396351303749994762600320946463204660826237570057858352419819198494028952402938741173921643706540568416726243785469986706642996364346678314022002596987673449407912026554386036201919964683365735440934605734375154143379435168701109819776189801;
            5'd5: xpb[122] = 1024'd111918211858719622355962496345590997840688992923994939687830287692689719273456972220957018204847497583186820148826945681585290734208422619829293704680550162288055844352913712139139397281262605175782982749989337464837324804366984083274437624966059762272559183022830432764694600961161382548240548843931118858334;
            5'd6: xpb[122] = 1024'd35048497683163753708115853690857651213068049808205380322890861179246146858301055537136364874090857652269664652626340070239097808377130876151024345603595361998714473567839480696863085384301361633891421213277413080713301085063663481557342294212688155313615096896102872893548298694250752644193706751416867042536;
            5'd7: xpb[122] = 1024'd82245479191732626459068138440938737330145533818151505086083289730779469780454277763330782757991892030795658563883227893471968723387059467027915111542971602643063777352336466592217012678857323813310057284952728542953638215981239652805225533142545997621490914183492371052508524501268755757265554485528209711069;
            5'd8: xpb[122] = 1024'd5375765016176757811221495786205390702524590702361945721143863217335897365298361079510129427235252099878503067682622282125775797555767723349645752466016802353722406567262235149940700781896080271418495748240804158829614496677919051088130202389174390662546828056764811181362222234358125853218712393013957895271;
            5'd9: xpb[122] = 1024'd52572746524745630562173780536286476819602074712308070484336291768869220287451583305704547311136286478404496978939510105358646712565696314226536518405393042998071710351759221045294628076452042450837131819916119621069951627595495222336013441319032232970422645344154309340322448041376128966290560127125300563804;
            5'd10: xpb[122] = 1024'd99769728033314503313126065286367562936679558722254195247528720320402543209604805531898965195037320856930490890196397928591517627575624905103427284344769283642421014136256206940648555371008004630255767891591435083310288758513071393583896680248890075278298462631543807499282673848394132079362407861236643232337;
            5'd11: xpb[122] = 1024'd22900013857758634665279422631634216309058615606464635882589293806958970794448888848078311864280680926013335393995792317245324701744333161425157925267814483353079643351181975498372243474046761088364206354879510699186265039209750791866801349495518468319354376504816247628136371581483502175315565768722391416539;
            5'd12: xpb[122] = 1024'd70096995366327507416231707381715302426136099616410760645781722358492293716602111074272729748181715304539329305252680140478195616754261752302048691207190723997428947135678961393726170768602723267782842426554826161426602170127326963114684588425376310627230193792205745787096597388501505288387413502833734085072;
            5'd13: xpb[122] = 1024'd117293976874896380167183992131796388543213583626356885408974150910025616638755333300467147632082749683065323216509567963711066531764190343178939457146566964641778250920175947289080098063158685447201478498230141623666939301044903134362567827355234152935106011079595243946056823195519508401459261236945076753605;
            5'd14: xpb[122] = 1024'd40424262699340511519337349477063041915592640510567326044034724396582044223599416616646494301326109752148167720308962352364873605932898599500670098069612164352436880135101715846803786166197441905309916961518217239542915581741582532645472496601862545976161924952867684074910520928608878497412419144430824937807;
            5'd15: xpb[122] = 1024'd87621244207909384270289634227144128032670124520513450807227152948115367145752638842840912185227144130674161631565850175597744520942827190377560864008988404996786183919598701742157713460753404084728553033193532701783252712659158703893355735531720388284037742240257182233870746735626881610484266878542167606340;
            5'd16: xpb[122] = 1024'd10751530032353515622442991572410781405049181404723891442287726434671794730596722159020258854470504199757006135365244564251551595111535446699291504932033604707444813134524470299881401563792160542836991496481608317659228993355838102176260404778348781325093656113529622362724444468716251706437424786027915790542;
            5'd17: xpb[122] = 1024'd57948511540922388373395276322491867522126665414670016205480154986205117652749944385214676738371538578283000046622132387484422510121464037576182270871409845351794116919021456195235328858348122722255627568156923779899566124273414273424143643708206623632969473400919120521684670275734254819509272520139258459075;
            5'd18: xpb[122] = 1024'd105145493049491261124347561072572953639204149424616140968672583537738440574903166611409094622272572956808993957879020210717293425131392628453073036810786085996143420703518442090589256152904084901674263639832239242139903255190990444672026882638064465940845290688308618680644896082752257932581120254250601127608;
            5'd19: xpb[122] = 1024'd28275778873935392476500918417839607011583206308826581603733157024294868159747249927588441291515933025891838461678414599371100499300100884774803677733831285706802049918444210648312944255942841359782702103120314858015879535887669842954931551884692858981901204561581058809498593815841628028534278161736349311810;
            5'd20: xpb[122] = 1024'd75472760382504265227453203167920693128660690318772706366925585575828191081900472153782859175416967404417832372935302422603971414310029475651694443673207526351151353702941196543666871550498803539201338174795630320256216666805246014202814790814550701289777021848970556968458819622859631141606125895847691980343;
            5'd21: xpb[122] = 1024'd122669741891073137978405487918001779245738174328718831130118014127361514004053694379977277059318001782943826284192190245836842329319958066528585209612583766995500657487438182439020798845054765718619974246470945782496553797722822185450698029744408543597652839136360055127419045429877634254677973629959034648876;
            5'd22: xpb[122] = 1024'd45800027715517269330558845263268432618117231212929271765178587613917941588897777696156623728561361852026670787991584634490649403488666322850315850535628966706159286702363950996744486948093522176728412709759021398372530078419501583733602698991036936638708753009632495256272743162967004350631131537444782833078;
            5'd23: xpb[122] = 1024'd92997009224086142081511130013349518735194715222875396528371016165451264511050999922351041612462396230552664699248472457723520318498594913727206616475005207350508590486860936892098414242649484356147048781434336860612867209337077754981485937920894778946584570297021993415232968969985007463702979271556125501611;
            5'd24: xpb[122] = 1024'd16127295048530273433664487358616172107573772107085837163431589652007692095895083238530388281705756299635509203047866846377327392667303170048937257398050407061167219701786705449822102345688240814255487244722412476488843490033757153264390607167523171987640484170294433544086666703074377559656137179041873685813;
            5'd25: xpb[122] = 1024'd63324276557099146184616772108697258224651256117031961926624018203541015018048305464724806165606790678161503114304754669610198307677231760925828023337426647705516523486283691345176029640244202993674123316397727938729180620951333324512273846097381014295516301457683931703046892510092380672727984913153216354346;
            5'd26: xpb[122] = 1024'd110521258065668018935569056858778344341728740126978086689816446755074337940201527690919224049507825056687497025561642492843069222687160351802718789276802888349865827270780677240529956934800165173092759388073043400969517751868909495760157085027238856603392118745073429862007118317110383785799832647264559022879;
            5'd27: xpb[122] = 1024'd33651543890112150287722414204044997714107797011188527324877020241630765525045611007098570718751185125770341529361036881496876296855868608124449430199848088060524456485706445798253645037838921631201197851361119016845494032565588894043061754273867249644448032618345869990860816050199753881752990554750307207081;
            5'd28: xpb[122] = 1024'd80848525398681023038674698954126083831185281021134652088069448793164088447198833233292988602652219504296335440617924704729747211865797199001340196139224328704873760270203431693607572332394883810619833923036434479085831163483165065290944993203725091952323849905735368149821041857217756994824838288861649875614;
            5'd29: xpb[122] = 1024'd3978811223125154390828056299392737203564337905345092723130022279720516032042916549472335271895579573379179944417319093383554286034505455323070837062269528415532389485129200251331260435433640268728272386324510094961807444179844463573849662450353484993379763779007808278674739590307127090777996196347398059816;
            5'd30: xpb[122] = 1024'd51175792731694027141780341049473823320641821915291217486322450831253838954196138775666753155796613951905173855674206916616425201044434046199961603001645769059881693269626186146685187729989602448146908457999825557202144575097420634821732901380211327301255581066397306437634965397325130203849843930458740728349;
            5'd31: xpb[122] = 1024'd98372774240262899892732625799554909437719305925237342249514879382787161876349361001861171039697648330431167766931094739849296116054362637076852368941022009704230997054123172042039115024545564627565544529675141019442481706014996806069616140310069169609131398353786804596595191204343133316921691664570083396882;
        endcase
    end

    always_comb begin
        case(flag[41][5:0])
            6'd0: xpb[123] = 1024'd0;
            6'd1: xpb[123] = 1024'd10751530032353515622442991572410781405049181404723891442287726434671794730596722159020258854470504199757006135365244564251551595111535446699291504932033604707444813134524470299881401563792160542836991496481608317659228993355838102176260404778348781325093656113529622362724444468716251706437424786027915790542;
            6'd2: xpb[123] = 1024'd21503060064707031244885983144821562810098362809447782884575452869343589461193444318040517708941008399514012270730489128503103190223070893398583009864067209414889626269048940599762803127584321085673982992963216635318457986711676204352520809556697562650187312227059244725448888937432503412874849572055831581084;
            6'd3: xpb[123] = 1024'd32254590097060546867328974717232344215147544214171674326863179304015384191790166477060776563411512599271018406095733692754654785334606340097874514796100814122334439403573410899644204691376481628510974489444824952977686980067514306528781214335046343975280968340588867088173333406148755119312274358083747371626;
            6'd4: xpb[123] = 1024'd43006120129414062489771966289643125620196725618895565769150905738687178922386888636081035417882016799028024541460978257006206380446141786797166019728134418829779252538097881199525606255168642171347965985926433270636915973423352408705041619113395125300374624454118489450897777874865006825749699144111663162168;
            6'd5: xpb[123] = 1024'd53757650161767578112214957862053907025245907023619457211438632173358973652983610795101294272352520998785030676826222821257757975557677233496457524660168023537224065672622351499407007818960802714184957482408041588296144966779190510881302023891743906625468280567648111813622222343581258532187123930139578952710;
            6'd6: xpb[123] = 1024'd64509180194121093734657949434464688430295088428343348653726358608030768383580332954121553126823025198542036812191467385509309570669212680195749029592201628244668878807146821799288409382752963257021948978889649905955373960135028613057562428670092687950561936681177734176346666812297510238624548716167494743252;
            6'd7: xpb[123] = 1024'd75260710226474609357100941006875469835344269833067240096014085042702563114177055113141811981293529398299042947556711949760861165780748126895040534524235232952113691941671292099169810946545123799858940475371258223614602953490866715233822833448441469275655592794707356539071111281013761945061973502195410533794;
            6'd8: xpb[123] = 1024'd86012240258828124979543932579286251240393451237791131538301811477374357844773777272162070835764033598056049082921956514012412760892283573594332039456268837659558505076195762399051212510337284342695931971852866541273831946846704817410083238226790250600749248908236978901795555749730013651499398288223326324336;
            6'd9: xpb[123] = 1024'd96763770291181640601986924151697032645442632642515022980589537912046152575370499431182329690234537797813055218287201078263964356003819020293623544388302442367003318210720232698932614074129444885532923468334474858933060940202542919586343643005139031925842905021766601264520000218446265357936823074251242114878;
            6'd10: xpb[123] = 1024'd107515300323535156224429915724107814050491814047238914422877264346717947305967221590202588544705041997570061353652445642515515951115354466992915049320336047074448131345244702998814015637921605428369914964816083176592289933558381021762604047783487813250936561135296223627244444687162517064374247860279157905420;
            6'd11: xpb[123] = 1024'd118266830355888671846872907296518595455540995451962805865164990781389742036563943749222847399175546197327067489017690206767067546226889913692206554252369651781892944479769173298695417201713765971206906461297691494251518926914219123938864452561836594576030217248825845989968889155878768770811672646307073695962;
            6'd12: xpb[123] = 1024'd4951664704117446070516971464114944115891749730951013179320862151084641429851526998228035038988376087640924216925441336439555300497205025836337934168072215555647083044722426260946579573988720792733700349392059965546387070049160453150146287656955926634303969948238410322586805550666387460130407605709395002173;
            6'd13: xpb[123] = 1024'd15703194736470961692959963036525725520940931135674904621608588585756436160448249157248293893458880287397930352290685900691106895608740472535629439100105820263091896179246896560827981137780881335570691845873668283205616063404998555326406692435304707959397626061768032685311250019382639166567832391737310792715;
            6'd14: xpb[123] = 1024'd26454724768824477315402954608936506925990112540398796063896315020428230891044971316268552747929384487154936487655930464942658490720275919234920944032139424970536709313771366860709382701573041878407683342355276600864845056760836657502667097213653489284491282175297655048035694488098890873005257177765226583257;
            6'd15: xpb[123] = 1024'd37206254801177992937845946181347288331039293945122687506184041455100025621641693475288811602399888686911942623021175029194210085831811365934212448964173029677981522448295837160590784265365202421244674838836884918524074050116674759678927501992002270609584938288827277410760138956815142579442681963793142373799;
            6'd16: xpb[123] = 1024'd47957784833531508560288937753758069736088475349846578948471767889771820352238415634309070456870392886668948758386419593445761680943346812633503953896206634385426335582820307460472185829157362964081666335318493236183303043472512861855187906770351051934678594402356899773484583425531394285880106749821058164341;
            6'd17: xpb[123] = 1024'd58709314865885024182731929326168851141137656754570470390759494324443615082835137793329329311340897086425954893751664157697313276054882259332795458828240239092871148717344777760353587392949523506918657831800101553842532036828350964031448311548699833259772250515886522136209027894247645992317531535848973954883;
            6'd18: xpb[123] = 1024'd69460844898238539805174920898579632546186838159294361833047220759115409813431859952349588165811401286182961029116908721948864871166417706032086963760273843800315961851869248060234988956741684049755649328281709871501761030184189066207708716327048614584865906629416144498933472362963897698754956321876889745425;
            6'd19: xpb[123] = 1024'd80212374930592055427617912470990413951236019564018253275334947193787204544028582111369847020281905485939967164482153286200416466277953152731378468692307448507760774986393718360116390520533844592592640824763318189160990023540027168383969121105397395909959562742945766861657916831680149405192381107904805535967;
            6'd20: xpb[123] = 1024'd90963904962945571050060904043401195356285200968742144717622673628458999274625304270390105874752409685696973299847397850451968061389488599430669973624341053215205588120918188659997792084326005135429632321244926506820219016895865270560229525883746177235053218856475389224382361300396401111629805893932721326509;
            6'd21: xpb[123] = 1024'd101715434995299086672503895615811976761334382373466036159910400063130794005222026429410364729222913885453979435212642414703519656501024046129961478556374657922650401255442658959879193648118165678266623817726534824479448010251703372736489930662094958560146874970005011587106805769112652818067230679960637117051;
            6'd22: xpb[123] = 1024'd112466965027652602294946887188222758166383563778189927602198126497802588735818748588430623583693418085210985570577886978955071251612559492829252983488408262630095214389967129259760595211910326221103615314208143142138677003607541474912750335440443739885240531083534633949831250237828904524504655465988552907593;
            6'd23: xpb[123] = 1024'd123218495060006117917389878760633539571432745182913819044485852932474383466415470747450882438163922284967991705943131543206622846724094939528544488420441867337540027524491599559641996775702486763940606810689751459797905996963379577089010740218792521210334187197064256312555694706545156230942080252016468698135;
            6'd24: xpb[123] = 1024'd9903329408234892141033942928229888231783499461902026358641724302169282859703053996456070077976752175281848433850882672879110600994410051672675868336144431111294166089444852521893159147977441585467400698784119931092774140098320906300292575313911853268607939896476820645173611101332774920260815211418790004346;
            6'd25: xpb[123] = 1024'd20654859440588407763476934500640669636832680866625917800929450736841077590299776155476328932447256375038854569216127237130662196105945498371967373268178035818738979223969322821774560711769602128304392195265728248752003133454159008476552980092260634593701596010006443007898055570049026626698239997446705794888;
            6'd26: xpb[123] = 1024'd31406389472941923385919926073051451041881862271349809243217177171512872320896498314496587786917760574795860704581371801382213791217480945071258878200211640526183792358493793121655962275561762671141383691747336566411232126809997110652813384870609415918795252123536065370622500038765278333135664783474621585430;
            6'd27: xpb[123] = 1024'd42157919505295439008362917645462232446931043676073700685504903606184667051493220473516846641388264774552866839946616365633765386329016391770550383132245245233628605493018263421537363839353923213978375188228944884070461120165835212829073789648958197243888908237065687733346944507481530039573089569502537375972;
            6'd28: xpb[123] = 1024'd52909449537648954630805909217873013851980225080797592127792630040856461782089942632537105495858768974309872975311860929885316981440551838469841888064278849941073418627542733721418765403146083756815366684710553201729690113521673315005334194427306978568982564350595310096071388976197781746010514355530453166514;
            6'd29: xpb[123] = 1024'd63660979570002470253248900790283795257029406485521483570080356475528256512686664791557364350329273174066879110677105494136868576552087285169133392996312454648518231762067204021300166966938244299652358181192161519388919106877511417181594599205655759894076220464124932458795833444914033452447939141558368957056;
            6'd30: xpb[123] = 1024'd74412509602355985875691892362694576662078587890245375012368082910200051243283386950577623204799777373823885246042350058388420171663622731868424897928346059355963044896591674321181568530730404842489349677673769837048148100233349519357855003984004541219169876577654554821520277913630285158885363927586284747598;
            6'd31: xpb[123] = 1024'd85164039634709501498134883935105358067127769294969266454655809344871845973880109109597882059270281573580891381407594622639971766775158178567716402860379664063407858031116144621062970094522565385326341174155378154707377093589187621534115408762353322544263532691184177184244722382346536865322788713614200538140;
            6'd32: xpb[123] = 1024'd95915569667063017120577875507516139472176950699693157896943535779543640704476831268618140913740785773337897516772839186891523361886693625267007907792413268770852671165640614920944371658314725928163332670636986472366606086945025723710375813540702103869357188804713799546969166851062788571760213499642116328682;
            6'd33: xpb[123] = 1024'd106667099699416532743020867079926920877226132104417049339231262214215435435073553427638399768211289973094903652138083751143074956998229071966299412724446873478297484300165085220825773222106886471000324167118594790025835080300863825886636218319050885194450844918243421909693611319779040278197638285670032119224;
            6'd34: xpb[123] = 1024'd117418629731770048365463858652337702282275313509140940781518988648887230165670275586658658622681794172851909787503328315394626552109764518665590917656480478185742297434689555520707174785899047013837315663600203107685064073656701928062896623097399666519544501031773044272418055788495291984635063071697947909766;
            6'd35: xpb[123] = 1024'd4103464079998822589107922819934050942626067788129148095674860018582129558957858835663846262494624063165766515411079445067114306380079630809722297572183041959496435999642808482958337158174001835364109551694571578979932216791643257274178458192518998577818253731185608605035972183282910673953798031100269215977;
            6'd36: xpb[123] = 1024'd14854994112352338211550914392344832347675249192853039537962586453253924289554580994684105116965128262922772650776324009318665901491615077509013802504216646666941249134167278782839738721966162378201101048176179896639161210147481359450438862970867779902911909844715230967760416651999162380391222817128185006519;
            6'd37: xpb[123] = 1024'd25606524144705853833993905964755613752724430597576930980250312887925719020151303153704363971435632462679778786141568573570217496603150524208305307436250251374386062268691749082721140285758322921038092544657788214298390203503319461626699267749216561228005565958244853330484861120715414086828647603156100797061;
            6'd38: xpb[123] = 1024'd36358054177059369456436897537166395157773612002300822422538039322597513750748025312724622825906136662436784921506813137821769091714685970907596812368283856081830875403216219382602541849550483463875084041139396531957619196859157563802959672527565342553099222071774475693209305589431665793266072389184016587603;
            6'd39: xpb[123] = 1024'd47109584209412885078879889109577176562822793407024713864825765757269308481344747471744881680376640862193791056872057702073320686826221417606888317300317460789275688537740689682483943413342644006712075537621004849616848190214995665979220077305914123878192878185304098055933750058147917499703497175211932378145;
            6'd40: xpb[123] = 1024'd57861114241766400701322880681987957967871974811748605307113492191941103211941469630765140534847145061950797192237302266324872281937756864306179822232351065496720501672265159982365344977134804549549067034102613167276077183570833768155480482084262905203286534298833720418658194526864169206140921961239848168687;
            6'd41: xpb[123] = 1024'd68612644274119916323765872254398739372921156216472496749401218626612897942538191789785399389317649261707803327602546830576423877049292311005471327164384670204165314806789630282246746540926965092386058530584221484935306176926671870331740886862611686528380190412363342781382638995580420912578346747267763959229;
            6'd42: xpb[123] = 1024'd79364174306473431946208863826809520777970337621196388191688945061284692673134913948805658243788153461464809462967791394827975472160827757704762832096418274911610127941314100582128148104719125635223050027065829802594535170282509972508001291640960467853473846525892965144107083464296672619015771533295679749771;
            6'd43: xpb[123] = 1024'd90115704338826947568651855399220302183019519025920279633976671495956487403731636107825917098258657661221815598333035959079527067272363204404054337028451879619054941075838570882009549668511286178060041523547438120253764163638348074684261696419309249178567502639422587506831527933012924325453196319323595540313;
            6'd44: xpb[123] = 1024'd100867234371180463191094846971631083588068700430644171076264397930628282134328358266846175952729161860978821733698280523331078662383898651103345841960485484326499754210363041181890951232303446720897033020029046437912993156994186176860522101197658030503661158752952209869555972401729176031890621105351511330855;
            6'd45: xpb[123] = 1024'd111618764403533978813537838544041864993117881835368062518552124365300076864925080425866434807199666060735827869063525087582630257495434097802637346892519089033944567344887511481772352796095607263734024516510654755572222150350024279036782505976006811828754814866481832232280416870445427738328045891379427121397;
            6'd46: xpb[123] = 1024'd122370294435887494435980830116452646398167063240091953960839850799971871595521802584886693661670170260492834004428769651834181852606969544501928851824552693741389380479411981781653754359887767806571016012992263073231451143705862381213042910754355593153848470980011454595004861339161679444765470677407342911939;
            6'd47: xpb[123] = 1024'd9055128784116268659624894284048995058517817519080161274995722169666770988809385833891881301483000150806690732336520781506669606877284656646060231740255257515143519044365234743904916732162722628097809901086631544526319286840803710424324745849474925212122223679424018927622777733949298134084205636809664218150;
            6'd48: xpb[123] = 1024'd19806658816469784282067885856459776463566998923804052717283448604338565719406107992912140155953504350563696867701765345758221201988820103345351736672288862222588332178889705043786318295954883170934801397568239862185548280196641812600585150627823706537215879792953641290347222202665549840521630422837580008692;
            6'd49: xpb[123] = 1024'd30558188848823299904510877428870557868616180328527944159571175039010360450002830151932399010424008550320703003067009910009772797100355550044643241604322466930033145313414175343667719859747043713771792894049848179844777273552479914776845555406172487862309535906483263653071666671381801546959055208865495799234;
            6'd50: xpb[123] = 1024'd41309718881176815526953869001281339273665361733251835601858901473682155180599552310952657864894512750077709138432254474261324392211890996743934746536356071637477958447938645643549121423539204256608784390531456497504006266908318016953105960184521269187403192020012886015796111140098053253396479994893411589776;
            6'd51: xpb[123] = 1024'd52061248913530331149396860573692120678714543137975727044146627908353949911196274469972916719365016949834715273797499038512875987323426443443226251468389676344922771582463115943430522987331364799445775887013064815163235260264156119129366364962870050512496848133542508378520555608814304959833904780921327380318;
            6'd52: xpb[123] = 1024'd62812778945883846771839852146102902083763724542699618486434354343025744641792996628993175573835521149591721409162743602764427582434961890142517756400423281052367584716987586243311924551123525342282767383494673132822464253619994221305626769741218831837590504247072130741245000077530556666271329566949243170860;
            6'd53: xpb[123] = 1024'd73564308978237362394282843718513683488812905947423509928722080777697539372389718788013434428306025349348727544527988167015979177546497336841809261332456885759812397851512056543193326114915685885119758879976281450481693246975832323481887174519567613162684160360601753103969444546246808372708754352977158961402;
            6'd54: xpb[123] = 1024'd84315839010590878016725835290924464893862087352147401371009807212369334102986440947033693282776529549105733679893232731267530772658032783541100766264490490467257210986036526843074727678707846427956750376457889768140922240331670425658147579297916394487777816474131375466693889014963060079146179139005074751944;
            6'd55: xpb[123] = 1024'd95067369042944393639168826863335246298911268756871292813297533647041128833583163106053952137247033748862739815258477295519082367769568230240392271196524095174702024120560997142956129242500006970793741872939498085800151233687508527834407984076265175812871472587660997829418333483679311785583603925032990542486;
            6'd56: xpb[123] = 1024'd105818899075297909261611818435746027703960450161595184255585260081712923564179885265074210991717537948619745950623721859770633962881103676939683776128557699882146837255085467442837530806292167513630733369421106403459380227043346630010668388854613957137965128701190620192142777952395563492021028711060906333028;
            6'd57: xpb[123] = 1024'd116570429107651424884054810008156809109009631566319075697872986516384718294776607424094469846188042148376752085988966424022185557992639123638975281060591304589591650389609937742718932370084328056467724865902714721118609220399184732186928793632962738463058784814720242554867222421111815198458453497088822123570;
            6'd58: xpb[123] = 1024'd3255263455880199107698874175753157769360385845307283012028857886079617688064190673099657486000872038690608813896717553694673312262954235783106660976293868363345788954563190704970094742359282877994518753997083192413477363534126061398210628728082070521332537514132806887485138815899433887777188456491143429781;
            6'd59: xpb[123] = 1024'd14006793488233714730141865748163939174409567250031174454316584320751412418660912832119916340471376238447614949261962117946224907374489682482398165908327473070790602089087661004851496306151443420831510250478691510072706356889964163574471033506430851846426193627662429250209583284615685594214613242519059220323;
            6'd60: xpb[123] = 1024'd24758323520587230352584857320574720579458748654755065896604310755423207149257634991140175194941880438204621084627206682197776502486025129181689670840361077778235415223612131304732897869943603963668501746960299827731935350245802265750731438284779633171519849741192051612934027753331937300652038028546975010865;
            6'd61: xpb[123] = 1024'd35509853552940745975027848892985501984507930059478957338892037190095001879854357150160434049412384637961627219992451246449328097597560575880981175772394682485680228358136601604614299433735764506505493243441908145391164343601640367926991843063128414496613505854721673975658472222048189007089462814574890801407;
            6'd62: xpb[123] = 1024'd46261383585294261597470840465396283389557111464202848781179763624766796610451079309180692903882888837718633355357695810700879692709096022580272680704428287193125041492661071904495700997527925049342484739923516463050393336957478470103252247841477195821707161968251296338382916690764440713526887600602806591949;
            6'd63: xpb[123] = 1024'd57012913617647777219913832037807064794606292868926740223467490059438591341047801468200951758353393037475639490722940374952431287820631469279564185636461891900569854627185542204377102561320085592179476236405124780709622330313316572279512652619825977146800818081780918701107361159480692419964312386630722382491;
        endcase
    end

    always_comb begin
        case(flag[41][11:6])
            6'd0: xpb[124] = 1024'd0;
            6'd1: xpb[124] = 1024'd67764443650001292842356823610217846199655474273650631665755216494110386071644523627221210612823897237232645626088184939203982882932166915978855690568495496608014667761710012504258504125112246135016467732886733098368851323669154674455773057398174758471894474195310541063831805628196944126401737172658638173033;
            6'd2: xpb[124] = 1024'd11462191615877844285914719815621259654612521421565579203378577923243876805979908344427350010990120165022141844718876443828901925023113497402551256120659952282338660953848807670886769058707286548722737857386226350373341797117412575946567545113120067676969044976504024097557083182465255235684784518691681861735;
            6'd3: xpb[124] = 1024'd79226635265879137128271543425839105854267995695216210869133794417354262877624431971648560623814017402254787470807061383032884807955280413381406946689155448890353328715558820175145273183819532683739205590272959448742193120786567250402340602511294826148863519171814565161388888810662199362086521691350320034768;
            6'd4: xpb[124] = 1024'd22924383231755688571829439631242519309225042843131158406757155846487753611959816688854700021980240330044283689437752887657803850046226994805102512241319904564677321907697615341773538117414573097445475714772452700746683594234825151893135090226240135353938089953008048195114166364930510471369569037383363723470;
            6'd5: xpb[124] = 1024'd90688826881756981414186263241460365508880517116781790072512372340598139683604340316075910634804137567276929315525937826861786732978393910783958202809815401172691989669407627846032042242526819232461943447659185799115534917903979826348908147624414893825832564148318589258945971993127454597771306210042001896503;
            6'd6: xpb[124] = 1024'd34386574847633532857744159446863778963837564264696737610135733769731630417939725033282050032970360495066425534156629331486705775069340492207653768361979856847015982861546423012660307176121859646168213572158679051120025391352237727839702635339360203030907134929512072292671249547395765707054353556075045585205;
            6'd7: xpb[124] = 1024'd102151018497634825700100983057081625163493038538347369275890950263842016489584248660503260645794257732299071160244814270690688658001507408186509458930475353455030650623256435516918811301234105781184681305045412149488876715021392402295475692737534961502801609124822613356503055175592709833456090728733683758238;
            6'd8: xpb[124] = 1024'd45848766463511377143658879262485038618450085686262316813514311692975507223919633377709400043960480660088567378875505775315607700092453989610205024482639809129354643815395230683547076234829146194890951429544905401493367188469650303786270180452480270707876179906016096390228332729861020942739138074766727446940;
            6'd9: xpb[124] = 1024'd113613210113512669986015702872702884818105559959912948479269528187085893295564157004930610656784377897321213004963690714519590583024620905589060715051135305737369311577105243187805580359941392329907419162431638499862218512138804978242043237850655029179770654101326637454060138358057965069140875247425365619973;
            6'd10: xpb[124] = 1024'd57310958079389221429573599078106298273062607107827896016892889616219384029899541722136750054950600825110709223594382219144509625115567487012756280603299761411693304769244038354433845293536432743613689286931131751866708985587062879732837725565600338384845224882520120487785415912326276178423922593458409308675;
            6'd11: xpb[124] = 1024'd1008706045265772873131495283509711728019654255742843554516251045352874764234926439342889453116823752900205442225073723769428667206514068436451846155464217086017297961382833521062110227131473157319959411430625003871199459035320781223632213280545647589919795663713603521510693466594587287706969939491452997377;
            6'd12: xpb[124] = 1024'd68773149695267065715488318893727557927675128529393475220271467539463260835879450066564100065940720990132851068313258662973411550138680984415307536723959713694031965723092846025320614352243719292336427144317358102240050782704475455679405270678720406061814269859024144585342499094791531414108707112150091170410;
            6'd13: xpb[124] = 1024'd12470897661143617159046215099130971382632175677308422757894828968596751570214834783770239464106943917922347286943950167598330592229627565839003102276124169368355958915231641191948879285838759706042697268816851354244541256152733357170199758393665715266888840640217627619067776649059842523391754458183134859112;
            6'd14: xpb[124] = 1024'd80235341311144910001403038709348817582287649950959054423650045462707137641859358410991450076930841155154992913032135106802313475161794481817858792844619665976370626676941653696207383410951005841059165001703584452613392579821888031625972815791840473738783314835528168682899582277256786649793491630841773032145;
            6'd15: xpb[124] = 1024'd23933089277021461444960934914752231037244697098874001961273406891840628376194743128197589475097064082944489131662826611427232517252741063241554358396784121650694619869080448862835648344546046254765435126203077704617883053270145933116767303506785782943857885616721651716624859831525097759076538976874816720847;
            6'd16: xpb[124] = 1024'd91697532927022754287317758524970077236900171372524633627028623385951014447839266755418800087920961320177134757751011550631215400184907979220410048965279618258709287630790461367094152469658292389781902859089810802986734376939300607572540360904960541415752359812032192780456665459722041885478276149533454893880;
            6'd17: xpb[124] = 1024'd35395280892899305730875654730373490691857218520439581164651984815084505182174651472624939486087184247966630976381703055256134442275854560644105614517444073933033280822929256533722417403253332803488172983589304054991224850387558509063334848619905850620826930593225675814181943013990352994761323495566498582582;
            6'd18: xpb[124] = 1024'd103159724542900598573232478340591336891512692794090212830407201309194891253819175099846150098911081485199276602469887994460117325208021476622961305085939570541047948584639269037980921528365578938504640716476037153360076174056713183519107906018080609092721404788536216878013748642187297121163060668225136755615;
            6'd19: xpb[124] = 1024'd46857472508777150016790374545994750346469739942005160368030562738328381988154559817052289497077304412988772821100579499085036367298968058046656870638104026215371941776778064204609186461960619352210910840975530405364566647504971085009902393733025918297795975569729699911739026196455608230446108014258180444317;
            6'd20: xpb[124] = 1024'd114621916158778442859147198156212596546125214215655792033785779232438768059799083444273500109901201650221418447188764438289019250231134974025512561206599522823386609538488076708867690587072865487227378573862263503733417971174125759465675451131200676769690449765040240975570831824652552356847845186916818617350;
            6'd21: xpb[124] = 1024'd58319664124654994302705094361616010001082261363570739571409140661572258794134468161479639508067424578010914665819455942913938292322081555449208126758763978497710602730626871875495955520667905900933648698361756755737908444622383660956469938846145985974765020546233724009296109378920863466130892532949862306052;
            6'd22: xpb[124] = 1024'd2017412090531545746262990567019423456039308511485687109032502090705749528469852878685778906233647505800410884450147447538857334413028136872903692310928434172034595922765667042124220454262946314639918822861250007742398918070641562447264426561091295179839591327427207043021386933189174575413939878982905994754;
            6'd23: xpb[124] = 1024'd69781855740532838588619814177237269655694782785136318774787718584816135600114376505906989519057544743033056510538332386742840217345195052851759382879423930780049263684475679546382724579375192449656386555747983106111250241739796236903037483959266053651734065522737748106853192561386118701815677051641544167787;
            6'd24: xpb[124] = 1024'd13479603706409390032177710382640683110651829933051266312411080013949626334449761223113128917223767670822552729169023891367759259436141634275454948431588386454373256876614474713010989512970232863362656680247476358115740715188054138393831971674211362856808636303931231140578470115654429811098724397674587856489;
            6'd25: xpb[124] = 1024'd81244047356410682874534533992858529310307304206701897978166296508060012406094284850334339530047664908055198355257208830571742142368308550254310639000083883062387924638324487217269493638082478998379124413134209456484592038857208812849605029072386121328703110499241772204410275743851373937500461570333226029522;
            6'd26: xpb[124] = 1024'd24941795322287234318092430198261942765264351354616845515789657937193503140429669567540478928213887835844694573887900335196661184459255131678006204552248338736711917830463282383897758571677519412085394537633702708489082512305466714340399516787331430533777681280435255238135553298119685046783508916366269718224;
            6'd27: xpb[124] = 1024'd92706238972288527160449253808479788964919825628267477181544874431303889212074193194761689541037785073077340199976085274400644067391422047656861895120743835344726585592173294888156262696789765547101862270520435806857933835974621388796172574185506189005672155475745796301967358926316629173185246089024907891257;
            6'd28: xpb[124] = 1024'd36403986938165078604007150013883202419876872776182424719168235860437379946409577911967828939204008000866836418606776779025563109482368629080557460672908291019050578784312090054784527630384805960808132395019929058862424309422879290286967061900451498210746726256939279335692636480584940282468293435057951579959;
            6'd29: xpb[124] = 1024'd104168430588166371446363973624101048619532347049833056384923452354547766018054101539189039552027905238099482044694961718229545992414535545059413151241403787627065246546022102559043031755497052095824600127906662157231275633092033964742740119298626256682641200452249820399524442108781884408870030607716589752992;
            6'd30: xpb[124] = 1024'd47866178554042922889921869829504462074489394197748003922546813783681256752389486256395178950194128165888978263325653222854465034505482126483108716793568243301389239738160897725671296689092092509530870252406155409235766106540291866233534607013571565887715771233443303433249719663050195518153077953749633441694;
            6'd31: xpb[124] = 1024'd115630622204044215732278693439722308274144868471398635588302030277791642824034009883616389563018025403121623889413838162058447917437649042461964407362063739909403907499870910229929800814204338644547337985292888507604617430209446540689307664411746324359610245428753844497081525291247139644554815126408271614727;
            6'd32: xpb[124] = 1024'd59328370169920767175836589645125721729101915619313583125925391706925133558369394600822528961184248330911120108044529666683366959528595623885659972914228195583727900692009705396558065747799379058253608109792381759609107903657704442180102152126691633564684816209947327530806802845515450753837862472441315303429;
            6'd33: xpb[124] = 1024'd3026118135797318619394485850529135184058962767228530663548753136058624292704779318028668359350471258700616326675221171308286001619542205309355538466392651258051893884148500563186330681394419471959878234291875011613598377105962343670896639841636942769759386991140810564532080399783761863120909818474358992131;
            6'd34: xpb[124] = 1024'd70790561785798611461751309460746981383714437040879162329303969630169010364349302945249878972174368495933261952763406110512268884551709121288211229034888147866066561645858513067444834806506665606976345967178608109982449700775117018126669697239811701241653861186451351628363886027980705989522646991132997165164;
            6'd35: xpb[124] = 1024'd14488309751675162905309205666150394838671484188794109866927331059302501098684687662456018370340591423722758171394097615137187926642655702711906794587052603540390554837997308234073099740101706020682616091678101361986940174223374919617464184954757010446728431967644834662089163582249017098805694337166040853866;
            6'd36: xpb[124] = 1024'd82252753401676455747666029276368241038326958462444741532682547553412887170329211289677228983164488660955403797482282554341170809574822618690762485155548100148405222599707320738331603865213952155699083824564834460355791497892529594073237242352931768918622906162955375725920969210445961225207431509824679026899;
            6'd37: xpb[124] = 1024'd25950501367553007191223925481771654493284005610359689070305908982546377904664596006883368381330711588744900016112974058966089851665769200114458050707712555822729215791846115904959868798808992569405353949064327712360281971340787495564031730067877078123697476944148858759646246764714272334490478855857722715601;
            6'd38: xpb[124] = 1024'd93714945017554300033580749091989500692939479884010320736061125476656763976309119634104578994154608825977545642201158998170072734597936116093313741276208052430743883553556128409218372923921238704421821681951060810729133295009942170019804787466051836595591951139459399823478052392911216460892216028516360888634;
            6'd39: xpb[124] = 1024'd37412692983430851477138645297392914147896527031925268273684486905790254710644504351310718392320831753767041860831850502794991776688882697517009306828372508105067876745694923575846637857516279118128091806450554062733623768458200071510599275180997145800666521920652882857203329947179527570175263374549404577336;
            6'd40: xpb[124] = 1024'd105177136633432144319495468907610760347552001305575899939439703399900640782289027978531929005144728990999687486920035441998974659621049613495864997396868004713082544507404936080105141982628525253144559539337287161102475092127354745966372332579171904272560996115963423921035135575376471696577000547208042750369;
            6'd41: xpb[124] = 1024'd48874884599308695763053365113014173802509048453490847477063064829034131516624412695738068403310951918789183705550726946623893701711996194919560562949032460387406537699543731246733406916223565666850829663836780413106965565575612647457166820294117213477635566897156906954760413129644782805860047893241086439071;
            6'd42: xpb[124] = 1024'd116639328249309988605410188723232020002164522727141479142818281323144517588268936322959279016134849156021829331638911885827876584644163110898416253517527956995421205461253743750991911041335811801867297396723513511475816889244767321912939877692291971949530041092467448018592218757841726932261785065899724612104;
            6'd43: xpb[124] = 1024'd60337076215186540048968084928635433457121569875056426680441642752278008322604321040165418414301072083811325550269603390452795626735109692322111819069692412669745198653392538917620175974930852215573567521223006763480307362693025223403734365407237281154604611873660931052317496312110038041544832411932768300806;
            6'd44: xpb[124] = 1024'd4034824181063091492525981134038846912078617022971374218065004181411499056939705757371557812467295011600821768900294895077714668826056273745807384621856868344069191845531334084248440908525892629279837645722500015484797836141283124894528853122182590359679182654854414086042773866378349150827879757965811989508;
            6'd45: xpb[124] = 1024'd71799267831064384334882804744256693111734091296622005883820220675521885128584229384592768425291192248833467394988479834281697551758223189724663075190352364952083859607241346588506945033638138764296305378609233113853649159810437799350301910520357348831573656850164955149874579494575293277229616930624450162541;
            6'd46: xpb[124] = 1024'd15497015796940935778440700949660106566691138444536953421443582104655375862919614101798907823457415176622963613619171338906616593849169771148358640742516820626407852799380141755135209967233179178002575503108726365858139633258695700841096398235302658036648227631358438183599857048843604386512664276657493851243;
            6'd47: xpb[124] = 1024'd83261459446942228620797524559877952766346612718187585087198798598765761934564137729020118436281312413855609239707356278110599476781336687127214331311012317234422520561090154259393714092345425313019043235995459464226990956927850375296869455633477416508542701826668979247431662677040548512914401449316132024276;
            6'd48: xpb[124] = 1024'd26959207412818780064355420765281366221303659866102532624822160027899252668899522446226257834447535341645105458338047782735518518872283268550909896863176772908746513753228949426021979025940465726725313360494952716231481430376108276787663943348422725713617272607862462281156940231308859622197448795349175712978;
            6'd49: xpb[124] = 1024'd94723651062820072906712244375499212420959134139753164290577376522009638740544046073447468447271432578877751084426232721939501401804450184529765587431672269516761181514938961930280483151052711861741781093381685814600332754045262951243437000746597484185511746803173003344988745859505803748599185968007813886011;
            6'd50: xpb[124] = 1024'd38421399028696624350270140580902625875916181287668111828200737951143129474879430790653607845437655506667247303056924226564420443895396765953461152983836725191085174707077757096908748084647752275448051217881179066604823227493520852734231488461542793390586317584366486378714023413774114857882233314040857574713;
            6'd51: xpb[124] = 1024'd106185842678697917192626964191120472075571655561318743493955954445253515546523954417874818458261552743899892929145109165768403326827563681932316843552332221799099842468787769601167252209759998410464518950767912164973674551162675527190004545859717551862480791779677027442545829041971058984283970486699495747746;
            6'd52: xpb[124] = 1024'd49883590644574468636184860396523885530528702709233691031579315874387006280859339135080957856427775671689389147775800670393322368918510263356012409104496677473423835660926564767795517143355038824170789075267405416978165024610933428680799033574662861067555362560870510476271106596239370093567017832732539436448;
            6'd53: xpb[124] = 1024'd117648034294575761478541684006741731730184176982884322697334532368497392352503862762302168469251672908922034773863985609597305251850677179334868099672992174081438503422636577272054021268467284959187256808154138515347016348280088103136572090972837619539449836756181051540102912224436314219968755005391177609481;
            6'd54: xpb[124] = 1024'd61345782260452312922099580212145145185141224130799270234957893797630883086839247479508307867417895836711530992494677114222224293941623760758563665225156629755762496614775372438682286202062325372893526932653631767351506821728346004627366578687782928744524407537374534573828189778704625329251802351424221298183;
            6'd55: xpb[124] = 1024'd5043530226328864365657476417548558640098271278714217772581255226764373821174632196714447265584118764501027211125368618847143336032570342182259230777321085430086489806914167605310551135657365786599797057153125019355997295176603906118161066402728237949598978318568017607553467332972936438534849697457264986885;
            6'd56: xpb[124] = 1024'd72807973876330157208014300027766404839753745552364849438336471720874759892819155823935657878408016001733672837213553558051126218964737258161114921345816582038101157568624180109569055260769611921616264790039858117724848618845758580573934123800902996421493452513878558671385272961169880564936586870115903159918;
            6'd57: xpb[124] = 1024'd16505721842206708651572196233169818294710792700279796975959833150008250627154540541141797276574238929523169055844245062676045261055683839584810486897981037712425150760762975276197320194364652335322534914539351369729339092294016482064728611515848305626568023295072041705110550515438191674219634216148946848620;
            6'd58: xpb[124] = 1024'd84270165492208001493929019843387664494366266973930428641715049644118636698799064168363007889398136166755814681932430001880028143987850755563666177466476534320439818522472987780455824319476898470339002647426084468098190415963171156520501668914023064098462497490382582768942356143635135800621371388807585021653;
            6'd59: xpb[124] = 1024'd27967913458084552937486916048791077949323314121845376179338411073252127433134448885569147287564359094545310900563121506504947186078797336987361743018640989994763811714611782947084089253071938884045272771925577720102680889411429058011296156628968373303537068271576065802667633697903446909904418734840628710355;
            6'd60: xpb[124] = 1024'd95732357108085845779843739659008924148978788395496007845093627567362513504778972512790357900388256331777956526651306445708930069010964252966217433587136486602778479476321795451342593378184185019061740504812310818471532213080583732467069214027143131775431542466886606866499439326100391036306155907499266883388;
            6'd61: xpb[124] = 1024'd39430105073962397223401635864412337603935835543410955382716988996496004239114357229996497298554479259567452745281997950333849111101910834389912999139300942277102472668460590617970858311779225432768010629311804070476022686528841633957863701742088440980506113248080089900224716880368702145589203253532310572090;
            6'd62: xpb[124] = 1024'd107194548723963690065758459474630183803591309817061587048472205490606390310758880857217707911378376496800098371370182889537831994034077750368768689707796438885117140430170603122229362436891471567784478362198537168844874010197996308413636759140263199452400587443390630964056522508565646271990940426190948745123;
            6'd63: xpb[124] = 1024'd50892296689840241509316355680033597258548356964976534586095566919739881045094265574423847309544599424589594590000874394162751036125024331792464255259960894559441133622309398288857627370486511981490748486698030420849364483646254209904431246855208508657475158224584113997781800062833957381273987772223992433825;
        endcase
    end

    always_comb begin
        case(flag[41][16:12])
            5'd0: xpb[125] = 1024'd0;
            5'd1: xpb[125] = 1024'd118656740339841534351673179290251443458203831238627166251850783413850267116738789201645057922368496661822240216089059333366733919057191247771319945828456391167455801384019410793116131495598758116507216219584763519218215807315408884360204304253383267129369632419894655061613605691030901507675724944882630606858;
            5'd2: xpb[125] = 1024'd113246784995558327304547431175688454171709235351518648375569711762723638896168439493275044630079319014201331024720625232154403997273162160987479766640581741401220928198467604248602023799680310511704234830782287192072070764409920995755430038823537084991919361425672252093120683308133169998232760063139666729385;
            5'd3: xpb[125] = 1024'd107836829651275120257421683061125464885214639464410130499288640111597010675598089784905031337790141366580421833352191130942074075489133074203639587452707091634986055012915797704087916103761862906901253441979810864925925721504433107150655773393690902854469090431449849124627760925235438488789795181396702851912;
            5'd4: xpb[125] = 1024'd102426874306991913210295934946562475598720043577301612623007568460470382455027740076535018045500963718959512641983757029729744153705103987419799408264832441868751181827363991159573808407843415302098272053177334537779780678598945218545881507963844720717018819437227446156134838542337706979346830299653738974439;
            5'd5: xpb[125] = 1024'd97016918962708706163170186831999486312225447690193094746726496809343754234457390368165004753211786071338603450615322928517414231921074900635959229076957792102516308641812184615059700711924967697295290664374858210633635635693457329941107242533998538579568548443005043187641916159439975469903865417910775096966;
            5'd6: xpb[125] = 1024'd91606963618425499116044438717436497025730851803084576870445425158217126013887040659794991460922608423717694259246888827305084310137045813852119049889083142336281435456260378070545593016006520092492309275572381883487490592787969441336332977104152356442118277448782640219148993776542243960460900536167811219493;
            5'd7: xpb[125] = 1024'd86197008274142292068918690602873507739236255915976058994164353507090497793316690951424978168633430776096785067878454726092754388353016727068278870701208492570046562270708571526031485320088072487689327886769905556341345549882481552731558711674306174304668006454560237250656071393644512451017935654424847342020;
            5'd8: xpb[125] = 1024'd80787052929859085021792942488310518452741660028867541117883281855963869572746341243054964876344253128475875876510020624880424466568987640284438691513333842803811689085156764981517377624169624882886346497967429229195200506976993664126784446244459992167217735460337834282163149010746780941574970772681883464547;
            5'd9: xpb[125] = 1024'd75377097585575877974667194373747529166247064141759023241602210204837241352175991534684951584055075480854966685141586523668094544784958553500598512325459193037576815899604958437003269928251177278083365109164952902049055464071505775522010180814613810029767464466115431313670226627849049432132005890938919587074;
            5'd10: xpb[125] = 1024'd69967142241292670927541446259184539879752468254650505365321138553710613131605641826314938291765897833234057493773152422455764623000929466716758333137584543271341942714053151892489162232332729673280383720362476574902910421166017886917235915384767627892317193471893028345177304244951317922689041009195955709601;
            5'd11: xpb[125] = 1024'd64557186897009463880415698144621550593257872367541987489040066902583984911035292117944924999476720185613148302404718321243434701216900379932918153949709893505107069528501345347975054536414282068477402331560000247756765378260529998312461649954921445754866922477670625376684381862053586413246076127452991832128;
            5'd12: xpb[125] = 1024'd59147231552726256833289950030058561306763276480433469612758995251457356690464942409574911707187542537992239111036284220031104779432871293149077974761835243738872196342949538803460946840495834463674420942757523920610620335355042109707687384525075263617416651483448222408191459479155854903803111245710027954655;
            5'd13: xpb[125] = 1024'd53737276208443049786164201915495572020268680593324951736477923600330728469894592701204898414898364890371329919667850118818774857648842206365237795573960593972637323157397732258946839144577386858871439553955047593464475292449554221102913119095229081479966380489225819439698537096258123394360146363967064077182;
            5'd14: xpb[125] = 1024'd48327320864159842739038453800932582733774084706216433860196851949204100249324242992834885122609187242750420728299416017606444935864813119581397616386085944206402449971845925714432731448658939254068458165152571266318330249544066332498138853665382899342516109495003416471205614713360391884917181482224100199709;
            5'd15: xpb[125] = 1024'd42917365519876635691912705686369593447279488819107915983915780298077472028753893284464871830320009595129511536930981916394115014080784032797557437198211294440167576786294119169918623752740491649265476776350094939172185206638578443893364588235536717205065838500781013502712692330462660375474216600481136322236;
            5'd16: xpb[125] = 1024'd37507410175593428644786957571806604160784892931999398107634708646950843808183543576094858538030831947508602345562547815181785092296754946013717258010336644673932703600742312625404516056822044044462495387547618612026040163733090555288590322805690535067615567506558610534219769947564928866031251718738172444763;
            5'd17: xpb[125] = 1024'd32097454831310221597661209457243614874290297044890880231353636995824215587613193867724845245741654299887693154194113713969455170512725859229877078822461994907697830415190506080890408360903596439659513998745142284879895120827602666683816057375844352930165296512336207565726847564667197356588286836995208567290;
            5'd18: xpb[125] = 1024'd26687499487027014550535461342680625587795701157782362355072565344697587367042844159354831953452476652266783962825679612757125248728696772446036899634587345141462957229638699536376300664985148834856532609942665957733750077922114778079041791945998170792715025518113804597233925181769465847145321955252244689817;
            5'd19: xpb[125] = 1024'd21277544142743807503409713228117636301301105270673844478791493693570959146472494450984818661163299004645874771457245511544795326944667685662196720446712695375228084044086892991862192969066701230053551221140189630587605035016626889474267526516151988655264754523891401628741002798871734337702357073509280812344;
            5'd20: xpb[125] = 1024'd15867588798460600456283965113554647014806509383565326602510422042444330925902144742614805368874121357024965580088811410332465405160638598878356541258838045608993210858535086447348085273148253625250569832337713303441459992111139000869493261086305806517814483529668998660248080415974002828259392191766316934871;
            5'd21: xpb[125] = 1024'd10457633454177393409158216998991657728311913496456808726229350391317702705331795034244792076584943709404056388720377309120135483376609512094516362070963395842758337672983279902833977577229806020447588443535236976295314949205651112264718995656459624380364212535446595691755158033076271318816427310023353057398;
            5'd22: xpb[125] = 1024'd5047678109894186362032468884428668441817317609348290849948278740191074484761445325874778784295766061783147197351943207907805561592580425310676182883088746076523464487431473358319869881311358415644607054732760649149169906300163223659944730226613442242913941541224192723262235650178539809373462428280389179925;
            5'd23: xpb[125] = 1024'd123704418449735720713705648174680111900021148847975457101799062154041341601500234527519836706664262723605387413441002541274539480649771673081996128711545137243979265871450884151436001376910116532151823274317524168367385713615572108020149034479996709372283573961118847784875841341209441317049187373163019786783;
            5'd24: xpb[125] = 1024'd118294463105452513666579900060117122613526552960866939225517990502914713380929884819149823414375085075984478222072568440062209558865742586298155949523670487477744392685899077606921893680991668927348841885515047841221240670710084219415374769050150527234833302966896444816382918958311709807606222491420055909310;
            5'd25: xpb[125] = 1024'd112884507761169306619454151945554133327031957073758421349236918851788085160359535110779810122085907428363569030704134338849879637081713499514315770335795837711509519500347271062407785985073221322545860496712571514075095627804596330810600503620304345097383031972674041847889996575413978298163257609677092031837;
            5'd26: xpb[125] = 1024'd107474552416886099572328403830991144040537361186649903472955847200661456939789185402409796829796729780742659839335700237637549715297684412730475591147921187945274646314795464517893678289154773717742879107910095186928950584899108442205826238190458162959932760978451638879397074192516246788720292727934128154364;
            5'd27: xpb[125] = 1024'd102064597072602892525202655716428154754042765299541385596674775549534828719218835694039783537507552133121750647967266136425219793513655325946635411960046538179039773129243657973379570593236326112939897719107618859782805541993620553601051972760611980822482489984229235910904151809618515279277327846191164276891;
            5'd28: xpb[125] = 1024'd96654641728319685478076907601865165467548169412432867720393703898408200498648485985669770245218374485500841456598832035212889871729626239162795232772171888412804899943691851428865462897317878508136916330305142532636660499088132664996277707330765798685032218990006832942411229426720783769834362964448200399418;
            5'd29: xpb[125] = 1024'd91244686384036478430951159487302176181053573525324349844112632247281572278078136277299756952929196837879932265230397934000559949945597152378955053584297238646570026758140044884351355201399430903333934941502666205490515456182644776391503441900919616547581947995784429973918307043823052260391398082705236521945;
            5'd30: xpb[125] = 1024'd85834731039753271383825411372739186894558977638215831967831560596154944057507786568929743660640019190259023073861963832788230028161568065595114874396422588880335153572588238339837247505480983298530953552700189878344370413277156887786729176471073434410131677001562027005425384660925320750948433200962272644472;
            5'd31: xpb[125] = 1024'd80424775695470064336699663258176197608064381751107314091550488945028315836937436860559730368350841542638113882493529731575900106377538978811274695208547939114100280387036431795323139809562535693727972163897713551198225370371668999181954911041227252272681406007339624036932462278027589241505468319219308766999;
        endcase
    end

    always_comb begin
        case(flag[42][5:0])
            6'd0: xpb[126] = 1024'd0;
            6'd1: xpb[126] = 1024'd37507410175593428644786957571806604160784892931999398107634708646950843808183543576094858538030831947508602345562547815181785092296754946013717258010336644673932703600742312625404516056822044044462495387547618612026040163733090555288590322805690535067615567506558610534219769947564928866031251718738172444763;
            6'd2: xpb[126] = 1024'd75014820351186857289573915143613208321569785863998796215269417293901687616367087152189717076061663895017204691125095630363570184593509892027434516020673289347865407201484625250809032113644088088924990775095237224052080327466181110577180645611381070135231135013117221068439539895129857732062503437476344889526;
            6'd3: xpb[126] = 1024'd112522230526780285934360872715419812482354678795998194322904125940852531424550630728284575614092495842525807036687643445545355276890264838041151774031009934021798110802226937876213548170466132133387486162642855836078120491199271665865770968417071605202846702519675831602659309842694786598093755156214517334289;
            6'd4: xpb[126] = 1024'd25962945018248973180348902882411983898441144602261908302406979522826479895425035394364362937465653480591259974792697826148076528345799449499708907025015537762040139833398033163987825035770970456539783941803234601739799804711465448189382721539532691003642366612117384106772551716331082447006317048327095294721;
            6'd5: xpb[126] = 1024'd63470355193842401825135860454218588059226037534261306410041688169777323703608578970459221475496485428099862320355245641329861620642554395513426165035352182435972843434140345789392341092593014501002279329350853213765839968444556003477973044345223226071257934118675994640992321663896011313037568767065267739484;
            6'd6: xpb[126] = 1024'd100977765369435830469922818026025192220010930466260704517676396816728167511792122546554080013527317375608464665917793456511646712939309341527143423045688827109905547034882658414796857149415058545464774716898471825791880132177646558766563367150913761138873501625234605175212091611460940179068820485803440184247;
            6'd7: xpb[126] = 1024'd14418479860904517715910848193017363636097396272524418497179250398702115982666527212633867336900475013673917604022847837114367964394843952985700556039694430850147576066053753702571134014719896868617072496058850591453559445689840341090175120273374846939669165717676157679325333485097236027981382377916018144679;
            6'd8: xpb[126] = 1024'd51925890036497946360697805764823967796882289204523816604813959045652959790850070788728725874931306961182519949585395652296153056691598898999417814050031075524080279666796066327975650071541940913079567883606469203479599609422930896378765443079065382007284733224234768213545103432662164894012634096654190589442;
            6'd9: xpb[126] = 1024'd89433300212091375005484763336630571957667182136523214712448667692603803599033614364823584412962138908691122295147943467477938148988353845013135072060367720198012983267538378953380166128363984957542063271154087815505639773156021451667355765884755917074900300730793378747764873380227093760043885815392363034205;
            6'd10: xpb[126] = 1024'd2874014703560062251472793503622743373753647942786928691951521274577752069908019030903371736335296546756575233252997848080659400443888456471692205054373323938255012298709474241154442993668823280694361050314466581167319086668215233990967519007217002875695964823234931251878115253863389608956447707504940994637;
            6'd11: xpb[126] = 1024'd40381424879153490896259751075429347534538540874786326799586229921528595878091562606998230274366128494265177578815545663262444492740643402485409463064709968612187715899451786866558959050490867325156856437862085193193359250401305789279557841812907537943311532329793541786097885201428318474987699426243113439400;
            6'd12: xpb[126] = 1024'd77888835054746919541046708647235951695323433806785724907220938568479439686275106183093088812396960441773779924378093478444229585037398348499126721075046613286120419500194099491963475107312911369619351825409703805219399414134396344568148164618598073010927099836352152320317655148993247341018951144981285884163;
            6'd13: xpb[126] = 1024'd115396245230340348185833666219042555856108326738785123014855647215430283494458649759187947350427792389282382269940641293626014677334153294512843979085383257960053123100936412117367991164134955414081847212957322417245439577867486899856738487424288608078542667342910762854537425096558176207050202863719458328926;
            6'd14: xpb[126] = 1024'd28836959721809035431821696386034727272194792545048836994358500797404231965333054425267734673800950027347835208045695674228735928789687905971401112079388861700295152132107507405142268029439793737234144992117701182907118891379680682180350240546749693879338331435352315358650666970194472055962764755832036289358;
            6'd15: xpb[126] = 1024'd66344369897402464076608653957841331432979685477048235101993209444355075773516598001362593211831781974856437553608243489410521021086442851985118370089725506374227855732849820030546784086261837781696640379665319794933159055112771237468940563352440228946953898941910925892870436917759400921994016474570208734121;
            6'd16: xpb[126] = 1024'd103851780072995892721395611529647935593764578409047633209627918091305919581700141577457451749862613922365039899170791304592306113383197797998835628100062151048160559333592132655951300143083881826159135767212938406959199218845861792757530886158130764014569466448469536427090206865324329788025268193308381178884;
            6'd17: xpb[126] = 1024'd17292494564464579967383641696640107009851044215311347189130771673279868052574546243537239073235771560430492837275845685195027364838732409457392761094067754788402588364763227943725577008388720149311433546373317172620878532358055575081142639280591849815365130540911088931203448738960625636937830085420959139316;
            6'd18: xpb[126] = 1024'd54799904740058008612170599268446711170635937147310745296765480320230711860758089819632097611266603507939095182838393500376812457135487355471110019104404399462335291965505540569130093065210764193773928933920935784646918696091146130369732962086282384882980698047469699465423218686525554502969081804159131584079;
            6'd19: xpb[126] = 1024'd92307314915651437256957556840253315331420830079310143404400188967181555668941633395726956149297435455447697528400941315558597549432242301484827277114741044136267995566247853194534609122032808238236424321468554396672958859824236685658323284891972919950596265554028309999642988634090483369000333522897304028842;
            6'd20: xpb[126] = 1024'd5748029407120124502945587007245486747507295885573857383903042549155504139816038061806743472670593093513150466505995696161318800887776912943384410108746647876510024597418948482308885987337646561388722100628933162334638173336430467981935038014434005751391929646469862503756230507726779217912895415009881989274;
            6'd21: xpb[126] = 1024'd43255439582713553147732544579052090908292188817573255491537751196106347947999581637901602010701425041021752812068543511343103893184531858957101668119083292550442728198161261107713402044159690605851217488176551774360678337069521023270525360820124540819007497153028473037976000455291708083944147133748054434037;
            6'd22: xpb[126] = 1024'd80762849758306981792519502150858695069077081749572653599172459843057191756183125213996460548732256988530355157631091326524888985481286804970818926129419937224375431798903573733117918100981734650313712875724170386386718500802611578559115683625815075886623064659587083572195770402856636949975398852486226878800;
            6'd23: xpb[126] = 1024'd118270259933900410437306459722665299229861974681572051706807168490008035564366668790091319086763088936038957503193639141706674077778041750984536184139756581898308135399645886358522434157803778694776208263271788998412758664535702133847706006431505610954238632166145694106415540350421565816006650571224399323563;
            6'd24: xpb[126] = 1024'd31710974425369097683294489889657470645948440487835765686310022071981984035241073456171106410136246574104410441298693522309395329233576362443093317133762185638550164430816981646296711023108617017928506042432167764074437978047895916171317759553966696755034296258587246610528782224057861664919212463336977283995;
            6'd25: xpb[126] = 1024'd69218384600962526328081447461464074806733333419835163793944730718932827843424617032265964948167078521613012786861241337491180421530331308456810575144098830312482868031559294271701227079930661062391001429979786376100478141780986471459908082359657231822649863765145857144748552171622790530950464182075149728758;
            6'd26: xpb[126] = 1024'd106725794776555954972868405033270678967518226351834561901579439365883671651608160608360823486197910469121615132423789152672965513827086254470527833154435474986415571632301606897105743136752705106853496817527404988126518305514077026748498405165347766890265431271704467678968322119187719396981715900813322173521;
            6'd27: xpb[126] = 1024'd20166509268024642218856435200262850383604692158098275881082292947857620122482565274440610809571068107187068070528843533275686765282620865929084966148441078726657600663472702184880020002057543430005794596687783753788197619026270809072110158287808852691061095364146020183081563992824015245894277792925900133953;
            6'd28: xpb[126] = 1024'd57673919443618070863643392772069454544389585090097673988717001594808463930666108850535469347601900054695670416091391348457471857579375811942802224158777723400590304264215014810284536058879587474468289984235402365814237782759361364360700481093499387758676662870704630717301333940388944111925529511664072578716;
            6'd29: xpb[126] = 1024'd95181329619211499508430350343876058705174478022097072096351710241759307738849652426630327885632732002204272761653939163639256949876130757956519482169114368074523007864957327435689052115701631518930785371783020977840277946492451919649290803899189922826292230377263241251521103887953872977956781230402245023479;
            6'd30: xpb[126] = 1024'd8622044110680186754418380510868230121260943828360786075854563823733256209724057092710115209005889640269725699758993544241978201331665369415076615163119971814765036896128422723463328981006469842083083150943399743501957260004645701972902557021651008627087894469704793755634345761590168826869343122514822983911;
            6'd31: xpb[126] = 1024'd46129454286273615399205338082674834282045836760360184183489272470684100017907600668804973747036721587778328045321541359423763293628420315428793873173456616488697740496870735348867845037828513886545578538491018355527997423737736257261492879827341543694703461976263404289854115709155097692900594841252995428674;
            6'd32: xpb[126] = 1024'd83636864461867044043992295654481438442830729692359582291123981117634943826091144244899832285067553535286930390884089174605548385925175261442511131183793261162630444097613047974272361094650557931008073926038636967554037587470826812550083202633032078762319029482822014824073885656720026558931846559991167873437;
            6'd33: xpb[126] = 1024'd121144274637460472688779253226288042603615622624358980398758689764585787634274687820994690823098385482795532736446636989787333478221930207456228389194129905836563147698355360599676877151472601975470569313586255579580077751203917367838673525438722613829934596989380625358293655604284955424963098278729340318200;
            6'd34: xpb[126] = 1024'd34584989128929159934767283393280214019702088430622694378261543346559736105149092487074478146471543120860985674551691370390054729677464818914785522188135509576805176729526455887451154016777440298622867092746634345241757064716111150162285278561183699630730261081822177862406897477921251273875660170841918278632;
            6'd35: xpb[126] = 1024'd72092399304522588579554240965086818180486981362622092485896251993510579913332636063169336684502375068369588020114239185571839821974219764928502780198472154250737880330268768512855670073599484343085362480294252957267797228449201705450875601366874234698345828588380788396626667425486180139906911889580090723395;
            6'd36: xpb[126] = 1024'd109599809480116017224341198536893422341271874294621490593530960640461423721516179639264195222533207015878190365676787000753624914270974710942220038208808798924670583931011081138260186130421528387547857867841871569293837392182292260739465924172564769765961396094939398930846437373051109005938163608318263168158;
            6'd37: xpb[126] = 1024'd23040523971584704470329228703885593757358340100885204573033814222435372192390584305343982545906364653943643303781841381356346165726509322400777171202814402664912612962182176426034462995726366710700155647002250334955516705694486043063077677295025855566757060187380951434959679246687404854850725500430841128590;
            6'd38: xpb[126] = 1024'd60547934147178133115116186275692197918143233032884602680668522869386216000574127881438841083937196601452245649344389196538131258023264268414494429213151047338845316562924489051438979052548410755162651034549868946981556869427576598351668000100716390634372627693939561969179449194252333720881977219169013573353;
            6'd39: xpb[126] = 1024'd98055344322771561759903143847498802078928125964884000788303231516337059808757671457533699621968028548960847994906937011719916350320019214428211687223487692012778020163666801676843495109370454799625146422097487559007597033160667153640258322906406925701988195200498172503399219141817262586913228937907186018116;
            6'd40: xpb[126] = 1024'd11496058814240249005891174014490973495014591771147714767806085098311008279632076123613486945341186187026300933011991392322637601775553825886768820217493295753020049194837896964617771974675293122777444201257866324669276346672860935963870076028868011502783859292939725007512461015453558435825790830019763978548;
            6'd41: xpb[126] = 1024'd49003468989833677650678131586297577655799484703147112875440793745261852087815619699708345483372018134534903278574539207504422694072308771900486078227829940426952752795580209590022288031497337167239939588805484936695316510405951491252460398834558546570399426799498335541732230963018487301857042548757936423311;
            6'd42: xpb[126] = 1024'd86510879165427106295465089158104181816584377635146510983075502392212695895999163275803204021402850082043505624137087022686207786369063717914203336238166585100885456396322522215426804088319381211702434976353103548721356674139042046541050721640249081638014994306056946075952000910583416167888294267496108868074;
            6'd43: xpb[126] = 1024'd124018289341020534940252046729910785977369270567145909090710211039163539704182706851898062559433682029552107969699634837867992878665818663927920594248503229774818159997064834840831320145141425256164930363900722160747396837872132601829641044445939616705630561812615556610171770858148345033919545986234281312837;
            6'd44: xpb[126] = 1024'd37459003832489222186240076896902957393455736373409623070213064621137488175057111517977849882806839667617560907804689218470714130121353275386477727242508833515060189028235930128605597010446263579317228143061100926409076151384326384153252797568400702506426225905057109114285012731784640882832107878346859273269;
            6'd45: xpb[126] = 1024'd74966414008082650831027034468709561554240629305409021177847773268088331983240655094072708420837671615126163253367237033652499222418108221400194985252845478188992892628978242754010113067268307623779723530608719538435116315117416939441843120374091237574041793411615719648504782679349569748863359597085031718032;
            6'd46: xpb[126] = 1024'd112473824183676079475813992040516165715025522237408419285482481915039175791424198670167566958868503562634765598929784848834284314714863167413912243263182122862925596229720555379414629124090351668242218918156338150461156478850507494730433443179781772641657360918174330182724552626914498614894611315823204162795;
            6'd47: xpb[126] = 1024'd25914538675144766721802022207508337131111988043672133264985335497013124262298603336247354282241661200700218537034839229437005566170397778872469376257187726603167625260891650667188905989395189991394516697316716916122835792362701277054045196302242858442453025010615882686837794500550794463807173207935782123227;
            6'd48: xpb[126] = 1024'd63421948850738195366588979779314941291896880975671531372620044143963968070482146912342212820272493148208820882597387044618790658467152724886186634267524371277100328861633963292593422046217234035857012084864335528148875956095791832342635519107933393510068592517174493221057564448115723329838424926673954567990;
            6'd49: xpb[126] = 1024'd100929359026331624011375937351121545452681773907670929480254752790914811878665690488437071358303325095717423228159934859800575750763907670899903892277861015951033032462376275917997938103039278080319507472411954140174916119828882387631225841913623928577684160023733103755277334395680652195869676645412127012753;
            6'd50: xpb[126] = 1024'd14370073517800311257363967518113716868768239713934643459757606372888760349540095154516858681676482733782876166264989240403297002219442282358461025271866619691275061493547371205772214968344116403471805251572332905836595433341076169954837595036085014378479824116174656259390576269316948044782238537524704973185;
            6'd51: xpb[126] = 1024'd51877483693393739902150925089920321029553132645934041567392315019839604157723638730611717219707314681291478511827537055585082094516197228372178283282203264365207765094289683831176731025166160447934300639119951517862635597074166725243427917841775549446095391622733266793610346216881876910813490256262877417948;
            6'd52: xpb[126] = 1024'd89384893868987168546937882661726925190338025577933439675027023666790447965907182306706575757738146628800080857390084870766867186812952174385895541292539909039140468695031996456581247081988204492396796026667570129888675760807257280532018240647466084513710959129291877327830116164446805776844741975001049862711;
            6'd53: xpb[126] = 1024'd2825608360455855792925912828719096606424491384197153654529877248764396436781586972786363081111304266865533795495139251369588438268486785844452674286545512779382497726203091744355523947293042815549093805827948895550355074319451062855629993769927170314506623221733429831943358038083101625757303867113627823143;
            6'd54: xpb[126] = 1024'd40333018536049284437712870400525700767209384316196551762164585895715240244965130548881221619142136214374136141057687066551373530565241731858169932296882157453315201326945404369760040004115086860011589193375567507576395238052541618144220316575617705382122190728292040366163127985648030491788555585851800267906;
            6'd55: xpb[126] = 1024'd77840428711642713082499827972332304927994277248195949869799294542666084053148674124976080157172968161882738486620234881733158622861996677871887190307218802127247904927687716995164556060937130904474084580923186119602435401785632173432810639381308240449737758234850650900382897933212959357819807304589972712669;
            6'd56: xpb[126] = 1024'd115347838887236141727286785544138909088779170180195347977434003189616927861332217701070938695203800109391340832182782696914943715158751623885604448317555446801180608528430029620569072117759174948936579968470804731628475565518722728721400962186998775517353325741409261434602667880777888223851059023328145157432;
            6'd57: xpb[126] = 1024'd28788553378704828973274815711131080504865635986459061956936856771590876332206622367150726018576957747456793770287837077517664966614286235344161581311561050541422637559601124908343348983064013272088877747631183497290154879030916511045012715309459861318148989833850813938715909754414184072763620915440723117864;
            6'd58: xpb[126] = 1024'd66295963554298257618061773282937684665650528918458460064571565418541720140390165943245584556607789694965396115850384892699450058911041181357878839321897695215355341160343437533747865039886057316551373135178802109316195042764007066333603038115150396385764557340409424472935679701979112938794872634178895562627;
            6'd59: xpb[126] = 1024'd103803373729891686262848730854744288826435421850457858172206274065492563948573709519340443094638621642473998461412932707881235151207796127371596097332234339889288044761085750159152381096708101361013868522726420721342235206497097621622193360920840931453380124846968035007155449649544041804826124352917068007390;
            6'd60: xpb[126] = 1024'd17244088221360373508836761021736460242521887656721572151709127647466512419448114185420230418011779280539451399517987088483956402663330738830153230326239943629530073792256845446926657962012939684166166301886799487003914520009291403945805114043302017254175788939409587511268691523180337653738686245029645967822;
            6'd61: xpb[126] = 1024'd54751498396953802153623718593543064403306780588720970259343836294417356227631657761515088956042611228048053745080534903665741494960085684843870488336576588303462777392999158072331174018834983728628661689434418099029954683742381959234395436848992552321791356445968198045488461470745266519769937963767818412585;
            6'd62: xpb[126] = 1024'd92258908572547230798410676165349668564091673520720368366978544941368200035815201337609947494073443175556656090643082718847526587256840630857587746346913232977395480993741470697735690075657027773091157076982036711055994847475472514522985759654683087389406923952526808579708231418310195385801189682505990857348;
            6'd63: xpb[126] = 1024'd5699623064015918044398706332341839980178139326984082346481398523342148506689606003689734817446600813622109028748137099450247838712375242316144879340918836717637510024912565985509966940961866096243454856142415476717674160987666296846597512777144173190202588044968361083821473291946491234713751574618568817780;
        endcase
    end

    always_comb begin
        case(flag[42][11:6])
            6'd0: xpb[127] = 1024'd0;
            6'd1: xpb[127] = 1024'd43207033239609346689185663904148444140963032258983480454116107170292992314873149579784593355477432761130711374310684914632032931009130188329862137351255481391570213625654878610914482997783910140705950243690034088743714324720756852135187835582834708257818155551526971618041243239511420100745003293356741262543;
            6'd2: xpb[127] = 1024'd86414066479218693378371327808296888281926064517966960908232214340585984629746299159569186710954865522261422748621369829264065862018260376659724274702510962783140427251309757221828965995567820281411900487380068177487428649441513704270375671165669416515636311103053943236082486479022840201490006586713482525086;
            6'd3: xpb[127] = 1024'd5554404034703298668758064307630899678190669651214757234216466445902081607310309829338708851774623973948984715474561309317034952186170230434426287037435403241019966307393418495113209801834524700807653122682862419866782123941373783440584937065274675506634563240463856824017201644605627285116320053444629303298;
            6'd4: xpb[127] = 1024'd48761437274312645357943728211779343819153701910198237688332573616195073922183459409123302207252056735079696089785246223949067883195300418764288424388690884632590179933048297106027692799618434841513603366372896508610496448662130635575772772648109383764452718791990828442058444884117047385861323346801370565841;
            6'd5: xpb[127] = 1024'd91968470513921992047129392115927787960116734169181718142448680786488066237056608988907895562729489496210407464095931138581100814204430607094150561739946366024160393558703175716942175797402344982219553610062930597354210773382887487710960608230944092022270874343517800060099688123628467486606326640158111828384;
            6'd6: xpb[127] = 1024'd11108808069406597337516128615261799356381339302429514468432932891804163214620619658677417703549247947897969430949122618634069904372340460868852574074870806482039932614786836990226419603669049401615306245365724839733564247882747566881169874130549351013269126480927713648034403289211254570232640106889258606596;
            6'd7: xpb[127] = 1024'd54315841309015944026701792519410243497344371561412994922549040062097155529493769238462011059026680709028680805259807533266102835381470649198714711426126287873610146240441715601140902601452959542321256489055758928477278572603504419016357709713384059271087282032454685266075646528722674670977643400245999869139;
            6'd8: xpb[127] = 1024'd97522874548625290715887456423558687638307403820396475376665147232390147844366918818246604414504113470159392179570492447898135766390600837528576848777381769265180359866096594212055385599236869683027206732745793017220992897324261271151545545296218767528905437583981656884116889768234094771722646693602741131682;
            6'd9: xpb[127] = 1024'd16663212104109896006274192922892699034572008953644271702649399337706244821930929488016126555323871921846954146423683927951104856558510691303278861112306209723059898922180255485339629405503574102422959368048587259600346371824121350321754811195824026519903689721391570472051604933816881855348960160333887909894;
            6'd10: xpb[127] = 1024'd59870245343719242695459856827041143175535041212627752156765506507999237136804079067800719910801304682977665520734368842583137787567640879633140998463561691114630112547835134096254112403287484243128909611738621348344060696544878202456942646778658734777721845272918542090092848173328301956093963453690629172437;
            6'd11: xpb[127] = 1024'd103077278583328589384645520731189587316498073471611232610881613678292229451677228647585313266278737444108376895045053757215170718576771067963003135814817172506200326173490012707168595401071394383834859855428655437087775021265635054592130482361493443035540000824445513708134091412839722056838966747047370434980;
            6'd12: xpb[127] = 1024'd22217616138813194675032257230523598712762678604859028936865865783608326429241239317354835407098495895795938861898245237268139808744680921737705148149741612964079865229573673980452839207338098803230612490731449679467128495765495133762339748261098702026538252961855427296068806578422509140465280213778517213192;
            6'd13: xpb[127] = 1024'd65424649378422541364217921134672042853725710863842509390981972953901318744114388897139428762575928656926650236208930151900172739753811110067567285500997094355650078855228552591367322205122008943936562734421483768210842820486251985897527583843933410284356408513382398914110049817933929241210283507135258475735;
            6'd14: xpb[127] = 1024'd108631682618031888053403585038820486994688743122825989845098080124194311058987538476924022118053361418057361610519615066532205670762941298397429422852252575747220292480883431202281805202905919084642512978111517856954557145207008838032715419426768118542174564064909370532151293057445349341955286800491999738278;
            6'd15: xpb[127] = 1024'd27772020173516493343790321538154498390953348256073786171082332229510408036551549146693544258873119869744923577372806546585174760930851152172131435187177016205099831536967092475566049009172623504038265613414312099333910619706868917202924685326373377533172816202319284120086008223028136425581600267223146516490;
            6'd16: xpb[127] = 1024'd70979053413125840032975985442302942531916380515057266625198439399803400351424698726478137614350552630875634951683491461217207691939981340501993572538432497596670045162621971086480532006956533644744215857104346188077624944427625769338112520909208085790990971753846255738127251462539556526326603560579887779033;
            6'd17: xpb[127] = 1024'd114186086652735186722161649346451386672879412774040747079314546570096392666297848306262730969827985392006346325994176375849240622949111528831855709889687978988240258788276849697395015004740443785450166100794380276821339269148382621473300356492042794048809127305373227356168494702050976627071606853936629041576;
            6'd18: xpb[127] = 1024'd33326424208219792012548385845785398069144017907288543405298798675412489643861858976032253110647743843693908292847367855902209713117021382606557722224612419446119797844360510970679258811007148204845918736097174519200692743648242700643509622391648053039807379442783140944103209867633763710697920320667775819788;
            6'd19: xpb[127] = 1024'd76533457447829138701734049749933842210107050166272023859414905845705481958735008555816846466125176604824619667158052770534242644126151570936419859575867900837690011470015389581593741808791058345551868979787208607944407068368999552778697457974482761297625534994310112562144453107145183811442923614024517082331;
            6'd20: xpb[127] = 1024'd119740490687438485390919713654082286351070082425255504313531013015998474273608158135601439821602609365955331041468737685166275575135281759266281996927123382229260225095670268192508224806574968486257819223477242696688121393089756404913885293557317469555443690545837084180185696346656603912187926907381258344874;
            6'd21: xpb[127] = 1024'd38880828242923090681306450153416297747334687558503300639515265121314571251172168805370961962422367817642893008321929165219244665303191613040984009262047822687139764151753929465792468612841672905653571858780036939067474867589616484084094559456922728546441942683246997768120411512239390995814240374112405123086;
            6'd22: xpb[127] = 1024'd82087861482532437370492114057564741888297719817486781093631372291607563566045318385155555317899800578773604382632614079851277596312321801370846146613303304078709977777408808076706951610625583046359522102470071027811189192310373336219282395039757436804260098234773969386161654751750811096559243667469146385629;
            6'd23: xpb[127] = 1024'd1228199038017042660878850556898753284562324950734577419615624396923660543609329054925077458719559030461166349485805559904246686480231655145548158948227744536589516833492469349991195416892287465755274737772865270190542666810233415389491660939362695795258350372183882974096369917333598180185557134200293163841;
            6'd24: xpb[127] = 1024'd44435232277626389350064514461047197425525357209718057873731731567216652858482478634709670814196991791591877723796490474536279617489361843475410296299483225928159730459147347960905678414676197606461224981462899358934256991530990267524679496522197404053076505923710854592137613156845018280930560427557034426384;
            6'd25: xpb[127] = 1024'd87642265517235736039250178365195641566488389468701538327847838737509645173355628214494264169674424552722589098107175389168312548498492031805272433650738707319729944084802226571820161412460107747167175225152933447677971316251747119659867332105032112310894661475237826210178856396356438381675563720913775688927;
            6'd26: xpb[127] = 1024'd6782603072720341329636914864529652962752994601949334653832090842825742150919638884263786310494183004410151064960366869221281638666401885579974445985663147777609483140885887845104405218726812166562927860455727690057324790751607198830076598004637371301892913612647739798113571561939225465301877187644922467139;
            6'd27: xpb[127] = 1024'd49989636312329688018822578768678097103716026860932815107948198013118734465792788464048379665971615765540862439271051783853314569675532073909836583336918629169179696766540766456018888216510722307268878104145761778801039115472364050965264433587472079559711069164174711416154814801450645566046880481001663729682;
            6'd28: xpb[127] = 1024'd93196669551939034708008242672826541244679059119916295562064305183411726780665938043832973021449048526671573813581736698485347500684662262239698720688174110560749910392195645066933371214294632447974828347835795867544753440193120903100452269170306787817529224715701683034196058040962065666791883774358404992225;
            6'd29: xpb[127] = 1024'd12337007107423639998394979172160552640943664253164091888048557288727823758229948713602495162268806978359135780434928178538316590852572116014400733023098551018629449448279306340217615020561336867370580983138590109924106914692980982270661535069912046808527476853111596622130773206544852750418197241089551770437;
            6'd30: xpb[127] = 1024'd55544040347032986687580643076308996781906696512147572342164664459020816073103098293387088517746239739489847154745613093170349521861702304344262870374354032410199663073934184951132098018345247008076531226828624198667821239413737834405849370652746755066345632404638568240172016446056272851163200534446293032980;
            6'd31: xpb[127] = 1024'd98751073586642333376766306980457440922869728771131052796280771629313808387976247873171681873223672500620558529056298007802382452870832492674125007725609513801769876699589063562046581016129157148782481470518658287411535564134494686541037206235581463324163787956165539858213259685567692951908203827803034295523;
            6'd32: xpb[127] = 1024'd17891411142126938667153043479791452319134333904378849122265023734629905365540258542941204014043430952308120495909489487855351543038742346448827020060533954259649415755672724835330824822395861568178234105821452529790889038634354765711246472135186722315162040093575453446147974851150480035534517294534181073735;
            6'd33: xpb[127] = 1024'd61098444381736285356338707383939896460097366163362329576381130904922897680413408122725797369520863713438831870220174402487384474047872534778689157411789435651219629381327603446245307820179771708884184349511486618534603363355111617846434307718021430572980195645102425064189218090661900136279520587890922336278;
            6'd34: xpb[127] = 1024'd104305477621345632045524371288088340601060398422345810030497238075215889995286557702510390724998296474569543244530859317119417405057002723108551294763044917042789843006982482057159790817963681849590134593201520707278317688075868469981622143300856138830798351196629396682230461330173320237024523881247663598821;
            6'd35: xpb[127] = 1024'd23445815176830237335911107787422351997325003555593606356481490180531986972850568372279912865818054926257105211384050797172386495224912576883253307097969357500669382063066143330444034624230386268985887228504314949657671162575728549151831409200461397821796603334039310270165176495756107320650837347978810377033;
            6'd36: xpb[127] = 1024'd66652848416439584025096771691570796138288035814577086810597597350824979287723717952064506221295487687387816585694735711804419426234042765213115444449224838892239595688721021941358517622014296409691837472194349038401385487296485401287019244783296106079614758885566281888206419735267527421395840641335551639576;
            6'd37: xpb[127] = 1024'd109859881656048930714282435595719240279251068073560567264713704521117971602596867531849099576772920448518527960005420626436452357243172953542977581800480320283809809314375900552273000619798206550397787715884383127145099812017242253422207080366130814337432914437093253506247662974778947522140843934692292902119;
            6'd38: xpb[127] = 1024'd29000219211533536004669172095053251675515673206808363590697956626434068580160878201618621717592678900206089926858612106489421447411082807317679594135404760741689348370459561825557244426064910969793540351187177369524453286517102332592416346265736073328431166574503167094182378140361734605767157401423439680331;
            6'd39: xpb[127] = 1024'd72207252451142882693854835999201695816478705465791844044814063796727060895034027781403215073070111661336801301169297021121454378420212995647541731486660242133259561996114440436471727423848821110499490594877211458268167611237859184727604181848570781586249322126030138712223621379873154706512160694780180942874;
            6'd40: xpb[127] = 1024'd115414285690752229383040499903350139957441737724775324498930170967020053209907177361187808428547544422467512675479981935753487309429343183977403868837915723524829775621769319047386210421632731251205440838567245547011881935958616036862792017431405489844067477677557110330264864619384574807257163988136922205417;
            6'd41: xpb[127] = 1024'd34554623246236834673427236402684151353706342858023120824914423072336150187471188030957330569367302874155074642333173415806456399597253037752105881172840163982709314677852980320670454227899435670601193473870039789391235410458476116033001283331010748835065729814967023918199579784967361890883477454868068983629;
            6'd42: xpb[127] = 1024'd77761656485846181362612900306832595494669375117006601279030530242629142502344337610741923924844735635285786016643858330438489330606383226081968018524095645374279528303507858931584937225683345811307143717560073878134949735179232968168189118913845457092883885366493995536240823024478781991628480748224810246172;
            6'd43: xpb[127] = 1024'd120968689725455528051798564210981039635632407375990081733146637412922134817217487190526517280322168396416497390954543245070522261615513414411830155875351126765849741929162737542499420223467255952013093961250107966878664059899989820303376954496680165350702040918020967154282066263990202092373484041581551508715;
            6'd44: xpb[127] = 1024'd40109027280940133342185300710315051031897012509237878059130889518238231794781497860296039421141926848104059357807734725123491351783423268186532168210275567223729280985246398815783664029733960371408846596552902209258017534399849899473586220396285424341700293055430880742216781429572989175999797508312698286927;
            6'd45: xpb[127] = 1024'd83316060520549480031370964614463495172860044768221358513246996688531224109654647440080632776619359609234770732118419639755524282792553456516394305561531048615299494610901277426698147027517870512114796840242936298001731859120606751608774055979120132599518448606957852360258024669084409276744800801669439549470;
            6'd46: xpb[127] = 1024'd2456398076034085321757701113797506569124649901469154839231248793847321087218658109850154917439118060922332698971611119808493372960463310291096317896455489073179033666984938699982390833784574931510549475545730540381085333620466830778983321878725391590516700744367765948192739834667196360371114268400586327682;
            6'd47: xpb[127] = 1024'd45663431315643432010943365017945950710087682160452635293347355964140313402091807689634748272916550822053044073282296034440526303969593498620958455247710970464749247292639817310896873831568485072216499719235764629124799658341223682914171157461560099848334856295894737566233983074178616461116117561757327590225;
            6'd48: xpb[127] = 1024'd88870464555252778700129028922094394851050714419436115747463463134433305716964957269419341628393983583183755447592980949072559234978723686950820592598966451856319460918294695921811356829352395212922449962925798717868513983061980535049358993044394808106153011847421709184275226313690036561861120855114068852768;
            6'd49: xpb[127] = 1024'd8010802110737383990515765421428406247315319552683912073447715239749402694528967939188863769213742034871317414446172429125528325146633540725522604933890892314198999974378357195095600635619099632318202598228592960247867457561840614219568258944000067097151263984831622772209941479272823645487434321845215630980;
            6'd50: xpb[127] = 1024'd51217835350346730679701429325576850388278351811667392527563822410042395009402117518973457124691174796002028788756857343757561256155763729055384742285146373705769213600033235806010083633403009773024152841918627048991581782282597466354756094526834775354969419536358594390251184718784243746232437615201956893523;
            6'd51: xpb[127] = 1024'd94424868589956077368887093229725294529241384070650872981679929580335387324275267098758050480168607557132740163067542258389594187164893917385246879636401855097339427225688114416924566631186919913730103085608661137735296107003354318489943930109669483612787575087885566008292427958295663846977440908558698156066;
            6'd52: xpb[127] = 1024'd13565206145440682659273829729059305925505989203898669307664181685651484301839277768527572620988366008820302129920733738442563277332803771159948891971326295555218966281771775690208810437453624333125855720911455380114649581503214397660153196009274742603785827225295479596227143123878450930603754375289844934278;
            6'd53: xpb[127] = 1024'd56772239385050029348459493633207750066469021462882149761780288855944476616712427348312165976465798769951013504231418653074596208341933959489811029322581776946789179907426654301123293435237534473831805964601489468858363906223971249795341031592109450861603982776822451214268386363389871031348757668646586196821;
            6'd54: xpb[127] = 1024'd99979272624659376037645157537356194207432053721865630215896396026237468931585576928096759331943231531081724878542103567706629139351064147819673166673837258338359393533081532912037776433021444614537756208291523557602078230944728101930528867174944159119422138328349422832309629602901291132093760962003327459364;
            6'd55: xpb[127] = 1024'd19119610180143981328031894036690205603696658855113426541880648131553565909149587597866281472762989982769286845395295047759598229518974001594375179008761698796238932589165194185322020239288149033933508843594317799981431705444588181100738133074549418110420390465759336420244344768484078215720074428734474237576;
            6'd56: xpb[127] = 1024'd62326643419753328017217557940838649744659691114096906995996755301846558224022737177650874828240422743899998219705979962391631160528104189924237316360017180187809146214820072796236503237072059174639459087284351888725146030165345033235925968657384126368238546017286308038285588007995498316465077722091215500119;
            6'd57: xpb[127] = 1024'd105533676659362674706403221844987093885622723373080387450112862472139550538895886757435468183717855505030709594016664877023664091537234378254099453711272661579379359840474951407150986234855969315345409330974385977468860354886101885371113804240218834626056701568813279656326831247506918417210081015447956762662;
            6'd58: xpb[127] = 1024'd24674014214847279996789958344321105281887328506328183776097114577455647516459897427204990324537613956718271560869856357076633181705144232028801466046197102037258898896558612680435230041122673734741161966277180219848213829385961964541323070139824093617054953706223193244261546413089705500836394482179103540874;
            6'd59: xpb[127] = 1024'd67881047454456626685975622248469549422850360765311664230213221747748639831333047006989583680015046717848982935180541271708666112714274420358663603397452583428829112522213491291349713038906583875447112209967214308591928154106718816676510905722658801874873109257750164862302789652601125601581397775535844803417;
            6'd60: xpb[127] = 1024'd111088080694065973375161286152617993563813393024295144684329328918041632146206196586774177035492479478979694309491226186340699043723404608688525740748708064820399326147868369902264196036690494016153062453657248397335642478827475668811698741305493510132691264809277136480344032892112545702326401068892586065960;
            6'd61: xpb[127] = 1024'd30228418249550578665548022651952004960077998157542941010313581023357729123770207256543699176312237930667256276344417666393668133891314462463227753083632505278278865203952031175548439842957198435548815088960042639714995953327335747981908007205098769123689516946687050068278748057695332785952714535623732844172;
            6'd62: xpb[127] = 1024'd73435451489159925354733686556100449101041030416526421464429688193650721438643356836328292531789670691797967650655102581025701064900444650793089890434887986669849078829606909786462922840741108576254765332650076728458710278048092600117095842787933477381507672498214021686319991297206752886697717828980474106715;
            6'd63: xpb[127] = 1024'd116642484728769272043919350460248893242004062675509901918545795363943713753516506416112885887267103452928679024965787495657733995909574839122952027786143468061419292455261788397377405838525018716960715576340110817202424602768849452252283678370768185639325828049740993304361234536718172987442721122337215369258;
        endcase
    end

    always_comb begin
        case(flag[42][16:12])
            5'd0: xpb[128] = 1024'd0;
            5'd1: xpb[128] = 1024'd35782822284253877334306086959582904638268667808757698244530047469259810731080517085882408028086861904616240991818978975710703086077484692897654040121067908519298831511345449670661649644791723136356468211642905059581778077268709531422492944270373444630324080187150906892295949702300960071069034589068362147470;
            5'd2: xpb[128] = 1024'd71565644568507754668612173919165809276537335617515396489060094938519621462161034171764816056173723809232481983637957951421406172154969385795308080242135817038597663022690899341323299289583446272712936423285810119163556154537419062844985888540746889260648160374301813784591899404601920142138069178136724294940;
            5'd3: xpb[128] = 1024'd107348466852761632002918260878748713914806003426273094733590142407779432193241551257647224084260585713848722975456936927132109258232454078692962120363203725557896494534036349011984948934375169409069404634928715178745334231806128594267478832811120333890972240561452720676887849106902880213207103767205086442410;
            5'd4: xpb[128] = 1024'd19064593452890767938425420433517185808376244109295108849988334812062347587012929433514560897689773309021814559818422468263748503468718437035456035467940593143504651475810581345016359387649686824115675238184380391962751458853941352724993207398264329254476417334486569539077270735275207267157448529647854105549;
            5'd5: xpb[128] = 1024'd54847415737144645272731507393100090446644911918052807094518382281322158318093446519396968925776635213638055551637401443974451589546203129933110075589008501662803482987156031015678009032441409960472143449827285451544529536122650884147486151668637773884800497521637476431373220437576167338226483118716216253019;
            5'd6: xpb[128] = 1024'd90630238021398522607037594352682995084913579726810505339048429750581969049173963605279376953863497118254296543456380419685154675623687822830764115710076410182102314498501480686339658677233133096828611661470190511126307613391360415569979095939011218515124577708788383323669170139877127409295517707784578400489;
            5'd7: xpb[128] = 1024'd2346364621527658542544753907451466978483820409832519455446622154864884442945341781146713767292684713427388127817865960816793920859952181173258030814813277767710471440275713019371069130507650511874882264725855724343724840439173174027493470526155213878628754481822232185858591768249454463245862470227346063628;
            5'd8: xpb[128] = 1024'd38129186905781535876850840867034371616752488218590217699976669624124695174025858867029121795379546618043629119636844936527497006937436874070912070935881186287009302951621162690032718775299373648231350476368760783925502917707882705449986414796528658508952834668973139078154541470550414534314897059295708211098;
            5'd9: xpb[128] = 1024'd73912009190035413211156927826617276255021156027347915944506717093384505905106375952911529823466408522659870111455823912238200093014921566968566111056949094806308134462966612360694368420091096784587818688011665843507280994976592236872479359066902103139276914856124045970450491172851374605383931648364070358568;
            5'd10: xpb[128] = 1024'd109694831474289290545463014786200180893289823836105614189036764562644316636186893038793937851553270427276111103274802887948903179092406259866220151178017003325606965974312062031356018064882819920944286899654570903089059072245301768294972303337275547769600995043274952862746440875152334676452966237432432506038;
            5'd11: xpb[128] = 1024'd21410958074418426480970174340968652786860064519127628305434956966927232029958271214661274664982458022449202687636288429080542424328670618208714066282753870911215122916086294364387428518157337335990557502910236116306476299293114526752486677924419543133105171816308801724935862503524661730403310999875200169177;
            5'd12: xpb[128] = 1024'd57193780358672303815276261300551557425128732327885326549965004436187042761038788300543682693069319927065443679455267404791245510406155311106368106403821779430513954427431744035049078162949060472347025714553141175888254376561824058174979622194792987763429252003459708617231812205825621801472345588943562316647;
            5'd13: xpb[128] = 1024'd92976602642926181149582348260134462063397400136643024794495051905446853492119305386426090721156181831681684671274246380501948596483640004004022146524889687949812785938777193705710727807740783608703493926196046235470032453830533589597472566465166432393753332190610615509527761908126581872541380178011924464117;
            5'd14: xpb[128] = 1024'd4692729243055317085089507814902933956967640819665038910893244309729768885890683562293427534585369426854776255635731921633587841719904362346516061629626555535420942880551426038742138261015301023749764529451711448687449680878346348054986941052310427757257508963644464371717183536498908926491724940454692127256;
            5'd15: xpb[128] = 1024'd40475551527309194419395594774485838595236308628422737155423291778989579616971200648175835562672231331471017247454710897344290927797389055244170101750694464054719774391896875709403787905807024160106232741094616508269227758147055879477479885322683872387581589150795371264013133238799868997560759529523054274726;
            5'd16: xpb[128] = 1024'd76258373811563071753701681734068743233504976437180435399953339248249390348051717734058243590759093236087258239273689873054994013874873748141824141871762372574018605903242325380065437550598747296462700952737521567851005835415765410899972829593057317017905669337946278156309082941100829068629794118591416422196;
            5'd17: xpb[128] = 1024'd112041196095816949088007768693651647871773644245938133644483386717509201079132234819940651618845955140703499231092668848765697099952358441039478181992830281093317437414587775050727087195390470432819169164380426627432783912684474942322465773863430761648229749525097185048605032643401789139698828707659778569666;
            5'd18: xpb[128] = 1024'd23757322695946085023514928248420119765343884928960147760881579121792116472903612995807988432275142735876590815454154389897336345188622799381972097097567148678925594356362007383758497648664987847865439767636091840650201139732287700779980148450574757011733926298131033910794454271774116193649173470102546232805;
            5'd19: xpb[128] = 1024'd59540144980199962357821015208003024403612552737717846005411626591051927203984130081690396460362004640492831807273133365608039431266107492279626137218635057198224425867707457054420147293456710984221907979278996900231979217000997232202473092720948201642058006485281940803090403974075076264718208059170908380275;
            5'd20: xpb[128] = 1024'd95322967264453839692127102167585929041881220546475544249941674060311737935064647167572804488448866545109072799092112341318742517343592185177280177339702965717523257379052906725081796938248434120578376190921901959813757294269706763624966036991321646272382086672432847695386353676376036335787242648239270527745;
            5'd21: xpb[128] = 1024'd7039093864582975627634261722354400935451461229497558366339866464594653328836025343440141301878054140282164383453597882450381762579856543519774092444439833303131414320827139058113207391522951535624646794177567173031174521317519522082480411578465641635886263445466696557575775304748363389737587410682038190884;
            5'd22: xpb[128] = 1024'd42821916148836852961940348681937305573720129038255256610869913933854464059916542429322549329964916044898405375272576858161084848657341236417428132565507741822430245832172588728774857036314674671981115005820472232612952598586229053504973355848839086266210343632617603449871725007049323460806621999750400338354;
            5'd23: xpb[128] = 1024'd78604738433090730296246435641520210211988796847012954855399961403114274790997059515204957358051777949514646367091555833871787934734825929315082172686575650341729077343518038399436506681106397808337583217463377292194730675854938584927466300119212530896534423819768510342167674709350283531875656588818762485824;
            5'd24: xpb[128] = 1024'd114387560717344607630552522601103114850257464655770653099930008872374085522077576601087365386138639854130887358910534809582491020812310622212736212807643558861027908854863488070098156325898120944694051429106282351776508753123648116349959244389585975526858504006919417234463624411651243602944691177887124633294;
            5'd25: xpb[128] = 1024'd26103687317473743566059682155871586743827705338792667216328201276657000915848954776954702199567827449303978943272020350714130266048574980555230127912380426446636065796637720403129566779172638359740322032361947564993925980171460874807473618976729970890362680779953266096653046040023570656895035940329892296433;
            5'd26: xpb[128] = 1024'd61886509601727620900365769115454491382096373147550365460858248745916811646929471862837110227654689353920219935090999326424833352126059673452884168033448334965934897307983170073791216423964361496096790244004852624575704057440170406229966563247103415520686760967104172988948995742324530727964070529398254443903;
            5'd27: xpb[128] = 1024'd97669331885981498234671856075037396020365040956308063705388296215176622378009988948719518255741551258536460926909978302135536438203544366350538208154516243485233728819328619744452866068756084632453258455647757684157482134708879937652459507517476860151010841154255079881244945444625490799033105118466616591373;
            5'd28: xpb[128] = 1024'd9385458486110634170179015629805867913935281639330077821786488619459537771781367124586855069170738853709552511271463843267175683439808724693032123259253111070841885761102852077484276522030602047499529058903422897374899361756692696109973882104620855514515017927288928743434367072997817852983449880909384254512;
            5'd29: xpb[128] = 1024'd45168280770364511504485102589388772552203949448087776066316536088719348502861884210469263097257600758325793503090442818977878769517293417590686163380321019590140717272448301748145926166822325183855997270546327956956677439025402227532466826374994300144839098114439835635730316775298777924052484469977746401982;
            5'd30: xpb[128] = 1024'd80951103054618388838791189548971677190472617256845474310846583557979159233942401296351671125344462662942034494909421794688581855594778110488340203501388928109439548783793751418807575811614048320212465482189233016538455516294111758954959770645367744775163178301590742528026266477599737995121519059046108549452;
            5'd31: xpb[128] = 1024'd116733925338872266173097276508554581828741285065603172555376631027238969965022918382234079153431324567558275486728400770399284941672262803385994243622456836628738380295139201089469225456405771456568933693832138076120233593562821290377452714915741189405487258488741649420322216179900698066190553648114470696922;
        endcase
    end

    always_comb begin
        case(flag[43][5:0])
            6'd0: xpb[129] = 1024'd0;
            6'd1: xpb[129] = 1024'd76258373811563071753701681734068743233504976437180435399953339248249390348051717734058243590759093236087258239273689873054994013874873748141824141871762372574018605903242325380065437550598747296462700952737521567851005835415765410899972829593057317017905669337946278156309082941100829068629794118591416422196;
            6'd2: xpb[129] = 1024'd28450051939001402108604436063323053722311525748625186671774823431521885358794296558101415966860512162731367071089886311530924186908527161728488158727193704214346537236913433422500635909680288871615204297087803289337650820610634048834967089502885184768991435261775498282511637808273025120140898410557238360061;
            6'd3: xpb[129] = 1024'd104708425750564473862306117797391796955816502185805622071728162679771275706846014292159659557619605398818625310363576184585918200783400909870312300598956076788365143140155758802566073460279036168077905249825324857188656656026399459734939919095942501786897104599721776438820720749373854188770692529148654782257;
            6'd4: xpb[129] = 1024'd56900103878002804217208872126646107444623051497250373343549646863043770717588593116202831933721024325462734142179772623061848373817054323456976317454387408428693074473826866845001271819360577743230408594175606578675301641221268097669934179005770369537982870523550996565023275616546050240281796821114476720122;
            6'd5: xpb[129] = 1024'd9091782005441134572111626455900417933429600808695124615371131046316265728331171940246004309822443252106842973995969061537778546850707737043640334309818740069021005807497974887436470178442119318382911938525888300161946626416136735604928438915598237289068636447380216691225830483718246291792901113080298657987;
            6'd6: xpb[129] = 1024'd85350155817004206325813308189969161166934577245875560015324470294565656076382889674304247900581536488194101213269658934592772560725581485185464476181581112643039611710740300267501907729040866614845612891263409868012952461831902146504901268508655554306974305785326494847534913424819075360422695231671715080183;
            6'd7: xpb[129] = 1024'd37541833944442536680716062519223471655741126557320311287145954477838151087125468498347420276682955414838210045085855373068702733759234898772128493037012444283367543044411408309937106088122408189998116235613691589499597447026770784439895528418483422058060071709155714973737468291991271411933799523637537018048;
            6'd8: xpb[129] = 1024'd113800207756005608434417744253292214889246102994500746687099293726087541435177186232405663867442048650925468284359545246123696747634108646913952634908774816857386148947653733690002543638721155486460817188351213157350603282442536195339868358011540739075965741047101993130046551233092100480563593642228953440244;
            6'd9: xpb[129] = 1024'd65991885883443938789320498582546525378052652305945497958920777909360036445919765056448836243543467577569577116175741684599626920667762060500616651764206148497714080281324841732437741997802697061613320532701494878837248267637404833274862617921368606827051506970931213256249106100264296532074697934194775378109;
            6'd10: xpb[129] = 1024'd18183564010882269144223252911800835866859201617390249230742262092632531456662343880492008619644886504213685947991938123075557093701415474087280668619637480138042011614995949774872940356884238636765823877051776600323893252832273471209856877831196474578137272894760433382451660967436492583585802226160597315974;
            6'd11: xpb[129] = 1024'd94441937822445340897924934645869579100364178054570684630695601340881921804714061614550252210403979740300944187265627996130551107576289222229104810491399852712060617518238275154938377907482985933228524829789298168174899088248038882109829707424253791596042942232706711538760743908537321652215596344752013738170;
            6'd12: xpb[129] = 1024'd46633615949883671252827688975123889589170727366015435902517085524154416815456640438593424586505398666945053019081824434606481280609942635815768827346831184352388548851909383197373576266564527508381028174139579889661544073442907520044823967334081659347128708156535931664963298775709517703726700636717835676035;
            6'd13: xpb[129] = 1024'd122891989761446743006529370709192632822675703803195871302470424772403807163508358172651668177264491903032311258355514307661475294484816383957592969218593556926407154755151708577439013817163274804843729126877101457512549908858672930944796796927138976365034377494482209821272381716810346772356494755309252098231;
            6'd14: xpb[129] = 1024'd75083667888885073361432125038446943311482253114640622574291908955676302174250936996694840553365910829676420090171710746137405467518469797544256986074024888566735086088822816619874212176244816379996232471227383178999194894053541568879791056836966844116120143418311429947474936583982542823867599047275074036096;
            6'd15: xpb[129] = 1024'd27275346016323403716334879367701253800288802426085373846113393138948797184993515820738012929467329756320528921987907184613335640552123211130921002929456220207063017422493924662309410535326357955148735815577664900485839879248410206814785316746794711867205909342140650073677491451154738875378703339240895973961;
            6'd16: xpb[129] = 1024'd103533719827886475470036561101769997033793778863265809246066732387198187533045233554796256520226422992407787161261597057668329654426996959272745144801218592781081623325736250042374848085925105251611436768315186468336845714664175617714758146339852028885111578680086928229986574392255567944008497457832312396157;
            6'd17: xpb[129] = 1024'd55725397955324805824939315431024307522600328174710560517888216570470682543787812378839428896327841919051895993077793496144259827460650372859409161656649924421409554659407358084810046445006646826763940112665468189823490699859044255649752406249679896636197344603916148356189129259427763995519601749798134334022;
            6'd18: xpb[129] = 1024'd7917076082763136179842069760278618011406877486155311789709700753743177554530391202882601272429260845696004824893989934620190000494303786446073178512081256061737485993078466127245244804088188401916443457015749911310135685053912893584746666159507764387283110527745368482391684126599960047030706041763956271887;
            6'd19: xpb[129] = 1024'd84175449894326207933543751494347361244911853923335747189663040001992567902582108936940844863188354081783263064167679807675184014369177534587897320383843628635756091896320791507310682354686935698379144409753271479161141520469678304484719495752565081405188779865691646638700767067700789115660500160355372694083;
            6'd20: xpb[129] = 1024'd36367128021764538288446505823601671733718403234780498461484524185265062913324687760984017239289773008427371895983876246151114187402830948174561337239274960276084023229991899549745880713768477273531647754103553200647786505664546942419713755662392949156274545789520866764903321934872985167171604452321194631948;
            6'd21: xpb[129] = 1024'd112625501833327610042148187557670414967223379671960933861437863433514453261376405495042260830048866244514630135257566119206108201277704696316385479111037332850102629133234224929811318264367224569994348706841074768498792341080312353319686585255450266174180215127467144921212404875973814235801398570912611054144;
            6'd22: xpb[129] = 1024'd64817179960765940397050941886924725456029928983405685133259347616786948272118984319085433206150285171158738967073762557682038374311358109903049495966468664490430560466905332972246516623448766145146852051191356489985437326275180991254680845165278133925265981051296365047414959743146010287312502862878432992009;
            6'd23: xpb[129] = 1024'd17008858088204270751953696216179035944836478294850436405080831800059443282861563143128605582251704097802847798889958996157968547345011523489713512821899996130758491800576441014681714982530307720299355395541638211472082311470049629189675105075106001676351746975125585173617514610318206338823607154844254929874;
            6'd24: xpb[129] = 1024'd93267231899767342505655377950247779178341454732030871805034171048308833630913280877186849173010797333890106038163648869212962561219885271631537654693662368704777097703818766394747152533129055016762056348279159779323088146885815040089647934668163318694257416313071863329926597551419035407453401273435671352070;
            6'd25: xpb[129] = 1024'd45458910027205672860558132279502089667148004043475623076855655231581328641655859701230021549112216260534214869979845307688892734253538685218201671549093700345105029037489874437182350892210596591914559692629441500809733132080683678024642194577991186445343182236901083456129152418591231458964505565401493289935;
            6'd26: xpb[129] = 1024'd121717283838768744614259814013570832900652980480656058476808994479830718989707577435288265139871309496621473109253535180743886748128412433360025813420856072919123634940732199817247788442809343888377260645366963068660738967496449088924615024171048503463248851574847361612438235359692060527594299683992909712131;
            6'd27: xpb[129] = 1024'd73908961966207074969162568342825143389459529792100809748630478663103214000450156259331437515972728423265581941069731619219816921162065846946689830276287404559451566274403307859682986801890885463529763989717244790147383952691317726859609284080876371214334617498676581738640790226864256579105403975958731649996;
            6'd28: xpb[129] = 1024'd26100640093645405324065322672079453878266079103545561020451962846375709011192735083374609892074147349909690772885928057695747094195719260533353847131718736199779497608074415902118185160972427038682267334067526511634028937886186364794603543990704238965420383422505801864843345094036452630616508267924553587861;
            6'd29: xpb[129] = 1024'd102359013905208477077767004406148197111771055540725996420405302094625099359244452817432853482833240585996949012159617930750741108070593008675177989003481108773798103511316741282183622711571174335144968286805048079485034773301951775694576373583761555983326052760452080021152428035137281699246302386515970010057;
            6'd30: xpb[129] = 1024'd54550692032646807432669758735402507600577604852170747692226786277897594369987031641476025858934659512641057843975814369226671281104246422261842005858912440414126034844987849324618821070652715910297471631155329800971679758496820413629570633493589423734411818684281300147354982902309477750757406678481791947922;
            6'd31: xpb[129] = 1024'd6742370160085137787572513064656818089384154163615498964048270461170089380729610465519198235036078439285166675792010807702601454137899835848506022714343772054453966178658957367054019429734257485449974975505611522458324743691689051564564893403417291485497584608110520273557537769481673802268510970447613885787;
            6'd32: xpb[129] = 1024'd83000743971648209541274194798725561322889130600795934364001609709419479728781328199577441825795171675372424915065700680757595468012773583990330164586106144628472572081901282747119456980333004781912675928243133090309330579107454462464537722996474608503403253946056798429866620710582502870898305089039030307983;
            6'd33: xpb[129] = 1024'd35192422099086539896176949127979871811695679912240685635823093892691974739523907023620614201896590602016533746881897119233525641046426997576994181441537476268800503415572390789554655339414546357065179272593414811795975564302323100399531982906302476254489019869886018556069175577754698922409409381004852245848;
            6'd34: xpb[129] = 1024'd111450795910649611649878630862048615045200656349421121035776433140941365087575624757678857792655683838103791986155586992288519654921300745718818323313299848842819109318814716169620092890013293653527880225330936379646981399718088511299504812499359793272394689207832296712378258518855527991039203499596268668044;
            6'd35: xpb[129] = 1024'd63642474038087942004781385191302925534007205660865872307597917324213860098318203581722030168757102764747900817971783430764449827954954159305482340168731180483147040652485824212055291249094835228680383569681218101133626384912957149234499072409187661023480455131661516838580813386027724042550307791562090605909;
            6'd36: xpb[129] = 1024'd15834152165526272359684139520557236022813754972310623579419401507486355109060782405765202544858521691392009649787979869240380000988607572892146357024162512123474971986156932254490489608176376803832886914031499822620271370107825787169493332319015528774566221055490736964783368253199920094061412083527912543774;
            6'd37: xpb[129] = 1024'd92092525977089344113385821254625979256318731409491058979372740755735745457112500139823446135617614927479267889061669742295374014863481321033970498895924884697493577889399257634555927158775124100295587866769021390471277205523591198069466161912072845792471890393437015121092451194300749162691206202119328965970;
            6'd38: xpb[129] = 1024'd44284204104527674468288575583880289745125280720935810251194224939008240467855078963866618511719033854123376720877866180771304187897134734620634515751356216337821509223070365676991125517856665675448091211119303111957922190718459836004460421821900713543557656317266235247295006061472945214202310494085150903835;
            6'd39: xpb[129] = 1024'd120542577916090746221990257317949032978630257158116245651147564187257630815906796697924862102478127090210634960151556053826298201772008482762458657623118588911840115126312691057056563068455412971910792163856824679808928026134225246904433251414958030561463325655212513403604089002573774282832104612676567326031;
            6'd40: xpb[129] = 1024'd72734256043529076576893011647203343467436806469560996922969048370530125826649375521968034478579546016854743791967752492302228374805661896349122674478549920552168046459983799099491761427536954547063295508207106401295573011329093884839427511324785898312549091579041733529806643869745970334343208904642389263896;
            6'd41: xpb[129] = 1024'd24925934170967406931795765976457653956243355781005748194790532553802620837391954346011206854680964943498852623783948930778158547839315309935786691333981252192495977793654907141926959786618496122215798852557388122782217996523962522774421771234613766063634857502870953656009198736918166385854313196608211201761;
            6'd42: xpb[129] = 1024'd101184307982530478685497447710526397189748332218186183594743871802052011185443672080069450445440058179586110863057638803833152561714189058077610833205743624766514583696897232521992397337217243418678499805294909690633223831939727933674394600827671083081540526840817231812318281678018995454484107315199627623957;
            6'd43: xpb[129] = 1024'd53375986109968809040400202039780707678554881529630934866565355985324506196186250904112622821541477106230219694873835242309082734747842471664274850061174956406842515030568340564427595696298784993831003149645191412119868817134596571609388860737498950832626292764646451938520836545191191505995211607165449561822;
            6'd44: xpb[129] = 1024'd5567664237407139395302956369035018167361430841075686138386840168597001206928829728155795197642896032874328526690031680785012907781495885250938866916606288047170446364239448606862794055380326568983506493995473133606513802329465209544383120647326818583712058688475672064723391412363387557506315899131271499687;
            6'd45: xpb[129] = 1024'd81826038048970211149004638103103761400866407278256121538340179416846391554980547462214038788401989268961586765963721553840006921656369633392763008788368660621189052267481773986928231605979073865446207446732994701457519637745230620444355950240384135601617728026421950221032474353464216626136110017722687921883;
            6'd46: xpb[129] = 1024'd34017716176408541503907392432358071889672956589700872810161663600118886565723126286257211164503408195605695597779917992315937094690023046979427025643799992261516983601152882029363429965060615440598710791083276422944164622940099258379350210150212003352703493950251170347235029220636412677647214309688509859748;
            6'd47: xpb[129] = 1024'd110276089987971613257609074166426815123177933026881308210115002848368276913774844020315454755262501431692953837053607865370931108564896795121251167515562364835535589504395207409428867515659362737061411743820797990795170458355864669279323039743269320370609163288197448503544112161737241746277008428279926281944;
            6'd48: xpb[129] = 1024'd62467768115409943612511828495681125611984482338326059481936487031640771924517422844358627131363920358337062668869804303846861281598550208707915184370993696475863520838066315451864065874740904312213915088171079712281815443550733307214317299653097188121694929212026668629746667028909437797788112720245748219809;
            6'd49: xpb[129] = 1024'd14659446242848273967414582824935436100791031649770810753757971214913266935260001668401799507465339284981171500686000742322791454632203622294579201226425028116191452171737423494299264233822445887366418432521361433768460428745601945149311559562925055872780695135855888755949221896081633849299217012211570157674;
            6'd50: xpb[129] = 1024'd90917820054411345721116264559004179334296008086951246153711310463162657283311719402460043098224432521068429739959690615377785468507077370436403343098187400690210058074979748874364701784421193183829119385258883001619466264161367356049284389155982372890686364473802166912258304837182462917929011130802986579870;
            6'd51: xpb[129] = 1024'd43109498181849676076019018888258489823102557398395997425532794646435152294054298226503215474325851447712538571775887053853715641540730784023067359953618732330537989408650856916799900143502734758981622729609164723106111249356235993984278649065810240641772130397631387038460859704354658969440115422768808517735;
            6'd52: xpb[129] = 1024'd119367871993412747829720700622327233056607533835576432825486133894684542642106015960561459065084944683799796811049576926908709655415604532164891501825381104904556595311893182296865337694101482055444323682346686290957117084772001404884251478658867557659677799735577665194769942645455488038069909541360224939931;
            6'd53: xpb[129] = 1024'd71559550120851078184623454951581543545414083147021184097307618077957037652848594784604631441186363610443905642865773365384639828449257945751555518680812436544884526645564290339300536053183023630596827026696968012443762069966870042819245738568695425410763565659406885320972497512627684089581013833326046877796;
            6'd54: xpb[129] = 1024'd23751228248289408539526209280835854034220632458465935369129102261229532663591173608647803817287782537088014474681969803860570001482911359338219535536243768185212457979235398381735734412264565205749330371047249733930407055161738680754239998478523293161849331583236105447175052379799880141092118125291868815661;
            6'd55: xpb[129] = 1024'd100009602059852480293227891014904597267725608895646370769082441509478923011642891342706047408046875773175272713955659676915564015357785107480043677408006140759231063882477723761801171962863312502212031323784771301781412890577504091654212828071580610179755000921182383603484135320900709209721912243883285237857;
            6'd56: xpb[129] = 1024'd52201280187290810648130645344158907756532158207091122040903925692751418022385470166749219784148294699819381545771856115391494188391438521066707694263437472399558995216148831804236370321944854077364534668135053023268057875772372729589207087981408477930840766845011603729686690188072905261233016535849107175722;
            6'd57: xpb[129] = 1024'd4392958314729141003033399673413218245338707518535873312725409876023913033128048990792392160249713626463490377588052553867424361425091934653371711118868804039886926549819939846671568681026395652517038012485334744754702860967241367524201347891236345681926532768840823855889245055245101312744120827814929113587;
            6'd58: xpb[129] = 1024'd80651332126292212756735081407481961478843683955716308712678749124273303381179766724850635751008806862550748616861742426922418375299965682795195852990631176613905532453062265226737006231625142948979738965222856312605708696383006778424174177484293662699832202106787102012198327996345930381373914946406345535783;
            6'd59: xpb[129] = 1024'd32843010253730543111637835736736271967650233267161059984500233307545798391922345548893808127110225789194857448677938865398348548333619096381859869846062508254233463786733373269172204590706684524132242309573138034092353681577875416359168437394121530450917968030616322138400882863518126432885019238372167473648;
            6'd60: xpb[129] = 1024'd109101384065293614865339517470805015201155209704341495384453572555795188739974063282952051717869319025282115687951628738453342562208492844523684011717824880828252069689975698649237642141305431820594943262310659601943359516993640827259141266987178847468823637368562600294709965804618955501514813356963583895844;
            6'd61: xpb[129] = 1024'd61293062192731945220242271800059325689961759015786246656275056739067683750716642106995224093970737951926224519767825176929272735242146258110348028573256212468580001023646806691672840500386973395747446606660941323430004502188509465194135526897006715219909403292391820420912520671791151553025917648929405833709;
            6'd62: xpb[129] = 1024'd13484740320170275575145026129313636178768308327230997928096540922340178761459220931038396470072156878570333351584021615405202908275799671697012045428687544108907932357317914734108038859468514970899949951011223044916649487383378103129129786806834582970995169216221040547115075538963347604537021940895227771574;
            6'd63: xpb[129] = 1024'd89743114131733347328846707863382379412273284764411433328049880170589569109510938665096640060831250114657591590857711488460196922150673419838836187300449916682926538260560240114173476410067262267362650903748744612767655322799143514029102616399891899988900838554167318703424158480064176673166816059486644193770;
        endcase
    end

    always_comb begin
        case(flag[43][11:6])
            6'd0: xpb[130] = 1024'd0;
            6'd1: xpb[130] = 1024'd41934792259171677683749462192636689901079834075856184599871364353862064120253517489139812436932669041301700422673907926936127095184326833425500204155881248323254469594231348156608674769148803842515154248099026334254300307994012151964096876309719767739986604477996538829626713347236372724677920351452466131635;
            6'd2: xpb[130] = 1024'd83869584518343355367498924385273379802159668151712369199742728707724128240507034978279624873865338082603400845347815853872254190368653666851000408311762496646508939188462696313217349538297607685030308496198052668508600615988024303928193752619439535479973208955993077659253426694472745449355840702904932263270;
            6'd3: xpb[130] = 1024'd1737681093390291652449459173095636958541075101832869671482237996609297023451413557404366096140332814461951860564230346229317444711760165721340487451312704036072734213122827132195785115929205806235265135909839156398540073761139682927312059245929853953139910019872558458773611967780485156915071227731803910574;
            6'd4: xpb[130] = 1024'd43672473352561969336198921365732326859620909177689054271353602350471361143704931046544178533073001855763652283238138273165444539896086999146840691607193952359327203807354175288804459885078009648750419384008865490652840381755151834891408935555649621693126514497869097288400325315016857881592991579184270042209;
            6'd5: xpb[130] = 1024'd85607265611733647019948383558369016760700743253545238871224966704333425263958448535683990970005670897065352705912046200101571635080413832572340895763075200682581673401585523445413134654226813491265573632107891824907140689749163986855505811865369389433113118975865636118027038662253230606270911930636736173844;
            6'd6: xpb[130] = 1024'd3475362186780583304898918346191273917082150203665739342964475993218594046902827114808732192280665628923903721128460692458634889423520331442680974902625408072145468426245654264391570231858411612470530271819678312797080147522279365854624118491859707906279820039745116917547223935560970313830142455463607821148;
            6'd7: xpb[130] = 1024'd45410154445952260988648380538827963818161984279521923942835840347080658167156344603948544629213334670225604143802368619394761984607847164868181179058506656395399938020477002421000245001007215454985684519918704647051380455516291517818720994801579475646266424517741655747173937282797343038508062806916073952783;
            6'd8: xpb[130] = 1024'd87344946705123938672397842731464653719241818355378108542707204700942722287409862093088357066146003711527304566476276546330889079792173998293681383214387904718654407614708350577608919770156019297500838768017730981305680763510303669782817871111299243386253028995738194576800650630033715763185983158368540084418;
            6'd9: xpb[130] = 1024'd5213043280170874957348377519286910875623225305498609014446713989827891070354240672213098288420998443385855581692691038687952334135280497164021462353938112108218202639368481396587355347787617418705795407729517469195620221283419048781936177737789561859419730059617675376320835903341455470745213683195411731722;
            6'd10: xpb[130] = 1024'd47147835539342552641097839711923600776703059381354793614318078343689955190607758161352910725353667484687556004366598965624079429319607330589521666509819360431472672233599829553196030116936421261220949655828543803449920529277431200746033054047509329599406334537614214205947549250577828195423134034647877863357;
            6'd11: xpb[130] = 1024'd89082627798514230324847301904560290677782893457210978214189442697552019310861275650492723162286336525989256427040506892560206524503934164015021870665700608754727141827831177709804704886085225103736103903927570137704220837271443352710129930357229097339392939015610753035574262597814200920101054386100343994992;
            6'd12: xpb[130] = 1024'd6950724373561166609797836692382547834164300407331478685928951986437188093805654229617464384561331257847807442256921384917269778847040662885361949805250816144290936852491308528783140463716823224941060543639356625594160295044558731709248236983719415812559640079490233835094447871121940627660284910927215642296;
            6'd13: xpb[130] = 1024'd48885516632732844293547298885019237735244134483187663285800316340299252214059171718757276821494000299149507864930829311853396874031367496310862153961132064467545406446722656685391815232865627067456214791738382959848460603038570883673345113293439183552546244557486772664721161218358313352338205262379681773931;
            6'd14: xpb[130] = 1024'd90820308891904521977296761077655927636323968559043847885671680694161316334312689207897089258426669340451208287604737238789523969215694329736362358117013312790799876040954004842000490002014430909971369039837409294102760911032583035637441989603158951292532849035483311494347874565594686077016125613832147905566;
            6'd15: xpb[130] = 1024'd8688405466951458262247295865478184792705375509164348357411189983046485117257067787021830480701664072309759302821151731146587223558800828606702437256563520180363671065614135660978925579646029031176325679549195781992700368805698414636560296229649269765699550099362792293868059838902425784575356138659019552870;
            6'd16: xpb[130] = 1024'd50623197726123135945996758058114874693785209585020532957282554336908549237510585276161642917634333113611459725495059658082714318743127662032202641412444768503618140659845483817587600348794832873691479927648222116247000676799710566600657172539369037505686154577359331123494773186138798509253276490111485684505;
            6'd17: xpb[130] = 1024'd92557989985294813629746220250751564594865043660876717557153918690770613357764102765301455354567002154913160148168967585018841413927454495457702845568326016826872610254076831974196275117943636716206634175747248450501300984793722718564754048849088805245672759055355869953121486533375171233931196841563951816140;
            6'd18: xpb[130] = 1024'd10426086560341749914696755038573821751246450610997218028893427979655782140708481344426196576841996886771711163385382077375904668270560994328042924707876224216436405278736962793174710695575234837411590815459034938391240442566838097563872355475579123718839460119235350752641671806682910941490427366390823463444;
            6'd19: xpb[130] = 1024'd52360878819513427598446217231210511652326284686853402628764792333517846260961998833566009013774665928073411586059290004312031763454887827753543128863757472539690874872968310949783385464724038679926745063558061272645540750560850249527969231785298891458826064597231889582268385153919283666168347717843289595079;
            6'd20: xpb[130] = 1024'd94295671078685105282195679423847201553406118762709587228636156687379910381215516322705821450707334969375112008733197931248158858639214661179043333019638720862945344467199659106392060233872842522441899311657087606899841058554862401492066108095018659198812669075228428411895098501155656390846268069295755726714;
            6'd21: xpb[130] = 1024'd12163767653732041567146214211669458709787525712830087700375665976265079164159894901830562672982329701233663023949612423605222112982321160049383412159188928252509139491859789925370495811504440643646855951368874094789780516327977780491184414721508977671979370139107909211415283774463396098405498594122627374018;
            6'd22: xpb[130] = 1024'd54098559912903719250895676404306148610867359788686272300247030330127143284413412390970375109914998742535363446623520350541349208166647993474883616315070176575763609086091138081979170580653244486162010199467900429044080824321989932455281291031228745411965974617104448041041997121699768823083418945575093505653;
            6'd23: xpb[130] = 1024'd96033352172075396934645138596942838511947193864542456900118394683989207404666929880110187546847667783837063869297428277477476303350974826900383820470951424899018078680322486238587845349802048328677164447566926763298381132316002084419378167340948513151952579095100986870668710468936141547761339297027559637288;
            6'd24: xpb[130] = 1024'd13901448747122333219595673384765095668328600814662957371857903972874376187611308459234928769122662515695614884513842769834539557694081325770723899610501632288581873704982617057566280927433646449882121087278713251188320590089117463418496473967438831625119280158980467670188895742243881255320569821854431284592;
            6'd25: xpb[130] = 1024'd55836241006294010903345135577401785569408434890519141971729268326736440307864825948374741206055331556997315307187750696770666652878408159196224103766382880611836343299213965214174955696582450292397275335377739585442620898083129615382593350277158599365105884636977006499815609089480253979998490173306897416227;
            6'd26: xpb[130] = 1024'd97771033265465688587094597770038475470488268966375326571600632680598504428118343437514553642988000598299015729861658623706793748062734992621724307922264128935090812893445313370783630465731254134912429583476765919696921206077141767346690226586878367105092489114973545329442322436716626704676410524759363547862;
            6'd27: xpb[130] = 1024'd15639129840512624872045132557860732626869675916495827043340141969483673211062722016639294865262995330157566745078073116063857002405841491492064387061814336324654607918105444189762066043362852256117386223188552407586860663850257146345808533213368685578259190178853026128962507710024366412235641049586235195166;
            6'd28: xpb[130] = 1024'd57573922099684302555794594750497422527949509992352011643211506323345737331316239505779107302195664371459267167751981042999984097590168324917564591217695584647909077512336792346370740812511656098632540471287578741841160971844269298309905409523088453318245794656849564958589221057260739136913561401038701326801;
            6'd29: xpb[130] = 1024'd99508714358855980239544056943134112429029344068208196243082870677207801451569756994918919739128333412760967590425888969936111192774495158343064795373576832971163547106568140502979415581660459941147694719386605076095461279838281450274002285832808221058232399134846103788215934404497111861591481752491167458436;
            6'd30: xpb[130] = 1024'd17376810933902916524494591730956369585410751018328696714822379966092970234514135574043660961403328144619518605642303462293174447117601657213404874513127040360727342131228271321957851159292058062352651359098391563985400737611396829273120592459298539531399100198725584587736119677804851569150712277318039105740;
            6'd31: xpb[130] = 1024'd59311603193074594208244053923593059486490585094184881314693744319955034354767653063183473398335997185921219028316211389229301542301928490638905078669008288683981811725459619478566525928440861904867805607197417898239701045605408981237217468769018307271385704676722123417362833025041224293828632628770505237375;
            6'd32: xpb[130] = 1024'd101246395452246271891993516116229749387570419170041065914565108673817098475021170552323285835268666227222919450990119316165428637486255324064405282824889537007236281319690967635175200697589665747382959855296444232494001353599421133201314345078738075011372309154718662246989546372277597018506552980222971369010;
            6'd33: xpb[130] = 1024'd19114492027293208176944050904052006543951826120161566386304617962702267257965549131448027057543660959081470466206533808522491891829361822934745361964439744396800076344351098454153636275221263868587916495008230720383940811372536512200432651705228393484539010218598143046509731645585336726065783505049843016314;
            6'd34: xpb[130] = 1024'd61049284286464885860693513096688696445031660196017750986175982316564331378219066620587839494476330000383170888880441735458618987013688656360245566120320992720054545938582446610762311044370067711103070743107257054638241119366548664164529528014948161224525614696594681876136444992821709450743703856502309147949;
            6'd35: xpb[130] = 1024'd102984076545636563544442975289325386346111494271873935586047346670426395498472584109727651931408999041684871311554349662394746082198015489785745770276202241043309015532813794767370985813518871553618224991206283388892541427360560816128626404324667928964512219174591220705763158340058082175421624207954775279584;
            6'd36: xpb[130] = 1024'd20852173120683499829393510077147643502492901221994436057786855959311564281416962688852393153683993773543422326770764154751809336541121988656085849415752448432872810557473925586349421391150469674823181630918069876782480885133676195127744710951158247437678920238470701505283343613365821882980854732781646926888;
            6'd37: xpb[130] = 1024'd62786965379855177513142972269784333403572735297850620657658220313173628401670480177992205590616662814845122749444672081687936431725448822081586053571633696756127280151705273742958096160299273517338335879017096211036781193127688347091841587260878015177665524716467240334910056960602194607658775084234113058523;
            6'd38: xpb[130] = 1024'd104721757639026855196892434462421023304652569373706805257529584667035692521923997667132018027549331856146823172118580008624063526909775655507086257727514945079381749745936621899566770929448077359853490127116122545291081501121700499055938463570597782917652129194463779164536770307838567332336695435686579190158;
            6'd39: xpb[130] = 1024'd22589854214073791481842969250243280461033976323827305729269093955920861304868376246256759249824326588005374187334994500981126781252882154377426336867065152468945544770596752718545206507079675481058446766827909033181020958894815878055056770197088101390818830258343259964056955581146307039895925960513450837462;
            6'd40: xpb[130] = 1024'd64524646473245469165592431442879970362113810399683490329140458309782925425121893735396571686756995629307074610008902427917253876437208987802926541022946400792200014364828100875153881276228479323573601014926935367435321266888828030019153646506807869130805434736339798793683668928382679764573846311965916969097;
            6'd41: xpb[130] = 1024'd106459438732417146849341893635516660263193644475539674929011822663644989545375411224536384123689664670608775032682810354853380971621535821228426745178827649115454483959059449031762556045377283166088755263025961701689621574882840181983250522816527636870792039214336337623310382275619052489251766663418383100732;
            6'd42: xpb[130] = 1024'd24327535307464083134292428423338917419575051425660175400751331952530158328319789803661125345964659402467326047899224847210444225964642320098766824318377856505018278983719579850740991623008881287293711902737748189579561032655955560982368829443017955343958740278215818422830567548926792196810997188245254748036;
            6'd43: xpb[130] = 1024'd66262327566635760818041890615975607320654885501516360000622696306392222448573307292800937782897328443769026470573132774146571321148969153524267028474259104828272748577950928007349666392157685129808866150836774523833861340649967712946465705752737723083945344756212357252457280896163164921488917539697720879671;
            6'd44: xpb[130] = 1024'd108197119825807438501791352808612297221734719577372544600494060660254286568826824781940750219829997485070726893247040701082698416333295986949767232630140353151527218172182276163958341161306488972324020398935800858088161648643979864910562582062457490823931949234208896082083994243399537646166837891150187011306;
            6'd45: xpb[130] = 1024'd26065216400854374786741887596434554378116126527493045072233569949139455351771203361065491442104992216929277908463455193439761670676402485820107311769690560541091013196842406982936776738938087093528977038647587345978101106417095243909680888688947809297098650298088376881604179516707277353726068415977058658610;
            6'd46: xpb[130] = 1024'd68000008660026052470491349789071244279195960603349229672104934303001519472024720850205303879037661258230978331137363120375888765860729319245607515925571808864345482791073755139545451508086890936044131286746613680232401414411107395873777764998667577037085254776084915711230892863943650078403988767429524790245;
            6'd47: xpb[130] = 1024'd109934800919197730154240811981707934180275794679205414271976298656863583592278238339345116315970330299532678753811271047312015861045056152671107720081453057187599952385305103296154126277235694778559285534845640014486701722405119547837874641308387344777071859254081454540857606211180022803081909118881990921880;
            6'd48: xpb[130] = 1024'd27802897494244666439191346769530191336657201629325914743715807945748752375222616918469857538245325031391229769027685539669079115388162651541447799221003264577163747409965234115132561854867292899764242174557426502376641180178234926836992947934877663250238560317960935340377791484487762510641139643708862569184;
            6'd49: xpb[130] = 1024'd69737689753416344122940808962166881237737035705182099343587172299610816495476134407609669975177994072692930191701593466605206210572489484966948003376884512900418217004196582271741236624016096742279396422656452836630941488172247078801089824244597430990225164795957474170004504831724135235319059995161328700819;
            6'd50: xpb[130] = 1024'd111672482012588021806690271154803571138816869781038283943458536653472880615729651896749482412110663113994630614375501393541333305756816318392448207532765761223672686598427930428349911393164900584794550670755479170885241796166259230765186700554317198730211769273954012999631218178960507959996980346613794832454;
            6'd51: xpb[130] = 1024'd29540578587634958091640805942625828295198276731158784415198045942358049398674030475874223634385657845853181629591915885898396560099922817262788286672315968613236481623088061247328346970796498705999507310467265658775181253939374609764305007180807517203378470337833493799151403452268247667556210871440666479758;
            6'd52: xpb[130] = 1024'd71475370846806635775390268135262518196278110807014969015069410296220113518927547965014036071318326887154882052265823812834523655284249650688288490828197216936490951217319409403937021739945302548514661558566291993029481561933386761728401883490527284943365074815830032628778116799504620392234131222893132611393;
            6'd53: xpb[130] = 1024'd113410163105978313459139730327899208097357944882871153614940774650082177639181065454153848508250995928456582474939731739770650750468576484113788694984078465259745420811550757560545696509094106391029815806665318327283781869927398913692498759800247052683351679293826571458404830146740993116912051574345598743028;
            6'd54: xpb[130] = 1024'd31278259681025249744090265115721465253739351832991654086680283938967346422125444033278589730525990660315133490156146232127714004811682982984128774123628672649309215836210888379524132086725704512234772446377104815173721327700514292691617066426737371156518380357706052257925015420048732824471282099172470390332;
            6'd55: xpb[130] = 1024'd73213051940196927427839727308358155154819185908847838686551648292829410542378961522418402167458659701616833912830054159063841099996009816409628978279509920972563685430442236536132806855874508354749926694476131149428021635694526444655713942736457138896504984835702591087551728767285105549149202450624936521967;
            6'd56: xpb[130] = 1024'd115147844199368605111589189500994845055899019984704023286423012646691474662632479011558214604391328742918534335503962085999968195180336649835129182435391169295818155024673584692741481625023312197265080942575157483682321943688538596619810819046176906636491589313699129917178442114521478273827122802077402653602;
            6'd57: xpb[130] = 1024'd33015940774415541396539724288817102212280426934824523758162521935576643445576857590682955826666323474777085350720376578357031449523443148705469261574941376685381950049333715511719917202654910318470037582286943971572261401461653975618929125672667225109658290377578610716698627387829217981386353326904274300906;
            6'd58: xpb[130] = 1024'd74950733033587219080289186481453792113360261010680708358033886289438707565830375079822768263598992516078785773394284505293158544707769982130969465730822625008636419643565063668328591971803714160985191830385970305826561709455666127583026001982386992849644894855575149546325340735065590706064273678356740432541;
            6'd59: xpb[130] = 1024'd116885525292758896764038648674090482014440095086536892957905250643300771686083892568962580700531661557380486196068192432229285639892096815556469669886703873331890889237796411824937266740952518003500346078484996640080862017449678279547122878292106760589631499333571688375952054082301963430742194029809206564176;
            6'd60: xpb[130] = 1024'd34753621867805833048989183461912739170821502036657393429644759932185940469028271148087321922806656289239037211284606924586348894235203314426809749026254080721454684262456542643915702318584116124705302718196783127970801475222793658546241184918597079062798200397451169175472239355609703138301424554636078211480;
            6'd61: xpb[130] = 1024'd76688414126977510732738645654549429071901336112513578029516124286048004589281788637227134359739325330540737633958514851522475989419530147852309953182135329044709153856687890800524377087732919967220456966295809462225101783216805810510338061228316846802784804875447708005098952702846075862979344906088544343115;
            6'd62: xpb[130] = 1024'd118623206386149188416488107847186118972981170188369762629387488639910068709535306126366946796671994371842438056632422778458603084603856981277810157338016577367963623450919238957133051856881723809735611214394835796479402091210817962474434937538036614542771409353444246834725666050082448587657265257541010474750;
            6'd63: xpb[130] = 1024'd36491302961196124701438642635008376129362577138490263101126997928795237492479684705491688018946989103700989071848837270815666338946963480148150236477566784757527418475579369776111487434513321930940567854106622284369341548983933341473553244164526933015938110417323727634245851323390188295216495782367882122054;
        endcase
    end

    always_comb begin
        case(flag[43][16:12])
            5'd0: xpb[131] = 1024'd0;
            5'd1: xpb[131] = 1024'd78426095220367802385188104827645066030442411214346447700998362282657301612733202194631500455879658145002689494522745197751793434131290313573650440633448033080781888069810717932720162203662125773455722102205648618623641856977945493437650120474246700755924714895320266463872564670626561019894416133820348253689;
            5'd2: xpb[131] = 1024'd32785494756610863371577282250475699316186395302957211273864869500337707888157265479247929697101641980562229581587996960924523027421360292592140756250565025227873101570050218527810085215807045825601246596024057390882922863734994213910321671265263952245029526376523474897638601267324489022670142441015102023047;
            5'd3: xpb[131] = 1024'd111211589976978665756765387078120765346628806517303658974863231782995009500890467673879430152981300125564919076110742158676316461552650606165791196884013058308654989639860936460530247419469171599056968698229706009506564720712939707347971791739510653000954241271843741361511165937951050042564558574835450276736;
            5'd4: xpb[131] = 1024'd65570989513221726743154564500951398632372790605914422547729739000675415776314530958495859394203283961124459163175993921849046054842720585184281512501130050455746203140100437055620170431614091651202493192048114781765845727469988427820643342530527904490059052753046949795277202534648978045340284882030204046094;
            5'd5: xpb[131] = 1024'd19930389049464787729543741923782031918116774694525186120596246218355822051738594243112288635425267796683999250241245685021775648132790564202771828118247042602837416640339937650710093443759011703348017685866523554025126734227037148293314893321545155979163864234250158229043239131346906048116011189224957815452;
            5'd6: xpb[131] = 1024'd98356484269832590114731846751427097948559185908871633821594608501013123664471796437743789091304925941686688744763990882773569082264080877776422268751695075683619304710150655583430255647421137476803739788072172172648768591204982641730965013795791856735088579129570424692915803801973467068010427323045306069141;
            5'd7: xpb[131] = 1024'd52715883806075651101121024174257731234303169997482397394461115718693529939895859722360218332526909777246228831829242645946298675554150856794912584368812067830710518210390156178520178659566057528949264281890580944908049597962031362203636564586809108224193390610773633126681840398671395070786153630240059838499;
            5'd8: xpb[131] = 1024'd7075283342318712087510201597088364520047154086093160967327622936373936215319923006976647573748893612805768918894494409119028268844220835813402899985929059977801731710629656773610101671710977581094788775708989717167330604719080082676308115377826359713298202091976841560447876995369323073561879937434813607857;
            5'd9: xpb[131] = 1024'd85501378562686514472698306424733430550489565300439608668325985219031237828053125201608148029628551757808458413417239606870821702975511149387053340619377093058583619780440374706330263875373103354550510877914638335790972461697025576113958235852073060469222916987297108024320441665995884093456296071255161861546;
            5'd10: xpb[131] = 1024'd39860778098929575459087483847564063836233549389050372241192492436711644103477188486224577270850535593367998500482491370043551296265581128405543656236494085205674833280679875301420186887518023406696035371733047108050253468454074296586629786643090311958327728468500316458086478262693812096232022378449915630904;
            5'd11: xpb[131] = 1024'd118286873319297377844275588675209129866675960603396819942190854719368945716210390680856077726730193738370687995005236567795344730396871441979194096869942118286456721350490593234140349091180149180151757473938695726673895325432019790024279907117337012714252443363820582921959042933320373116126438512270263884593;
            5'd12: xpb[131] = 1024'd72646272855540438830664766098039763152419944692007583515057361937049351991634453965472506967952177573930228082070488330968074323686941420997684412487059110433547934850730093829230272103325069232297281967757104498933176332189068510496951457908354264203357254845023791355725079530018301118902164819465017653951;
            5'd13: xpb[131] = 1024'd27005672391783499817053943520870396438163928780618347087923869154729758267058517250088936209174161409489768169135740094140803916977011400016174728104176102580639148350969594424320195115469989284442806461575513271192457338946117230969623008699371515692462066326226999789491116126716229121677891126659771423309;
            5'd14: xpb[131] = 1024'd105431767612151302202242048348515462468606339994964794788922231437387059879791719444720436665053819554492457663658485291892597351108301713589825168737624135661421036420780312357040357319132115057898528563781161889816099195924062724407273129173618216448386781221547266253363680797342790141572307260480119676998;
            5'd15: xpb[131] = 1024'd59791167148394363188631225771346095754350324083575558361788738655067466155215782729336865906275803390051997750723737055065326944398371692608315484354741127808512249921019812952130280331277035110044053057599570662075380202681111444879944679964635467937491592702750474687129717394040718144348033567674873446356;
            5'd16: xpb[131] = 1024'd14150566684637424175020403194176729040094308172186321934655245872747872430639846013953295147497787225611537837788988818238056537688441671626805799971858119955603463421259313547220203343421955162189577551417979434334661209438160165352616230755652719426596404183953683120895753990738646147123759874869627215714;
            5'd17: xpb[131] = 1024'd92576661905005226560208508021821795070536719386532769635653608155405174043373048208584795603377445370614227332311734015989849971819731985200456240605306153036385351491070031479940365547084080935645299653623628052958303066416105658790266351229899420182521119079273949584768318661365207167018176008689975469403;
            5'd18: xpb[131] = 1024'd46936061441248287546597685444652428356280703475143533208520115373085580318797111493201224844599429206173767419376985779162579565109801964218946556222423145183476564991309532075030288559229000987790824147442036825217584073173154379262937902020916671671625930560477158018534355258063135169793902315884729238761;
            5'd19: xpb[131] = 1024'd1295460977491348532986862867483061642024687563754296781386622590765986594221174777817654085821413041733307506442237542335309158399871943237436871839540137330567778491549032670120211571373921039936348641260445597476865079930203099735609452811933923160730742041680366452300391854761063172569628623079483008119;
            5'd20: xpb[131] = 1024'd79721556197859150918174967695128127672467098778100744482384984873423288206954376972449154541701071186735997000964982740087102592531162256811087312472988170411349666561359750602840373775036046813392070743466094216100506936908148593173259573286180623916655456937000632916172956525387624192464044756899831261808;
            5'd21: xpb[131] = 1024'd34080955734102211904564145117958760958211082866711508055251492091103694482378440257065583782923055022295537088030234503259832185821232235829577628090105162558440880061599251197930296787180966865537595237284502988359787943665197313645931124077197875405760268418203841349938993122085552195239771064094585031166;
            5'd22: xpb[131] = 1024'd112507050954470014289752249945603826988653494081057955756249854373760996095111642451697084238802713167298226582552979701011625619952522549403228068723553195639222768131409969130650458990843092638993317339490151606983429800643142807083581244551444576161684983313524107813811557792712113215134187197914933284855;
            5'd23: xpb[131] = 1024'd66866450490713075276141427368434460274397478169668719329116361591441402370535705736313513480024697002857766669618231464184355213242592528421718384340670187786313981631649469725740382002988012691138841833308560379242710807400191527556252795342461827650789794794727316247577594389410041217909913505109687054213;
            5'd24: xpb[131] = 1024'd21225850026956136262530604791265093560141462258279482901982868809121808645959769020929942721246680838417306756683483227357084806532662507440208699957787179933405195131888970320830305015132932743284366327126969151501991814157240248028924346133479079139894606275930524681343630986107969220685639812304440823571;
            5'd25: xpb[131] = 1024'd99651945247323938647718709618910159590583873472625930602981231091779110258692971215561443177126338983419996251206228425108878240663952821013859140591235213014187083201699688253550467218795058516740088429332617770125633671135185741466574466607725779895819321171250791145216195656734530240580055946124789077260;
            5'd26: xpb[131] = 1024'd54011344783566999634107887041740792876327857561236694175847738309459516534117034500177872418348322818979536338271480188281607833954022800032349456208352205161278296701939188848640390230939978568885612923151026542384914677892234461939246017398743031384924132652453999578982232253432458243355782253319542846618;
            5'd27: xpb[131] = 1024'd8370744319810060620497064464571426162071841649847457748714245527139922809541097784794301659570306654539076425336731951454337427244092779050839771825469197308369510202178689443730313243084898621031137416969435314644195684649283182411917568189760282874028944133657208012748268850130386246131508560514296615976;
            5'd28: xpb[131] = 1024'd86796839540177863005685169292216492192514252864193905449712607809797224422274299979425802115449964799541765919859477149206130861375383092624490212458917230389151398271989407376450475446747024394486859519175083933267837541627228675849567688664006983629953659028977474476620833520756947266025924694334644869665;
            5'd29: xpb[131] = 1024'd41156239076420923992074346715047125478258236952804669022579115027477630697698363264042231356671948635101306006924728912378860454665453071642980528076034222536242611772228907971540398458891944446632384012993492705527118548384277396322239239455024235119058470510180682910386870117454875268801651001529398639023;
            5'd30: xpb[131] = 1024'd119582334296788726377262451542692191508700648167151116723577477310134932310431565458673731812551606780103995501447474110130653888796743385216630968709482255617024499842039625904260560662554070220088106115199141324150760405362222889759889359929270935874983185405500949374259434788081436288696067135349746892712;
            5'd31: xpb[131] = 1024'd73941733833031787363651628965522824794444632255761880296443984527815338585855628743290161053773590615663535588512725873303383482086813364235121284326599247764115713342279126499350483674698990272233630609017550096410041412119271610232560910720288187364087996886704157808025471384779364291471793442544500662070;
        endcase
    end

    always_comb begin
        case(flag[44][5:0])
            6'd0: xpb[132] = 1024'd0;
            6'd1: xpb[132] = 1024'd14150566684637424175020403194176729040094308172186321934655245872747872430639846013953295147497787225611537837788988818238056537688441671626805799971858119955603463421259313547220203343421955162189577551417979434334661209438160165352616230755652719426596404183953683120895753990738646147123759874869627215714;
            6'd2: xpb[132] = 1024'd28301133369274848350040806388353458080188616344372643869310491745495744861279692027906590294995574451223075675577977636476113075376883343253611599943716239911206926842518627094440406686843910324379155102835958868669322418876320330705232461511305438853192808367907366241791507981477292294247519749739254431428;
            6'd3: xpb[132] = 1024'd42451700053912272525061209582530187120282924516558965803965737618243617291919538041859885442493361676834613513366966454714169613065325014880417399915574359866810390263777940641660610030265865486568732654253938303003983628314480496057848692266958158279789212551861049362687261972215938441371279624608881647142;
            6'd4: xpb[132] = 1024'd56602266738549696700081612776706916160377232688745287738620983490991489722559384055813180589991148902446151351155955272952226150753766686507223199887432479822413853685037254188880813373687820648758310205671917737338644837752640661410464923022610877706385616735814732483583015962954584588495039499478508862856;
            6'd5: xpb[132] = 1024'd70752833423187120875102015970883645200471540860931609673276229363739362153199230069766475737488936128057689188944944091190282688442208358134028999859290599778017317106296567736101016717109775810947887757089897171673306047190800826763081153778263597132982020919768415604478769953693230735618799374348136078570;
            6'd6: xpb[132] = 1024'd84903400107824545050122419165060374240565849033117931607931475236487234583839076083719770884986723353669227026733932909428339226130650029760834799831148719733620780527555881283321220060531730973137465308507876606007967256628960992115697384533916316559578425103722098725374523944431876882742559249217763294284;
            6'd7: xpb[132] = 1024'd99053966792461969225142822359237103280660157205304253542586721109235107014478922097673066032484510579280764864522921727666395763819091701387640599803006839689224243948815194830541423403953686135327042859925856040342628466067121157468313615289569035986174829287675781846270277935170523029866319124087390509998;
            6'd8: xpb[132] = 1024'd113204533477099393400163225553413832320754465377490575477241966981982979445118768111626361179982297804892302702311910545904452301507533373014446399774864959644827707370074508377761626747375641297516620411343835474677289675505281322820929846045221755412771233471629464967166031925909169176990078998957017725712;
            6'd9: xpb[132] = 1024'd3288404477612076176384701342776128616150346423941213283765357789753956538449475215564585112822410721060691132643405929563444998354754710086092074730392038666740496221762604587351590899280390738396000354374575062647590034722544715208567507117645025572547734241466090057955257842719182306995149047201050457095;
            6'd10: xpb[132] = 1024'd17438971162249500351405104536952857656244654596127535218420603662501828969089321229517880260320197946672228970432394747801501536043196381712897874702250158622343959643021918134571794242702345900585577905792554496982251244160704880561183737873297744999144138425419773178851011833457828454118908922070677672809;
            6'd11: xpb[132] = 1024'd31589537846886924526425507731129586696338962768313857153075849535249701399729167243471175407817985172283766808221383566039558073731638053339703674674108278577947423064281231681791997586124301062775155457210533931316912453598865045913799968628950464425740542609373456299746765824196474601242668796940304888523;
            6'd12: xpb[132] = 1024'd45740104531524348701445910925306315736433270940500179087731095407997573830369013257424470555315772397895304646010372384277614611420079724966509474645966398533550886485540545229012200929546256224964733008628513365651573663037025211266416199384603183852336946793327139420642519814935120748366428671809932104237;
            6'd13: xpb[132] = 1024'd59890671216161772876466314119483044776527579112686501022386341280745446261008859271377765702813559623506842483799361202515671149108521396593315274617824518489154349906799858776232404272968211387154310560046492799986234872475185376619032430140255903278933350977280822541538273805673766895490188546679559319951;
            6'd14: xpb[132] = 1024'd74041237900799197051486717313659773816621887284872822957041587153493318691648705285331060850311346849118380321588350020753727686796963068220121074589682638444757813328059172323452607616390166549343888111464472234320896081913345541971648660895908622705529755161234505662434027796412413042613948421549186535665;
            6'd15: xpb[132] = 1024'd88191804585436621226507120507836502856716195457059144891696833026241191122288551299284355997809134074729918159377338838991784224485404739846926874561540758400361276749318485870672810959812121711533465662882451668655557291351505707324264891651561342132126159345188188783329781787151059189737708296418813751379;
            6'd16: xpb[132] = 1024'd102342371270074045401527523702013231896810503629245466826352078898989063552928397313237651145306921300341455997166327657229840762173846411473732674533398878355964740170577799417893014303234076873723043214300431102990218500789665872676881122407214061558722563529141871904225535777889705336861468171288440967093;
            6'd17: xpb[132] = 1024'd116492937954711469576547926896189960936904811801431788761007324771736935983568243327190946292804708525952993834955316475467897299862288083100538474505256998311568203591837112965113217646656032035912620765718410537324879710227826038029497353162866780985318967713095555025121289768628351483985228046158068182807;
            6'd18: xpb[132] = 1024'd6576808955224152352769402685552257232300692847882426567530715579507913076898950431129170225644821442121382265286811859126889996709509420172184149460784077333480992443525209174703181798560781476792000708749150125295180069445089430417135014235290051145095468482932180115910515685438364613990298094402100914190;
            6'd19: xpb[132] = 1024'd20727375639861576527789805879728986272395001020068748502185961452255785507538796445082465373142608667732920103075800677364946534397951091798989949432642197289084455864784522721923385141982736638981578260167129559629841278883249595769751244990942770571691872666885863236806269676177010761114057969271728129904;
            6'd20: xpb[132] = 1024'd34877942324499000702810209073905715312489309192255070436841207325003657938178642459035760520640395893344457940864789495603003072086392763425795749404500317244687919286043836269143588485404691801171155811585108993964502488321409761122367475746595489998288276850839546357702023666915656908237817844141355345618;
            6'd21: xpb[132] = 1024'd49028509009136424877830612268082444352583617364441392371496453197751530368818488472989055668138183118955995778653778313841059609774834435052601549376358437200291382707303149816363791828826646963360733363003088428299163697759569926474983706502248209424884681034793229478597777657654303055361577719010982561332;
            6'd22: xpb[132] = 1024'd63179075693773849052851015462259173392677925536627714306151699070499402799458334486942350815635970344567533616442767132079116147463276106679407349348216557155894846128562463363583995172248602125550310914421067862633824907197730091827599937257900928851481085218746912599493531648392949202485337593880609777046;
            6'd23: xpb[132] = 1024'd77329642378411273227871418656435902432772233708814036240806944943247275230098180500895645963133757570179071454231755950317172685151717778306213149320074677111498309549821776910804198515670557287739888465839047296968486116635890257180216168013553648278077489402700595720389285639131595349609097468750236992760;
            6'd24: xpb[132] = 1024'd91480209063048697402891821850612631472866541881000358175462190815995147660738026514848941110631544795790609292020744768555229222840159449933018949291932797067101772971081090458024401859092512449929466017257026731303147326074050422532832398769206367704673893586654278841285039629870241496732857343619864208474;
            6'd25: xpb[132] = 1024'd105630775747686121577912225044789360512960850053186680110117436688743020091377872528802236258129332021402147129809733586793285760528601121559824749263790917022705236392340404005244605202514467612119043568675006165637808535512210587885448629524859087131270297770607961962180793620608887643856617218489491424188;
            6'd26: xpb[132] = 1024'd119781342432323545752932628238966089553055158225373002044772682561490892522017718542755531405627119247013684967598722405031342298217042793186630549235649036978308699813599717552464808545936422774308621120092985599972469744950370753238064860280511806557866701954561645083076547611347533790980377093359118639902;
            6'd27: xpb[132] = 1024'd9865213432836228529154104028328385848451039271823639851296073369261869615348425646693755338467232163182073397930217788690334995064264130258276224191176116000221488665287813762054772697841172215188001063123725187942770104167634145625702521352935076717643202724398270173865773528157546920985447141603151371285;
            6'd28: xpb[132] = 1024'd24015780117473652704174507222505114888545347444009961785951319242009742045988271660647050485965019388793611235719206606928391532752705801885082024163034235955824952086547127309274976041263127377377578614541704622277431313605794310978318752108587796144239606908351953294761527518896193068109207016472778586999;
            6'd29: xpb[132] = 1024'd38166346802111076879194910416681843928639655616196283720606565114757614476628117674600345633462806614405149073508195425166448070441147473511887824134892355911428415507806440856495179384685082539567156165959684056612092523043954476330934982864240515570836011092305636415657281509634839215232966891342405802713;
            6'd30: xpb[132] = 1024'd52316913486748501054215313610858572968733963788382605655261810987505486907267963688553640780960593840016686911297184243404504608129589145138693624106750475867031878929065754403715382728107037701756733717377663490946753732482114641683551213619893234997432415276259319536553035500373485362356726766212033018427;
            6'd31: xpb[132] = 1024'd66467480171385925229235716805035302008828271960568927589917056860253359337907809702506935928458381065628224749086173061642561145818030816765499424078608595822635342350325067950935586071528992863946311268795642925281414941920274807036167444375545954424028819460213002657448789491112131509480486641081660234141;
            6'd32: xpb[132] = 1024'd80618046856023349404256119999212031048922580132755249524572302733001231768547655716460231075956168291239762586875161879880617683506472488392305224050466715778238805771584381498155789414950948026135888820213622359616076151358434972388783675131198673850625223644166685778344543481850777656604246515951287449855;
            6'd33: xpb[132] = 1024'd94768613540660773579276523193388760089016888304941571459227548605749104199187501730413526223453955516851300424664150698118674221194914160019111024022324835733842269192843695045375992758372903188325466371631601793950737360796595137741399905886851393277221627828120368899240297472589423803728006390820914665569;
            6'd34: xpb[132] = 1024'd108919180225298197754296926387565489129111196477127893393882794478496976629827347744366821370951742742462838262453139516356730758883355831645916823994182955689445732614103008592596196101794858350515043923049581228285398570234755303094016136642504112703818032012074052020136051463328069950851766265690541881283;
            6'd35: xpb[132] = 1024'd123069746909935621929317329581742218169205504649314215328538040351244849060467193758320116518449529968074376100242128334594787296571797503272722623966041075645049196035362322139816399445216813512704621474467560662620059779672915468446632367398156832130414436196027735141031805454066716097975526140560169096997;
            6'd36: xpb[132] = 1024'd13153617910448304705538805371104514464601385695764853135061431159015826153797900862258340451289642884242764530573623718253779993419018840344368298921568154666961984887050418349406363597121562953584001417498300250590360138890178860834270028470580102290190936965864360231821031370876729227980596188804201828380;
            6'd37: xpb[132] = 1024'd27304184595085728880559208565281243504695693867951175069716677031763698584437746876211635598787430109854302368362612536491836531107460511971174098893426274622565448308309731896626566940543518115773578968916279684925021348328339026186886259226232821716787341149818043352716785361615375375104356063673829044094;
            6'd38: xpb[132] = 1024'd41454751279723153055579611759457972544790002040137497004371922904511571015077592890164930746285217335465840206151601354729893068795902183597979898865284394578168911729569045443846770283965473277963156520334259119259682557766499191539502489981885541143383745333771726473612539352354021522228115938543456259808;
            6'd39: xpb[132] = 1024'd55605317964360577230600014953634701584884310212323818939027168777259443445717438904118225893783004561077378043940590172967949606484343855224785698837142514533772375150828358991066973627387428440152734071752238553594343767204659356892118720737538260569980149517725409594508293343092667669351875813413083475522;
            6'd40: xpb[132] = 1024'd69755884648998001405620418147811430624978618384510140873682414650007315876357284918071521041280791786688915881729578991206006144172785526851591498809000634489375838572087672538287176970809383602342311623170217987929004976642819522244734951493190979996576553701679092715404047333831313816475635688282710691236;
            6'd41: xpb[132] = 1024'd83906451333635425580640821341988159665072926556696462808337660522755188306997130932024816188778579012300453719518567809444062681861227198478397298780858754444979301993346986085507380314231338764531889174588197422263666186080979687597351182248843699423172957885632775836299801324569959963599395563152337906950;
            6'd42: xpb[132] = 1024'd98057018018272849755661224536164888705167234728882784742992906395503060737636976945978111336276366237911991557307556627682119219549668870105203098752716874400582765414606299632727583657653293926721466726006176856598327395519139852949967413004496418849769362069586458957195555315308606110723155438021965122664;
            6'd43: xpb[132] = 1024'd112207584702910273930681627730341617745261542901069106677648152268250933168276822959931406483774153463523529395096545445920175757238110541732008898724574994356186228835865613179947787001075249088911044277424156290932988604957300018302583643760149138276365766253540142078091309306047252257846915312891592338378;
            6'd44: xpb[132] = 1024'd2291455703422956706903103519703914040657423947519744484171543076021910261607530063869630416614266379691917825428040829579168454085331878803654573680102073378099017687553709389537751152979998529790424220454895878903288964174563410690221304832572408436142267023376767168880535222857265387851985361135625069761;
            6'd45: xpb[132] = 1024'd16442022388060380881923506713880643080751732119706066418826788948769782692247376077822925564112053605303455663217029647817224991773773550430460373651960193333702481108813022936757954496401953691980001771872875313237950173612723576042837535588225127862738671207330450289776289213595911534975745236005252285475;
            6'd46: xpb[132] = 1024'd30592589072697805056943909908057372120846040291892388353482034821517655122887222091776220711609840830914993501006018466055281529462215222057266173623818313289305944530072336483978157839823908854169579323290854747572611383050883741395453766343877847289335075391284133410672043204334557682099505110874879501189;
            6'd47: xpb[132] = 1024'd44743155757335229231964313102234101160940348464078710288137280694265527553527068105729515859107628056526531338795007284293338067150656893684071973595676433244909407951331650031198361183245864016359156874708834181907272592489043906748069997099530566715931479575237816531567797195073203829223264985744506716903;
            6'd48: xpb[132] = 1024'd58893722441972653406984716296410830201034656636265032222792526567013399984166914119682811006605415282138069176583996102531394604839098565310877773567534553200512871372590963578418564526667819178548734426126813616241933801927204072100686227855183286142527883759191499652463551185811849976347024860614133932617;
            6'd49: xpb[132] = 1024'd73044289126610077582005119490587559241128964808451354157447772439761272414806760133636106154103202507749607014372984920769451142527540236937683573539392673156116334793850277125638767870089774340738311977544793050576595011365364237453302458610836005569124287943145182773359305176550496123470784735483761148331;
            6'd50: xpb[132] = 1024'd87194855811247501757025522684764288281223272980637676092103018312509144845446606147589401301600989733361144852161973739007507680215981908564489373511250793111719798215109590672858971213511729502927889528962772484911256220803524402805918689366488724995720692127098865894255059167289142270594544610353388364045;
            6'd51: xpb[132] = 1024'd101345422495884925932045925878941017321317581152823998026758264185257017276086452161542696449098776958972682689950962557245564217904423580191295173483108913067323261636368904220079174556933684665117467080380751919245917430241684568158534920122141444422317096311052549015150813158027788417718304485223015579759;
            6'd52: xpb[132] = 1024'd115495989180522350107066329073117746361411889325010319961413510058004889706726298175495991596596564184584220527739951375483620755592865251818100973454967033022926725057628217767299377900355639827307044631798731353580578639679844733511151150877794163848913500495006232136046567148766434564842064360092642795473;
            6'd53: xpb[132] = 1024'd5579860181035032883287804862480042656807770371460957767936900865775866800057005279434215529436677100752608958071446759142613452440086588889746648410494112044839513909316313976889342052260389268186424574829470941550878998897108125898788811950217434008690001264842857226835793065576447694847134408336675526856;
            6'd54: xpb[132] = 1024'd19730426865672457058308208056656771696902078543647279702592146738523739230696851293387510676934464326364146795860435577380669990128528260516552448382352232000442977330575627524109545395682344430376002126247450375885540208335268291251405042705870153435286405448796540347731547056315093841970894283206302742570;
            6'd55: xpb[132] = 1024'd33880993550309881233328611250833500736996386715833601637247392611271611661336697307340805824432251551975684633649424395618726527816969932143358248354210351956046440751834941071329748739104299592565579677665429810220201417773428456604021273461522872861882809632750223468627301047053739989094654158075929958284;
            6'd56: xpb[132] = 1024'd48031560234947305408349014445010229777090694888019923571902638484019484091976543321294100971930038777587222471438413213856783065505411603770164048326068471911649904173094254618549952082526254754755157229083409244554862627211588621956637504217175592288479213816703906589523055037792386136218414032945557173998;
            6'd57: xpb[132] = 1024'd62182126919584729583369417639186958817185003060206245506557884356767356522616389335247396119427826003198760309227402032094839603193853275396969848297926591867253367594353568165770155425948209916944734780501388678889523836649748787309253734972828311715075618000657589710418809028531032283342173907815184389712;
            6'd58: xpb[132] = 1024'd76332693604222153758389820833363687857279311232392567441213130229515228953256235349200691266925613228810298147016390850332896140882294947023775648269784711822856831015612881712990358769370165079134312331919368113224185046087908952661869965728481031141672022184611272831314563019269678430465933782684811605426;
            6'd59: xpb[132] = 1024'd90483260288859577933410224027540416897373619404578889375868376102263101383896081363153986414423400454421835984805379668570952678570736618650581448241642831778460294436872195260210562112792120241323889883337347547558846255526069118014486196484133750568268426368564955952210317010008324577589693657554438821140;
            6'd60: xpb[132] = 1024'd104633826973497002108430627221717145937467927576765211310523621975010973814535927377107281561921187680033373822594368486809009216259178290277387248213500951734063757858131508807430765456214075403513467434755326981893507464964229283367102427239786469994864830552518639073106071000746970724713453532424066036854;
            6'd61: xpb[132] = 1024'd118784393658134426283451030415893874977562235748951533245178867847758846245175773391060576709418974905644911660383357305047065753947619961904193048185359071689667221279390822354650968799636030565703044986173306416228168674402389448719718657995439189421461234736472322194001824991485616871837213407293693252568;
            6'd62: xpb[132] = 1024'd8868264658647109059672506205256171272958116795402171051702258655529823338506480494998800642259087821813300090714852688706058450794841298975838723140886150711580010131078918564240932951540780006582424929204046004198469033619652841107356319067862459581237735506308947284791050908295630001842283455537725983951;
            6'd63: xpb[132] = 1024'd23018831343284533234692909399432900313052424967588492986357504528277695769146326508952095789756875047424837928503841506944114988483282970602644523112744270667183473552338232111461136294962735168772002480622025438533130243057813006459972549823515179007834139690262630405686804899034276148966043330407353199665;
        endcase
    end

    always_comb begin
        case(flag[44][11:6])
            6'd0: xpb[133] = 1024'd0;
            6'd1: xpb[133] = 1024'd37169398027921957409713312593609629353146733139774814921012750401025568199786172522905390937254662273036375766292830325182171526171724642229450323084602390622786936973597545658681339638384690330961580032040004872867791452495973171812588780579167898434430543874216313526582558889772922296089803205276980415379;
            6'd2: xpb[133] = 1024'd74338796055843914819426625187219258706293466279549629842025500802051136399572345045810781874509324546072751532585660650364343052343449284458900646169204781245573873947195091317362679276769380661923160064080009745735582904991946343625177561158335796868861087748432627053165117779545844592179606410553960830758;
            6'd3: xpb[133] = 1024'd111508194083765872229139937780828888059440199419324444763038251203076704599358517568716172811763986819109127298878490975546514578515173926688350969253807171868360810920792636976044018915154070992884740096120014618603374357487919515437766341737503695303291631622648940579747676669318766888269409615830941246137;
            6'd4: xpb[133] = 1024'd24610896427563088240054322969624084667888505433363575555919146539125377461835551181606492534360974782702353657713827866149622263845678234362641167322078521557457073324818965297095119362021555602536122519772779645106804959762995914285376552633442144470902272082748196076223707485163056167240522994482327177185;
            6'd5: xpb[133] = 1024'd61780294455485045649767635563233714021035238573138390476931896940150945661621723704511883471615637055738729424006658191331793790017402876592091490406680912180244010298416510955776459000406245933497702551812784517974596412258969086097965333212610042905332815956964509602806266374935978463330326199759307592564;
            6'd6: xpb[133] = 1024'd98949692483407003059480948156843343374181971712913205397944647341176513861407896227417274408870299328775105190299488516513965316189127518821541813491283302803030947272014056614457798638790936264459282583852789390842387864754942257910554113791777941339763359831180823129388825264708900759420129405036288007943;
            6'd7: xpb[133] = 1024'd12052394827204219070395333345638539982630277726952336190825542677225186723884929840307594131467287292368331549134825407117073001519631826495832011559554652492127209676040384935508899085658420874110665007505554417345818467030018656758164324687716390507374000291280078625864856080553190038391242783687673938991;
            6'd8: xpb[133] = 1024'd49221792855126176480108645939248169335777010866727151111838293078250754923671102363212985068721949565404707315427655732299244527691356468725282334644157043114914146649637930594190238724043111205072245039545559290213609919525991828570753105266884288941804544165496392152447414970326112334481045988964654354370;
            6'd9: xpb[133] = 1024'd86391190883048133889821958532857798688923744006501966032851043479276323123457274886118376005976611838441083081720486057481416053863081110954732657728759433737701083623235476252871578362427801536033825071585564163081401372021965000383341885846052187376235088039712705679029973860099034630570849194241634769749;
            6'd10: xpb[133] = 1024'd123560588910970091299535271126467428042070477146276780953863793880301891323243447409023766943231274111477458848013316382663587580034805753184182980813361824360488020596833021911552918000812491866995405103625569035949192824517938172195930666425220085810665631913929019205612532749871956926660652399518615185128;
            6'd11: xpb[133] = 1024'd36663291254767307310449656315262624650518783160315911746744689216350564185720481021914086665828262075070685206848653273266695265365310060858473178881633174049584283000859350232604018447679976476646787527278334062452623426793014571043540877321158534978276272374028274702088563565716246205631765778170001116176;
            6'd12: xpb[133] = 1024'd73832689282689264720162968908872254003665516300090726667757439617376132385506653544819477603082924348107060973141483598448866791537034703087923501966235564672371219974456895891285358086064666807608367559318338935320414879288987742856129657900326433412706816248244588228671122455489168501721568983446981531555;
            6'd13: xpb[133] = 1024'd111002087310611222129876281502481883356812249439865541588770190018401700585292826067724868540337586621143436739434313923631038317708759345317373825050837955295158156948054441549966697724449357138569947591358343808188206331784960914668718438479494331847137360122460901755253681345262090797811372188723961946934;
            6'd14: xpb[133] = 1024'd24104789654408438140790666691277079965260555453904672381651085354450373447769859680615188262934574584736663098269650814234146003039263652991664023119109304984254419352080769871017798171316841748221330015011108834691636934060037313516328649375432781014748000582560157251729712161106380076782485567375347877982;
            6'd15: xpb[133] = 1024'd61274187682330395550503979284886709318407288593679487302663835755475941647556032203520579200189236857773038864562481139416317529210988295221114346203711695607041356325678315529699137809701532079182910047051113707559428386556010485328917429954600679449178544456776470778312271050879302372872288772652328293361;
            6'd16: xpb[133] = 1024'd98443585710252352960217291878496338671554021733454302223676586156501509847342204726425970137443899130809414630855311464598489055382712937450564669288314086229828293299275861188380477448086222410144490079091118580427219839051983657141506210533768577883609088330992784304894829940652224668962091977929308708740;
            6'd17: xpb[133] = 1024'd11546288054049568971131677067291535280002327747493433016557481492550182709819238339316289860040887094402640989690648355201596740713217245124854867356585435918924555703302189509431577894953707019795872502743883606930650441327060055989116421429707027051219728791092039801370860756496513947933205356580694639788;
            6'd18: xpb[133] = 1024'd48715686081971526380844989660901164633149060887268247937570231893575750909605410862221680797295549367439016755983478680383768266884941887354305190441187826541711492676899735168112917533338397350757452534783888479798441893823033227801705202008874925485650272665308353327953419646269436244023008561857675055167;
            6'd19: xpb[133] = 1024'd85885084109893483790558302254510793986295794027043062858582982294601319109391583385127071734550211640475392522276309005565939793056666529583755513525790217164498429650497280826794257171723087681719032566823893352666233346319006399614293982588042823920080816539524666854535978536042358540112811767134655470546;
            6'd20: xpb[133] = 1024'd123054482137815441200271614848120423339442527166817877779595732695626887309177755908032462671804873913511768288569139330748111319228391171813205836610392607787285366624094826485475596810107778012680612598863898225534024798814979571426882763167210722354511360413740980381118537425815280836202614972411635885925;
            6'd21: xpb[133] = 1024'd36157184481612657211186000036915619947890833180857008572476628031675560171654789520922782394401861877104994647404476221351219004558895479487496034678663957476381629028121154806526697256975262622331995022516663252037455401090055970274492974063149171522122000873840235877594568241659570115173728351063021816973;
            6'd22: xpb[133] = 1024'd73326582509534614620899312630525249301037566320631823493489378432701128371440962043828173331656524150141370413697306546533390530730620121716946357763266348099168566001718700465208036895359952953293575054556668124905246853586029142087081754642317069956552544748056549404177127131432492411263531556340002232352;
            6'd23: xpb[133] = 1024'd110495980537456572030612625224134878654184299460406638414502128833726696571227134566733564268911186423177746179990136871715562056902344763946396680847868738721955502975316246123889376533744643284255155086596672997773038306082002313899670535221484968390983088622272862930759686021205414707353334761616982647731;
            6'd24: xpb[133] = 1024'd23598682881253788041527010412930075262632605474445769207383024169775369433704168179623883991508174386770972538825473762318669742232849071620686878916140088411051765379342574444940476980612127893906537510249438024276468908357078712747280746117423417558593729082372118427235716837049703986324448140268368578779;
            6'd25: xpb[133] = 1024'd60768080909175745451240323006539704615779338614220584128395774570800937633490340702529274928762836659807348305118304087500841268404573713850137202000742479033838702352940120103621816618996818224868117542289442897144260360853051884559869526696591315993024272956588431953818275726822626282414251345545348994158;
            6'd26: xpb[133] = 1024'd97937478937097702860953635600149333968926071753995399049408524971826505833276513225434665866017498932843724071411134412683012794576298356079587525085344869656625639326537665762303156257381508555829697574329447770012051813349025056372458307275759214427454816830804745480400834616595548578504054550822329409537;
            6'd27: xpb[133] = 1024'd11040181280894918871868020788944530577374377768034529842289420307875178695753546838324985588614486896436950430246471303286120479906802663753877723153616219345721901730563994083354256704248993165481079997982212796515482415624101455220068518171697663595065457290904000976876865432439837857475167929473715340585;
            6'd28: xpb[133] = 1024'd48209579308816876281581333382554159930521110907809344763302170708900746895539719361230376525869149169473326196539301628468292006078527305983328046238218609968508838704161539742035596342633683496442660030022217669383273868120074627032657298750865562029496001165120314503459424322212760153564971134750695755964;
            6'd29: xpb[133] = 1024'd85378977336738833691294645976163789283667844047584159684314921109926315095325891884135767463123811442509701962832131953650463532250251948212778369322821000591295775677759085400716935981018373827404240062062222542251065320616047798845246079330033460463926545039336628030041983211985682449654774340027676171343;
            6'd30: xpb[133] = 1024'd122548375364660791101007958569773418636814577187358974605327671510951883295112064407041158400378473715546077729124962278832635058421976590442228692407423391214082712651356631059398275619403064158365820094102227415118856773112020970657834859909201358898357088913552941556624542101758604745744577545304656586722;
            6'd31: xpb[133] = 1024'd35651077708458007111922343758568615245262883201398105398208566847000556157589098019931478122975461679139304087960299169435742743752480898116518890475694740903178975055382959380449376066270548768017202517754992441622287375387097369505445070805139808065967729373652197053100572917602894024715690923956042517770;
            6'd32: xpb[133] = 1024'd72820475736379964521635656352178244598409616341172920319221317248026124357375270542836869060230123952175679854253129494617914269924205540345969213560297131525965912028980505039130715704655239098978782549794997314490078827883070541318033851384307706500398273247868510579683131807375816320805494129233022933149;
            6'd33: xpb[133] = 1024'd109989873764301921931348968945787873951556349480947735240234067649051692557161443065742259997484786225212055620545959819800085796095930182575419536644899522148752849002578050697812055343039929429940362581835002187357870280379043713130622631963475604934828817122084824106265690697148738616895297334510003348528;
            6'd34: xpb[133] = 1024'd23092576108099137942263354134583070560004655494986866033114962985100365419638476678632579720081774188805281979381296710403193481426434490249709734713170871837849111406604379018863155789907414039591745005487767213861300882654120111978232842859414054102439457582184079602741721512993027895866410713161389279576;
            6'd35: xpb[133] = 1024'd60261974136021095351976666728192699913151388634761680954127713386125933619424649201537970657336436461841657745674127035585365007598159132479160057797773262460636048380201924677544495428292104370553325037527772086729092335150093283790821623438581952536870001456400393129324280402765950191956213918438369694955;
            6'd36: xpb[133] = 1024'd97431372163943052761689979321802329266298121774536495875140463787151501819210821724443361594591098734878033511966957360767536533769883774708610380882375653083422985353799470336225835066676794701514905069567776959596883787646066455603410404017749850971300545330616706655906839292538872488046017123715350110334;
            6'd37: xpb[133] = 1024'd10534074507740268772604364510597525874746427788575626668021359123200174681687855337333681317188086698471259870802294251370644219100388082382900578950647002772519247757825798657276935513544279311166287493220541986100314389921142854451020614913688300138911185790715962152382870108383161767017130502366736041382;
            6'd38: xpb[133] = 1024'd47703472535662226182317677104207155227893160928350441589034109524225742881474027860239072254442748971507635637095124576552815745272112724612350902035249393395306184731423344315958275151928969642127867525260546858968105842417116026263609395492856198573341729664932275678965428998156084063106933707643716456761;
            6'd39: xpb[133] = 1024'd84872870563584183592030989697816784581039894068125256510046859925251311081260200383144463191697411244544011403387954901734987271443837366841801225119851784018093121705020889974639614790313659973089447557300551731835897294913089198076198176072024097007772273539148589205547987887929006359196736912920696872140;
            6'd40: xpb[133] = 1024'd122042268591506141001744302291426413934186627207900071431059610326276879281046372906049854128952073517580387169680785226917158797615562009071251548204454174640880058678618435633320954428698350304051027589340556604703688747409062369888786956651191995442202817413364902732130546777701928655286540118197677287519;
            6'd41: xpb[133] = 1024'd35144970935303357012658687480221610542634933221939202223940505662325552143523406518940173851549061481173613528516122117520266482946066316745541746272725524329976321082644763954372054875565834913702410012993321631207119349684138768736397167547130444609813457873464158228606577593546217934257653496849063218567;
            6'd42: xpb[133] = 1024'd72314368963225314422372000073831239895781666361714017144953256063351120343309579041845564788803723754209989294808952442702438009117790958974992069357327914952763258056242309613053394513950525244663990045033326504074910802180111940548985948126298343044244001747680471755189136483319140230347456702126043633946;
            6'd43: xpb[133] = 1024'd109483766991147271832085312667440869248928399501488832065966006464376688543095751564750955726058386027246365061101782767884609535289515601204442392441930305575550195029839855271734734152335215575625570077073331376942702254676085112361574728705466241478674545621896785281771695373092062526437259907403024049325;
            6'd44: xpb[133] = 1024'd22586469334944487842999697856236065857376705515527962858846901800425361405572785177641275448655373990839591419937119658487717220620019908878732590510201655264646457433866183592785834599202700185276952500726096403446132856951161511209184939601404690646285186081996040778247726188936351805408373286054409980373;
            6'd45: xpb[133] = 1024'd59755867362866445252713010449845695210523438655302777779859652201450929605358957700546666385910036263875967186229949983669888746791744551108182913594804045887433394407463729251467174237587390516238532532766101276313924309447134683021773720180572589080715729956212354304830285078709274101498176491331390395752;
            6'd46: xpb[133] = 1024'd96925265390788402662426323043455324563670171795077592700872402602476497805145130223452057323164698536912342952522780308852060272963469193337633236679406436510220331381061274910148513875972080847200112564806106149181715761943107854834362500759740487515146273830428667831412843968482196397587979696608370811131;
            6'd47: xpb[133] = 1024'd10027967734585618673340708232250521172118477809116723493753297938525170667622163836342377045761686500505569311358117199455167958293973501011923434747677786199316593785087603231199614322839565456851494988458871175685146364218184253681972711655678936682756914290527923327888874784326485676559093075259756742179;
            6'd48: xpb[133] = 1024'd47197365762507576083054020825860150525265210948891538414766048339550738867408336359247767983016348773541945077650947524637339484465698143241373757832280176822103530758685148889880953961224255787813075020498876048552937816714157425494561492234846835117187458164744236854471433674099407972648896280536737157558;
            6'd49: xpb[133] = 1024'd84366763790429533492767333419469779878411944088666353335778798740576307067194508882153158920271011046578320843943777849819511010637422785470824080916882567444890467732282694548562293599608946118774655052538880921420729269210130597307150272814014733551618002038960550381053992563872330268738699485813717572937;
            6'd50: xpb[133] = 1024'd121536161818351490902480646013079409231558677228441168256791549141601875266980681405058549857525673319614696610236608175001682536809147427700274404001484958067677404705880240207243633237993636449736235084578885794288520721706103769119739053393182631986048545913176863907636551453645252564828502691090697988316;
            6'd51: xpb[133] = 1024'd34638864162148706913395031201874605840006983242480299049672444477650548129457715017948869580122661283207922969071945065604790222139651735374564602069756307756773667109906568528294733684861121059387617508231650820791951323981180167967349264289121081153659186373276119404112582269489541843799616069742083919364;
            6'd52: xpb[133] = 1024'd71808262190070664323108343795484235193153716382255113970685194878676116329243887540854260517377323556244298735364775390786961748311376377604014925154358698379560604083504114186976073323245811390349197540271655693659742776477153339779938044868288979588089730247492432930695141159262464139889419275019064334743;
            6'd53: xpb[133] = 1024'd108977660217992621732821656389093864546300449522029928891697945279701684529030060063759651454631985829280674501657605715969133274483101019833465248238961089002347541057101659845657412961630501721310777572311660566527534228973126511592526825447456878022520274121708746457277700049035386435979222480296044750122;
            6'd54: xpb[133] = 1024'd22080362561789837743736041577889061154748755536069059684578840615750357391507093676649971177228973792873900860492942606572240959813605327507755446307232438691443803461127988166708513408497986330962159995964425593030964831248202910440137036343395327190130914581808001953753730864879675714950335858947430681170;
            6'd55: xpb[133] = 1024'd59249760589711795153449354171498690507895488675843874605591591016775925591293266199555362114483636065910276626785772931754412485985329969737205769391834829314230740434725533825389853046882676661923740028004430465898756283744176082252725816922563225624561458456024315480336289754652598011040139064224411096549;
            6'd56: xpb[133] = 1024'd96419158617633752563162666765108319861042221815618689526604341417801493791079438722460753051738298338946652393078603256936584012157054611966656092476437219937017677408323079484071192685267366992885320060044435338766547736240149254065314597501731124058992002330240629006918848644425520307129942269501391511928;
            6'd57: xpb[133] = 1024'd9521860961430968574077051953903516469490527829657820319485236753850166653556472335351072774335286302539878751913940147539691697487558919640946290544708569626113939812349407805122293132134851602536702483697200365269978338515225652912924808397669573226602642790339884503394879460269809586101055648152777442976;
            6'd58: xpb[133] = 1024'd46691258989352925983790364547513145822637260969432635240497987154875734853342644858256463711589948575576254518206770472721863223659283561870396613629310960248900876785946953463803632770519541933498282515737205238137769791011198824725513588976837471661033186664556198029977438350042731882190858853429757858355;
            6'd59: xpb[133] = 1024'd83860657017274883393503677141122775175783994109207450161510737555901303053128817381161854648844610848612630284499600797904034749831008204099846936713913350871687813759544499122484972408904232264459862547777210111005561243507171996538102369556005370095463730538772511556559997239815654178280662058706738273734;
            6'd60: xpb[133] = 1024'd121030055045196840803216989734732404528930727248982265082523487956926871252914989904067245586099273121649006050792431123086206276002732846329297259798515741494474750733142044781166312047288922595421442579817214983873352696003145168350691150135173268529894274412988825083142556129588576474370465263983718689113;
            6'd61: xpb[133] = 1024'd34132757388994056814131374923527601137379033263021395875404383292975544115392023516957565308696261085242232409627768013689313961333237154003587457866787091183571013137168373102217412494156407205072825003469980010376783298278221567198301361031111717697504914873088080579618586945432865753341578642635104620161;
            6'd62: xpb[133] = 1024'd71302155416916014223844687517137230490525766402796210796417133694001112315178196039862956245950923358278608175920598338871485487504961796233037780951389481806357950110765918760898752132541097536034405035509984883244574750774194739010890141610279616131935458747304394106201145835205788049431381847912085035540;
            6'd63: xpb[133] = 1024'd108471553444837971633558000110746859843672499542571025717429884095026680514964368562768347183205585631314983942213428664053657013676686438462488104035991872429144887084363464419580091770925787866995985067549989756112366203270167910823478922189447514566366002621520707632783704724978710345521185053189065450919;
        endcase
    end

    always_comb begin
        case(flag[44][16:12])
            5'd0: xpb[134] = 1024'd0;
            5'd1: xpb[134] = 1024'd21574255788635187644472385299542056452120805556610156510310779431075353377441402175658666905802573594908210301048765554656764699007190746136778302104263222118241149488389792740631192217793272476647367491202754782615796805545244309671089133085385963733976643081619963129259735540822999624492298431840451381967;
            5'd2: xpb[134] = 1024'd43148511577270375288944770599084112904241611113220313020621558862150706754882804351317333811605147189816420602097531109313529398014381492273556604208526444236482298976779585481262384435586544953294734982405509565231593611090488619342178266170771927467953286163239926258519471081645999248984596863680902763934;
            5'd3: xpb[134] = 1024'd64722767365905562933417155898626169356362416669830469530932338293226060132324206526976000717407720784724630903146296663970294097021572238410334906312789666354723448465169378221893576653379817429942102473608264347847390416635732929013267399256157891201929929244859889387779206622468998873476895295521354145901;
            5'd4: xpb[134] = 1024'd86297023154540750577889541198168225808483222226440626041243117724301413509765608702634667623210294379632841204195062218627058796028762984547113208417052888472964597953559170962524768871173089906589469964811019130463187222180977238684356532341543854935906572326479852517038942163291998497969193727361805527868;
            5'd5: xpb[134] = 1024'd107871278943175938222361926497710282260604027783050782551553897155376766887207010878293334529012867974541051505243827773283823495035953730683891510521316110591205747441948963703155961088966362383236837456013773913078984027726221548355445665426929818669883215408099815646298677704114998122461492159202256909835;
            5'd6: xpb[134] = 1024'd5378839047686384468035384392437905968026406213925254933732821521475224927339274143936930220157767260006112398835099893361524353201924142265509687609248291775756222360767539106156914115242429138574007338829288849330419983050569085061556228829086333137039955075602720745451885171009364729835100764417113807471;
            5'd7: xpb[134] = 1024'd26953094836321572112507769691979962420147211770535411444043600952550578304780676319595597125960340854914322699883865448018289052209114888402287989713511513893997371849157331846788106333035701615221374830032043631946216788595813394732645361914472296871016598157222683874711620711832364354327399196257565189438;
            5'd8: xpb[134] = 1024'd48527350624956759756980154991522018872268017327145567954354380383625931682222078495254264031762914449822533000932631002675053751216305634539066291817774736012238521337547124587419298550828974091868742321234798414562013594141057704403734494999858260604993241238842647003971356252655363978819697628098016571405;
            5'd9: xpb[134] = 1024'd70101606413591947401452540291064075324388822883755724464665159814701285059663480670912930937565488044730743301981396557331818450223496380675844593922037958130479670825936917328050490768622246568516109812437553197177810399686302014074823628085244224338969884320462610133231091793478363603311996059938467953372;
            5'd10: xpb[134] = 1024'd91675862202227135045924925590606131776509628440365880974975939245776638437104882846571597843368061639638953603030162111988583149230687126812622896026301180248720820314326710068681682986415519045163477303640307979793607205231546323745912761170630188072946527402082573262490827334301363227804294491778919335339;
            5'd11: xpb[134] = 1024'd113250117990862322690397310890148188228630433996976037485286718676851991814546285022230264749170635234547163904078927666645347848237877872949401198130564402366961969802716502809312875204208791521810844794843062762409404010776790633417001894256016151806923170483702536391750562875124362852296592923619370717306;
            5'd12: xpb[134] = 1024'd10757678095372768936070768784875811936052812427850509867465643042950449854678548287873860440315534520012224797670199786723048706403848284531019375218496583551512444721535078212313828230484858277148014677658577698660839966101138170123112457658172666274079910151205441490903770342018729459670201528834227614942;
            5'd13: xpb[134] = 1024'd32331933884007956580543154084417868388173617984460666377776422474025803232119950463532527346118108114920435098718965341379813405411039030667797677322759805669753594209924870952945020448278130753795382168861332481276636771646382479794201590743558630008056553232825404620163505882841729084162499960674678996909;
            5'd14: xpb[134] = 1024'd53906189672643144225015539383959924840294423541070822888087201905101156609561352639191194251920681709828645399767730896036578104418229776804575979427023027787994743698314663693576212666071403230442749660064087263892433577191626789465290723828944593742033196314445367749423241423664728708654798392515130378876;
            5'd15: xpb[134] = 1024'd75480445461278331869487924683501981292415229097680979398397981336176509987002754814849861157723255304736855700816496450693342803425420522941354281531286249906235893186704456434207404883864675707090117151266842046508230382736871099136379856914330557476009839396065330878682976964487728333147096824355581760843;
            5'd16: xpb[134] = 1024'd97054701249913519513960309983044037744536034654291135908708760767251863364444156990508528063525828899645066001865262005350107502432611269078132583635549472024477042675094249174838597101657948183737484642469596829124027188282115408807468989999716521209986482477685294007942712505310727957639395256196033142810;
            5'd17: xpb[134] = 1024'd118628957038548707158432695282586094196656840210901292419019540198327216741885559166167194969328402494553276302914027560006872201439802015214910885739812694142718192163484041915469789319451220660384852133672351611739823993827359718478558123085102484943963125559305257137202448046133727582131693688036484524777;
            5'd18: xpb[134] = 1024'd16136517143059153404106153177313717904079218641775764801198464564425674782017822431810790660473301780018337196505299680084573059605772426796529062827744875327268667082302617318470742345727287415722022016487866547991259949151707255184668686487258999411119865226808162236355655513028094189505302293251341422413;
            5'd19: xpb[134] = 1024'd37710772931694341048578538476855774356200024198385921311509243995501028159459224607469457566275875374926547497554065234741337758612963172933307364932008097445509816570692410059101934563520559892369389507690621330607056754696951564855757819572644963145096508308428125365615391053851093813997600725091792804380;
            5'd20: xpb[134] = 1024'd59285028720329528693050923776397830808320829754996077821820023426576381536900626783128124472078448969834757798602830789398102457620153919070085667036271319563750966059082202799733126781313832369016756998893376113222853560242195874526846952658030926879073151390048088494875126594674093438489899156932244186347;
            5'd21: xpb[134] = 1024'd80859284508964716337523309075939887260441635311606234332130802857651734914342028958786791377881022564742968099651596344054867156627344665206863969140534541681992115547471995540364318999107104845664124490096130895838650365787440184197936085743416890613049794471668051624134862135497093062982197588772695568314;
            5'd22: xpb[134] = 1024'd102433540297599903981995694375481943712562440868216390842441582288727088291783431134445458283683596159651178400700361898711631855634535411343642271244797763800233265035861788280995511216900377322311491981298885678454447171332684493869025218828802854347026437553288014753394597676320092687474496020613146950281;
            5'd23: xpb[134] = 1024'd124007796086235091626468079675024000164683246424826547352752361719802441669224833310104125189486169754559388701749127453368396554641726157480420573349060985918474414524251581021626703434693649798958859472501640461070243976877928803540114351914188818081003080634907977882654333217143092311966794452453598332248;
            5'd24: xpb[134] = 1024'd21515356190745537872141537569751623872105624855701019734931286085900899709357096575747720880631069040024449595340399573446097412807696569062038750436993167103024889443070156424627656460969716554296029355317155397321679932202276340246224915316345332548159820302410882981807540684037458919340403057668455229884;
            5'd25: xpb[134] = 1024'd43089611979380725516613922869293680324226430412311176245242065516976253086798498751406387786433642634932659896389165128102862111814887315198817052541256389221266038931459949165258848678762989030943396846519910179937476737747520649917314048401731296282136463384030846111067276224860458543832701489508906611851;
            5'd26: xpb[134] = 1024'd64663867768015913161086308168835736776347235968921332755552844948051606464239900927065054692236216229840870197437930682759626810822078061335595354645519611339507188419849741905890040896556261507590764337722664962553273543292764959588403181487117260016113106465650809240327011765683458168324999921349357993818;
            5'd27: xpb[134] = 1024'd86238123556651100805558693468377793228468041525531489265863624379126959841681303102723721598038789824749080498486696237416391509829268807472373656749782833457748337908239534646521233114349533984238131828925419745169070348838009269259492314572503223750089749547270772369586747306506457792817298353189809375785;
            5'd28: xpb[134] = 1024'd107812379345286288450031078767919849680588847082141645776174403810202313219122705278382388503841363419657290799535461792073156208836459553609151958854046055575989487396629327387152425332142806460885499320128174527784867154383253578930581447657889187484066392628890735498846482847329457417309596785030260757752;
            5'd29: xpb[134] = 1024'd5319939449796734695704536662647473388011225513016118158353328176300771259254968544025984194986262705122351693126733912150857067002429965190770135941978236760539962315447902790153378358418873216222669202943689464036303109707601115636692011060045701951223132296393640597999690314223824024683205390245117655388;
            5'd30: xpb[134] = 1024'd26894195238431922340176921962189529840132031069626274668664107607376124636696370719684651100788836300030561994175499466807621766009620711327548438046241458878781111803837695530784570576212145692870036694146444246652099915252845425307781144145431665685199775378013603727259425855046823649175503822085569037355;
            5'd31: xpb[134] = 1024'd48468451027067109984649307261731586292252836626236431178974887038451478014137772895343318006591409894938772295224265021464386465016811457464326740150504680997022261292227488271415762794005418169517404185349199029267896720798089734978870277230817629419176418459633566856519161395869823273667802253926020419322;
        endcase
    end

    always_comb begin
        case(flag[45][5:0])
            6'd0: xpb[135] = 1024'd0;
            6'd1: xpb[135] = 1024'd97054701249913519513960309983044037744536034654291135908708760767251863364444156990508528063525828899645066001865262005350107502432611269078132583635549472024477042675094249174838597101657948183737484642469596829124027188282115408807468989999716521209986482477685294007942712505310727957639395256196033142810;
            6'd2: xpb[135] = 1024'd70042706815702297629121692561273642744373642182846587689285666469526831391579175071001984912393983489846982596273030576121151164024002203601105042254767903115263410780617281012046955011798690646164771676551953811883693526343334044649959410316203593153153061541253529985778896936692822898160100685766471801289;
            6'd3: xpb[135] = 1024'd43030712381491075744283075139503247744211249711402039469862572171801799418714193151495441761262138080048899190680799146892194825615393138124077500873986334206049778886140312849255312921939433108592058710634310794643359864404552680492449830632690665096319640604821765963615081368074917838680806115336910459768;
            6'd4: xpb[135] = 1024'd16018717947279853859444457717732852744048857239957491250439477874076767445849211231988898610130292670250815785088567717663238487206784072647049959493204765296836146991663344686463670832080175571019345744716667777403026202465771316334940250949177737039486219668390001941451265799457012779201511544907349118247;
            6'd5: xpb[135] = 1024'd113073419197193373373404767700776890488584891894248627159148238641328630810293368222497426673656121569895881786953829723013345989639395341725182543128754237321313189666757593861302267933738123754756830387186264606527053390747886725142409240948894258249472702146075295949393978304767740736840906801103382261057;
            6'd6: xpb[135] = 1024'd86061424762982151488566150279006495488422499422804078939725144343603598837428386302990883522524276160097798381361598293784389651230786276248155001747972668412099557772280625698510625843878866217184117421268621589286719728809105360984899661265381330192639281209643531927230162736149835677361612230673820919536;
            6'd7: xpb[135] = 1024'd59049430328770929603727532857236100488260106951359530720302050045878566864563404383484340371392430750299714975769366864555433312822177210771127460367191099502885925877803657535718983754019608679611404455350978572046386066870323996827390081581868402135805860273211767905066347167531930617882317660244259578015;
            6'd8: xpb[135] = 1024'd32037435894559707718888915435465705488097714479914982500878955748153534891698422463977797220260585340501631570177135435326476974413568145294099918986409530593672293983326689372927341664160351142038691489433335554806052404931542632669880501898355474078972439336780003882902531598914025558403023089814698236494;
            6'd9: xpb[135] = 1024'd5025441460348485834050298013695310487935322008470434281455861450428502918833440544471254069128739930703548164584904006097520636004959079817072377605627961684458662088849721210135699574301093604465978523515692537565718742992761268512370922214842546022139018400348239860738716030296120498923728519385136894973;
            6'd10: xpb[135] = 1024'd102080142710262005348010607996739348232471356662761570190164622217680366283277597534979782132654568830348614166450166011447628138437570348895204961241177433708935704763943970384974296675959041788203463165985289366689745931274876677319839912214559067232125500878033533868681428535606848456563123775581170037783;
            6'd11: xpb[135] = 1024'd75068148276050783463171990574968953232308964191317021970741527919955334310412615615473238981522723420550530760857934582218671800028961283418177419860395864799722072869467002222182654586099784250630750200067646349449412269336095313162330332531046139175292079941601769846517612966988943397083829205151608696262;
            6'd12: xpb[135] = 1024'd48056153841839561578333373153198558232146571719872473751318433622230302337547633695966695830390878010752447355265703152989715461620352217941149878479614295890508440974990034059391012496240526713058037234150003332209078607397313949004820752847533211118458659005170005824353797398371038337604534634722047354741;
            6'd13: xpb[135] = 1024'd21044159407628339693494755731428163231984179248427925531895339324505270364682651776460152679259032600954363949673471723760759123211743152464122337098832726981294809080513065896599370406381269175485324268232360314968744945458532584847311173164020283061625238068738241802189981829753133278125240064292486013220;
            6'd14: xpb[135] = 1024'd118098860657541859207455065714472200976520213902719061440604100091757133729126808766968680742784861500599429951538733729110866625644354421542254920734382199005771851755607315071437967508039217359222808910701957144092772133740647993654780163163736804271611720546423535810132694335063861235764635320488519156030;
            6'd15: xpb[135] = 1024'd91086866223330637322616448292701805976357821431274513221181005794032101756261826847462137591653016090801346545946502299881910287235745356065227379353600630096558219861130346908646325418179959821650095944784314126852438471801866629497270583480223876214778299609991771787968878766445956176285340750058957814509;
            6'd16: xpb[135] = 1024'd64074871789119415437777830870931410976195428959829965001757911496307069783396844927955594440521170681003263140354270870652953948827136290588199837972819061187344587966653378745854683328320702284077382978866671109612104809863085265339761003796710948157944878673560007765805063197828051116806046179629396472988;
            6'd17: xpb[135] = 1024'd37062877354908193552939213449161015976033036488385416782334817198582037810531863008449051289389325271205179734762039441423997610418527225111172296592037492278130956072176410583063041238461444746504670012949028092371771147924303901182251424113198020101111457737128243743641247629210146057326751609199835131467;
            6'd18: xpb[135] = 1024'd10050882920696971668100596027390620975870644016940868562911722900857005837666881088942508138257479861407096329169808012195041272009918159634144755211255923368917324177699442420271399148602187208931957047031385075131437485985522537024741844429685092044278036800696479721477432060592240997847457038770273789946;
            6'd19: xpb[135] = 1024'd107105584170610491182060906010434658720406678671232004471620483668108869202111038079451036201783308761052162331035070017545148774442529428712277338846805395393394366852793691595109996250260135392669441689500981904255464674267637945832210834429401613254264519278381773729420144565902968955486852294966306932756;
            6'd20: xpb[135] = 1024'd80093589736399269297222288588664263720244286199787456252197389370383837229246056159944493050651463351254078925442838588316192436033920363235249797466023826484180734958316723432318354160400877855096728723583338887015131012328856581674701254745888685197431098341950009707256328997285063896007557724536745591235;
            6'd21: xpb[135] = 1024'd53081595302188047412383671166893868720081893728342908032774295072658805256381074240437949899519617941455995519850607159087236097625311297758222256085242257574967103063839755269526712070541620317524015757665695869774797350390075217517191675062375757140597677405518245685092513428667158836528263154107184249714;
            6'd22: xpb[135] = 1024'd26069600867976825527545053745123473719919501256898359813351200774933773283516092320931406748387772531657912114258375729858279759216702232281194714704460688665753471169362787106735069980682362779951302791748052852534463688451293853359682095378862829083764256469086481662928697860049253777048968583677622908193;
            6'd23: xpb[135] = 1024'd123124302117890345041505363728167511464455535911189495722059961542185636647960249311439934811913601431302978116123637735208387261649313501359327298340010160690230513844457036281573667082340310963688787434217649681658490876733409262167151085378579350293750738946771775670871410365359981734688363839873656051003;
            6'd24: xpb[135] = 1024'd96112307683679123156666746306397116464293143439744947502636867244460604675095267391933391660781756021504894710531406305979430923240704435882299756959228591781016881949980068118782024992481053426116074468300006664418157214794627898009641505695066422236917318010340011648707594796742076675209069269444094709482;
            6'd25: xpb[135] = 1024'd69100313249467901271828128884626721464130750968300399283213772946735572702230285472426848509649910611706811304939174876750474584832095370405272215578447022871803250055503099955990382902621795888543361502382363647177823552855846533852131926011553494180083897073908247626543779228124171615729774699014533367961;
            6'd26: xpb[135] = 1024'd42088318815256679386989511462856326463968358496855851063790678649010540729365303552920305358518065201908727899346943447521518246423486304928244674197665453962589618161026131793198740812762538350970648536464720629937489890917065169694622346328040566123250476137476483604379963659506266556250480128584972026440;
            6'd27: xpb[135] = 1024'd15076324381045457502150894041085931463805966025411302844367584351285508756500321633413762207386219792110644493754712018292561908014877239451217132816883885053375986266549163630407098722903280813397935570547077612697156228978283805537112766644527638066417055201044719582216148090888361496771185558155410684919;
            6'd28: xpb[135] = 1024'd112131025630958977016111204024129969208342000679702438753076345118537372120944478623922290270912048691755710495619974023642669410447488508529349716452433357077853028941643412805245695824561228997135420213016674441821183417260399214344581756644244159276403537678730013590158860596199089454410580814351443827729;
            6'd29: xpb[135] = 1024'd85119031196747755131272586602359574208179608208257890533653250820812340148079496704415747119780203281957627090027742594413713072038879443052322175071651788168639397047166444642454053734701971459562707247099031424580849755321617850187072176960731231219570116742298249567995045027581184394931286243921882486208;
            6'd30: xpb[135] = 1024'd58107036762536533246433969180589179208017215736813342314230156523087308175214514784909203968648357872159543684435511165184756733630270377575294633690870219259425765152689476479662411644842713921989994281181388407340516093382836486029562597277218303162736695805866485545831229458963279335451991673492321144687;
            6'd31: xpb[135] = 1024'd31095042328325311361595351758818784207854823265368794094807062225362276202349532865402660817516512462361460278843279735955800395221661312098267092310088650350212133258212508316870769554983456384417281315263745390100182431444055121872053017593705375105903274869434721523667413890345374275972697103062759803166;
            6'd32: xpb[135] = 1024'd4083047894114089476756734337048389207692430793924245875383967927637244229484550945896117666384667052563376873251048306726844056813052246621239550929307081440998501363735540154079127465124198846844568349346102372859848769505273757714543437910192447049069853933002957501503598321727469216493402532633198461645;
            6'd33: xpb[135] = 1024'd101137749144027608990717044320092426952228465448215381784092728694889107593928707936404645729910495952208442875116310312076951559245663515699372134564856553465475544038829789328917724566782147030582052991815699201983875957787389166522012427909908968259056336410688251509446310827038197174132797788829231604455;
            6'd34: xpb[135] = 1024'd74125754709816387105878426898322031952066072976770833564669634397164075621063726016898102578778650542410359469524078882847995220837054450222344593184074984556261912144352821166126082476922889493009340025898056184743542295848607802364502848226396040202222915474256487487282495258420292114653503218399670262934;
            6'd35: xpb[135] = 1024'd47113760275605165221039809476551636951903680505326285345246540099439043648198744097391559427646805132612276063931847453619038882428445384745317051803293415647048280249875853003334440387063631955436627059980413167503208633909826438206993268542883112145389494537824723465118679689802387055174208647970108921413;
            6'd36: xpb[135] = 1024'd20101765841393943336201192054781241951741288033881737125823445801714011675333762177885016276514959722814192658339616024390082544019836319268289510422511846737834648355398884840542798297204374417863914094062770150262874971971045074049483688859370184088556073601392959442954864121184481995694914077540547579892;
            6'd37: xpb[135] = 1024'd117156467091307462850161502037825279696277322688172873034532206568965875039777919168393544340040788622459258660204878029740190046452447588346422094058061318762311691030493134015381395398862322601601398736532366979386902160253160482856952678859086705298542556079078253450897576626495209953334309333736580722702;
            6'd38: xpb[135] = 1024'd90144472657096240965322884616054884696114930216728324815109112271240843066912937248887001188908943212661175254612646600511233708043838522869394552677279749853098059136016165852589753309003065064028685770614723962146568498314379118699443099175573777241709135142646489428733761057877304893855014763307019381181;
            6'd39: xpb[135] = 1024'd63132478222885019080484267194284489695952537745283776595686017973515811094047955329380458037777097802863091849020415171282277369635229457392367011296498180943884427241539197689798111219143807526455972804697080944906234836375597754541933519492060849184875714206214725406569945489259399834375720192877458039660;
            6'd40: xpb[135] = 1024'd36120483788673797195645649772514094695790145273839228376262923675790779121182973409873914886645252393065008443428183742053321031226620391915339469915716612034670795347062229527006469129284549988883259838779437927665901174436816390384423939808547921128042293269782961384406129920641494774896425622447896698139;
            6'd41: xpb[135] = 1024'd9108489354462575310807032350743699695627752802394680156839829378065747148317991490367371735513406983266925037835952312824364692818011326438311928534935043125457163452585261364214827039425292451310546872861794910425567512498035026226914360125034993071208872333351197362242314352023589715417131052018335356618;
            6'd42: xpb[135] = 1024'd106163190604376094824767342333787737440163787456685816065548590145317610512762148480875899799039235882911991039701214318174472195250622595516444512170484515149934206127679510539053424141083240635048031515331391739549594700780150435034383350124751514281195354811036491370185026857334317673056526308214368499428;
            6'd43: xpb[135] = 1024'd79151196170164872939928724912017342440001394985241267846125495847592578539897166561369356647907390473113907634108982888945515856842013530039416970789702946240720574233202542376261782051223983097475318549413748722309261038841369070876873770441238586224361933874604727348021211288716412613577231737784807157907;
            6'd44: xpb[135] = 1024'd52139201735953651055090107490246947439839002513796719626702401549867546567032184641862813496775545063315824228516751459716559518433404464562389429408921377331506942338725574213470139961364725559902605583496105705068927376902587706719364190757725658167528512938172963325857395720098507554097937167355245816386;
            6'd45: xpb[135] = 1024'd25127207301742429170251490068476552439676610042352171407279307252142514594167202722356270345643699653517740822924520030487603180024795399085361888028139808422293310444248606050678497871505468022329892617578462687828593714963806342561854611074212730110695092001741199303693580151480602494618642596925684474865;
            6'd46: xpb[135] = 1024'd122181908551655948684211800051520590184212644696643307315988068019394377958611359712864798409169528553162806824789782035837710682457406668163494471663689280446770353119342855225517094973163416206067377260048059516952620903245921751369323601073929251320681574479426493311636292656791330452258037853121717617675;
            6'd47: xpb[135] = 1024'd95169914117444726799373182629750195184050252225198759096564973721669345985746377793358255258037683143364723419197550606608754344048797602686466930282907711537556721224865887062725452883304158668494664294130416499712287241307140387211814021390416323263848153542994729289472477088173425392778743282692156276154;
            6'd48: xpb[135] = 1024'd68157919683233504914534565207979800183887859753754210877141879423944314012881395873851712106905837733566640013605319177379798005640188537209439388902126142628343089330388918899933810793444901130921951328212773482471953579368359023054304441706903395207014732606562965267308661519555520333299448712262594934633;
            6'd49: xpb[135] = 1024'd41145925249022283029695947786209405183725467282309662657718785126219282040016413954345168955773992323768556608013087748150841667231579471732411847521344573719129457435911950737142168703585643593349238362295130465231619917429577658896794862023390467150181311670131201245144845950937615273820154141833033593112;
            6'd50: xpb[135] = 1024'd14133930814811061144857330364439010183563074810865114438295690828494250067151432034838625804642146913970473202420856318921885328822970406255384306140563004809915825541434982574350526613726386055776525396377487447991286255490796294739285282339877539093347890733699437222981030382319710214340859571403472251591;
            6'd51: xpb[135] = 1024'd111188632064724580658817640347483047928099109465156250347004451595746113431595589025347153868167975813615539204286118324271992831255581675333516889776112476834392868216529231749189123715384334239514010038847084277115313443772911703546754272339594060303334373211384731230923742887630438171980254827599505394401;
            6'd52: xpb[135] = 1024'd84176637630513358773979022925712652927936716993711702127581357298021081458730607105840610717036130403817455798693886895043036492846972609856489348395330907925179236322052263586397481625525076701941297072929441259874979781834130339389244692656081132246500952274952967208759927319012533112500960257169944052880;
            6'd53: xpb[135] = 1024'd57164643196302136889140405503942257927774324522267153908158263000296049485865625186334067565904284994019372393101655465814080154438363544379461807014549339015965604427575295423605839535665819164368584107011798242634646119895348975231735112972568204189667531338521203186596111750394628053021665686740382711359;
            6'd54: xpb[135] = 1024'd30152648762090915004301788082171862927611932050822605688735168702571017513000643266827524414772439584221288987509424036585123816029754478902434265633767770106751972533098327260814197445806561626795871141094155225394312457956567611074225533289055276132834110402089439164432296181776722993542371116310821369838;
            6'd55: xpb[135] = 1024'd3140654327879693119463170660401467927449539579378057469312074404845985540135661347320981263640594174423205581917192607356167477621145413425406724252986201197538340638621359098022555355947304089223158175176512208153978796017786246916715953605542348076000689465657675142268480613158817934063076545881260028317;
            6'd56: xpb[135] = 1024'd100195355577793212633423480643445505671985574233669193378020835172097848904579818337829509327166423074068271583782454612706274980053756682503539307888535673222015383313715608272861152457605252272960642817646109037278005984299901655724184943605258869285987171943342969150211193118469545891702471802077293171127;
            6'd57: xpb[135] = 1024'd73183361143581990748584863221675110671823181762224645158597740874372816931714836418322966176034577664270188178190223183477318641645147617026511766507754104312801751419238640110069510367745994735387929851728466020037672322361120291566675363921745941229153751006911205128047377549851640832223177231647731829606;
            6'd58: xpb[135] = 1024'd46171366709370768863746245799904715671660789290780096939174646576647784958849854498816423024902732254472104772597991754248362303236538551549484225126972535403588119524761671947277868277886737197815216885810823002797338660422338927409165784238233013172320330070479441105883561981233735772743882661218170488085;
            6'd59: xpb[135] = 1024'd19159372275159546978907628378134320671498396819335548719751552278922752985984872579309879873770886844674021367005760325019405964827929486072456683746190966494374487630284703784486226188027479660242503919893179985557004998483557563251656204554720085115486909134047677083719746412615830713264588090788609146564;
            6'd60: xpb[135] = 1024'd116214073525073066492867938361178358416034431473626684628460313046174616350429029569818407937296715744319087368871022330369513467260540755150589267381740438518851530305378952959324823289685427843979988562362776814681032186765672972059125194554436606325473391611732971091662458917926558670903983346984642289374;
            6'd61: xpb[135] = 1024'd89202079090861844608029320939407963415872039002182136409037218748449584377564047650311864786164870334521003963278790901140557128851931689673561726000958869609637898410901984796533181199826170306407275596445133797440698524826891607901615614870923678268639970675301207069498643349308653611424688776555080947853;
            6'd62: xpb[135] = 1024'd62190084656650622723190703517637568415709646530737588189614124450724552404699065730805321635033024924722920557686559471911600790443322624196534184620177300700424266516425016633741539109966912768834562630527490780200364862888110243744106035187410750211806549738869443047334827780690748551945394206125519606332;
            6'd63: xpb[135] = 1024'd35178090222439400838352086095867173415547254059293039970191030152999520431834083811298778483901179514924837152094328042682644452034713558719506643239395731791210634621948048470949897020107655231261849664609847762960031200949328879586596455503897822154973128802437679025171012212072843492466099635695958264811;
        endcase
    end

    always_comb begin
        case(flag[45][11:6])
            6'd0: xpb[136] = 1024'd0;
            6'd1: xpb[136] = 1024'd8166095788228178953513468674096778415384861587848491750767935855274488458969101891792235332769334105126753746502096613453688113626104493242479101858614162881997002727471080308158254930248397693689136698692204745719697539010547515429086875820384894098139707866005915003007196643454938432986805065266396923290;
            6'd2: xpb[136] = 1024'd16332191576456357907026937348193556830769723175696983501535871710548976917938203783584470665538668210253507493004193226907376227252208986484958203717228325763994005454942160616316509860496795387378273397384409491439395078021095030858173751640769788196279415732011830006014393286909876865973610130532793846580;
            6'd3: xpb[136] = 1024'd24498287364684536860540406022290335246154584763545475252303807565823465376907305675376705998308002315380261239506289840361064340878313479727437305575842488645991008182413240924474764790745193081067410096076614237159092617031642546287260627461154682294419123598017745009021589930364815298960415195799190769870;
            6'd4: xpb[136] = 1024'd32664383152912715814053874696387113661539446351393967003071743421097953835876407567168941331077336420507014986008386453814752454504417972969916407434456651527988010909884321232633019720993590774756546794768818982878790156042190061716347503281539576392558831464023660012028786573819753731947220261065587693160;
            6'd5: xpb[136] = 1024'd40830478941140894767567343370483892076924307939242458753839679276372442294845509458961176663846670525633768732510483067268440568130522466212395509293070814409985013637355401540791274651241988468445683493461023728598487695052737577145434379101924470490698539330029575015035983217274692164934025326331984616450;
            6'd6: xpb[136] = 1024'd48996574729369073721080812044580670492309169527090950504607615131646930753814611350753411996616004630760522479012579680722128681756626959454874611151684977291982016364826481848949529581490386162134820192153228474318185234063285092574521254922309364588838247196035490018043179860729630597920830391598381539740;
            6'd7: xpb[136] = 1024'd57162670517597252674594280718677448907694031114939442255375550986921419212783713242545647329385338735887276225514676294175816795382731452697353713010299140173979019092297562157107784511738783855823956890845433220037882773073832608003608130742694258686977955062041405021050376504184569030907635456864778463030;
            6'd8: xpb[136] = 1024'd65328766305825431628107749392774227323078892702787934006143486842195907671752815134337882662154672841014029972016772907629504909008835945939832814868913303055976021819768642465266039441987181549513093589537637965757580312084380123432695006563079152785117662928047320024057573147639507463894440522131175386320;
            6'd9: xpb[136] = 1024'd73494862094053610581621218066871005738463754290636425756911422697470396130721917026130117994924006946140783718518869521083193022634940439182311916727527465937973024547239722773424294372235579243202230288229842711477277851094927638861781882383464046883257370794053235027064769791094445896881245587397572309610;
            6'd10: xpb[136] = 1024'd81660957882281789535134686740967784153848615878484917507679358552744884589691018917922353327693341051267537465020966134536881136261044932424791018586141628819970027274710803081582549302483976936891366986922047457196975390105475154290868758203848940981397078660059150030071966434549384329868050652663969232900;
            6'd11: xpb[136] = 1024'd89827053670509968488648155415064562569233477466333409258447294408019373048660120809714588660462675156394291211523062747990569249887149425667270120444755791701967030002181883389740804232732374630580503685614252202916672929116022669719955634024233835079536786526065065033079163078004322762854855717930366156190;
            6'd12: xpb[136] = 1024'd97993149458738147442161624089161340984618339054181901009215230263293861507629222701506823993232009261521044958025159361444257363513253918909749222303369954583964032729652963697899059162980772324269640384306456948636370468126570185149042509844618729177676494392070980036086359721459261195841660783196763079480;
            6'd13: xpb[136] = 1024'd106159245246966326395675092763258119400003200642030392759983166118568349966598324593299059326001343366647798704527255974897945477139358412152228324161984117465961035457124044006057314093229170017958777082998661694356068007137117700578129385665003623275816202258076895039093556364914199628828465848463160002770;
            6'd14: xpb[136] = 1024'd114325341035194505349188561437354897815388062229878884510751101973842838425567426485091294658770677471774552451029352588351633590765462905394707426020598280347958038184595124314215569023477567711647913781690866440075765546147665216007216261485388517373955910124082810042100753008369138061815270913729556926060;
            6'd15: xpb[136] = 1024'd122491436823422684302702030111451676230772923817727376261519037829117326884536528376883529991540011576901306197531449201805321704391567398637186527879212443229955040912066204622373823953725965405337050480383071185795463085158212731436303137305773411472095617990088725045107949651824076494802075978995953849350;
            6'd16: xpb[136] = 1024'd6590836927526121857416571380734021901459358279840183884155118619414920006196491358660694109651671372584910536576052380679945977176451557324505504721495565178261369069966067592901839692457157377715989570688036085150799773947863473900411443442928856303415422441977582018008618221350381910670191217636756288309;
            6'd17: xpb[136] = 1024'd14756932715754300810930040054830800316844219867688675634923054474689408465165593250452929442421005477711664283078148994133634090802556050566984606580109728060258371797437147901060094622705555071405126269380240830870497312958410989329498319263313750401555130307983497021015814864805320343656996282903153211599;
            6'd18: xpb[136] = 1024'd22923028503982479764443508728927578732229081455537167385690990329963896924134695142245164775190339582838418029580245607587322204428660543809463708438723890942255374524908228209218349552953952765094262968072445576590194851968958504758585195083698644499694838173989412024023011508260258776643801348169550134889;
            6'd19: xpb[136] = 1024'd31089124292210658717956977403024357147613943043385659136458926185238385383103797034037400107959673687965171776082342221041010318054765037051942810297338053824252377252379308517376604483202350458783399666764650322309892390979506020187672070904083538597834546039995327027030208151715197209630606413435947058179;
            6'd20: xpb[136] = 1024'd39255220080438837671470446077121135562998804631234150887226862040512873842072898925829635440729007793091925522584438834494698431680869530294421912155952216706249379979850388825534859413450748152472536365456855068029589929990053535616758946724468432695974253906001242030037404795170135642617411478702343981469;
            6'd21: xpb[136] = 1024'd47421315868667016624983914751217913978383666219082642637994797895787362301042000817621870773498341898218679269086535447948386545306974023536901014014566379588246382707321469133693114343699145846161673064149059813749287469000601051045845822544853326794113961772007157033044601438625074075604216543968740904759;
            6'd22: xpb[136] = 1024'd55587411656895195578497383425314692393768527806931134388762733751061850760011102709414106106267676003345433015588632061402074658933078516779380115873180542470243385434792549441851369273947543539850809762841264559468985008011148566474932698365238220892253669638013072036051798082080012508591021609235137828049;
            6'd23: xpb[136] = 1024'd63753507445123374532010852099411470809153389394779626139530669606336339218980204601206341439037010108472186762090728674855762772559183010021859217731794705352240388162263629750009624204195941233539946461533469305188682547021696081904019574185623114990393377504018987039058994725534950941577826674501534751339;
            6'd24: xpb[136] = 1024'd71919603233351553485524320773508249224538250982628117890298605461610827677949306492998576771806344213598940508592825288309450886185287503264338319590408868234237390889734710058167879134444338927229083160225674050908380086032243597333106450006008009088533085370024902042066191368989889374564631739767931674629;
            6'd25: xpb[136] = 1024'd80085699021579732439037789447605027639923112570476609641066541316885316136918408384790812104575678318725694255094921901763138999811391996506817421449023031116234393617205790366326134064692736620918219858917878796628077625042791112762193325826392903186672793236030817045073388012444827807551436805034328597919;
            6'd26: xpb[136] = 1024'd88251794809807911392551258121701806055307974158325101391834477172159804595887510276583047437345012423852448001597018515216827113437496489749296523307637193998231396344676870674484388994941134314607356557610083542347775164053338628191280201646777797284812501102036732048080584655899766240538241870300725521209;
            6'd27: xpb[136] = 1024'd96417890598036090346064726795798584470692835746173593142602413027434293054856612168375282770114346528979201748099115128670515227063600982991775625166251356880228399072147950982642643925189532008296493256302288288067472703063886143620367077467162691382952208968042647051087781299354704673525046935567122444499;
            6'd28: xpb[136] = 1024'd104583986386264269299578195469895362886077697334022084893370348882708781513825714060167518102883680634105955494601211742124203340689705476234254727024865519762225401799619031290800898855437929701985629954994493033787170242074433659049453953287547585481091916834048562054094977942809643106511852000833519367789;
            6'd29: xpb[136] = 1024'd112750082174492448253091664143992141301462558921870576644138284737983269972794815951959753435653014739232709241103308355577891454315809969476733828883479682644222404527090111598959153785686327395674766653686697779506867781084981174478540829107932479579231624700054477057102174586264581539498657066099916291079;
            6'd30: xpb[136] = 1024'd120916177962720627206605132818088919716847420509719068394906220593257758431763917843751988768422348844359462987605404969031579567941914462719212930742093845526219407254561191907117408715934725089363903352378902525226565320095528689907627704928317373677371332566060392060109371229719519972485462131366313214369;
            6'd31: xpb[136] = 1024'd5015578066824064761319674087371265387533854971831876017542301383555351553423880825529152886534008640043067326650008147906203840726798621406531907584376967474525735412461054877645424454665917061742842442683867424581902008885179432371736011065472818508691137017949249033010039799245825388353577370007115653328;
            6'd32: xpb[136] = 1024'd13181673855052243714833142761468043802918716559680367768310237238829840012392982717321388219303342745169821073152104761359891954352903114649011009442991130356522738139932135185803679384914314755431979141376072170301599547895726947800822886885857712606830844883955164036017236442700763821340382435273512576618;
            6'd33: xpb[136] = 1024'd21347769643280422668346611435564822218303578147528859519078173094104328471362084609113623552072676850296574819654201374813580067979007607891490111301605293238519740867403215493961934315162712449121115840068276916021297086906274463229909762706242606704970552749961079039024433086155702254327187500539909499908;
            6'd34: xpb[136] = 1024'd29513865431508601621860080109661600633688439735377351269846108949378816930331186500905858884842010955423328566156297988267268181605112101133969213160219456120516743594874295802120189245411110142810252538760481661740994625916821978658996638526627500803110260615966994042031629729610640687313992565806306423198;
            6'd35: xpb[136] = 1024'd37679961219736780575373548783758379049073301323225843020614044804653305389300288392698094217611345060550082312658394601720956295231216594376448315018833619002513746322345376110278444175659507836499389237452686407460692164927369494088083514347012394901249968481972909045038826373065579120300797631072703346488;
            6'd36: xpb[136] = 1024'd45846057007964959528887017457855157464458162911074334771381980659927793848269390284490329550380679165676836059160491215174644408857321087618927416877447781884510749049816456418436699105907905530188525936144891153180389703937917009517170390167397288999389676347978824048046023016520517553287602696339100269778;
            6'd37: xpb[136] = 1024'd54012152796193138482400486131951935879843024498922826522149916515202282307238492176282564883150013270803589805662587828628332522483425580861406518736061944766507751777287536726594954036156303223877662634837095898900087242948464524946257265987782183097529384213984739051053219659975455986274407761605497193068;
            6'd38: xpb[136] = 1024'd62178248584421317435913954806048714295227886086771318272917852370476770766207594068074800215919347375930343552164684442082020636109530074103885620594676107648504754504758617034753208966404700917566799333529300644619784781959012040375344141808167077195669092079990654054060416303430394419261212826871894116358;
            6'd39: xpb[136] = 1024'd70344344372649496389427423480145492710612747674619810023685788225751259225176695959867035548688681481057097298666781055535708749735634567346364722453290270530501757232229697342911463896653098611255936032221505390339482320969559555804431017628551971293808799945996569057067612946885332852248017892138291039648;
            6'd40: xpb[136] = 1024'd78510440160877675342940892154242271125997609262468301774453724081025747684145797851659270881458015586183851045168877668989396863361739060588843824311904433412498759959700777651069718826901496304945072730913710136059179859980107071233517893448936865391948507812002484060074809590340271285234822957404687962938;
            6'd41: xpb[136] = 1024'd86676535949105854296454360828339049541382470850316793525221659936300236143114899743451506214227349691310604791670974282443084976987843553831322926170518596294495762687171857959227973757149893998634209429605914881778877398990654586662604769269321759490088215678008399063082006233795209718221628022671084886228;
            6'd42: xpb[136] = 1024'd94842631737334033249967829502435827956767332438165285275989595791574724602084001635243741546996683796437358538173070895896773090613948047073802028029132759176492765414642938267386228687398291692323346128298119627498574938001202102091691645089706653588227923544014314066089202877250148151208433087937481809518;
            6'd43: xpb[136] = 1024'd103008727525562212203481298176532606372152194026013777026757531646849213061053103527035976879766017901564112284675167509350461204240052540316281129887746922058489768142114018575544483617646689386012482826990324373218272477011749617520778520910091547686367631410020229069096399520705086584195238153203878732808;
            6'd44: xpb[136] = 1024'd111174823313790391156994766850629384787537055613862268777525467502123701520022205418828212212535352006690866031177264122804149317866157033558760231746361084940486770869585098883702738547895087079701619525682529118937970016022297132949865396730476441784507339276026144072103596164160025017182043218470275656098;
            6'd45: xpb[136] = 1024'd119340919102018570110508235524726163202921917201710760528293403357398189978991307310620447545304686111817619777679360736257837431492261526801239333604975247822483773597056179191860993478143484773390756224374733864657667555032844648378952272550861335882647047142032059075110792807614963450168848283736672579388;
            6'd46: xpb[136] = 1024'd3440319206122007665222776794008508873608351663823568150929484147695783100651270292397611663416345907501224116723963915132461704277145685488558310447258369770790101754956042162389009216874676745769695314679698764013004243822495390843060578688016780713966851593920916048011461377141268866036963522377475018347;
            6'd47: xpb[136] = 1024'd11606414994350186618736245468105287288993213251672059901697420002970271559620372184189846996185680012627977863226060528586149817903250178731037412305872532652787104482427122470547264147123074439458832013371903509732701782833042906272147454508401674812106559459926831051018658020596207299023768587643871941637;
            6'd48: xpb[136] = 1024'd19772510782578365572249714142202065704378074839520551652465355858244760018589474075982082328955014117754731609728157142039837931529354671973516514164486695534784107209898202778705519077371472133147968712064108255452399321843590421701234330328786568910246267325932746054025854664051145732010573652910268864927;
            6'd49: xpb[136] = 1024'd27938606570806544525763182816298844119762936427369043403233291713519248477558575967774317661724348222881485356230253755493526045155459165215995616023100858416781109937369283086863774007619869826837105410756313001172096860854137937130321206149171463008385975191938661057033051307506084164997378718176665788217;
            6'd50: xpb[136] = 1024'd36104702359034723479276651490395622535147798015217535154001227568793736936527677859566552994493682328008239102732350368947214158781563658458474717881715021298778112664840363395022028937868267520526242109448517746891794399864685452559408081969556357106525683057944576060040247950961022597984183783443062711507;
            6'd51: xpb[136] = 1024'd44270798147262902432790120164492400950532659603066026904769163424068225395496779751358788327263016433134992849234446982400902272407668151700953819740329184180775115392311443703180283868116665214215378808140722492611491938875232967988494957789941251204665390923950491063047444594415961030970988848709459634797;
            6'd52: xpb[136] = 1024'd52436893935491081386303588838589179365917521190914518655537099279342713854465881643151023660032350538261746595736543595854590386033772644943432921598943347062772118119782524011338538798365062907904515506832927238331189477885780483417581833610326145302805098789956406066054641237870899463957793913975856558087;
            6'd53: xpb[136] = 1024'd60602989723719260339817057512685957781302382778763010406305035134617202313434983534943258992801684643388500342238640209308278499659877138185912023457557509944769120847253604319496793728613460601593652205525131984050887016896327998846668709430711039400944806655962321069061837881325837896944598979242253481377;
            6'd54: xpb[136] = 1024'd68769085511947439293330526186782736196687244366611502157072970989891690772404085426735494325571018748515254088740736822761966613285981631428391125316171672826766123574724684627655048658861858295282788904217336729770584555906875514275755585251095933499084514521968236072069034524780776329931404044508650404667;
            6'd55: xpb[136] = 1024'd76935181300175618246843994860879514612072105954459993907840906845166179231373187318527729658340352853642007835242833436215654726912086124670870227174785835708763126302195764935813303589110255988971925602909541475490282094917423029704842461071480827597224222387974151075076231168235714762918209109775047327957;
            6'd56: xpb[136] = 1024'd85101277088403797200357463534976293027456967542308485658608842700440667690342289210319964991109686958768761581744930049669342840538190617913349329033399998590760129029666845243971558519358653682661062301601746221209979633927970545133929336891865721695363930253980066078083427811690653195905014175041444251247;
            6'd57: xpb[136] = 1024'd93267372876631976153870932209073071442841829130156977409376778555715156149311391102112200323879021063895515328247026663123030954164295111155828430892014161472757131757137925552129813449607051376350199000293950966929677172938518060563016212712250615793503638119985981081090624455145591628891819240307841174537;
            6'd58: xpb[136] = 1024'd101433468664860155107384400883169849858226690718005469160144714410989644608280492993904435656648355169022269074749123276576719067790399604398307532750628324354754134484609005860288068379855449070039335698986155712649374711949065575992103088532635509891643345985991896084097821098600530061878624305574238097827;
            6'd59: xpb[136] = 1024'd109599564453088334060897869557266628273611552305853960910912650266264133067249594885696670989417689274149022821251219890030407181416504097640786634609242487236751137212080086168446323310103846763728472397678360458369072250959613091421189964353020403989783053851997811087105017742055468494865429370840635021117;
            6'd60: xpb[136] = 1024'd117765660241316513014411338231363406688996413893702452661680586121538621526218696777488906322187023379275776567753316503484095295042608590883265736467856650118748139939551166476604578240352244457417609096370565204088769789970160606850276840173405298087922761718003726090112214385510406927852234436107031944407;
            6'd61: xpb[136] = 1024'd1865060345419950569125879500645752359682848355815260284316666911836214647878659759266070440298683174959380906797919682358719567827492749570584713310139772067054468097451029447132593979083436429796548186675530103444106478759811349314385146310560742919242566169892583063012882955036712343720349674747834383366;
            6'd62: xpb[136] = 1024'd10031156133648129522639348174742530775067709943663752035084602767110703106847761651058305773068017280086134653300016295812407681453597242813063815168753934949051470824922109755290848909331834123485684885367734849163804017770358864743472022130945637017382274035898498066020079598491650776707154740014231306656;
            6'd63: xpb[136] = 1024'd18197251921876308476152816848839309190452571531512243785852538622385191565816863542850541105837351385212888399802112909266095795079701736055542917027368097831048473552393190063449103839580231817174821584059939594883501556780906380172558897951330531115521981901904413069027276241946589209693959805280628229946;
        endcase
    end

    always_comb begin
        case(flag[45][16:12])
            5'd0: xpb[137] = 1024'd0;
            5'd1: xpb[137] = 1024'd26363347710104487429666285522936087605837433119360735536620474477659680024785965434642776438606685490339642146304209522719783908705806229298022018885982260713045476279864270371607358769828629510863958282752144340603199095791453895601645773771715425213661689767910328072034472885401527642680764870547025153236;
            5'd2: xpb[137] = 1024'd52726695420208974859332571045872175211674866238721471073240948955319360049571930869285552877213370980679284292608419045439567817411612458596044037771964521426090952559728540743214717539657259021727916565504288681206398191582907791203291547543430850427323379535820656144068945770803055285361529741094050306472;
            5'd3: xpb[137] = 1024'd79090043130313462288998856568808262817512299358082206609861423432979040074357896303928329315820056471018926438912628568159351726117418687894066056657946782139136428839592811114822076309485888532591874848256433021809597287374361686804937321315146275640985069303730984216103418656204582928042294611641075459708;
            5'd4: xpb[137] = 1024'd105453390840417949718665142091744350423349732477442942146481897910638720099143861738571105754426741961358568585216838090879135634823224917192088075543929042852181905119457081486429435079314518043455833131008577362412796383165815582406583095086861700854646759071641312288137891541606110570723059482188100612944;
            5'd5: xpb[137] = 1024'd7750042866397695749532500209866005284488738471067993554970517323321504786620688263198810978375753142255061324063554179019855702687810811934949969413580262631536706829750134520406554657625941833009593805373481856651634628736372705043250299175347676801488545425434582330065836353079005196285134526109531281849;
            5'd6: xpb[137] = 1024'd34113390576502183179198785732802092890326171590428729091590991800981184811406653697841587416982438632594703470367763701739639611393617041232971988299562523344582183109614404892013913427454571343873552088125626197254833724527826600644896072947063102015150235193344910402100309238480532838965899396656556435085;
            5'd7: xpb[137] = 1024'd60476738286606670608865071255738180496163604709789464628211466278640864836192619132484363855589124122934345616671973224459423520099423270530994007185544784057627659389478675263621272197283200854737510370877770537858032820319280496246541846718778527228811924961255238474134782123882060481646664267203581588321;
            5'd8: xpb[137] = 1024'd86840085996711158038531356778674268102001037829150200164831940756300544860978584567127140294195809613273987762976182747179207428805229499829016026071527044770673135669342945635228630967111830365601468653629914878461231916110734391848187620490493952442473614729165566546169255009283588124327429137750606741557;
            5'd9: xpb[137] = 1024'd113203433706815645468197642301610355707838470948510935701452415233960224885764550001769916732802495103613629909280392269898991337511035729127038044957509305483718611949207216006835989736940459876465426936382059219064431011902188287449833394262209377656135304497075894618203727894685115767008194008297631894793;
            5'd10: xpb[137] = 1024'd15500085732795391499065000419732010568977476942135987109941034646643009573241376526397621956751506284510122648127108358039711405375621623869899938827160525263073413659500269040813109315251883666019187610746963713303269257472745410086500598350695353602977090850869164660131672706158010392570269052219062563698;
            5'd11: xpb[137] = 1024'd41863433442899878928731285942668098174814910061496722646561509124302689598027341961040398395358191774849764794431317880759495314081427853167921957713142785976118889939364539412420468085080513176883145893499108053906468353264199305688146372122410778816638780618779492732166145591559538035251033922766087716934;
            5'd12: xpb[137] = 1024'd68226781153004366358397571465604185780652343180857458183181983601962369622813307395683174833964877265189406940735527403479279222787234082465943976599125046689164366219228809784027826854909142687747104176251252394509667449055653201289792145894126204030300470386689820804200618476961065677931798793313112870170;
            5'd13: xpb[137] = 1024'd94590128863108853788063856988540273386489776300218193719802458079622049647599272830325951272571562755529049087039736926199063131493040311763965995485107307402209842499093080155635185624737772198611062459003396735112866544847107096891437919665841629243962160154600148876235091362362593320612563663860138023406;
            5'd14: xpb[137] = 1024'd120953476573213341217730142511476360992327209419578929256422932557281729672385238264968727711178248245868691233343946448918847040198846541061988014371089568115255318778957350527242544394566401709475020741755541075716065640638560992493083693437557054457623849922510476948269564247764120963293328534407163176642;
            5'd15: xpb[137] = 1024'd23250128599193087248597500629598015853466215413203980664911551969964514359862064789596432935127259426765183972190662537059567108063432435804849908240740787894610120489250403561219663972877825499028781416120445569954903886209118115129750897526043030404465636276303746990197509059237015588855403578328593845547;
            5'd16: xpb[137] = 1024'd49613476309297574678263786152534103459303648532564716201532026447624194384648030224239209373733944917104826118494872059779351016769238665102871927126723048607655596769114673932827022742706455009892739698872589910558102982000572010731396671297758455618127326044214075062231981944638543231536168448875618998783;
            5'd17: xpb[137] = 1024'd75976824019402062107930071675470191065141081651925451738152500925283874409433995658881985812340630407444468264799081582499134925475044894400893946012705309320701073048978944304434381512535084520756697981624734251161302077792025906333042445069473880831789015812124403134266454830040070874216933319422644152019;
            5'd18: xpb[137] = 1024'd102340171729506549537596357198406278670978514771286187274772975402943554434219961093524762250947315897784110411103291105218918834180851123698915964898687570033746549328843214676041740282363714031620656264376878591764501173583479801934688218841189306045450705580034731206300927715441598516897698189969669305255;
            5'd19: xpb[137] = 1024'd4636823755486295568463715316527933532117520764911238683261594815626339121696787618152467474896327078680603149950007193359638902045437018441777858768338789813101351039136267710018859860675137821174416938741783086003339419154036924571355422929675281992292491933828001248228872526914493142459773233891099974160;
            5'd20: xpb[137] = 1024'd31000171465590782998130000839464021137954953884271974219882069293286019146482753052795243913503012569020245296254216716079422810751243247739799877654321050526146827319000538081626218630503767332038375221493927426606538514945490820173001196701390707205954181701738329320263345412316020785140538104438125127396;
            5'd21: xpb[137] = 1024'd57363519175695270427796286362400108743792387003632709756502543770945699171268718487438020352109698059359887442558426238799206719457049477037821896540303311239192303598864808453233577400332396842902333504246071767209737610736944715774646970473106132419615871469648657392297818297717548427821302974985150280632;
            5'd22: xpb[137] = 1024'd83726866885799757857462571885336196349629820122993445293123018248605379196054683922080796790716383549699529588862635761518990628162855706335843915426285571952237779878729078824840936170161026353766291786998216107812936706528398611376292744244821557633277561237558985464332291183119076070502067845532175433868;
            5'd23: xpb[137] = 1024'd110090214595904245287128857408272283955467253242354180829743492726265059220840649356723573229323069040039171735166845284238774536868661935633865934312267832665283256158593349196448294939989655864630250069750360448416135802319852506977938518016536982846939251005469313536366764068520603713182832716079200587104;
            5'd24: xpb[137] = 1024'd12386866621883991317996215526393938816606259235979232238232112138947843908317475881351278453272080220935664474013561372379494604733247830376727828181919052444638057868886402230425414518301079654184010744115264942654974047890409629614605722105022958793781037359262583578294708879993498338744907760000631256009;
            5'd25: xpb[137] = 1024'd38750214331988478747662501049330026422443692355339967774852586616607523933103441315994054891878765711275306620317770895099278513439054059674749847067901313157683534148750672602032773288129709165047969026867409283258173143681863525216251495876738384007442727127172911650329181765395025981425672630547656409245;
            5'd26: xpb[137] = 1024'd65113562042092966177328786572266114028281125474700703311473061094267203957889406750636831330485451201614948766621980417819062422144860288972771865953883573870729010428614942973640132057958338675911927309619553623861372239473317420817897269648453809221104416895083239722363654650796553624106437501094681562481;
            5'd27: xpb[137] = 1024'd91476909752197453606995072095202201634118558594061438848093535571926883982675372185279607769092136691954590912926189940538846330850666518270793884839865834583774486708479213345247490827786968186775885592371697964464571335264771316419543043420169234434766106662993567794398127536198081266787202371641706715717;
            5'd28: xpb[137] = 1024'd117840257462301941036661357618138289239955991713422174384714010049586564007461337619922384207698822182294233059230399463258630239556472747568815903725848095296819962988343483716854849597615597697639843875123842305067770431056225212021188817191884659648427796430903895866432600421599608909467967242188731868953;
            5'd29: xpb[137] = 1024'd20136909488281687067528715736259944101094997707047225793202629462269348694938164144550089431647833363190725798077115551399350307421058642311677797595499315076174764698636536750831969175927021487193604549488746799306608676626782334657856021280370635595269582784697165908360545233072503535030042286110162537858;
            5'd30: xpb[137] = 1024'd46500257198386174497195001259196031706932430826407961329823103939929028719724129579192865870254518853530367944381325074119134216126864871609699816481481575789220240978500807122439327945755650998057562832240891139909807772418236230259501795052086060808931272552607493980395018118474031177710807156657187691094;
            5'd31: xpb[137] = 1024'd72863604908490661926861286782132119312769863945768696866443578417588708744510095013835642308861204343870010090685534596838918124832671100907721835367463836502265717258365077494046686715584280508921521114993035480513006868209690125861147568823801486022592962320517822052429491003875558820391572027204212844330;
        endcase
    end

    always_comb begin
        case(flag[46][5:0])
            6'd0: xpb[138] = 1024'd0;
            6'd1: xpb[138] = 1024'd49613476309297574678263786152534103459303648532564716201532026447624194384648030224239209373733944917104826118494872059779351016769238665102871927126723048607655596769114673932827022742706455009892739698872589910558102982000572010731396671297758455618127326044214075062231981944638543231536168448875618998783;
            6'd2: xpb[138] = 1024'd99226952618595149356527572305068206918607297065129432403064052895248388769296060448478418747467889834209652236989744119558702033538477330205743854253446097215311193538229347865654045485412910019785479397745179821116205964001144021462793342595516911236254652088428150124463963889277086463072336897751237997566;
            6'd3: xpb[138] = 1024'd24773733243767982635992431052787877633212518471958464476464224277895687816634951762702556906544160441871328948027122744758989209466495660753455656363838104889276115737772804460850829036602159308368021488230529885309948095780819259229211444210045917587562074718525167156589417759986996677489815520001262512018;
            6'd4: xpb[138] = 1024'd74387209553065557314256217205321981092516167004523180677996250725519882201282981986941766280278105358976155066521994804538340226235734325856327583490561153496931712506887478393677851779308614318260761187103119795868051077781391269960608115507804373205689400762739242218821399704625539909025983968876881510801;
            6'd5: xpb[138] = 1024'd124000685862363131992520003357856084551819815537087896879528277173144076585931012211180975654012050276080981185016866864317691243004972990959199510617284202104587309276002152326504874522015069328153500885975709706426154059781963280692004786805562828823816726806953317281053381649264083140562152417752500509584;
            6'd6: xpb[138] = 1024'd49547466487535965271984862105575755266425036943916928952928448555791375633269903525405113813088320883742657896054245489517978418932991321506911312727676209778552231475545608921701658073204318616736042976461059770619896191561638518458422888420091835175124149437050334313178835519973993354979631040002525024036;
            6'd7: xpb[138] = 1024'd99160942796833539950248648258109858725728685476481645154460475003415570017917933749644323186822265800847484014549117549297329435702229986609783239854399258386207828244660282854528680815910773626628782675333649681177999173562210529189819559717850290793251475481264409375410817464612536586515799488878144022819;
            6'd8: xpb[138] = 1024'd24707723422006373229713507005829529440333906883310677227860646386062869065256825063868461345898536408509160725586496174497616611630248317157495041964791266060172750444203739449725464367100022915211324765818999745371741305341885766956237661332379297144558898111361426407536271335322446800933278111128168537271;
            6'd9: xpb[138] = 1024'd74321199731303947907977293158363632899637555415875393429392672833687063449904855288107670719632481325613986844081368234276967628399486982260366969091514314667828347213318413382552487109806477925104064464691589655929844287342457777687634332630137752762686224155575501469768253279960990032469446560003787536054;
            6'd10: xpb[138] = 1024'd123934676040601522586241079310897736358941203948440109630924699281311257834552885512346880093366426242718812962576240294056318645168725647363238896218237363275483943982433087315379509852512932934996804163564179566487947269343029788419031003927896208380813550199789576532000235224599533264005615008879406534837;
            6'd11: xpb[138] = 1024'd49481456665774355865705938058617407073546425355269141704324870663958556881891776826571018252442696850380489673613618919256605821096743977910950698328629370949448866181976543910576293403702182223579346254049529630681689401122705026185449105542425214732120972829886593564125689095309443478423093631129431049289;
            6'd12: xpb[138] = 1024'd99094932975071930543969724211151510532850073887833857905856897111582751266539807050810227626176641767485315792108490979035956837865982643013822625455352419557104462951091217843403316146408637233472085952922119541239792383123277036916845776840183670350248298874100668626357671039947986709959262080005050048072;
            6'd13: xpb[138] = 1024'd24641713600244763823434582958871181247455295294662889979257068494230050313878698365034365785252912375146992503145869604236244013794000973561534427565744427231069385150634674438600099697597886522054628043407469605433534514902952274683263878454712676701555721504197685658483124910657896924376740702255074562524;
            6'd14: xpb[138] = 1024'd74255189909542338501698369111405284706758943827227606180789094941854244698526728589273575158986857292251818621640741664015595030563239638664406354692467475838724981919749348371427122440304341531947367742280059515991637496903524285414660549752471132319683047548411760720715106855296440155912909151130693561307;
            6'd15: xpb[138] = 1024'd123868666218839913179962155263939388166062592359792322382321121389478439083174758813512784532720802209356644740135613723794946047332478303767278281819190524446380578688864022304254145183010796541840107441152649426549740478904096296146057221050229587937810373592625835782947088799934983387449077600006312560090;
            6'd16: xpb[138] = 1024'd49415446844012746459427014011659058880667813766621354455721292772125738130513650127736922691797072817018321451172992348995233223260496634314990083929582532120345500888407478899450928734200045830422649531637999490743482610683771533912475322664758594289117796222722852815072542670644893601866556222256337074542;
            6'd17: xpb[138] = 1024'd99028923153310321137690800164193162339971462299186070657253319219749932515161680351976132065531017734123147569667864408774584240029735299417862011056305580728001097657522152832277951476906500840315389230510589401301585592684343544643871993962517049907245122266936927877304524615283436833402724671131956073325;
            6'd18: xpb[138] = 1024'd24575703778483154417155658911912833054576683706015102730653490602397231562500571666200270224607288341784824280705243033974871415957753629965573813166697588401966019857065609427474735028095750128897931320995939465495327724464018782410290095577046056258552544897033944909429978485993347047820203293381980587777;
            6'd19: xpb[138] = 1024'd74189180087780729095419445064446936513880332238579818932185517050021425947148601890439479598341233258889650399200115093754222432726992295068445740293420637009621616626180283360301757770802205138790671019868529376053430706464590793141686766874804511876679870941248019971661960430631890279356371742257599586560;
            6'd20: xpb[138] = 1024'd123802656397078303773683231216981039973183980771144535133717543497645620331796632114678688972075178175994476517694987153533573449496230960171317667420143685617277213395294957293128780513508660148683410718741119286611533688465162803873083438172562967494807196985462095033893942375270433510892540191133218585343;
            6'd21: xpb[138] = 1024'd49349437022251137053148089964700710687789202177973567207117714880292919379135523428902827131151448783656153228732365778733860625424249290719029469530535693291242135594838413888325564064697909437265952809226469350805275820244838041639501539787091973846114619615559112066019396245980343725310018813383243099795;
            6'd22: xpb[138] = 1024'd98962913331548711731411876117234814147092850710538283408649741327917113763783553653142036504885393700760979347227237838513211642193487955821901396657258741898897732363953087821152586807404364447158692508099059261363378802245410052370898211084850429464241945659773187128251378190618886956846187262258862098578;
            6'd23: xpb[138] = 1024'd24509693956721545010876734864954484861698072117367315482049912710564412811122444967366174663961664308422656058264616463713498818121506286369613198767650749572862654563496544416349370358593613735741234598584409325557120934025085290137316312699379435815549368289870204160376832061328797171263665884508886613030;
            6'd24: xpb[138] = 1024'd74123170266019119689140521017488588321001720649932031683581939158188607195770475191605384037695609225527482176759488523492849834890744951472485125894373798180518251332611218349176393101300068745633974297456999236115223916025657300868712983997137891433676694334084279222608814005967340402799834333384505611813;
            6'd25: xpb[138] = 1024'd123736646575316694367404307170022691780305369182496747885113965605812801580418505415844593411429554142632308295254360583272200851659983616575357053021096846788173848101725892282003415844006523755526713996329589146673326898026229311600109655294896347051804020378298354284840795950605883634336002782260124610596;
            6'd26: xpb[138] = 1024'd49283427200489527646869165917742362494910590589325779958514136988460100627757396730068731570505824750293985006291739208472488027588001947123068855131488854462138770301269348877200199395195773044109256086814939210867069029805904549366527756909425353403111443008395371316966249821315793848753481404510149125048;
            6'd27: xpb[138] = 1024'd98896903509787102325132952070276465954214239121890496160046163436084295012405426954307940944239769667398811124786611268251839044357240612225940782258211903069794367070384022810027222137902228054001995785687529121425172011806476560097924428207183809021238769052609446379198231765954337080289649853385768123831;
            6'd28: xpb[138] = 1024'd24443684134959935604597810817996136668819460528719528233446334818731594059744318268532079103316040275060487835823989893452126220285258942773652584368603910743759289269927479405224005689091477342584537876172879185618914143586151797864342529821712815372546191682706463411323685636664247294707128475635792638283;
            6'd29: xpb[138] = 1024'd74057160444257510282861596970530240128123109061284244434978361266355788444392348492771288477049985192165313954318861953231477237054497607876524511495326959351414886039042153338051028431797932352477277575045469096177017125586723808595739201119471270990673517726920538473555667581302790526243296924511411637066;
            6'd30: xpb[138] = 1024'd123670636753555084961125383123064343587426757593848960636510387713979982829040378717010497850783930109270140072813734013010828253823736272979396438622050007959070482808156827270878051174504387362370017273918059006735120107587295819327135872417229726608800843771134613535787649525941333757779465373387030635849;
            6'd31: xpb[138] = 1024'd49217417378727918240590241870784014302031979000677992709910559096627281876379270031234636009860200716931816783851112638211115429751754603527108240732442015633035405007700283866074834725693636650952559364403409070928862239366971057093553974031758732960108266401231630567913103396651243972196943995637055150301;
            6'd32: xpb[138] = 1024'd98830893688025492918854028023318117761335627533242708911442585544251476261027300255473845383594145634036642902345984697990466446520993268629980167859165064240691001776814957798901857468400091660845299063275998981486965221367543067824950645329517188578235592445445705630145085341289787203733112444512674149084;
            6'd33: xpb[138] = 1024'd24377674313198326198318886771037788475940848940071740984842756926898775308366191569697983542670416241698319613383363323190753622449011599177691969969557071914655923976358414394098641019589340949427841153761349045680707353147218305591368746944046194929543015075542722662270539211999697418150591066762698663536;
            6'd34: xpb[138] = 1024'd73991150622495900876582672923571891935244497472636457186374783374522969693014221793937192916404361158803145731878235382970104639218250264280563897096280120522311520745473088326925663762295795959320580852633938956238810335147790316322765418241804650547670341119756797724502521156638240649686759515638317662319;
            6'd35: xpb[138] = 1024'd123604626931793475554846459076105995394548146005201173387906809822147164077662252018176402290138306075907971850373107442749455655987488929383435824223003169129967117514587762259752686505002250969213320551506528866796913317148362327054162089539563106165797667163970872786734503101276783881222927964513936661102;
            6'd36: xpb[138] = 1024'd49151407556966308834311317823825666109153367412030205461306981204794463125001143332400540449214576683569648561410486067949742831915507259931147626333395176803932039714131218854949470056191500257795862641991878930990655448928037564820580191154092112517105089794067889818859956971986694095640406586763961175554;
            6'd37: xpb[138] = 1024'd98764883866263883512575103976359769568457015944594921662839007652418657509649173556639749822948521600674474679905358127729093848684745925034019553460118225411587636483245892787776492798897955267688602340864468841548758430928609575551976862451850568135232415838281964881091938916625237327176575035639580174337;
            6'd38: xpb[138] = 1024'd24311664491436716792039962724079440283062237351423953736239179035065956556988064870863887982024792208336151390942736752929381024612764255581731355570510233085552558682789349382973276350087204556271144431349818905742500562708284813318394964066379574486539838468378981913217392787335147541594053657889604688789;
            6'd39: xpb[138] = 1024'd73925140800734291470303748876613543742365885883988669937771205482690150941636095095103097355758737125440977509437608812708732041382002920684603282697233281693208155451904023315800299092793659566163884130222408816300603544708856824049791635364138030104667164512593056975449374731973690773130222106765223687572;
            6'd40: xpb[138] = 1024'd123538617110031866148567535029147647201669534416553386139303231930314345326284125319342306729492682042545803627932480872488083058151241585787475209823956330300863752221018697248627321835500114576056623829094998726858706526709428834781188306661896485722794490556807132037681356676612234004666390555640842686355;
            6'd41: xpb[138] = 1024'd49085397735204699428032393776867317916274755823382418212703403312961644373623016633566444888568952650207480338969859497688370234079259916335187011934348337974828674420562153843824105386689363864639165919580348791052448658489104072547606408276425492074101913186904149069806810547322144219083869177890867200807;
            6'd42: xpb[138] = 1024'd98698874044502274106296179929401421375578404355947134414235429760585838758271046857805654262302897567312306457464731557467721250848498581438058939061071386582484271189676827776651128129395818874531905618452938701610551640489676083279003079574183947692229239231118224132038792491960687450620037626766486199590;
            6'd43: xpb[138] = 1024'd24245654669675107385761038677121092090183625762776166487635601143233137805609938172029792421379168174973983168502110182668008426776516911985770741171463394256449193389220284371847911680585068163114447708938288765804293772269351321045421181188712954043536661861215241164164246362670597665037516249016510714042;
            6'd44: xpb[138] = 1024'd73859130978972682064024824829655195549487274295340882689167627590857332190257968396269001795113113092078809286996982242447359443545755577088642668298186442864104790158334958304674934423291523173007187407810878676362396754269923331776817852486471409661663987905429316226396228307309140896573684697892129712825;
            6'd45: xpb[138] = 1024'd123472607288270256742288610982189299008790922827905598890699654038481526574905998620508211168847058009183635405491854302226710460314994242191514595424909491471760386927449632237501957165997978182899927106683468586920499736270495342508214523784229865279791313949643391288628210251947684128109853146767748711608;
            6'd46: xpb[138] = 1024'd49019387913443090021753469729908969723396144234734630964099825421128825622244889934732349327923328616845312116529232927426997636243012572739226397535301499145725309126993088832698740717187227471482469197168818651114241868050170580274632625398758871631098736579740408320753664122657594342527331769017773226060;
            6'd47: xpb[138] = 1024'd98632864222740664700017255882443073182699792767299347165631851868753020006892920158971558701657273533950138235024104987206348653012251237842098324662024547753380905896107762765525763459893682481375208896041408561672344850050742591006029296696517327249226062623954483382985646067296137574063500217893392224843;
            6'd48: xpb[138] = 1024'd24179644847913497979482114630162743897305014174128379239032023251400319054231811473195696860733544141611814946061483612406635828940269568389810126772416555427345828095651219360722547011082931769957750986526758625866086981830417828772447398311046333600533485254051500415111099938006047788480978840143416739295;
            6'd49: xpb[138] = 1024'd73793121157211072657745900782696847356608662706693095440564049699024513438879841697434906234467489058716641064556355672185986845709508233492682053899139604035001424864765893293549569753789386779850490685399348536424189963830989839503844069608804789218660811298265575477343081882644591020017147289019035738078;
            6'd50: xpb[138] = 1024'd123406597466508647336009686935230950815912311239257811642096076146648707823527871921674115608201433975821467183051227731965337862478746898595553981025862652642657021633880567226376592496495841789743230384271938446982292945831561850235240740906563244836788137342479650539575063827283134251553315737894654736861;
            6'd51: xpb[138] = 1024'd48953378091681480615474545682950621530517532646086843715496247529296006870866763235898253767277704583483143894088606357165625038406765229143265783136254660316621943833424023821573376047685091078325772474757288511176035077611237088001658842521092251188095559972576667571700517697993044465970794360144679251313;
            6'd52: xpb[138] = 1024'd98566854400979055293738331835484724989821181178651559917028273976920201255514793460137463141011649500587970012583478416944976055176003894246137710262977708924277540602538697754400398790391546088218512173629878421734138059611809098733055513818850706806222886016790742633932499642631587697506962809020298250096;
            6'd53: xpb[138] = 1024'd24113635026151888573203190583204395704426402585480591990428445359567500302853684774361601300087920108249646723620857042145263231104022224793849512373369716598242462802082154349597182341580795376801054264115228485927880191391484336499473615433379713157530308646887759666057953513341497911924441431270322764548;
            6'd54: xpb[138] = 1024'd73727111335449463251466976735738499163730051118045308191960471807191694687501714998600810673821865025354472842115729101924614247873260889896721439500092765205898059571196828282424205084287250386693793962987818396485983173392056347230870286731138168775657634691101834728289935457980041143460609880145941763331;
            6'd55: xpb[138] = 1024'd123340587644747037929730762888272602623033699650610024393492498254815889072149745222840020047555809942459298960610601161703965264642499554999593366626815813813553656340311502215251227826993705396586533661860408307044086155392628357962266958028896624393784960735315909790521917402618584374996778329021560762114;
            6'd56: xpb[138] = 1024'd48887368269919871209195621635992273337638921057439056466892669637463188119488636537064158206632080550120975671647979786904252440570517885547305168737207821487518578539854958810448011378182954685169075752345758371237828287172303595728685059643425630745092383365412926822647371273328494589414256951271585276566;
            6'd57: xpb[138] = 1024'd98500844579217445887459407788526376796942569590003772668424696085087382504136666761303367580366025467225801790142851846683603457339756550650177095863930870095174175308969632743275034120889409695061815451218348281795931269172875606460081730941184086363219709409627001884879353217967037820950425400147204275349;
            6'd58: xpb[138] = 1024'd24047625204390279166924266536246047511547790996832804741824867467734681551475558075527505739442296074887478501180230471883890633267774881197888897974322877769139097508513089338471817672078658983644357541703698345989673400952550844226499832555713092714527132039724018917004807088676948035367904022397228789801;
            6'd59: xpb[138] = 1024'd73661101513687853845188052688780150970851439529397520943356893915358875936123588299766715113176240991992304619675102531663241650037013546300760825101045926376794694277627763271298840414785113993537097240576288256547776382953122854957896503853471548332654458083938093979236789033315491266904072471272847788584;
            6'd60: xpb[138] = 1024'd123274577822985428523451838841314254430155088061962237144888920362983070320771618524005924486910185909097130738169974591442592666806252211403632752227768974984450291046742437204125863157491569003429836939448878167105879364953694865689293175151230003950781784128152169041468770977954034498440240920148466787367;
            6'd61: xpb[138] = 1024'd48821358448158261802916697589033925144760309468791269218289091745630369368110509838230062645986456516758807449207353216642879842734270541951344554338160982658415213246285893799322646708680818292012379029934228231299621496733370103455711276765759010302089206758249186073594224848663944712857719542398491301819;
            6'd62: xpb[138] = 1024'd98434834757455836481180483741568028604063958001355985419821118193254563752758540062469272019720401433863633567702225276422230859503509207054216481464884031266070810015400567732149669451387273301905118728806818141857724478733942114187107948063517465920216532802463261135826206793302487944393887991274110300602;
            6'd63: xpb[138] = 1024'd23981615382628669760645342489287699318669179408185017493221289575901862800097431376693410178796672041525310278739603901622518035431527537601928283575276038940035732214944024327346453002576522590487660819292168206051466610513617351953526049678046472271523955432560278167951660664012398158811366613524134815054;
        endcase
    end

    always_comb begin
        case(flag[46][11:6])
            6'd0: xpb[139] = 1024'd0;
            6'd1: xpb[139] = 1024'd73595091691926244438909128641821802777972827940749733694753316023526057184745461600932619552530616958630136397234475961401869052200766202704800210701999087547691328984058698260173475745282977600380400518164758116609569592514189362684922720975804927889651281476774353230183642608650941390347535062399753813837;
            6'd2: xpb[139] = 1024'd23123487699727747479019329878829172811247228755763783261374776982075219032181784291850167890403559607817123387011458488224674263560312070854440296387667134161691983398546179182716712299048749479450603427942276386854778334807481952404866872268380406512482659539431648430260757143373249763576380298173913143343;
            6'd3: xpb[139] = 1024'd96718579391653991917928458520650975589220056696513516956128093005601276216927245892782787442934176566447259784245934449626543315761078273559240507089666221709383312382604877442890188044331727079831003946107034503464347927321671315089789593244185334402133941016206001660444399752024191153923915360573666957180;
            6'd4: xpb[139] = 1024'd46246975399455494958038659757658345622494457511527566522749553964150438064363568583700335780807119215634246774022916976449348527120624141708880592775334268323383966797092358365433424598097498958901206855884552773709556669614963904809733744536760813024965319078863296860521514286746499527152760596347826286686;
            6'd5: xpb[139] = 1024'd119842067091381739396947788399480148400467285452277300217502869987676495249109030184632955333337736174264383171257392937851217579321390344413680803477333355871075295781151056625606900343380476559281607374049310890319126262129153267494656465512565740914616600555637650090705156895397440917500295658747580100523;
            6'd6: xpb[139] = 1024'd69370463099183242437057989636487518433741686267291349784124330946225657096545352875550503671210678823451370161034375464674022790680936212563320889163001402485075950195638537548150136897146248438351810283826829160564335004422445857214600616805141219537447978618294945290782271430119749290729140894521739430029;
            6'd7: xpb[139] = 1024'd18898859106984745477168190873494888467016087082305399350745791904774818943981675566468052009083621472638357150811357991496828002040482080712960974848669449099076604610126018470693373450912020317422013193604347430809543746715738446934544768097716698160279356680952240490859385964842057663957986130295898759535;
            6'd8: xpb[139] = 1024'd92493950798910989916077319515316691244988915023055133045499107928300876128727137167400671561614238431268493548045833952898697054241248283417761185550668536646767933594184716730866849196194997917802413711769105547419113339229927809619467489073521626049930638157726593721043028573492999054305521192695652573372;
            6'd9: xpb[139] = 1024'd42022346806712492956187520752324061278263315838069182612120568886850037976163459858318219899487181080455480537822816479721502265600794151567401271236336583260768588008672197653410085749960769796872616621546623817664322081523220399339411640366097104672762016220383888921120143108215307427534366428469811902878;
            6'd10: xpb[139] = 1024'd115617438498638737395096649394145864056236143778818916306873884910376095160908921459250839452017798039085616935057292441123371317801560354272201481938335670808459916992730895913583561495243747397253017139711381934273891674037409762024334361341902032562413297697158242151303785716866248817881901490869565716715;
            6'd11: xpb[139] = 1024'd65145834506440240435206850631153234089510544593832965873495345868925257008345244150168387789890740688272603924834274967946176529161106222421841567624003717422460571407218376836126798049009519276323220049488900204519100416330702351744278512634477511185244675759815537351380900251588557191110746726643725046221;
            6'd12: xpb[139] = 1024'd14674230514241743475317051868160604122784945408847015440116806827474418855781566841085936127763683337459590914611257494768981740520652090571481653309671764036461225821705857758670034602775291155393422959266418474764309158623994941464222663927052989808076053822472832551458014786310865564339591962417884375727;
            6'd13: xpb[139] = 1024'd88269322206167987914226180509982406900757773349596749134870122851000476040527028442018555680294300296089727311845733456170850792721418293276281864011670851584152554805764556018843510348058268755773823477431176591373878751138184304149145384902857917697727335299247185781641657394961806954687127024817638189564;
            6'd14: xpb[139] = 1024'd37797718213969490954336381746989776934032174164610798701491583809549637887963351132936104018167242945276714301622715982993656004080964161425921949697338898198153209220252036941386746901824040634844026387208694861619087493431476893869089536195433396320558713361904480981718771929684115327915972260591797519070;
            6'd15: xpb[139] = 1024'd111392809905895735393245510388811579712005002105360532396244899833075695072708812733868723570697859903906850698857191944395525056281730364130722160399337985745844538204310735201560222647107018235224426905373452978228657085945666256554012257171238324210209994838678834211902414538335056718263507322991551332907;
            6'd16: xpb[139] = 1024'd60921205913697238433355711625818949745279402920374581962866360791624856920145135424786271908570802553093837688634174471218330267641276232280362246085006032359845192618798216124103459200872790114294629815150971248473865828238958846273956408463813802833041372901336129411979529073057365091492352558765710662413;
            6'd17: xpb[139] = 1024'd10449601921498741473465912862826319778553803735388631529487821750174018767581458115703820246443745202280824678411156998041135479000822100430002331770674078973845847033285697046646695754638561993364832724928489518719074570532251435993900559756389281455872750963993424612056643607779673464721197794539869991919;
            6'd18: xpb[139] = 1024'd84044693613424985912375041504648122556526631676138365224241137773700075952326919716636439798974362160910961075645632959443004531201588303134802542472673166521537176017344395306820171499921539593745233243093247635328644163046440798678823280732194209345524032440767777842240286216430614855068732856939623805756;
            6'd19: xpb[139] = 1024'd33573089621226488952485242741655492589801032491152414790862598732249237799763242407553988136847304810097948065422615486265809742561134171284442628158341213135537830431831876229363408053687311472815436152870765905573852905339733388398767432024769687968355410503425073042317400751152923228297578092713783135262;
            6'd20: xpb[139] = 1024'd107168181313152733391394371383477295367773860431902148485615914755775294984508704008486607689377921768728084462657091447667678794761900373989242838860340300683229159415890574489536883798970289073195836671035524022183422497853922751083690153000574615858006691980199426272501043359803864618645113155113536949099;
            6'd21: xpb[139] = 1024'd56696577320954236431504572620484665401048261246916198052237375714324456831945026699404156027250864417915071452434073974490484006121446242138882924546008347297229813830378055412080120352736060952266039580813042292428631240147215340803634304293150094480838070042856721472578157894526172991873958390887696278605;
            6'd22: xpb[139] = 1024'd6224973328755739471614773857492035434322662061930247618858836672873618679381349390321704365123807067102058442211056501313289217480992110288523010231676393911230468244865536334623356906501832831336242490590560562673839982440507930523578455585725573103669448105514016672655272429248481365102803626661855608111;
            6'd23: xpb[139] = 1024'd79820065020681983910523902499313838212295490002679981313612152696399675864126810991254323917654424025732194839445532462715158269681758312993323220933675481458921797228924234594796832651784810431716643008755318679283409574954697293208501176561530500993320729582288369902838915037899422755450338689061609421948;
            6'd24: xpb[139] = 1024'd29348461028483486950634103736321208245569890817694030880233613654948837711563133682171872255527366674919181829222514989537963481041304181142963306619343528072922451643411715517340069205550582310786845918532836949528618317247989882928445327854105979616152107644945665102916029572621731128679183924835768751454;
            6'd25: xpb[139] = 1024'd102943552720409731389543232378143011023542718758443764574986929678474894896308595283104491808057983633549318226456990950939832533242070383847763517321342615620613780627470413777513544950833559911167246436697595066138187909762179245613368048829910907505803389121720018333099672181272672519026718987235522565291;
            6'd26: xpb[139] = 1024'd52471948728211234429653433615150381056817119573457814141608390637024056743744917974022040145930926282736305216233973477762637744601616251997403603007010662234614435041957894700056781504599331790237449346475113336383396652055471835333312200122486386128634767184377313533176786715994980892255564223009681894797;
            6'd27: xpb[139] = 1024'd2000344736012737469763634852157751090091520388471863708229851595573218591181240664939588483803868931923292206010956004585442955961162120147043688692678708848615089456445375622600018058365103669307652256252631606628605394348764425053256351415061864751466145247034608733253901250717289265484409458783841224303;
            6'd28: xpb[139] = 1024'd75595436427938981908672763493979553868064348329221597402983167619099275775926702265872208036334485890553428603245431965987312008161928322851843899394677796396306418440504073882773493803648081269688052774417389723238174986862953787738179072390866792641117426723808961963437543859368230655831944521183595038140;
            6'd29: xpb[139] = 1024'd25123832435740484948782964730986923901338749144235646969604628577648437623363024956789756374207428539740415593022414492810117219521474191001483985080345843010307072854991554805316730357413853148758255684194907993483383729156246377458123223683442271263948804786466257163514658394090539029060789756957754367646;
            6'd30: xpb[139] = 1024'd98718924127666729387692093372808726679311577084985380664357944601174494808108486557722375926738045498370551990256890454211986271722240393706284195782344930557998401839050253065490206102696830749138656202359666110092953321670435740143045944659247199153600086263240610393698301002741480419408324819357508181483;
            6'd31: xpb[139] = 1024'd48247320135468232427802294609816096712585977899999430230979405559723656655544809248639924264610988147557538980033872981034791483081786261855924281468012977171999056253537733988033442656462602628208859112137184380338162063963728329862990095951822677776431464325897905593775415537463788792637170055131667510989;
            6'd32: xpb[139] = 1024'd121842411827394476866711423251637899490558805840749163925732721583249713840290270849572543817141605106187675377268348942436660535282552464560724492170012064719690385237596432248206918401745580228589259630301942496947731656477917692547912816927627605666082745802672258823959058146114730182984705117531421324826;
            6'd33: xpb[139] = 1024'd71370807835195979906821624488645269523833206655763213492354182541798875687726593540490092155014547755374662367045331469259465746642098332710364577855680111333691039652083913170750154955511352107659462540079460767192940398771210282267856968220203084288914123865329554024036172680837038556213550353305580654332;
            6'd34: xpb[139] = 1024'd20899203842997482946931825725652639557107607470777263058975643500348037535162916231407640492887490404561649356822313996082270958001644200860004663541348157947691694066571394093293391509277123986729665449856979037438149141064502871987801119512778562911745501927986849224113287215559346929442395589079739983838;
            6'd35: xpb[139] = 1024'd94494295534923727385840954367474442335080435411526996753728959523874094719908377832340260045418107363191785754056789957484140010202410403564804874243347245495383023050630092353466867254560101587110065968021737154047718733578692234672723840488583490801396783404761202454296929824210288319789930651479493797675;
            6'd36: xpb[139] = 1024'd44022691542725230425951155604481812368354836226541046320350420482423256567344700523257808383291050012378772743833772484306945221561956271714444959929015292109383677465117573276010103808325873466180268877799255424292927475871984824392667991781158969424228161467418497654374044358932596693018775887253653127181;
            6'd37: xpb[139] = 1024'd117617783234651474864860284246303615146327664167290780015103736505949313752090162124190427935821666971008909141068248445708814273762722474419245170631014379657075006449176271536183579553608851066560669395964013540902497068386174187077590712756963897313879442944192850884557686967583538083366310949653406941018;
            6'd38: xpb[139] = 1024'd67146179242452977904970485483310985179602064982304829581725197464498475599526484815107976273694609620195896130845230972531619485122268342568885256316682426271075660863663752458726816107374622945630872305741531811147705810679466776797534864049539375936710821006850146084634801502305846456595156185427566270524;
            6'd39: xpb[139] = 1024'd16674575250254480945080686720318355212876465797318879148346658423047637446962807506025524611567552269382883120622213499354424696481814210718525342002350472885076315278151233381270052661140394824701075215519050081392914552972759366517479015342114854559542199069507441284711916037028154829824001421201725600030;
            6'd40: xpb[139] = 1024'd90269666942180725383989815362140157990849293738068612843099974446573694631708269106958144164098169228013019517856689460756293748682580413423325552704349560432767644262209931641443528406423372425081475733683808198002484145486948729202401736317919782449193480546281794514895558645679096220171536483601479413867;
            6'd41: xpb[139] = 1024'd39798062949982228424100016599147528024123694553082662409721435405122856479144591797875692501971111877200006507633671987579098960042126281572965638390017607046768298676697412563986764960189144304151678643461326468247692887780241318922345887610495261072024858608939089714972673180401404593400381719375638743373;
            6'd42: xpb[139] = 1024'd113393154641908472863009145240969330802096522493832396104474751428648913663890053398808312054501728835830142904868147948980968012242892484277765849092016694594459627660756110824160240705472121904532079161626084584857262480294430681607268608586300188961676140085713442945156315789052345983747916781775392557210;
            6'd43: xpb[139] = 1024'd62921550649709975903119346477976700835370923308846445671096212387198075511326376089725860392374671485017129894645130475803773223602438352427405934777684741208460282075243591746703477259237893783602282071403602855102471222587723271327212759878875667584507518148370738145233430323774654356976762017549551886716;
            6'd44: xpb[139] = 1024'd12449946657511478943229547714984070868645324123860495237717673345747237358762698780643408730247614134204116884422113002626578434961984220577046020463352787822460936489731072669246713813003665662672484981181121125347679964881015861047156911171451146207338896211028033345310544858496962730205607253323711216222;
            6'd45: xpb[139] = 1024'd86045038349437723382138676356805873646618152064610228932470989369273294543508160381576028282778231092834253281656588964028447487162750423281846231165351875370152265473789770929420189558286643263052885499345879241957249557395205223732079632147256074096990177687802386575494187467147904120553142315723465030059;
            6'd46: xpb[139] = 1024'd35573434357239226422248877593813243679892552879624278499092450327822456390944483072493576620651173742021240271433571490851252698522296291431486316851019921984152919888277251851963426112052415142123088409123397512202458299688497813452023783439831552719821555750459681775571302001870212493781987551497624359565;
            6'd47: xpb[139] = 1024'd109168526049165470861158006235635046457865380820374012193845766351348513575689944673426196173181790700651376668668047452253121750723062494136286527553019009531844248872335950112136901857335392742503488927288155628812027892202687176136946504415636480609472837227234035005754944610521153884129522613897378173402;
            6'd48: xpb[139] = 1024'd58696922056966973901268207472642416491139781635388061760467227309897675423126267364343744511054733349838363658445029979075926962082608362285926613238687056145844903286823431034680138411101164621573691837065673899057236634495979765856890655708211959232304215289891330205832059145243462257358367849671537502908;
            6'd49: xpb[139] = 1024'd8225318064768476941378408709649786524414182450402111327088688268446837270562590055261292848927675999025350648222012505898732173442154230435566698924355102759845557701310911957223374964866936500643894746843192169302445376789272355576834807000787437855135593352548625405909173679965770630587213085445696832414;
            6'd50: xpb[139] = 1024'd81820409756694721380287537351471589302387010391151845021842004291972894455308051656193912401458292957655487045456488467300601225642920433140366909626354190307536886685369610217396850710149914101024295265007950285912014969303461718261757527976592365744786874829322978636092816288616712020934748147845450646251;
            6'd51: xpb[139] = 1024'd31348805764496224420397738588478959335661411206165894588463465250522056302744374347111460739331235606842474035233470994123406437002466301290006995312022236921537541099857091139940087263915685980094498174785468556157223711596754307981701679269167844367618252891980273836169930823339020394163593383619609975757;
            6'd52: xpb[139] = 1024'd104943897456422468859306867230300762113634239146915628283216781274048113487489835948044080291861852565472610432467946955525275489203232503994807206014021324469228870083915789400113563009198663580474898692950226672766793304110943670666624400244972772257269534368754627066353573431989961784511128446019363789594;
            6'd53: xpb[139] = 1024'd54472293464223971899417068467308132146908639961929677849838242232597275334926158638961628629734795214659597422244929482348080700562778372144447291699689371083229524498403270322656799562964435459545101602727744943012002046404236260386568551537548250880100912431411922266430687966712270157739973681793523119100;
            6'd54: xpb[139] = 1024'd4000689472025474939527269704315502180183040776943727416459703191146437182362481329879176967607737863846584412021912009170885911922324240294087377385357417697230178912890751245200036116730207338615304512505263213257210788697528850106512702830123729502932290494069217466507802501434578530968818917567682448606;
            6'd55: xpb[139] = 1024'd77595781163951719378436398346137304958155868717693461111213019214672494367107942930811796520138354822476720809256387970572754964123090442998887588087356505244921507896949449505373511862013184938995705030670021329866780381211718212791435423805928657392583571970843570696691445110085519921316353979967436262443;
            6'd56: xpb[139] = 1024'd27124177171753222418546599583144674991430269532707510677834480173221656214544265621729344858011297471663707799033370497395560175482636311148527673773024551858922162311436930427916748415778956818065907940447539600111989123505010802511379575098504136015414950033500865896768559644807828294545199215741595591949;
            6'd57: xpb[139] = 1024'd100719268863679466857455728224966477769403097473457244372587796196747713399289727222661964410541914430293844196267846458797429227683402513853327884475023639406613491295495628688090224161061934418446308458612297716721558716019200165196302296074309063905066231510275219126952202253458769684892734278141349405786;
            6'd58: xpb[139] = 1024'd50247664871480969897565929461973847802677498288471293939209257155296875246726049913579512748414857079480831186044828985620234439042948382002967970160691686020614145709983109610633460714827706297516511368389815986966767458312492754916246447366884542527897609572932514327029316788181078058121579513915508735292;
            6'd59: xpb[139] = 1024'd123842756563407214336475058103795650580650326229221027633962573178822932431471511514512132300945474038110967583279304947022103491243714584707768180862690773568305474694041807870806936460110683897896911886554574103576337050826682117601169168342689470417548891049706867557212959396832019448469114576315262549129;
            6'd60: xpb[139] = 1024'd73371152571208717376585259340803020613924727044235077200584034137372094278907834205429680638818416687297954573056287473844908702603260452857408266548358820182306129108529288793350173013876455776967114796332092373821545793119974707321113319635264949040380269112364162757290073931554327821697959812089421878635;
            6'd61: xpb[139] = 1024'd22899548579010220416695460577810390647199127859249126767205495095921256126344156896347228976691359336484941562833270000667713913962806321007048352234026866796306783523016769715893409567642227656037317706109610644066754535413267297041057470927840427663211647175021457957367188466276636194926805047863581208141;
            6'd62: xpb[139] = 1024'd96494640270936464855604589219632193425171955799998860461958811119447313311089618497279848529221976295115077960067745962069582966163572523711848562936025954343998112507075467976066885312925205256417718224274368760676324127927456659725980191903645355552862928651795811187550831074927577585274340110263335021978;
            6'd63: xpb[139] = 1024'd46023036278737967895714790456639563458446356615012910028580272077996475158525941188197396867094918944302064949844728488892388177523118391861488648621694000957998766921562948898610121866690977135487921134051887030921532870220749249445924343196220834175694306714453106387627945609649885958503185346037494351484;
        endcase
    end

    always_comb begin
        case(flag[46][16:12])
            5'd0: xpb[140] = 1024'd0;
            5'd1: xpb[140] = 1024'd119618127970664212334623919098461366236419184555762643723333588101522532343271402789130016419625535902932201347079204450294257229723884594566288859323693088505690095905621647158783597611973954735868321652216645147531102462734938612130847064172025762065345588191227459617811588218300827348850720408437248165321;
            5'd2: xpb[140] = 1024'd115169560257203683270448910792108299728139941985789603318535321138068169349233666668244961624593397496421253286700915466009450618606548854577417593631055136077689517241672076979936956032430703750426445696046050448697844075248980451296715558660822074863871272968337861205516648362673021680582750990248901846311;
            5'd3: xpb[140] = 1024'd110720992543743154206273902485755233219860699415816562913737054174613806355195930547359906829561259089910305226322626481724644007489213114588546327938417183649688938577722506801090314452887452764984569739875455749864585687763022290462584053149618387662396957745448262793221708507045216012314781572060555527301;
            5'd4: xpb[140] = 1024'd106272424830282625142098894179402166711581456845843522508938787211159443361158194426474852034529120683399357165944337497439837396371877374599675062245779231221688359913772936622243672873344201779542693783704861051031327300277064129628452547638414700460922642522558664380926768651417410344046812153872209208291;
            5'd5: xpb[140] = 1024'd101823857116822096077923885873049100203302214275870482104140520247705080367120458305589797239496982276888409105566048513155030785254541634610803796553141278793687781249823366443397031293800950794100817827534266352198068912791105968794321042127211013259448327299669065968631828795789604675778842735683862889281;
            5'd6: xpb[140] = 1024'd97375289403361567013748877566696033695022971705897441699342253284250717373082722184704742444464843870377461045187759528870224174137205894621932530860503326365687202585873796264550389714257699808658941871363671653364810525305147807960189536616007326057974012076779467556336888940161799007510873317495516570271;
            5'd7: xpb[140] = 1024'd92926721689901037949573869260342967186743729135924401294543986320796354379044986063819687649432705463866512984809470544585417563019870154633061265167865373937686623921924226085703748134714448823217065915193076954531552137819189647126058031104803638856499696853889869144041949084533993339242903899307170251261;
            5'd8: xpb[140] = 1024'd88478153976440508885398860953989900678464486565951360889745719357341991385007249942934632854400567057355564924431181560300610951902534414644189999475227421509686045257974655906857106555171197837775189959022482255698293750333231486291926525593599951655025381631000270731747009228906187670974934481118823932251;
            5'd9: xpb[140] = 1024'd84029586262979979821223852647636834170185243995978320484947452393887628390969513822049578059368428650844616864052892576015804340785198674655318733782589469081685466594025085728010464975627946852333314002851887556865035362847273325457795020082396264453551066408110672319452069373278382002706965062930477613241;
            5'd10: xpb[140] = 1024'd79581018549519450757048844341283767661906001426005280080149185430433265396931777701164523264336290244333668803674603591730997729667862934666447468089951516653684887930075515549163823396084695866891438046681292858031776975361315164623663514571192577252076751185221073907157129517650576334438995644742131294231;
            5'd11: xpb[140] = 1024'd75132450836058921692873836034930701153626758856032239675350918466978902402894041580279468469304151837822720743296314607446191118550527194677576202397313564225684309266125945370317181816541444881449562090510698159198518587875357003789532009059988890050602435962331475494862189662022770666171026226553784975221;
            5'd12: xpb[140] = 1024'd70683883122598392628698827728577634645347516286059199270552651503524539408856305459394413674272013431311772682918025623161384507433191454688704936704675611797683730602176375191470540236998193896007686134340103460365260200389398842955400503548785202849128120739441877082567249806394964997903056808365438656211;
            5'd13: xpb[140] = 1024'd66235315409137863564523819422224568137068273716086158865754384540070176414818569338509358879239875024800824622539736638876577896315855714699833671012037659369683151938226805012623898657454942910565810178169508761532001812903440682121268998037581515647653805516552278670272309950767159329635087390177092337201;
            5'd14: xpb[140] = 1024'd61786747695677334500348811115871501628789031146113118460956117576615813420780833217624304084207736618289876562161447654591771285198519974710962405319399706941682573274277234833777257077911691925123934221998914062698743425417482521287137492526377828446179490293662680257977370095139353661367117971988746018191;
            5'd15: xpb[140] = 1024'd57338179982216805436173802809518435120509788576140078056157850613161450426743097096739249289175598211778928501783158670306964674081184234722091139626761754513681994610327664654930615498368440939682058265828319363865485037931524360453005987015174141244705175070773081845682430239511547993099148553800399699181;
            5'd16: xpb[140] = 1024'd52889612268756276371998794503165368612230546006167037651359583649707087432705360975854194494143459805267980441404869686022158062963848494733219873934123802085681415946378094476083973918825189954240182309657724665032226650445566199618874481503970454043230859847883483433387490383883742324831179135612053380171;
            5'd17: xpb[140] = 1024'd48441044555295747307823786196812302103951303436193997246561316686252724438667624854969139699111321398757032381026580701737351451846512754744348608241485849657680837282428524297237332339281938968798306353487129966198968262959608038784742975992766766841756544624993885021092550528255936656563209717423707061161;
            5'd18: xpb[140] = 1024'd43992476841835218243648777890459235595672060866220956841763049722798361444629888734084084904079182992246084320648291717452544840729177014755477342548847897229680258618478954118390690759738687983356430397316535267365709875473649877950611470481563079640282229402104286608797610672628130988295240299235360742151;
            5'd19: xpb[140] = 1024'd39543909128374689179473769584106169087392818296247916436964782759343998450592152613199030109047044585735136260270002733167738229611841274766606076856209944801679679954529383939544049180195436997914554441145940568532451487987691717116479964970359392438807914179214688196502670817000325320027270881047014423141;
            5'd20: xpb[140] = 1024'd35095341414914160115298761277753102579113575726274876032166515795889635456554416492313975314014906179224188199891713748882931618494505534777734811163571992373679101290579813760697407600652186012472678484975345869699193100501733556282348459459155705237333598956325089784207730961372519651759301462858668104131;
            5'd21: xpb[140] = 1024'd30646773701453631051123752971400036070834333156301835627368248832435272462516680371428920518982767772713240139513424764598125007377169794788863545470934039945678522626630243581850766021108935027030802528804751170865934713015775395448216953947952018035859283733435491371912791105744713983491332044670321785121;
            5'd22: xpb[140] = 1024'd26198205987993101986948744665046969562555090586328795222569981868980909468478944250543865723950629366202292079135135780313318396259834054799992279778296087517677943962680673403004124441565684041588926572634156472032676325529817234614085448436748330834384968510545892959617851250116908315223362626481975466111;
            5'd23: xpb[140] = 1024'd21749638274532572922773736358693903054275848016355754817771714905526546474441208129658810928918490959691344018756846796028511785142498314811121014085658135089677365298731103224157482862022433056147050616463561773199417938043859073779953942925544643632910653287656294547322911394489102646955393208293629147101;
            5'd24: xpb[140] = 1024'd17301070561072043858598728052340836545996605446382714412973447942072183480403472008773756133886352553180395958378557811743705174025162574822249748393020182661676786634781533045310841282479182070705174660292967074366159550557900912945822437414340956431436338064766696135027971538861296978687423790105282828091;
            5'd25: xpb[140] = 1024'd12852502847611514794423719745987770037717362876409674008175180978617820486365735887888701338854214146669447898000268827458898562907826834833378482700382230233676207970831962866464199702935931085263298704122372375532901163071942752111690931903137269229962022841877097722733031683233491310419454371916936509081;
            5'd26: xpb[140] = 1024'd8403935134150985730248711439634703529438120306436633603376914015163457492327999767003646543822075740158499837621979843174091951790491094844507217007744277805675629306882392687617558123392680099821422747951777676699642775585984591277559426391933582028487707618987499310438091827605685642151484953728590190071;
            5'd27: xpb[140] = 1024'd3955367420690456666073703133281637021158877736463593198578647051709094498290263646118591748789937333647551777243690858889285340673155354855635951315106325377675050642932822508770916543849429114379546791781182977866384388100026430443427920880729894827013392396097900898143151971977879973883515535540243871061;
            5'd28: xpb[140] = 1024'd123573495391354669000697622231743003257578062292226236921912235153231626841561666435248608168415473236579753124322895309183542570397039949421924810638799413883365146548554469667554514155823383850247868443997828125397486850834965042574274985052755656892358980587325360515954740190278707322734235943977492036382;
            5'd29: xpb[140] = 1024'd119124927677894139936522613925389936749298819722253196517113968189777263847523930314363553373383334830068805063944606324898735959279704209433053544946161461455364567884604899488707872576280132864805992487827233426564228463349006881740143479541551969690884665364435762103659800334650901654466266525789145717372;
            5'd30: xpb[140] = 1024'd114676359964433610872347605619036870241019577152280156112315701226322900853486194193478498578351196423557857003566317340613929348162368469444182279253523509027363989220655329309861230996736881879364116531656638727730970075863048720906011974030348282489410350141546163691364860479023095986198297107600799398362;
            5'd31: xpb[140] = 1024'd110227792250973081808172597312683803732740334582307115707517434262868537859448458072593443783319058017046908943188028356329122737045032729455311013560885556599363410556705759131014589417193630893922240575486044028897711688377090560071880468519144595287936034918656565279069920623395290317930327689412453079352;
        endcase
    end

    always_comb begin
        case(flag[47][5:0])
            6'd0: xpb[141] = 1024'd0;
            6'd1: xpb[141] = 1024'd52889612268756276371998794503165368612230546006167037651359583649707087432705360975854194494143459805267980441404869686022158062963848494733219873934123802085681415946378094476083973918825189954240182309657724665032226650445566199618874481503970454043230859847883483433387490383883742324831179135612053380171;
            6'd2: xpb[141] = 1024'd105779224537512552743997589006330737224461092012334075302719167299414174865410721951708388988286919610535960882809739372044316125927696989466439747868247604171362831892756188952167947837650379908480364619315449330064453300891132399237748963007940908086461719695766966866774980767767484649662358271224106760342;
            6'd3: xpb[141] = 1024'd34602141122144087717197456104681673091993210892765428825946895884144366960806944017547512267772705106360791916757115623487410348050325149644499496786040365323353573269563066090621682564958364141410349320585934148732319101115801825891644874828681912862872676129533392270055943077722593957374847580210565656182;
            6'd4: xpb[141] = 1024'd87491753390900364089196250607847041704223756898932466477306479533851454393512304993401706761916164911628772358161985309509568411014173644377719370720164167409034989215941160566705656483783554095650531630243658813764545751561368025510519356332652366906103535977416875703443433461606336282206026715822619036353;
            6'd5: xpb[141] = 1024'd16314669975531899062396117706197977571755875779363820000534208118581646488908527059240830041401950407453603392109361560952662633136801804555779119637956928561025730592748037705159391211091538328580516331514143632432411551786037452164415268153393371682514492411183301106724395771561445589918516024809077932193;
            6'd6: xpb[141] = 1024'd69204282244288175434394912209363346183986421785530857651893791768288733921613888035095024535545410212721583833514231246974820696100650299288998993572080730646707146539126132181243365129916728282820698641171868297464638202231603651783289749657363825725745352259066784540111886155445187914749695160421131312364;
            6'd7: xpb[141] = 1024'd122093894513044451806393706712528714796216967791697895303253375417995821354319249010949219029688870017989564274919100932996978759064498794022218867506204532732388562485504226657327339048741918237060880950829592962496864852677169851402164231161334279768976212106950267973499376539328930239580874296033184692535;
            6'd8: xpb[141] = 1024'd50916811097675986779593573810879650663749086672129248826481104002726013449715471076788342309174655513814395308866477184440072981187126954200278616423997293884379303862311103795781073776049902469990865652100077781164730652901839278056060142982075284545387168540716693376780338849284039547293363605019643588375;
            6'd9: xpb[141] = 1024'd103806423366432263151592368314045019275979632678296286477840687652433100882420832052642536803318115319082375750271346870462231044150975448933498490358121095970060719808689198271865047694875092424231047961757802446196957303347405477674934624486045738588618028388600176810167829233167781872124542740631696968546;
            6'd10: xpb[141] = 1024'd32629339951063798124792235412395955143511751558727640001068416237163292977817054118481660082803900814907206784218723121905325266273603609111558239275913857122051461185496075410318782422183076657161032663028287264864823103572074904328830536306786743365028984822366602213448791543122891179837032049618155864386;
            6'd11: xpb[141] = 1024'd85518952219820074496791029915561323755742297564894677652427999886870380410522415094335854576947360620175187225623592807927483329237452103844778113210037659207732877131874169886402756341008266611401214972686011929897049754017641103947705017810757197408259844670250085646836281927006633504668211185230209244557;
            6'd12: xpb[141] = 1024'd14341868804451609469990897013912259623274416445326031175655728471600572505918637160174977856433146116000018259570969059370577551360080264022837862127830420359723618508681047024856491068316250844331199673956496748564915554242310530601600929631498202184670801104016511050117244236961742812380700494216668140397;
            6'd13: xpb[141] = 1024'd67231481073207885841989691517077628235504962451493068827015312121307659938623998136029172350576605921267998700975838745392735614323928758756057736061954222445405034455059141500940464987141440798571381983614221413597142204687876730220475411135468656227901660951899994483504734620845485137211879629828721520568;
            6'd14: xpb[141] = 1024'd120121093341964162213988486020242996847735508457660106478374895771014747371329359111883366844720065726535979142380708431414893677287777253489277609996078024531086450401437235977024438905966630752811564293271946078629368855133442929839349892639439110271132520799783477916892225004729227462043058765440774900739;
            6'd15: xpb[141] = 1024'd48944009926595697187188353118593932715267627338091460001602624355744939466725581177722490124205851222360810176328084682857987899410405413667337358913870785683077191778244113115478173633274614985741548994542430897297234655358112356493245804460180115047543477233549903320173187314684336769755548074427233796579;
            6'd16: xpb[141] = 1024'd101833622195351973559187147621759301327498173344258497652962208005452026899430942153576684618349311027628790617732954368880145962374253908400557232847994587768758607724622207591562147552099804939981731304200155562329461305803678556112120285964150569090774337081433386753560677698568079094586727210039287176750;
            6'd17: xpb[141] = 1024'd30656538779983508532387014720110237195030292224689851176189936590182218994827164219415807897835096523453621651680330620323240184496882068578616981765787348920749349101429084730015882279407789172911716005470640380997327106028347982766016197784891573867185293515199812156841640008523188402299216519025746072590;
            6'd18: xpb[141] = 1024'd83546151048739784904385809223275605807260838230856888827549520239889306427532525195270002391978556328721602093085200306345398247460730563311836855699911151006430765047807179206099856198232979127151898315128365046029553756473914182384890679288862027910416153363083295590229130392406930727130395654637799452761;
            6'd19: xpb[141] = 1024'd12369067633371319877585676321626541674792957111288242350777248824619498522928747261109125671464341824546433127032576557788492469583358723489896604617703912158421506424614056344553590925540963360081883016398849864697419556698583609038786591109603032686827109796849720993510092702362040034842884963624258348601;
            6'd20: xpb[141] = 1024'd65258679902127596249584470824791910287023503117455280002136832474326585955634108236963320165607801629814413568437446243810650532547207218223116478551827714244102922370992150820637564844366153314322065326056574529729646207144149808657661072613573486730057969644733204426897583086245782359674064099236311728772;
            6'd21: xpb[141] = 1024'd118148292170883872621583265327957278899254049123622317653496416124033673388339469212817514659751261435082394009842315929832808595511055712956336352485951516329784338317370245296721538763191343268562247635714299194761872857589716008276535554117543940773288829492616687860285073470129524684505243234848365108943;
            6'd22: xpb[141] = 1024'd46971208755515407594783132426308214766786168004053671176724144708763865483735691278656637939237046930907225043789692181275902817633683873134396101403744277481775079694177122435175273490499327501492232336984784013429738657814385434930431465938284945549699785926383113263566035780084633992217732543834824004783;
            6'd23: xpb[141] = 1024'd99860821024271683966781926929473583379016714010220708828083728358470952916441052254510832433380506736175205485194561867298060880597532367867615975337868079567456495640555216911259247409324517455732414646642508678461965308259951634549305947442255399592930645774266596696953526163968376317048911679446877384954;
            6'd24: xpb[141] = 1024'd28683737608903218939981794027824519246548832890652062351311456943201145011837274320349955712866292232000036519141938118741155102720160528045675724255660840719447237017362094049712982136632501688662399347912993497129831108484621061203201859262996404369341602208033022100234488473923485624761400988433336280794;
            6'd25: xpb[141] = 1024'd81573349877659495311980588530989887858779378896819100002671040592908232444542635296204150207009752037268016960546807804763313165684009022778895598189784642805128652963740188525796956055457691642902581657570718162162057758930187260822076340766966858412572462055916505533621978857807227949592580124045389660965;
            6'd26: xpb[141] = 1024'd10396266462291030285180455629340823726311497777250453525898769177638424539938857362043273486495537533092847994494184056206407387806637182956955347107577403957119394340547065664250690782765675875832566358841202980829923559154856687475972252587707863188983418489682930936902941167762337257305069433031848556805;
            6'd27: xpb[141] = 1024'd63285878731047306657179250132506192338542043783417491177258352827345511972644218337897467980638997338360828435899053742228565450770485677690175221041701206042800810286925160140334664701590865830072748668498927645862150209600422887094846734091678317232214278337566414370290431551646079582136248568643901936976;
            6'd28: xpb[141] = 1024'd116175490999803583029178044635671560950772589789584528828617936477052599405349579313751662474782457143628808877303923428250723513734334172423395094975825008128482226233303254616418638620416055784312930978156652310894376860045989086713721215595648771275445138185449897803677921935529821906967427704255955317147;
            6'd29: xpb[141] = 1024'd44998407584435118002377911734022496818304708670015882351845665061782791500745801379590785754268242639453639911251299679693817735856962332601454843893617769280472967610110131754872373347724040017242915679427137129562242660270658513367617127416389776051856094619216323206958884245484931214679917013242414212987;
            6'd30: xpb[141] = 1024'd97888019853191394374376706237187865430535254676182920003205248711489878933451162355444980248411702444721620352656169365715975798820810827334674717827741571366154383556488226230956347266549229971483097989084861794594469310716224712986491608920360230095086954467099806640346374629368673539511096148854467593158;
            6'd31: xpb[141] = 1024'd26710936437822929347576573335538801298067373556614273526432977296220071028847384421284103527897487940546451386603545617159070020943438987512734466745534332518145124933295103369410081993857214204413082690355346613262335110940894139640387520741101234871497910900866232043627336939323782847223585457840926488998;
            6'd32: xpb[141] = 1024'd79600548706579205719575367838704169910297919562781311177792560945927158461552745397138298022040947745814431828008415303181228083907287482245954340679658134603826540879673197845494055912682404158653265000013071278294561761386460339259262002245071688914728770748749715477014827323207525172054764593452979869169;
            6'd33: xpb[141] = 1024'd8423465291210740692775234937055105777830038443212664701020289530657350556948967462977421301526733241639262861955791554624322306029915642424014089597450895755817282256480074983947790639990388391583249701283556096962427561611129765913157914065812693691139727182516140880295789633162634479767253902439438765009;
            6'd34: xpb[141] = 1024'd61313077559967017064774029440220474390060584449379702352379873180364437989654328438831615795670193046907243303360661240646480368993764137157233963531574697841498698202858169460031764558815578345823432010941280761994654212056695965532032395569783147734370587030399624313683280017046376804598433038051492145180;
            6'd35: xpb[141] = 1024'd114202689828723293436772823943385843002291130455546740003739456830071525422359689414685810289813652852175223744765530926668638431957612631890453837465698499927180114149236263936115738477640768300063614320599005427026880862502262165150906877073753601777601446878283107747070770400930119129429612173663545525351;
            6'd36: xpb[141] = 1024'd43025606413354828409972691041736778869823249335978093526967185414801717517755911480524933569299438348000054778712907178111732654080240792068513586383491261079170855526043141074569473204948752532993599021869490245694746662726931591804802788894494606554012403312049533150351732710885228437142101482650004421191;
            6'd37: xpb[141] = 1024'd95915218682111104781971485544902147482053795342145131178326769064508804950461272456379128063442898153268035220117776864133890717044089286801733460317615063164852271472421235550653447123773942487233781331527214910726973313172497791423677270398465060597243263159933016583739223094768970761973280618262057801362;
            6'd38: xpb[141] = 1024'd24738135266742639755171352643253083349585914222576484701554497649238997045857494522218251342928683649092866254065153115576984939166717446979793209235407824316843012849228112689107181851081926720163766032797699729394839113397167218077573182219206065373654219593699441987020185404724080069685769927248516697202;
            6'd39: xpb[141] = 1024'd77627747535498916127170147146418451961816460228743522352914081298946084478562855498072445837072143454360846695470022801599143002130565941713013083169531626402524428795606207165191155769907116674403948342455424394427065763842733417696447663723176519416885079441582925420407675788607822394516949062860570077373;
            6'd40: xpb[141] = 1024'd6450664120130451100370014244769387829348579109174875876141809883676276573959077563911569116557928950185677729417399053042237224253194101891072832087324387554515170172413084303644890497215100907333933043725909213094931564067402844350343575543917524193296035875349350823688638098562931702229438371847028973213;
            6'd41: xpb[141] = 1024'd59340276388886727472368808747934756441579125115341913527501393533383364006664438539765763610701388755453658170822268739064395287217042596624292706021448189640196586118791178779728864416040290861574115353383633878127158214512969043969218057047887978236526895723232834257076128482446674027060617507459082353384;
            6'd42: xpb[141] = 1024'd112229888657643003844367603251100125053809671121508951178860977183090451439369799515619958104844848560721638612227138425086553350180891091357512579955571991725878002065169273255812838334865480815814297663041358543159384864958535243588092538551858432279757755571116317690463618866330416351891796643071135733555;
            6'd43: xpb[141] = 1024'd41052805242274538817567470349451060921341790001940304702088705767820643534766021581459081384330634056546469646174514676529647572303519251535572328873364752877868743441976150394266573062173465048744282364311843361827250665183204670241988450372599437056168712004882743093744581176285525659604285952057594629395;
            6'd44: xpb[141] = 1024'd93942417511030815189566264852616429533572336008107342353448289417527730967471382557313275878474093861814450087579384362551805635267367746268792202807488554963550159388354244870350546980998655002984464673969568026859477315628770869860862931876569891099399571852766226527132071560169267984435465087669648009566;
            6'd45: xpb[141] = 1024'd22765334095662350162766131950967365401104454888538695876676018002257923062867604623152399157959879357639281121526760613994899857389995906446851951725281316115540900765161122008804281708306639235914449375240052845527343115853440296514758843697310895875810528286532651930413033870124377292147954396656106905406;
            6'd46: xpb[141] = 1024'd75654946364418626534764926454132734013335000894705733528035601651965010495572965599006593652103339162907261562931630300017057920353844401180071825659405118201222316711539216484888255627131829190154631684897777510559569766299006496133633325201281349919041388134416135363800524254008119616979133532268160285577;
            6'd47: xpb[141] = 1024'd4477862949050161507964793552483669880867119775137087051263330236695202590969187664845716931589124658732092596879006551460152142476472561358131574577197879353213058088346093623341990354439813423084616386168262329227435566523675922787529237022022354695452344568182560767081486563963228924691622841254619181417;
            6'd48: xpb[141] = 1024'd57367475217806437879963588055649038493097665781304124702622913886402290023674548640699911425732584464000073038283876237482310205440321056091351448511321681438894474034724188099425964273265003377324798695825986994259662216969242122406403718525992808738683204416066044200468976947846971249522801976866672561588;
            6'd49: xpb[141] = 1024'd110257087486562714251962382558814407105328211787471162353982497536109377456379909616554105919876044269268053479688745923504468268404169550824571322445445483524575889981102282575509938192090193331564981005483711659291888867414808322025278200029963262781914064263949527633856467331730713574353981112478725941759;
            6'd50: xpb[141] = 1024'd39080004071194249225162249657165342972860330667902515877210226120839569551776131682393229199361829765092884513636122174947562490526797711002631071363238244676566631357909159713963672919398177564494965706754196477959754667639477748679174111850704267558325020697715953037137429641685822882066470421465184837599;
            6'd51: xpb[141] = 1024'd91969616339950525597161044160330711585090876674069553528569809770546656984481492658247423693505289570360864955040991860969720553490646205735850945297362046762248047304287254190047646838223367518735148016411921142991981318085043948298048593354674721601555880545599436470524920025569565206897649557077238217770;
            6'd52: xpb[141] = 1024'd20792532924582060570360911258681647452622995554500907051797538355276849079877714724086546972991075066185695988988368112412814775613274365913910694215154807914238788681094131328501381565531351751665132717682405961659847118309713374951944505175415726377966836979365861873805882335524674514610138866063697113610;
            6'd53: xpb[141] = 1024'd73682145193338336942359705761847016064853541560667944703157122004983936512583075699940741467134534871453676430393237798434972838577122860647130568149278609999920204627472225804585355484356541705905315027340130626692073768755279574570818986679386180421197696827249345307193372719408416839441318001675750493781;
            6'd54: xpb[141] = 1024'd2505061777969871915559572860197951932385660441099298226384850589714128607979297765779864746620320367278507464340614049878067060699751020825190317067071371151910946004279102943039090211664525938835299728610615445359939568979949001224714898500127185197608653261015770710474335029363526147153807310662209389621;
            6'd55: xpb[141] = 1024'd55394674046726148287558367363363320544616206447266335877744434239421216040684658741634059240763780172546487905745483735900225123663599515558410191001195173237592361950657197419123064130489715893075482038268340110392166219425515200843589380004097639240839513108899254143861825413247268471984986446274262769792;
            6'd56: xpb[141] = 1024'd108284286315482424659557161866528689156846752453433373529104017889128303473390019717488253734907239977814468347150353421922383186627448010291630064935318975323273777897035291895207038049314905847315664347926064775424392869871081400462463861508068093284070372956782737577249315797131010796816165581886316149963;
            6'd57: xpb[141] = 1024'd37107202900113959632757028964879625024378871333864727052331746473858495568786241783327377014393025473639299381097729673365477408750076170469689813853111736475264519273842169033660772776622890080245649049196549594092258670095750827116359773328809098060481329390549162980530278107086120104528654890872775045803;
            6'd58: xpb[141] = 1024'd89996815168870236004755823468044993636609417340031764703691330123565583001491602759181571508536485278907279822502599359387635471713924665202909687787235538560945935220220263509744746695448080034485831358854274259124485320541317026735234254832779552103712189238432646413917768490969862429359834026484828425974;
            6'd59: xpb[141] = 1024'd18819731753501770977955690566395929504141536220463118226919058708295775096887824825020694788022270774732110856449975610830729693836552825380969436705028299712936676597027140648198481422756064267415816060124759077792351120765986453389130166653520556880123145672199071817198730800924971737072323335471287321814;
            6'd60: xpb[141] = 1024'd71709344022258047349954485069561298116372082226630155878278642358002862529593185800874889282165730580000091297854845296852887756800401320114189310639152101798618092543405235124282455341581254221655998369782483742824577771211552653008004648157491010923354005520082555250586221184808714061903502471083340701985;
            6'd61: xpb[141] = 1024'd532260606889582323154352167912233983904201107061509401506370942733054624989407866714012561651516075824922331802221548295981978923029480292249059556944862950608833920212112262736190068889238454585983071052968561492443571436222079661900559978232015699764961953848980653867183494763823369615991780069799597825;
            6'd62: xpb[141] = 1024'd53421872875645858695153146671077602596134747113228547052865954592440142057694768842568207055794975881092902773207091234318140041886877975025468933491068665036290249866590206738820163987714428408826165380710693226524670221881788279280775041482202469742995821801732464087254673878647565694447170915681852977996;
            6'd63: xpb[141] = 1024'd106311485144402135067151941174242971208365293119395584704225538242147229490400129818422401549938435686360883214611960920340298104850726469758688807425192467121971665812968301214904137906539618363066347690368417891556896872327354478899649522986172923786226681649615947520642164262531308019278350051293906358167;
        endcase
    end

    always_comb begin
        case(flag[47][11:6])
            6'd0: xpb[142] = 1024'd0;
            6'd1: xpb[142] = 1024'd35134401729033670040351808272593907075897411999826938227453266826877421585796351884261524829424221182185714248559337171783392326973354629936748556342985228273962407189775178353357872633847602595996332391638902710224762672552023905553545434806913928562637638083382372923923126572486417326990839360280365254007;
            6'd2: xpb[142] = 1024'd70268803458067340080703616545187814151794823999653876454906533653754843171592703768523049658848442364371428497118674343566784653946709259873497112685970456547924814379550356706715745267695205191992664783277805420449525345104047811107090869613827857125275276166764745847846253144972834653981678720560730508014;
            6'd3: xpb[142] = 1024'd105403205187101010121055424817781721227692235999480814682359800480632264757389055652784574488272663546557142745678011515350176980920063889810245669028955684821887221569325535060073617901542807787988997174916708130674288017656071716660636304420741785687912914250147118771769379717459251980972518080841095762021;
            6'd4: xpb[142] = 1024'd16470911232009938762608305685561195558891220873572068781681212242532791005876268627031028103039210419299707586779855252554505467052198185191834100355609872162158954189529496075801251343873204662675131958168370994534689839987198849249203169544426264983730648919412433665585978216017036290844667614495866531697;
            6'd5: xpb[142] = 1024'd51605312961043608802960113958155102634788632873399007009134479069410212591672620511292552932463431601485421835339192424337897794025552815128582656698595100436121361379304674429159123977720807258671464349807273704759452512539222754802748604351340193546368287002794806589509104788503453617835506974776231785704;
            6'd6: xpb[142] = 1024'd86739714690077278843311922230749009710686044873225945236587745896287634177468972395554077761887652783671136083898529596121290120998907445065331213041580328710083768569079852782516996611568409854667796741446176414984215185091246660356294039158254122109005925086177179513432231360989870944826346335056597039711;
            6'd7: xpb[142] = 1024'd121874116419110948883663730503342916786583456873052883464041012723165055763265324279815602591311873965856850332457866767904682447972262075002079769384565556984046175758855031135874869245416012450664129133085079125208977857643270565909839473965168050671643563169559552437355357933476288271817185695336962293718;
            6'd8: xpb[142] = 1024'd32941822464019877525216611371122391117782441747144137563362424485065582011752537254062056206078420838599415173559710505109010934104396370383668200711219744324317908379058992151602502687746409325350263916336741989069379679974397698498406339088852529967461297838824867331171956432034072581689335228991733063394;
            6'd9: xpb[142] = 1024'd68076224193053547565568419643716298193679853746971075790815691311943003597548889138323581035502642020785129422119047676892403261077751000320416757054204972598280315568834170504960375321594011921346596307975644699294142352526421604051951773895766458530098935922207240255095083004520489908680174589272098317401;
            6'd10: xpb[142] = 1024'd103210625922087217605920227916310205269577265746798014018268958138820425183345241022585105864926863202970843670678384848675795588051105630257165313397190200872242722758609348858318247955441614517342928699614547409518905025078445509605497208702680387092736574005589613179018209577006907235671013949552463571408;
            6'd11: xpb[142] = 1024'd14278331966996146247473108784089679600776250620889268117590369900720951431832453996831559479693410075713408511780228585880124074183239925638753744723844388212514455378813309874045881397772011392029063482866210273379306847409572642194064073826364866388554308674854928072834808075564691545543163483207234341084;
            6'd12: xpb[142] = 1024'd49412733696029816287824917056683586676673662620716206345043636727598373017628805881093084309117631257899122760339565757663516401156594555575502301066829616486476862568588488227403754031619613988025395874505112983604069519961596547747609508633278794951191946758237300996757934648051108872534002843487599595091;
            6'd13: xpb[142] = 1024'd84547135425063486328176725329277493752571074620543144572496903554475794603425157765354609138541852440084837008898902929446908728129949185512250857409814844760439269758363666580761626665467216584021728266144015693828832192513620453301154943440192723513829584841619673920681061220537526199524842203767964849098;
            6'd14: xpb[142] = 1024'd119681537154097156368528533601871400828468486620370082799950170381353216189221509649616133967966073622270551257458240101230301055103303815448999413752800073034401676948138844934119499299314819180018060657782918404053594865065644358854700378247106652076467222925002046844604187793023943526515681564048330103105;
            6'd15: xpb[142] = 1024'd30749243199006085010081414469650875159667471494461336899271582143253742437708722623862587582732620495013116098560083838434629541235438110830587845079454260374673409568342805949847132741645216054704195441034581267913996687396771491443267243370791131372284957594267361738420786291581727836387831097703100872781;
            6'd16: xpb[142] = 1024'd65883644928039755050433222742244782235564883494288275126724848970131164023505074508124112412156841677198830347119421010218021868208792740767336401422439488648635816758117984303205005375492818650700527832673483978138759359948795396996812678177705059934922595677649734662343912864068145163378670457983466126788;
            6'd17: xpb[142] = 1024'd101018046657073425090785031014838689311462295494115213354178115797008585609301426392385637241581062859384544595678758182001414195182147370704084957765424716922598223947893162656562878009340421246696860224312386688363522032500819302550358112984618988497560233761032107586267039436554562490369509818263831380795;
            6'd18: xpb[142] = 1024'd12085752701982353732337911882618163642661280368206467453499527558909111857788639366632090856347609732127109436780601919205742681314281666085673389092078904262869956568097123672290511451670818121382995007564049552223923854831946435138924978108303467793377968430297422480083637935112346800241659351918602150471;
            6'd19: xpb[142] = 1024'd47220154431016023772689720155212070718558692368033405680952794385786533443584991250893615685771830914312823685339939090989135008287636296022421945435064132536832363757872302025648384085518420717379327399202952262448686527383970340692470412915217396356015606513679795404006764507598764127232498712198967404478;
            6'd20: xpb[142] = 1024'd82354556160049693813041528427805977794456104367860343908406061212663955029381343135155140515196052096498537933899276262772527335260990925959170501778049360810794770947647480379006256719366023313375659790841854972673449199935994246246015847722131324918653244597062168327929891080085181454223338072479332658485;
            6'd21: xpb[142] = 1024'd117488957889083363853393336700399884870353516367687282135859328039541376615177695019416665344620273278684252182458613434555919662234345555895919058121034589084757178137422658732364129353213625909371992182480757682898211872488018151799561282529045253481290882680444541251853017652571598781214177432759697912492;
            6'd22: xpb[142] = 1024'd28556663933992292494946217568179359201552501241778536235180739801441902863664907993663118959386820151426817023560457171760248148366479851277507489447688776425028910757626619748091762795544022784058126965732420546758613694819145284388128147652729732777108617349709856145669616151129383091086326966414468682168;
            6'd23: xpb[142] = 1024'd63691065663025962535298025840773266277449913241605474462634006628319324449461259877924643788811041333612531272119794343543640475339834481214256045790674004698991317947401798101449635429391625380054459357371323256983376367371169189941673582459643661339746255433092229069592742723615800418077166326694833936175;
            6'd24: xpb[142] = 1024'd98825467392059632575649834113367173353347325241432412690087273455196746035257611762186168618235262515798245520679131515327032802313189111151004602133659232972953725137176976454807508063239227976050791749010225967208139039923193095495219017266557589902383893516474601993515869296102217745068005686975199190182;
            6'd25: xpb[142] = 1024'd9893173436968561217202714981146647684546310115523666789408685217097272283744824736432622233001809388540810361780975252531361288445323406532593033460313420313225457757380937470535141505569624850736926532261888831068540862254320228083785882390242069198201628185739916887332467794660002054940155220629969959858;
            6'd26: xpb[142] = 1024'd45027575166002231257554523253740554760443722115350605016861952043974693869541176620694147062426030570726524610340312424314753615418678036469341589803298648587187864947156115823893014139417227446733258923900791541293303534806344133637331317197155997760839266269122289811255594367146419381930994580910335213865;
            6'd27: xpb[142] = 1024'd80161976895035901297906331526334461836341134115177543244315218870852115455337528504955671891850251752912238858899649596098145942392032666406090146146283876861150272136931294177250886773264830042729591315539694251518066207358368039190876752004069926323476904352504662735178720939632836708921833941190700467872;
            6'd28: xpb[142] = 1024'd115296378624069571338258139798928368912238546115004481471768485697729537041133880389217196721274472935097953107458986767881538269365387296342838702489269105135112679326706472530608759407112432638725923707178596961742828879910391944744422186810983854886114542435887035659101847512119254035912673301471065721879;
            6'd29: xpb[142] = 1024'd26364084668978499979811020666707843243437530989095735571089897459630063289621093363463650336041019807840517948560830505085866755497521591724427133815923292475384411946910433546336392849442829513412058490430259825603230702241519077332989051934668334181932277105152350552918446010677038345784822835125836491555;
            6'd30: xpb[142] = 1024'd61498486398012170020162828939301750319334942988922673798543164286507484875417445247725175165465240990026232197120167676869259082470876221661175690158908520749346819136685611899694265483290432109408390882069162535827993374793542982886534486741582262744569915188534723476841572583163455672775662195406201745562;
            6'd31: xpb[142] = 1024'd96632888127045840060514637211895657395232354988749612025996431113384906461213797131986699994889462172211946445679504848652651409444230851597924246501893749023309226326460790253052138117138034705404723273708065246052756047345566888440079921548496191307207553271917096400764699155649872999766501555686566999569;
            6'd32: xpb[142] = 1024'd7700594171954768702067518079675131726431339862840866125317842875285432709701010106233153609656009044954511286781348585856979895576365146979512677828547936363580958946664751268779771559468431580090858056959728109913157869676694021028646786672180670603025287941182411294581297654207657309638651089341337769245;
            6'd33: xpb[142] = 1024'd42834995900988438742419326352269038802328751862667804352771109702162854295497361990494678439080230227140225535340685757640372222549719776916261234171533164637543366136439929622137644193316034176087190448598630820137920542228717926582192221479094599165662926024564784218504424226694074636629490449621703023252;
            6'd34: xpb[142] = 1024'd77969397630022108782771134624862945878226163862494742580224376529040275881293713874756203268504451409325939783900022929423764549523074406853009790514518392911505773326215107975495516827163636772083522840237533530362683214780741832135737656286008527728300564107947157142427550799180491963620329809902068277259;
            6'd35: xpb[142] = 1024'd113103799359055778823122942897456852954123575862321680807677643355917697467090065759017728097928672591511654032459360101207156876496429036789758346857503621185468180515990286328853389461011239368079855231876436240587445887332765737689283091092922456290938202191329530066350677371666909290611169170182433531266;
            6'd36: xpb[142] = 1024'd24171505403964707464675823765236327285322560736412934906999055117818223715577278733264181712695219464254218873561203838411485362628563332171346778184157808525739913136194247344581022903341636242765990015128099104447847709663892870277849956216606935586755936860594844960167275870224693600483318703837204300942;
            6'd37: xpb[142] = 1024'd59305907132998377505027632037830234361219972736239873134452321944695645301373630617525706542119440646439933122120541010194877689601917962108095334527143036799702320325969425697938895537189238838762322406767001814672610382215916775831395391023520864149393574943977217884090402442711110927474158064117569554949;
            6'd38: xpb[142] = 1024'd94440308862032047545379440310424141437117384736066811361905588771573066887169982501787231371543661828625647370679878181978270016575272592044843890870128265073664727515744604051296768171036841434758654798405904524897373054767940681384940825830434792712031213027359590808013529015197528254464997424397934808956;
            6'd39: xpb[142] = 1024'd5508014906940976186932321178203615768316369610158065461227000533473593135657195476033684986310208701368212211781721919182598502707406887426432322196782452413936460135948565067024401613367238309444789581657567388757774877099067813973507690954119272007848947696624905701830127513755312564337146958052705578632;
            6'd40: xpb[142] = 1024'd40642416635974646227284129450797522844213781609985003688680267360351014721453547360295209815734429883553926460341059090965990829680761517363180878539767680687898867325723743420382274247214840905441121973296470098982537549651091719527053125761033200570486585780007278625753254086241729891327986318333070832639;
            6'd41: xpb[142] = 1024'd75776818365008316267635937723391429920111193609811941916133534187228436307249899244556734645158651065739640708900396262749383156654116147299929434882752908961861274515498921773740146881062443501437454364935372809207300222203115625080598560567947129133124223863389651549676380658728147218318825678613436086646;
            6'd42: xpb[142] = 1024'd110911220094041986307987745995985336996008605609638880143586801014105857893046251128818259474582872247925354957459733434532775483627470777236677991225738137235823681705274100127098019514910046097433786756574275519432062894755139530634143995374861057695761861946772024473599507231214564545309665038893801340653;
            6'd43: xpb[142] = 1024'd21978926138950914949540626863764811327207590483730134242908212776006384141533464103064713089349419120667919798561577171737103969759605072618266422552392324576095414325478061142825652957240442972119921539825938383292464717086266663222710860498545536991579596616037339367416105729772348855181814572548572110329;
            6'd44: xpb[142] = 1024'd57113327867984584989892435136358718403105002483557072470361479602883805727329815987326237918773640302853634047120914343520496296732959702555014978895377552850057821515253239496183525591088045568116253931464841093517227389638290568776256295305459465554217234699419712291339232302258766182172653932828937364336;
            6'd45: xpb[142] = 1024'd92247729597018255030244243408952625479002414483384010697814746429761227313126167871587762748197861485039348295680251515303888623706314332491763535238362781124020228705028417849541398224935648164112586323103743803741990062190314474329801730112373394116854872782802085215262358874745183509163493293109302618343;
            6'd46: xpb[142] = 1024'd3315435641927183671797124276732099810201399357475264797136158191661753561613380845834216362964408357781913136782095252508217109838448627873351966565016968464291961325232378865269031667266045038798721106355406667602391884521441606918368595236057873412672607452067400109078957373302967819035642826764073388019;
            6'd47: xpb[142] = 1024'd38449837370960853712148932549326006886098811357302203024589425018539175147409732730095741192388629539967627385341432424291609436811803257810100522908002196738254368515007557218626904301113647634795053497994309377827154557073465512471914030042971801975310245535449773033002083945789385146026482187044438642026;
            6'd48: xpb[142] = 1024'd73584239099994523752500740821919913961996223357129141252042691845416596733206084614357266021812850722153341633900769596075001763785157887746849079250987425012216775704782735571984776934961250230791385889633212088051917229625489418025459464849885730537947883618832145956925210518275802473017321547324803896033;
            6'd49: xpb[142] = 1024'd108718640829028193792852549094513821037893635356956079479495958672294018319002436498618790851237071904339055882460106767858394090758512517683597635593972653286179182894557913925342649568808852826787718281272114798276679902177513323579004899656799659100585521702214518880848337090762219800008160907605169150040;
            6'd50: xpb[142] = 1024'd19786346873937122434405429962293295369092620231047333578817370434194544567489649472865244466003618777081620723561950505062722576890646813065186066920626840626450915514761874941070283011139249701473853064523777662137081724508640456167571764780484138396403256371479833774664935589320004109880310441259939919716;
            6'd51: xpb[142] = 1024'd54920748602970792474757238234887202444990032230874271806270637261071966153286001357126769295427839959267334972121287676846114903864001443001934623263612068900413322704537053294428155644986852297470185456162680372361844397060664361721117199587398066959040894454862206698588062161806421436871149801540305173723;
            6'd52: xpb[142] = 1024'd90055150332004462515109046507481109520887444230701210033723904087949387739082353241388294124852061141453049220680624848629507230837356072938683179606597297174375729894312231647786028278834454893466517847801583082586607069612688267274662634394311995521678532538244579622511188734292838763861989161820670427730;
            6'd53: xpb[142] = 1024'd1122856376913391156661927375260583852086429104792464133045315849849913987569566215634747739618608014195614061782468585833835716969490368320271610933251484514647462514516192663513661721164851768152652631053245946447008891943815399863229499517996474817496267207509894516327787232850623073734138695475441197406;
            6'd54: xpb[142] = 1024'd36257258105947061197013735647854490927983841104619402360498582676727335573365918099896272569042829196381328310341805757617228043942844998257020167276236712788609869704291371016871534355012454364148985022692148656671771564495839305416774934324910403380133905290892267440250913805337040400724978055755806451413;
            6'd55: xpb[142] = 1024'd71391659834980731237365543920448398003881253104446340587951849503604757159162269984157797398467050378567042558901142929400620370916199628193768723619221941062572276894066549370229406988860056960145317414331051366896534237047863210970320369131824331942771543374274640364174040377823457727715817416036171705420;
            6'd56: xpb[142] = 1024'd106526061564014401277717352193042305079778665104273278815405116330482178744958621868419322227891271560752756807460480101184012697889554258130517279962207169336534684083841727723587279622707659556141649805969954077121296909599887116523865803938738260505409181457657013288097166950309875054706656776316536959427;
            6'd57: xpb[142] = 1024'd17593767608923329919270233060821779410977649978364532914726528092382704993445834842665775842657818433495321648562323838388341184021688553512105711288861356676806416704045688739314913065038056430827784589221616940981698731931014249112432669062422739801226916126922328181913765448867659364578806309971307729103;
            6'd58: xpb[142] = 1024'd52728169337956999959622041333415686486875061978191471142179794919260126579242186726927300672082039615681035897121661010171733510995043183448854267631846584950768823893820867092672785698885659026824116980860519651206461404483038154665978103869336668363864554210304701105836892021354076691569645670251672983110;
            6'd59: xpb[142] = 1024'd87862571066990669999973849606009593562772473978018409369633061746137548165038538611188825501506260797866750145680998181955125837968397813385602823974831813224731231083596045446030658332733261622820449372499422361431224077035062060219523538676250596926502192293687074029760018593840494018560485030532038237117;
            6'd60: xpb[142] = 1024'd122996972796024340040325657878603500638669885977845347597086328573014969750834890495450350330930481980052464394240335353738518164941752443322351380317817041498693638273371223799388530966580864218816781764138325071655986749587085965773068973483164525489139830377069446953683145166326911345551324390812403491124;
            6'd61: xpb[142] = 1024'd34064678840933268681878538746382974969868870851936601696407740334915495999322103469696803945697028852795029235342179090942846651073886738703939811644471228838965370893575184815116164408911261093502916547389987935516388571918213098361635838606849004784957565046334761847499743664884695655423473924467174260800;
            6'd62: xpb[142] = 1024'd69199080569966938722230347018976882045766282851763539923861007161792917585118455353958328775121250034980743483901516262726238978047241368640688367987456457112927778083350363168474037042758863689499248939028890645741151244470237003915181273413762933347595203129717134771422870237371112982414313284747539514807;
            6'd63: xpb[142] = 1024'd104333482299000608762582155291570789121663694851590478151314273988670339170914807238219853604545471217166457732460853434509631305020595998577436924330441685386890185273125541521831909676606466285495581330667793355965913917022260909468726708220676861910232841213099507695345996809857530309405152645027904768814;
        endcase
    end

    always_comb begin
        case(flag[47][16:12])
            5'd0: xpb[143] = 1024'd0;
            5'd1: xpb[143] = 1024'd15401188343909537404135036159350263452862679725681732250635685750570865419402020212466307219312018089909022573562697171713959791152730293959025355657095872727161917893329502537559543118936863160181716113919456219826315739353388042057293573344361341206050575882364822589162595308415314619277302178682675538490;
            5'd2: xpb[143] = 1024'd30802376687819074808270072318700526905725359451363464501271371501141730838804040424932614438624036179818045147125394343427919582305460587918050711314191745454323835786659005075119086237873726320363432227838912439652631478706776084114587146688722682412101151764729645178325190616830629238554604357365351076980;
            5'd3: xpb[143] = 1024'd46203565031728612212405108478050790358588039177045196751907057251712596258206060637398921657936054269727067720688091515141879373458190881877076066971287618181485753679988507612678629356810589480545148341758368659478947218060164126171880720033084023618151727647094467767487785925245943857831906536048026615470;
            5'd4: xpb[143] = 1024'd61604753375638149616540144637401053811450718902726929002542743002283461677608080849865228877248072359636090294250788686855839164610921175836101422628383490908647671573318010150238172475747452640726864455677824879305262957413552168229174293377445364824202303529459290356650381233661258477109208714730702153960;
            5'd5: xpb[143] = 1024'd77005941719547687020675180796751317264313398628408661253178428752854327097010101062331536096560090449545112867813485858569798955763651469795126778285479363635809589466647512687797715594684315800908580569597281099131578696766940210286467866721806706030252879411824112945812976542076573096386510893413377692450;
            5'd6: xpb[143] = 1024'd92407130063457224424810216956101580717176078354090393503814114503425192516412121274797843315872108539454135441376183030283758746916381763754152133942575236362971507359977015225357258713621178961090296683516737318957894436120328252343761440066168047236303455294188935534975571850491887715663813072096053230940;
            5'd7: xpb[143] = 1024'd107808318407366761828945253115451844170038758079772125754449800253996057935814141487264150535184126629363158014938880201997718538069112057713177489599671109090133425253306517762916801832558042121272012797436193538784210175473716294401055013410529388442354031176553758124138167158907202334941115250778728769430;
            5'd8: xpb[143] = 1024'd123209506751276299233080289274802107622901437805453858005085486004566923355216161699730457754496144719272180588501577373711678329221842351672202845256766981817295343146636020300476344951494905281453728911355649758610525914827104336458348586754890729648404607058918580713300762467322516954218417429461404307920;
            5'd9: xpb[143] = 1024'd14543999411061095238416398029337938331065690405399906127589316690160893437309043002181693759150488499738053754606781110846574279533352311076068075897531813610766586470394305500405648878914562720325247416887866132072480803959595605550663590416022621587635279527166345272356829701809198556377029781518485362079;
            5'd10: xpb[143] = 1024'd29945187754970632642551434188688201783928370131081638378225002440731758856711063214648000978462506589647076328169478282560534070686082605035093431554627686337928504363723808037965191997851425880506963530807322351898796543312983647607957163760383962793685855409531167861519425010224513175654331960201160900569;
            5'd11: xpb[143] = 1024'd45346376098880170046686470348038465236791049856763370628860688191302624276113083427114308197774524679556098901732175454274493861838812898994118787211723559065090422257053310575524735116788289040688679644726778571725112282666371689665250737104745303999736431291895990450682020318639827794931634138883836439059;
            5'd12: xpb[143] = 1024'd60747564442789707450821506507388728689653729582445102879496373941873489695515103639580615417086542769465121475294872625988453652991543192953144142868819431792252340150382813113084278235725152200870395758646234791551428022019759731722544310449106645205787007174260813039844615627055142414208936317566511977549;
            5'd13: xpb[143] = 1024'd76148752786699244854956542666738992142516409308126835130132059692444355114917123852046922636398560859374144048857569797702413444144273486912169498525915304519414258043712315650643821354662015361052111872565691011377743761373147773779837883793467986411837583056625635629007210935470457033486238496249187516039;
            5'd14: xpb[143] = 1024'd91549941130608782259091578826089255595379089033808567380767745443015220534319144064513229855710578949283166622420266969416373235297003780871194854183011177246576175937041818188203364473598878521233827986485147231204059500726535815837131457137829327617888158938990458218169806243885771652763540674931863054529;
            5'd15: xpb[143] = 1024'd106951129474518319663226614985439519048241768759490299631403431193586085953721164276979537075022597039192189195982964141130333026449734074830220209840107049973738093830371320725762907592535741681415544100404603451030375240079923857894425030482190668823938734821355280807332401552301086272040842853614538593019;
            5'd16: xpb[143] = 1024'd122352317818427857067361651144789782501104448485172031882039116944156951373123184489445844294334615129101211769545661312844292817602464368789245565497202922700900011723700823263322450711472604841597260214324059670856690979433311899951718603826552010029989310703720103396494996860716400891318145032297214131509;
            5'd17: xpb[143] = 1024'd13686810478212653072697759899325613209268701085118080004542947629750921455216065791897080298988958909567084935650865049979188767913974328193110796137967754494371255047459108463251754638892262280468778719856276044318645868565803169044033607487683901969219983171967867955551064095203082493476757384354295185668;
            5'd18: xpb[143] = 1024'd29087998822122190476832796058675876662131380810799812255178633380321786874618086004363387518300976999476107509213562221693148559066704622152136151795063627221533172940788611000811297757829125440650494833775732264144961607919191211101327180832045243175270559054332690544713659403618397112754059563036970724158;
            5'd19: xpb[143] = 1024'd44489187166031727880967832218026140114994060536481544505814319130892652294020106216829694737612995089385130082776259393407108350219434916111161507452159499948695090834118113538370840876765988600832210947695188483971277347272579253158620754176406584381321134936697513133876254712033711732031361741719646262648;
            5'd20: xpb[143] = 1024'd59890375509941265285102868377376403567856740262163276756450004881463517713422126429296001956925013179294152656338956565121068141372165210070186863109255372675857008727447616075930383995702851761013927061614644703797593086625967295215914327520767925587371710819062335723038850020449026351308663920402321801138;
            5'd21: xpb[143] = 1024'd75291563853850802689237904536726667020719419987845009007085690632034383132824146641762309176237031269203175229901653736835027932524895504029212218766351245403018926620777118613489927114639714921195643175534100923623908825979355337273207900865129266793422286701427158312201445328864340970585966099084997339628;
            5'd22: xpb[143] = 1024'd90692752197760340093372940696076930473582099713526741257721376382605248552226166854228616395549049359112197803464350908548987723677625797988237574423447118130180844514106621151049470233576578081377359289453557143450224565332743379330501474209490607999472862583791980901364040637279655589863268277767672878118;
            5'd23: xpb[143] = 1024'd106093940541669877497507976855427193926444779439208473508357062133176113971628187066694923614861067449021220377027048080262947514830356091947262930080542990857342762407436123688609013352513441241559075403373013363276540304686131421387795047553851949205523438466156803490526635945694970209140570456450348416608;
            5'd24: xpb[143] = 1024'd121495128885579414901643013014777457379307459164890205758992747883746979391030207279161230834173085538930242950589745251976907305983086385906288285737638863584504680300765626226168556471450304401740791517292469583102856044039519463445088620898213290411574014348521626079689231254110284828417872635133023955098;
            5'd25: xpb[143] = 1024'd12829621545364210906979121769313288087471711764836253881496578569340949473123088581612466838827429319396116116694948989111803256294596345310153516378403695377975923624523911426097860398869961840612310022824685956564810933172010732537403624559345182350804686816769390638745298488596966430576484987190105009257;
            5'd26: xpb[143] = 1024'd28230809889273748311114157928663551540334391490517986132132264319911814892525108794078774058139447409305138690257646160825763047447326639269178872035499568105137841517853413963657403517806825000794026136744142176391126672525398774594697197903706523556855262699134213227907893797012281049853787165872780547747;
            5'd27: xpb[143] = 1024'd43631998233183285715249194088013814993197071216199718382767950070482680311927129006545081277451465499214161263820343332539722838600056933228204227692595440832299759411182916501216946636743688160975742250663598396217442411878786816651990771248067864762905838581499035817070489105427595669131089344555456086237;
            5'd28: xpb[143] = 1024'd59033186577092823119384230247364078446059750941881450633403635821053545731329149219011388496763483589123183837383040504253682629752787227187229583349691313559461677304512419038776489755680551321157458364583054616043758151232174858709284344592429205968956414463863858406233084413842910288408391523238131624727;
            5'd29: xpb[143] = 1024'd74434374921002360523519266406714341898922430667563182884039321571624411150731169431477695716075501679032206410945737675967642420905517521146254939006787186286623595197841921576336032874617414481339174478502510835870073890585562900766577917936790547175006990346228680995395679722258224907685693701920807163217;
            5'd30: xpb[143] = 1024'd89835563264911897927654302566064605351785110393244915134675007322195276570133189643944002935387519768941228984508434847681602212058247815105280294663883059013785513091171424113895575993554277641520890592421967055696389629938950942823871491281151888381057566228593503584558275030673539526962995880603482701707;
            5'd31: xpb[143] = 1024'd105236751608821435331789338725414868804647790118926647385310693072766141989535209856410310154699537858850251558071132019395562003210978109064305650320978931740947430984500926651455119112491140801702606706341423275522705369292338984881165064625513229587108142110958326173720870339088854146240298059286158240197;
        endcase
    end

    always_comb begin
        case(flag[48][5:0])
            6'd0: xpb[144] = 1024'd0;
            6'd1: xpb[144] = 1024'd122352317818427857067361651144789782501104448485172031882039116944156951373123184489445844294334615129101211769545661312844292817602464368789245565497202922700900011723700823263322450711472604841597260214324059670856690979433311899951718603826552010029989310703720103396494996860716400891318145032297214131509;
            6'd2: xpb[144] = 1024'd120637939952730972735924374884765132257510469844608379635946378823337007408937230068876617374011555948759274131633829191109521794363708403023331005978074804468109348877830429189014662231428003961884322820260879495349021108645727026938458637969874570793158717993323148762883465647504168765517600237968833778687;
            6'd3: xpb[144] = 1024'd118923562087034088404487098624740482013916491204044727389853640702517063444751275648307390453688496768417336493721997069374750771124952437257416446458946686235318686031960035114706873751383403082171385426197699319841351237858142153925198672113197131556328125282926194129271934434291936639717055443640453425865;
            6'd4: xpb[144] = 1024'd117209184221337204073049822364715831770322512563481075143760902581697119480565321227738163533365437588075398855810164947639979747886196471491501886939818568002528023186089641040399085271338802202458448032134519144333681367070557280911938706256519692319497532572529239495660403221079704513916510649312073073043;
            6'd5: xpb[144] = 1024'd115494806355640319741612546104691181526728533922917422897668164460877175516379366807168936613042378407733461217898332825905208724647440505725587327420690449769737360340219246966091296791294201322745510638071338968826011496282972407898678740399842253082666939862132284862048872007867472388115965854983692720221;
            6'd6: xpb[144] = 1024'd113780428489943435410175269844666531283134555282353770651575426340057231552193412386599709692719319227391523579986500704170437701408684539959672767901562331536946697494348852891783508311249600443032573244008158793318341625495387534885418774543164813845836347151735330228437340794655240262315421060655312367399;
            6'd7: xpb[144] = 1024'd112066050624246551078737993584641881039540576641790118405482688219237287588007457966030482772396260047049585942074668582435666678169928574193758208382434213304156034648478458817475719831204999563319635849944978617810671754707802661872158808686487374609005754441338375594825809581443008136514876266326932014577;
            6'd8: xpb[144] = 1024'd110351672758549666747300717324617230795946598001226466159389950098417343623821503545461255852073200866707648304162836460700895654931172608427843648863306095071365371802608064743167931351160398683606698455881798442303001883920217788858898842829809935372175161730941420961214278368230776010714331471998551661755;
            6'd9: xpb[144] = 1024'd108637294892852782415863441064592580552352619360662813913297211977597399659635549124892028931750141686365710666251004338966124631692416642661929089344177976838574708956737670668860142871115797803893761061818618266795332013132632915845638876973132496135344569020544466327602747155018543884913786677670171308933;
            6'd10: xpb[144] = 1024'd106922917027155898084426164804567930308758640720099161667204473856777455695449594704322802011427082506023773028339172217231353608453660676896014529825049858605784046110867276594552354391071196924180823667755438091287662142345048042832378911116455056898513976310147511693991215941806311759113241883341790956111;
            6'd11: xpb[144] = 1024'd105208539161459013752988888544543280065164662079535509421111735735957511731263640283753575091104023325681835390427340095496582585214904711130099970305921740372993383264996882520244565911026596044467886273692257915779992271557463169819118945259777617661683383599750557060379684728594079633312697089013410603289;
            6'd12: xpb[144] = 1024'd103494161295762129421551612284518629821570683438971857175018997615137567767077685863184348170780964145339897752515507973761811561976148745364185410786793622140202720419126488445936777430981995164754948879629077740272322400769878296805858979403100178424852790889353602426768153515381847507512152294685030250467;
            6'd13: xpb[144] = 1024'd101779783430065245090114336024493979577976704798408204928926259494317623802891731442615121250457904964997960114603675852027040538737392779598270851267665503907412057573256094371628988950937394285042011485565897564764652529982293423792599013546422739188022198178956647793156622302169615381711607500356649897645;
            6'd14: xpb[144] = 1024'd100065405564368360758677059764469329334382726157844552682833521373497679838705777022045894330134845784656022476691843730292269515498636813832356291748537385674621394727385700297321200470892793405329074091502717389256982659194708550779339047689745299951191605468559693159545091088957383255911062706028269544823;
            6'd15: xpb[144] = 1024'd98351027698671476427239783504444679090788747517280900436740783252677735874519822601476667409811786604314084838780011608557498492259880848066441732229409267441830731881515306223013411990848192525616136697439537213749312788407123677766079081833067860714361012758162738525933559875745151130110517911699889192001;
            6'd16: xpb[144] = 1024'd96636649832974592095802507244420028847194768876717248190648045131857791910333868180907440489488727423972147200868179486822727469021124882300527172710281149209040069035644912148705623510803591645903199303376357038241642917619538804752819115976390421477530420047765783892322028662532919004309973117371508839179;
            6'd17: xpb[144] = 1024'd94922271967277707764365230984395378603600790236153595944555307011037847946147913760338213569165668243630209562956347365087956445782368916534612613191153030976249406189774518074397835030758990766190261909313176862733973046831953931739559150119712982240699827337368829258710497449320686878509428323043128486357;
            6'd18: xpb[144] = 1024'd93207894101580823432927954724370728360006811595589943698462568890217903981961959339768986648842609063288271925044515243353185422543612950768698053672024912743458743343904124000090046550714389886477324515249996687226303176044369058726299184263035543003869234626971874625098966236108454752708883528714748133535;
            6'd19: xpb[144] = 1024'd91493516235883939101490678464346078116412832955026291452369830769397960017776004919199759728519549882946334287132683121618414399304856985002783494152896794510668080498033729925782258070669789006764387121186816511718633305256784185713039218406358103767038641916574919991487435022896222626908338734386367780713;
            6'd20: xpb[144] = 1024'd89779138370187054770053402204321427872818854314462639206277092648578016053590050498630532808196490702604396649220850999883643376066101019236868934633768676277877417652163335851474469590625188127051449727123636336210963434469199312699779252549680664530208049206177965357875903809683990501107793940057987427891;
            6'd21: xpb[144] = 1024'd88064760504490170438616125944296777629224875673898986960184354527758072089404096078061305887873431522262459011309018878148872352827345053470954375114640558045086754806292941777166681110580587247338512333060456160703293563681614439686519286693003225293377456495781010724264372596471758375307249145729607075069;
            6'd22: xpb[144] = 1024'd86350382638793286107178849684272127385630897033335334714091616406938128125218141657492078967550372341920521373397186756414101329588589087705039815595512439812296091960422547702858892630535986367625574938997275985195623692894029566673259320836325786056546863785384056090652841383259526249506704351401226722247;
            6'd23: xpb[144] = 1024'd84636004773096401775741573424247477142036918392771682467998878286118184161032187236922852047227313161578583735485354634679330306349833121939125256076384321579505429114552153628551104150491385487912637544934095809687953822106444693659999354979648346819716271074987101457041310170047294123706159557072846369425;
            6'd24: xpb[144] = 1024'd82921626907399517444304297164222826898442939752208030221906140165298240196846232816353625126904253981236646097573522512944559283111077156173210696557256203346714766268681759554243315670446784608199700150870915634180283951318859820646739389122970907582885678364590146823429778956835061997905614762744466016603;
            6'd25: xpb[144] = 1024'd81207249041702633112867020904198176654848961111644377975813402044478296232660278395784398206581194800894708459661690391209788259872321190407296137038128085113924103422811365479935527190402183728486762756807735458672614080531274947633479423266293468346055085654193192189818247743622829872105069968416085663781;
            6'd26: xpb[144] = 1024'd79492871176005748781429744644173526411254982471080725729720663923658352268474323975215171286258135620552770821749858269475017236633565224641381577518999966881133440576940971405627738710357582848773825362744555283164944209743690074620219457409616029109224492943796237556206716530410597746304525174087705310959;
            6'd27: xpb[144] = 1024'd77778493310308864449992468384148876167661003830517073483627925802838408304288369554645944365935076440210833183838026147740246213394809258875467017999871848648342777731070577331319950230312981969060887968681375107657274338956105201606959491552938589872393900233399282922595185317198365620503980379759324958137;
            6'd28: xpb[144] = 1024'd76064115444611980118555192124124225924067025189953421237535187682018464340102415134076717445612017259868895545926194026005475190156053293109552458480743730415552114885200183257012161750268381089347950574618194932149604468168520328593699525696261150635563307523002328288983654103986133494703435585430944605315;
            6'd29: xpb[144] = 1024'd74349737578915095787117915864099575680473046549389768991442449561198520375916460713507490525288958079526957908014361904270704166917297327343637898961615612182761452039329789182704373270223780209635013180555014756641934597380935455580439559839583711398732714812605373655372122890773901368902890791102564252493;
            6'd30: xpb[144] = 1024'd72635359713218211455680639604074925436879067908826116745349711440378576411730506292938263604965898899185020270102529782535933143678541361577723339442487493949970789193459395108396584790179179329922075786491834581134264726593350582567179593982906272161902122102208419021760591677561669243102345996774183899671;
            6'd31: xpb[144] = 1024'd70920981847521327124243363344050275193285089268262464499256973319558632447544551872369036684642839718843082632190697660801162120439785395811808779923359375717180126347589001034088796310134578450209138392428654405626594855805765709553919628126228832925071529391811464388149060464349437117301801202445803546849;
            6'd32: xpb[144] = 1024'd69206603981824442792806087084025624949691110627698812253164235198738688483358597451799809764319780538501144994278865539066391097201029430045894220404231257484389463501718606959781007830089977570496200998365474230118924985018180836540659662269551393688240936681414509754537529251137204991501256408117423194027;
            6'd33: xpb[144] = 1024'd67492226116127558461368810824000974706097131987135160007071497077918744519172643031230582843996721358159207356367033417331620073962273464279979660885103139251598800655848212885473219350045376690783263604302294054611255114230595963527399696412873954451410343971017555120925998037924972865700711613789042841205;
            6'd34: xpb[144] = 1024'd65777848250430674129931534563976324462503153346571507760978758957098800554986688610661355923673662177817269718455201295596849050723517498514065101365975021018808137809977818811165430870000775811070326210239113879103585243443011090514139730556196515214579751260620600487314466824712740739900166819460662488383;
            6'd35: xpb[144] = 1024'd64063470384733789798494258303951674218909174706007855514886020836278856590800734190092129003350602997475332080543369173862078027484761532748150541846846902786017474964107424736857642389956174931357388816175933703595915372655426217500879764699519075977749158550223645853702935611500508614099622025132282135561;
            6'd36: xpb[144] = 1024'd62349092519036905467056982043927023975315196065444203268793282715458912626614779769522902083027543817133394442631537052127307004246005566982235982327718784553226812118237030662549853909911574051644451422112753528088245501867841344487619798842841636740918565839826691220091404398288276488299077230803901782739;
            6'd37: xpb[144] = 1024'd60634714653340021135619705783902373731721217424880551022700544594638968662428825348953675162704484636791456804719704930392535981007249601216321422808590666320436149272366636588242065429866973171931514028049573352580575631080256471474359832986164197504087973129429736586479873185076044362498532436475521429917;
            6'd38: xpb[144] = 1024'd58920336787643136804182429523877723488127238784316898776607806473819024698242870928384448242381425456449519166807872808657764957768493635450406863289462548087645486426496242513934276949822372292218576633986393177072905760292671598461099867129486758267257380419032781952868341971863812236697987642147141077095;
            6'd39: xpb[144] = 1024'd57205958921946252472745153263853073244533260143753246530515068352999080734056916507815221322058366276107581528896040686922993934529737669684492303770334429854854823580625848439626488469777771412505639239923213001565235889505086725447839901272809319030426787708635827319256810758651580110897442847818760724273;
            6'd40: xpb[144] = 1024'd55491581056249368141307877003828423000939281503189594284422330232179136769870962087245994401735307095765643890984208565188222911290981703918577744251206311622064160734755454365318699989733170532792701845860032826057566018717501852434579935416131879793596194998238872685645279545439347985096898053490380371451;
            6'd41: xpb[144] = 1024'd53777203190552483809870600743803772757345302862625942038329592111359192805685007666676767481412247915423706253072376443453451888052225738152663184732078193389273497888885060291010911509688569653079764451796852650549896147929916979421319969559454440556765602287841918052033748332227115859296353259162000018629;
            6'd42: xpb[144] = 1024'd52062825324855599478433324483779122513751324222062289792236853990539248841499053246107540561089188735081768615160544321718680864813469772386748625212950075156482835043014666216703123029643968773366827057733672475042226277142332106408060003702777001319935009577444963418422217119014883733495808464833619665807;
            6'd43: xpb[144] = 1024'd50348447459158715146996048223754472270157345581498637546144115869719304877313098825538313640766129554739830977248712199983909841574713806620834065693821956923692172197144272142395334549599367893653889663670492299534556406354747233394800037846099562083104416867048008784810685905802651607695263670505239312985;
            6'd44: xpb[144] = 1024'd48634069593461830815558771963729822026563366940934985300051377748899360913127144404969086720443070374397893339336880078249138818335957840854919506174693838690901509351273878068087546069554767013940952269607312124026886535567162360381540071989422122846273824156651054151199154692590419481894718876176858960163;
            6'd45: xpb[144] = 1024'd46919691727764946484121495703705171782969388300371333053958639628079416948941189984399859800120011194055955701425047956514367795097201875089004946655565720458110846505403483993779757589510166134228014875544131948519216664779577487368280106132744683609443231446254099517587623479378187356094174081848478607341;
            6'd46: xpb[144] = 1024'd45205313862068062152684219443680521539375409659807680807865901507259472984755235563830632879796952013714018063513215834779596771858445909323090387136437602225320183659533089919471969109465565254515077481480951773011546793991992614355020140276067244372612638735857144883976092266165955230293629287520098254519;
            6'd47: xpb[144] = 1024'd43490935996371177821246943183655871295781431019244028561773163386439529020569281143261405959473892833372080425601383713044825748619689943557175827617309483992529520813662695845164180629420964374802140087417771597503876923204407741341760174419389805135782046025460190250364561052953723104493084493191717901697;
            6'd48: xpb[144] = 1024'd41776558130674293489809666923631221052187452378680376315680425265619585056383326722692179039150833653030142787689551591310054725380933977791261268098181365759738857967792301770856392149376363495089202693354591421996207052416822868328500208562712365898951453315063235616753029839741490978692539698863337548875;
            6'd49: xpb[144] = 1024'd40062180264977409158372390663606570808593473738116724069587687144799641092197372302122952118827774472688205149777719469575283702142178012025346708579053247526948195121921907696548603669331762615376265299291411246488537181629237995315240242706034926662120860604666280983141498626529258852891994904534957196053;
            6'd50: xpb[144] = 1024'd38347802399280524826935114403581920564999495097553071823494949023979697128011417881553725198504715292346267511865887347840512678903422046259432149059925129294157532276051513622240815189287161735663327905228231070980867310841653122301980276849357487425290267894269326349529967413317026727091450110206576843231;
            6'd51: xpb[144] = 1024'd36633424533583640495497838143557270321405516456989419577402210903159753163825463460984498278181656112004329873954055226105741655664666080493517589540797011061366869430181119547933026709242560855950390511165050895473197440054068249288720310992680048188459675183872371715918436200104794601290905315878196490409;
            6'd52: xpb[144] = 1024'd34919046667886756164060561883532620077811537816425767331309472782339809199639509040415271357858596931662392236042223104370970632425910114727603030021668892828576206584310725473625238229197959976237453117101870719965527569266483376275460345136002608951629082473475417082306904986892562475490360521549816137587;
            6'd53: xpb[144] = 1024'd33204668802189871832623285623507969834217559175862115085216734661519865235453554619846044437535537751320454598130390982636199609187154148961688470502540774595785543738440331399317449749153359096524515723038690544457857698478898503262200379279325169714798489763078462448695373773680330349689815727221435784765;
            6'd54: xpb[144] = 1024'd31490290936492987501186009363483319590623580535298462839123996540699921271267600199276817517212478570978516960218558860901428585948398183195773910983412656362994880892569937325009661269108758216811578328975510368950187827691313630248940413422647730477967897052681507815083842560468098223889270932893055431943;
            6'd55: xpb[144] = 1024'd29775913070796103169748733103458669347029601894734810593031258419879977307081645778707590596889419390636579322306726739166657562709642217429859351464284538130204218046699543250701872789064157337098640934912330193442517956903728757235680447565970291241137304342284553181472311347255866098088726138564675079121;
            6'd56: xpb[144] = 1024'd28061535205099218838311456843434019103435623254171158346938520299060033342895691358138363676566360210294641684394894617431886539470886251663944791945156419897413555200829149176394084309019556457385703540849150017934848086116143884222420481709292852004306711631887598547860780134043633972288181344236294726299;
            6'd57: xpb[144] = 1024'd26347157339402334506874180583409368859841644613607506100845782178240089378709736937569136756243301029952704046483062495697115516232130285898030232426028301664622892354958755102086295828974955577672766146785969842427178215328559011209160515852615412767476118921490643914249248920831401846487636549907914373477;
            6'd58: xpb[144] = 1024'd24632779473705450175436904323384718616247665973043853854753044057420145414523782516999909835920241849610766408571230373962344492993374320132115672906900183431832229509088361027778507348930354697959828752722789666919508344540974138195900549995937973530645526211093689280637717707619169720687091755579534020655;
            6'd59: xpb[144] = 1024'd22918401608008565843999628063360068372653687332480201608660305936600201450337828096430682915597182669268828770659398252227573469754618354366201113387772065199041566663217966953470718868885753818246891358659609491411838473753389265182640584139260534293814933500696734647026186494406937594886546961251153667833;
            6'd60: xpb[144] = 1024'd21204023742311681512562351803335418129059708691916549362567567815780257486151873675861455995274123488926891132747566130492802446515862388600286553868643946966250903817347572879162930388841152938533953964596429315904168602965804392169380618282583095056984340790299780013414655281194705469086002166922773315011;
            6'd61: xpb[144] = 1024'd19489645876614797181125075543310767885465730051352897116474829694960313521965919255292229074951064308584953494835734008758031423277106422834371994349515828733460240971477178804855141908796552058821016570533249140396498732178219519156120652425905655820153748079902825379803124067982473343285457372594392962189;
            6'd62: xpb[144] = 1024'd17775268010917912849687799283286117641871751410789244870382091574140369557779964834723002154628005128243015856923901887023260400038350457068457434830387710500669578125606784730547353428751951179108079176470068964888828861390634646142860686569228216583323155369505870746191592854770241217484912578266012609367;
            6'd63: xpb[144] = 1024'd16060890145221028518250523023261467398277772770225592624289353453320425593594010414153775234304945947901078219012069765288489376799594491302542875311259592267878915279736390656239564948707350299395141782406888789381158990603049773129600720712550777346492562659108916112580061641558009091684367783937632256545;
        endcase
    end

    always_comb begin
        case(flag[48][11:6])
            6'd0: xpb[145] = 1024'd0;
            6'd1: xpb[145] = 1024'd14346512279524144186813246763236817154683794129661940378196615332500481629408055993584548313981886767559140581100237643553718353560838525536628315792131474035088252433865996581931776468662749419682204388343708613873489119815464900116340754855873338109661969948711961478968530428345776965883822989609251903723;
            6'd2: xpb[145] = 1024'd28693024559048288373626493526473634309367588259323880756393230665000963258816111987169096627963773535118281162200475287107436707121677051073256631584262948070176504867731993163863552937325498839364408776687417227746978239630929800232681509711746676219323939897423922957937060856691553931767645979218503807446;
            6'd3: xpb[145] = 1024'd43039536838572432560439740289710451464051382388985821134589845997501444888224167980753644941945660302677421743300712930661155060682515576609884947376394422105264757301597989745795329405988248259046613165031125841620467359446394700349022264567620014328985909846135884436905591285037330897651468968827755711169;
            6'd4: xpb[145] = 1024'd57386049118096576747252987052947268618735176518647761512786461330001926517632223974338193255927547070236562324400950574214873414243354102146513263168525896140353009735463986327727105874650997678728817553374834455493956479261859600465363019423493352438647879794847845915874121713383107863535291958437007614892;
            6'd5: xpb[145] = 1024'd71732561397620720934066233816184085773418970648309701890983076662502408147040279967922741569909433837795702905501188217768591767804192627683141578960657370175441262169329982909658882343313747098411021941718543069367445599077324500581703774279366690548309849743559807394842652141728884829419114948046259518615;
            6'd6: xpb[145] = 1024'd86079073677144865120879480579420902928102764777971642269179691995002889776448335961507289883891320605354843486601425861322310121365031153219769894752788844210529514603195979491590658811976496518093226330062251683240934718892789400698044529135240028657971819692271768873811182570074661795302937937655511422338;
            6'd7: xpb[145] = 1024'd100425585956669009307692727342657720082786558907633582647376307327503371405856391955091838197873207372913984067701663504876028474925869678756398210544920318245617767037061976073522435280639245937775430718405960297114423838708254300814385283991113366767633789640983730352779712998420438761186760927264763326061;
            6'd8: xpb[145] = 1024'd114772098236193153494505974105894537237470353037295523025572922660003853035264447948676386511855094140473124648801901148429746828486708204293026526337051792280706019470927972655454211749301995357457635106749668910987912958523719200930726038846986704877295759589695691831748243426766215727070583916874015229784;
            6'd9: xpb[145] = 1024'd5051914831592556282520293464316921647455720041221779275637682927527439327363365032245863611179306598589115822444645357404401341206326395274494717112852225382103597335222751899755749026447539055829641886706137678497041228118287328082088224019630593720137826124290595280610245781183359675835717079857672649176;
            6'd10: xpb[145] = 1024'd19398427111116700469333540227553738802139514170883719653834298260027920956771421025830411925161193366148256403544883000958119694767164920811123032904983699417191849769088748481687525495110288475511846275049846292370530347933752228198428978875503931829799796073002556759578776209529136641719540069466924552899;
            6'd11: xpb[145] = 1024'd33744939390640844656146786990790555956823308300545660032030913592528402586179477019414960239143080133707396984645120644511838048328003446347751348697115173452280102202954745063619301963773037895194050663393554906244019467749217128314769733731377269939461766021714518238547306637874913607603363059076176456622;
            6'd12: xpb[145] = 1024'd48091451670164988842960033754027373111507102430207600410227528925028884215587533012999508553124966901266537565745358288065556401888841971884379664489246647487368354636820741645551078432435787314876255051737263520117508587564682028431110488587250608049123735970426479717515837066220690573487186048685428360345;
            6'd13: xpb[145] = 1024'd62437963949689133029773280517264190266190896559869540788424144257529365844995589006584056867106853668825678146845595931619274755449680497421007980281378121522456607070686738227482854901098536734558459440080972133990997707380146928547451243443123946158785705919138441196484367494566467539371009038294680264068;
            6'd14: xpb[145] = 1024'd76784476229213277216586527280501007420874690689531481166620759590029847474403645000168605181088740436384818727945833575172993109010519022957636296073509595557544859504552734809414631369761286154240663828424680747864486827195611828663791998298997284268447675867850402675452897922912244505254832027903932167791;
            6'd15: xpb[145] = 1024'd91130988508737421403399774043737824575558484819193421544817374922530329103811700993753153495070627203943959309046071218726711462571357548494264611865641069592633111938418731391346407838424035573922868216768389361737975947011076728780132753154870622378109645816562364154421428351258021471138655017513184071514;
            6'd16: xpb[145] = 1024'd105477500788261565590213020806974641730242278948855361923013990255030810733219756987337701809052513971503099890146308862280429816132196074030892927657772543627721364372284727973278184307086784993605072605112097975611465066826541628896473508010743960487771615765274325633389958779603798437022478007122435975237;
            6'd17: xpb[145] = 1024'd119824013067785709777026267570211458884926073078517302301210605587531292362627812980922250123034400739062240471246546505834148169693034599567521243449904017662809616806150724555209960775749534413287276993455806589484954186642006529012814262866617298597433585713986287112358489207949575402906300996731687878960;
            6'd18: xpb[145] = 1024'd10103829663185112565040586928633843294911440082443558551275365855054878654726730064491727222358613197178231644889290714808802682412652790548989434225704450764207194670445503799511498052895078111659283773412275356994082456236574656164176448039261187440275652248581190561220491562366719351671434159715345298352;
            6'd19: xpb[145] = 1024'd24450341942709256751853833691870660449595234212105498929471981187555360284134786058076275536340499964737372225989528358362521035973491316085617750017835924799295447104311500381443274521557827531341488161755983970867571576052039556280517202895134525549937622197293152040189021990712496317555257149324597202075;
            6'd20: xpb[145] = 1024'd38796854222233400938667080455107477604279028341767439307668596520055841913542842051660823850322386732296512807089766001916239389534329841622246065809967398834383699538177496963375050990220576951023692550099692584741060695867504456396857957751007863659599592146005113519157552419058273283439080138933849105798;
            6'd21: xpb[145] = 1024'd53143366501757545125480327218344294758962822471429379685865211852556323542950898045245372164304273499855653388190003645469957743095168367158874381602098872869471951972043493545306827458883326370705896938443401198614549815682969356513198712606881201769261562094717074998126082847404050249322903128543101009521;
            6'd22: xpb[145] = 1024'd67489878781281689312293573981581111913646616601091320064061827185056805172358954038829920478286160267414793969290241289023676096656006892695502697394230346904560204405909490127238603927546075790388101326787109812488038935498434256629539467462754539878923532043429036477094613275749827215206726118152352913244;
            6'd23: xpb[145] = 1024'd81836391060805833499106820744817929068330410730753260442258442517557286801767010032414468792268047034973934550390478932577394450216845418232131013186361820939648456839775486709170380396208825210070305715130818426361528055313899156745880222318627877988585501992140997956063143704095604181090549107761604816967;
            6'd24: xpb[145] = 1024'd96182903340329977685920067508054746223014204860415200820455057850057768431175066025999017106249933802533075131490716576131112803777683943768759328978493294974736709273641483291102156864871574629752510103474527040235017175129364056862220977174501216098247471940852959435031674132441381146974372097370856720690;
            6'd25: xpb[145] = 1024'd110529415619854121872733314271291563377697998990077141198651673182558250060583122019583565420231820570092215712590954219684831157338522469305387644770624769009824961707507479873033933333534324049434714491818235654108506294944828956978561732030374554207909441889564920914000204560787158112858195086980108624413;
            6'd26: xpb[145] = 1024'd809232215253524660747633629713947787683365994003397448716433450081836352682039103153042519556033028208206886233698428659485670058140660286855835546425202111222539571802259117335470610679867747806721271774704421617634564539397084129923917203018443050751508424159824362862206915204302061623328249963766043805;
            6'd27: xpb[145] = 1024'd15155744494777668847560880392950764942367160123665337826913048782582317982090095096737590833537919795767347467333936072213204023618979185823484151338556676146310792005668255699267247079342617167488925660118413035491123684354861984246264672058891781160413478372871785841830737343550079027507151239573017947528;
            6'd28: xpb[145] = 1024'd29502256774301813034374127156187582097050954253327278205109664115082799611498151090322139147519806563326488048434173715766922377179817711360112467130688150181399044439534252281199023548005366587171130048462121649364612804170326884362605426914765119270075448321583747320799267771895855993390974229182269851251;
            6'd29: xpb[145] = 1024'd43848769053825957221187373919424399251734748382989218583306279447583281240906207083906687461501693330885628629534411359320640730740656236896740782922819624216487296873400248863130800016668116006853334436805830263238101923985791784478946181770638457379737418270295708799767798200241632959274797218791521754974;
            6'd30: xpb[145] = 1024'd58195281333350101408000620682661216406418542512651158961502894780083762870314263077491235775483580098444769210634649002874359084301494762433369098714951098251575549307266245445062576485330865426535538825149538877111591043801256684595286936626511795489399388219007670278736328628587409925158620208400773658697;
            6'd31: xpb[145] = 1024'd72541793612874245594813867445898033561102336642313099339699510112584244499722319071075784089465466866003909791734886646428077437862333287969997414507082572286663801741132242026994352953993614846217743213493247490985080163616721584711627691482385133599061358167719631757704859056933186891042443198010025562420;
            6'd32: xpb[145] = 1024'd86888305892398389781627114209134850715786130771975039717896125445084726129130375064660332403447353633563050372835124289981795791423171813506625730299214046321752054174998238608926129422656364265899947601836956104858569283432186484827968446338258471708723328116431593236673389485278963856926266187619277466143;
            6'd33: xpb[145] = 1024'd101234818171922533968440360972371667870469924901636980096092740777585207758538431058244880717429240401122190953935361933535514144984010339043254046091345520356840306608864235190857905891319113685582151990180664718732058403247651384944309201194131809818385298065143554715641919913624740822810089177228529369866;
            6'd34: xpb[145] = 1024'd115581330451446678155253607735608485025153719031298920474289356110085689387946487051829429031411127168681331535035599577089232498544848864579882361883476994391928559042730231772789682359981863105264356378524373332605547523063116285060649956050005147928047268013855516194610450341970517788693912166837781273589;
            6'd35: xpb[145] = 1024'd5861147046846080943267927094030869435139086035225176724354116377609275680045404135398906130735339626797322708678343786063887011264467055561350552659277427493326136907025011017091219637127406803636363158480842100114675792657684412212012141222649036770889334548450419643472452696387661737459045329821438692981;
            6'd36: xpb[145] = 1024'd20207659326370225130081173857267686589822880164887117102550731710109757309453460128983454444717226394356463289778581429617605364825305581097978868451408901528414389340891007599022996105790156223318567546824550713988164912473149312328352896078522374880551304497162381122440983124733438703342868319430690596704;
            6'd37: xpb[145] = 1024'd34554171605894369316894420620504503744506674294549057480747347042610238938861516122568002758699113161915603870878819073171323718386144106634607184243540375563502641774757004180954772574452905643000771935168259327861654032288614212444693650934395712990213274445874342601409513553079215669226691309039942500427;
            6'd38: xpb[145] = 1024'd48900683885418513503707667383741320899190468424210997858943962375110720568269572116152551072680999929474744451979056716725042071946982632171235500035671849598590894208623000762886549043115655062682976323511967941735143152104079112561034405790269051099875244394586304080378043981424992635110514298649194404150;
            6'd39: xpb[145] = 1024'd63247196164942657690520914146978138053874262553872938237140577707611202197677628109737099386662886697033885033079294360278760425507821157707863815827803323633679146642488997344818325511778404482365180711855676555608632271919544012677375160646142389209537214343298265559346574409770769600994337288258446307873;
            6'd40: xpb[145] = 1024'd77593708444466801877334160910214955208558056683534878615337193040111683827085684103321647700644773464593025614179532003832478779068659683244492131619934797668767399076354993926750101980441153902047385100199385169482121391735008912793715915502015727319199184292010227038315104838116546566878160277867698211596;
            6'd41: xpb[145] = 1024'd91940220723990946064147407673451772363241850813196818993533808372612165456493740096906196014626660232152166195279769647386197132629498208781120447412066271703855651510220990508681878449103903321729589488543093783355610511550473812910056670357889065428861154240722188517283635266462323532761983267476950115319;
            6'd42: xpb[145] = 1024'd106286733003515090250960654436688589517925644942858759371730423705112647085901796090490744328608546999711306776380007290939915486190336734317748763204197745738943903944086987090613654917766652741411793876886802397229099631365938713026397425213762403538523124189434149996252165694808100498645806257086202019042;
            6'd43: xpb[145] = 1024'd120633245283039234437773901199925406672609439072520699749927039037613128715309852084075292642590433767270447357480244934493633839751175259854377078996329219774032156377952983672545431386429402161093998265230511011102588751181403613142738180069635741648185094138146111475220696123153877464529629246695453922765;
            6'd44: xpb[145] = 1024'd10913061878438637225788220558347791082594806076446955999991799305136715007408769167644769741914646225386438531122989143468288352470793450835845269772129652875429734242247762916846968663574945859466005045186979778611717020775971740294100365242279630491027160672741014924082698477571021413294762409679111342157;
            6'd45: xpb[145] = 1024'd25259574157962781412601467321584608237278600206108896378188414637637196636816825161229318055896532992945579112223226787022006706031631976372473585564261126910517986676113759498778745132237695279148209433530688392485206140591436640410441120098152968600689130621452976403051228905916798379178585399288363245880;
            6'd46: xpb[145] = 1024'd39606086437486925599414714084821425391962394335770836756385029970137678266224881154813866369878419760504719693323464430575725059592470501909101901356392600945606239109979756080710521600900444698830413821874397006358695260406901540526781874954026306710351100570164937882019759334262575345062408388897615149603;
            6'd47: xpb[145] = 1024'd53952598717011069786227960848058242546646188465432777134581645302638159895632937148398414683860306528063860274423702074129443413153309027445730217148524074980694491543845752662642298069563194118512618210218105620232184380222366440643122629809899644820013070518876899360988289762608352310946231378506867053326;
            6'd48: xpb[145] = 1024'd68299110996535213973041207611295059701329982595094717512778260635138641525040993141982962997842193295623000855523939717683161766714147552982358532940655549015782743977711749244574074538225943538194822598561814234105673500037831340759463384665772982929675040467588860839956820190954129276830054368116118957049;
            6'd49: xpb[145] = 1024'd82645623276059358159854454374531876856013776724756657890974875967639123154449049135567511311824080063182141436624177361236880120274986078518986848732787023050870996411577745826505851006888692957877026986905522847979162619853296240875804139521646321039337010416300822318925350619299906242713877357725370860772;
            6'd50: xpb[145] = 1024'd96992135555583502346667701137768694010697570854418598269171491300139604783857105129152059625805966830741282017724415004790598473835824604055615164524918497085959248845443742408437627475551442377559231375249231461852651739668761140992144894377519659148998980365012783797893881047645683208597700347334622764495;
            6'd51: xpb[145] = 1024'd111338647835107646533480947901005511165381364984080538647368106632640086413265161122736607939787853598300422598824652648344316827396663129592243480317049971121047501279309738990369403944214191797241435763592940075726140859484226041108485649233392997258660950313724745276862411475991460174481523336943874668218;
            6'd52: xpb[145] = 1024'd1618464430507049321495267259427895575366731988006794897432866900163672705364078206306085039112066056416413772467396857318971340116281320573711671092850404222445079143604518234670941221359735495613442543549408843235269129078794168259847834406036886101503016848319648725724413830408604123246656499927532087610;
            6'd53: xpb[145] = 1024'd15964976710031193508308514022664712730050526117668735275629482232664154334772134199890633353093952823975554353567634500872689693677119846110339986884981878257533331577470514816602717690022484915295646931893117457108758248894259068376188589261910224211164986797031610204692944258754381089130479489536783991333;
            6'd54: xpb[145] = 1024'd30311488989555337695121760785901529884734320247330675653826097565164635964180190193475181667075839591534694934667872144426408047237958371646968302677113352292621584011336511398534494158685234334977851320236826070982247368709723968492529344117783562320826956745743571683661474687100158055014302479146035895056;
            6'd55: xpb[145] = 1024'd44658001269079481881935007549138347039418114376992616032022712897665117593588246187059729981057726359093835515768109787980126400798796897183596618469244826327709836445202507980466270627347983754660055708580534684855736488525188868608870098973656900430488926694455533162630005115445935020898125468755287798779;
            6'd56: xpb[145] = 1024'd59004513548603626068748254312375164194101908506654556410219328230165599222996302180644278295039613126652976096868347431533844754359635422720224934261376300362798088879068504562398047096010733174342260096924243298729225608340653768725210853829530238540150896643167494641598535543791711986781948458364539702502;
            6'd57: xpb[145] = 1024'd73351025828127770255561501075611981348785702636316496788415943562666080852404358174228826609021499894212116677968585075087563107920473948256853250053507774397886341312934501144329823564673482594024464485267951912602714728156118668841551608685403576649812866591879456120567065972137488952665771447973791606225;
            6'd58: xpb[145] = 1024'd87697538107651914442374747838848798503469496765978437166612558895166562481812414167813374923003386661771257259068822718641281461481312473793481565845639248432974593746800497726261600033336232013706668873611660526476203847971583568957892363541276914759474836540591417599535596400483265918549594437583043509948;
            6'd59: xpb[145] = 1024'd102044050387176058629187994602085615658153290895640377544809174227667044111220470161397923236985273429330397840169060362194999815042150999330109881637770722468062846180666494308193376501998981433388873261955369140349692967787048469074233118397150252869136806489303379078504126828829042884433417427192295413671;
            6'd60: xpb[145] = 1024'd116390562666700202816001241365322432812837085025302317923005789560167525740628526154982471550967160196889538421269298005748718168602989524866738197429902196503151098614532490890125152970661730853071077650299077754223182087602513369190573873253023590978798776438015340557472657257174819850317240416801547317394;
            6'd61: xpb[145] = 1024'd6670379262099605604015560723744817222822452029228574173070549827691112032727443238551948650291372655005529594912042214723372681322607715848206388205702629604548676478827270134426690247807274551443084430255546521732310357197081496341936058425667479821640842972610244006334659611591963799082373579785204736786;
            6'd62: xpb[145] = 1024'd21016891541623749790828807486981634377506246158890514551267165160191593662135499232136496964273259422564670176012279858277091034883446241384834703997834103639636928912693266716358466716470023971125288818599255135605799477012546396458276813281540817931302812921322205485303190039937740764966196569394456640509;
            6'd63: xpb[145] = 1024'd35363403821147893977642054250218451532190040288552454929463780492692075291543555225721045278255146190123810757112517501830809388444284766921463019789965577674725181346559263298290243185132773390807493206942963749479288596828011296574617568137414156040964782870034166964271720468283517730850019559003708544232;
        endcase
    end

    always_comb begin
        case(flag[48][16:12])
            5'd0: xpb[146] = 1024'd0;
            5'd1: xpb[146] = 1024'd49709916100672038164455301013455268686873834418214395307660395825192556920951611219305593592237032957682951338212755145384527742005123292458091335582097051709813433780425259880222019653795522810489697595286672363352777716643476196690958322993287494150626752818746128443240250896629294696733842548612960447955;
            5'd2: xpb[146] = 1024'd99419832201344076328910602026910537373747668836428790615320791650385113841903222438611187184474065915365902676425510290769055484010246584916182671164194103419626867560850519760444039307591045620979395190573344726705555433286952393381916645986574988301253505637492256886480501793258589393467685097225920895910;
            5'd3: xpb[146] = 1024'd25063052617891373094566975635551373315923076128907501794849332410600775425545694747901709562053424563605704607180772001574519385174149542819113881729960114195749626771704562303035819769869362710158895177472777243693972299709531817107896399296633033185060355042121327299614224615959251073082837819213286859534;
            5'd4: xpb[146] = 1024'd74772968718563411259022276649006642002796910547121897102509728235793332346497305967207303154290457521288655945393527146959047127179272835277205217312057165905563060552129822183257839423664885520648592772759449607046750016353008013798854722289920527335687107860867455742854475512588545769816680367826247307489;
            5'd5: xpb[146] = 1024'd416189135110708024678650257647477944972317839600608282038268996008993930139778276497825531869816169528457876148788857764511028343175793180136427877823176681685819762983864725849619885943202609828092759658882124035166882775587437524834475599978572219493957265496526155988198335289207449431833089813613271113;
            5'd6: xpb[146] = 1024'd50126105235782746189133951271102746631846152257815003589698664821201550851091389495803419124106849127211409214361544003149038770348299085638227763459920228391499253543409124606071639539738725420317790354945554487387944599419063634215792798593266066370120710084242654599228449231918502146165675638426573719068;
            5'd7: xpb[146] = 1024'd99836021336454784353589252284558015318719986676029398897359060646394107772043000715109012716343882084894360552574299148533566512353422378096319099042017280101312687323834384486293659193534248230807487950232226850740722316062539830906751121586553560520747462902988783042468700128547796842899518187039534167023;
            5'd8: xpb[146] = 1024'd25479241753002081119245625893198851260895393968508110076887601406609769355685473024399535093923240733134162483329560859339030413517325335999250309607783290877435446534688427028885439655812565319986987937131659367729139182485119254632730874896611605404554312307617853455602422951248458522514670909026900130647;
            5'd9: xpb[146] = 1024'd75189157853674119283700926906654119947769228386722505384547997231802326276637084243705128686160273690817113821542316004723558155522448628457341645189880342587248880315113686909107459309608088130476685532418331731081916899128595451323689197889899099555181065126363981898842673847877753219248513457639860578602;
            5'd10: xpb[146] = 1024'd832378270221416049357300515294955889944635679201216564076537992017987860279556552995651063739632339056915752297577715529022056686351586360272855755646353363371639525967729451699239771886405219656185519317764248070333765551174875049668951199957144438987914530993052311976396670578414898863666179627226542226;
            5'd11: xpb[146] = 1024'd50542294370893454213812601528750224576818470097415611871736933817210544781231167772301244655976665296739867090510332860913549798691474878818364191337743405073185073306392989331921259425681928030145883114604436611423111482194651071740627274193244638589614667349739180755216647567207709595597508728240186990181;
            5'd12: xpb[146] = 1024'd100252210471565492378267902542205493263692304515630007179397329642403101702182778991606838248213698254422818428723088006298077540696598171276455526919840456782998507086818249212143279079477450840635580709891108974775889198838127268431585597186532132740241420168485309198456898463837004292331351276853147438136;
            5'd13: xpb[146] = 1024'd25895430888112789143924276150846329205867711808108718358925870402618763285825251300897360625793056902662620359478349717103541441860501129179386737485606467559121266297672291754735059541755767929815080696790541491764306065260706692157565350496590177624048269573114379611590621286537665971946503998840513401760;
            5'd14: xpb[146] = 1024'd75605346988784827308379577164301597892741546226323113666586266227811320206776862520202954218030089860345571697691104862488069183865624421637478073067703519268934700078097551634957079195551290740304778292077213855117083781904182888848523673489877671774675022391860508054830872183166960668680346547453473849715;
            5'd15: xpb[146] = 1024'd1248567405332124074035950772942433834916953518801824846114806988026981790419334829493476595609448508585373628446366573293533085029527379540409283633469530045057459288951594177548859657829607829484278278976646372105500648326762312574503426799935716658481871796489578467964595005867622348295499269440839813339;
            5'd16: xpb[146] = 1024'd50958483506004162238491251786397702521790787937016220153775202813219538711370946048799070187846481466268324966659121718678060827034650671998500619215566581754870893069376854057770879311625130639973975874263318735458278364970238509265461749793223210809108624615235706911204845902496917045029341818053800261294;
            5'd17: xpb[146] = 1024'd100668399606676200402946552799852971208664622355230615461435598638412095632322557268104663780083514423951276304871876864062588569039773964456591954797663633464684326849802113937992898965420653450463673469549991098811056081613714705956420072786510704959735377433981835354445096799126211741763184366666760709249;
            5'd18: xpb[146] = 1024'd26311620023223497168602926408493807150840029647709326640964139398627757215965029577395186157662873072191078235627138574868052470203676922359523165363429644240807086060656156480584679427698970539643173456449423615799472948036294129682399826096568749843542226838610905767578819621826873421378337088654126672873;
            5'd19: xpb[146] = 1024'd76021536123895535333058227421949075837713864065923721948624535223820314136916640796700779749899906029874029573839893720252580212208800214817614500945526695950620519841081416360806699081494493350132871051736095979152250664679770326373358149089856243994168979657357034210819070518456168118112179637267087120828;
            5'd20: xpb[146] = 1024'd1664756540442832098714601030589911779889271358402433128153075984035975720559113105991302127479264678113831504595155431058044113372703172720545711511292706726743279051935458903398479543772810439312371038635528496140667531102349750099337902399914288877975829061986104623952793341156829797727332359254453084452;
            5'd21: xpb[146] = 1024'd51374672641114870263169902044045180466763105776616828435813471809228532641510724325296895719716297635796782842807910576442571855377826465178637047093389758436556712832360718783620499197568333249802068633922200859493445247745825946790296225393201783028602581880732233067193044237786124494461174907867413532407;
            5'd22: xpb[146] = 1024'd101084588741786908427625203057500449153636940194831223743473867634421089562462335544602489311953330593479734181020665721827099597382949757636728382675486810146370146612785978663842518851363856060291766229208873222846222964389302143481254548386489277179229334699478361510433295134415419191195017456480373980362;
            5'd23: xpb[146] = 1024'd26727809158334205193281576666141285095812347487309934923002408394636751146104807853893011689532689241719536111775927432632563498546852715539659593241252820922492905823640021206434299313642173149471266216108305739834639830811881567207234301696547322063036184104107431923567017957116080870810170178467739943986;
            5'd24: xpb[146] = 1024'd76437725259006243357736877679596553782686181905524330230662804219829308067056419073198605281769722199402487449988682578017091240551976007997750928823349872632306339604065281086656318967437695959960963811394978103187417547455357763898192624689834816213662936922853560366807268853745375567544012727080700391941;
            5'd25: xpb[146] = 1024'd2080945675553540123393251288237389724861589198003041410191344980044969650698891382489127659349080847642289380743944288822555141715878965900682139389115883408429098814919323629248099429716013049140463798294410620175834413877937187624172377999892861097469786327482630779940991676446037247159165449068066355565;
            5'd26: xpb[146] = 1024'd51790861776225578287848552301692658411735423616217436717851740805237526571650502601794721251586113805325240718956699434207082883721002258358773474971212935118242532595344583509470119083511535859630161393581082983528612130521413384315130700993180355248096539146228759223181242573075331943893007997681026803520;
            5'd27: xpb[146] = 1024'd101500777876897616452303853315147927098609258034431832025512136630430083492602113821100314843823146763008192057169454579591610625726125550816864810553309986828055966375769843389692138737307058670119858988867755346881389847164889581006089023986467849398723291964974887666421493469704626640626850546293987251475;
            5'd28: xpb[146] = 1024'd27143998293444913217960226923788763040784665326910543205040677390645745076244586130390837221402505411247993987924716290397074526890028508719796021119075997604178725586623885932283919199585375759299358975767187863869806713587469004732068777296525894282530141369603958079555216292405288320242003268281353215099;
            5'd29: xpb[146] = 1024'd76853914394116951382415527937244031727658499745124938512701073215838301997196197349696430813639538368930945326137471435781602268895151801177887356701173049313992159367049145812505938853380898569789056571053860227222584430230945201423027100289813388433156894188350086522795467189034583016975845816894313663054;
            5'd30: xpb[146] = 1024'd2497134810664248148071901545884867669833907037603649692229613976053963580838669658986953191218897017170747256892733146587066170059054759080818567266939060090114918577903188355097719315659215658968556557953292744211001296653524625149006853599871433316963743592979156935929190011735244696590998538881679626678;
            5'd31: xpb[146] = 1024'd52207050911336286312527202559340136356707741455818044999890009801246520501790280878292546783455929974853698595105488291971593912064178051538909902849036111799928352358328448235319738969454738469458254153239965107563779013297000821839965176593158927467590496411725285379169440908364539393324841087494640074633;
        endcase
    end

    always_comb begin
        case(flag[49][5:0])
            6'd0: xpb[147] = 1024'd0;
            6'd1: xpb[147] = 1024'd50958483506004162238491251786397702521790787937016220153775202813219538711370946048799070187846481466268324966659121718678060827034650671998500619215566581754870893069376854057770879311625130639973975874263318735458278364970238509265461749793223210809108624615235706911204845902496917045029341818053800261294;
            6'd2: xpb[147] = 1024'd101916967012008324476982503572795405043581575874032440307550405626439077422741892097598140375692962932536649933318243437356121654069301343997001238431133163509741786138753708115541758623250261279947951748526637470916556729940477018530923499586446421618217249230471413822409691804993834090058683636107600522588;
            6'd3: xpb[147] = 1024'd28808754833887745316674827954378674820673936685312976333193753374681720796803699236382139348881770089361825492519871721455118640262731681440341732630368704330922004638559344835682398743358186198611730014402716360010474244689818754831406679696440183160505970431590062703508009633562118117969335627535806299551;
            6'd4: xpb[147] = 1024'd79767238339891907555166079740776377342464724622329196486968956187901259508174645285181209536728251555630150459178993440133179467297382353438842351845935286085792897707936198893453278054983316838585705888666035095468752609660057264096868429489663393969614595046825769614712855536059035162998677445589606560845;
            6'd5: xpb[147] = 1024'd6659026161771328394858404122359647119557085433609732512612303936143902882236452423965208509917058712455326018380621724232176453490812690882182846045170826906973116207741835613593918175091241757249484154542113984562670124409399000397351609599657155511903316247944418495811173364627319190909329437017812337808;
            6'd6: xpb[147] = 1024'd57617509667775490633349655908757349641347873370625952666387506749363441593607398472764278697763540178723650985039743442910237280525463362880683465260737408661844009277118689671364797486716372397223460028805432720020948489379637509662813359392880366321011940863180125407016019267124236235938671255071612599102;
            6'd7: xpb[147] = 1024'd108575993173779652871840907695155052163138661307642172820162709562582980304978344521563348885610021644991975951698865161588298107560114034879184084476303990416714902346495543729135676798341503037197435903068751455479226854349876018928275109186103577130120565478415832318220865169621153280968013073125412860396;
            6'd8: xpb[147] = 1024'd35467780995659073711533232076738321940231022118922708845806057310825623679040151660347347858798828801817151510900493445687295093753544372322524578675539531237895120846301180449276316918449427955861214168944830344573144369099217755228758289296097338672409286679534481199319182998189437308878665064553618637359;
            6'd9: xpb[147] = 1024'd86426264501663235950024483863136024462021810055938928999581260124045162390411097709146418046645310268085476477559615164365355920788195044321025197891106112992766013915678034507047196230074558595835190043208149080031422734069456264494220039089320549481517911294770188110524028900686354353908006882607418898653;
            6'd10: xpb[147] = 1024'd13318052323542656789716808244719294239114170867219465025224607872287805764472904847930417019834117424910652036761243448464352906981625381764365692090341653813946232415483671227187836350182483514498968309084227969125340248818798000794703219199314311023806632495888836991622346729254638381818658874035624675616;
            6'd11: xpb[147] = 1024'd64276535829546819028208060031116996760904958804235685178999810685507344475843850896729487207680598891178977003420365167142413734016276053762866311305908235568817125484860525284958715661807614154472944183347546704583618613789036510060164968992537521832915257111124543902827192631751555426848000692089424936910;
            6'd12: xpb[147] = 1024'd115235019335550981266699311817514699282695746741251905332775013498726883187214796945528557395527080357447301970079486885820474561050926725761366930521474817323688018554237379342729594973432744794446920057610865440041896978759275019325626718785760732642023881726360250814032038534248472471877342510143225198204;
            6'd13: xpb[147] = 1024'd42126807157430402106391636199097969059788107552532441358418361246969526561276604084312556368715887514272477529281115169919471547244357063204707424720710358144868237054043016062870235093540669713110698323486944329135814493508616755626109898895754494184312602927478899695130356362816756499787994501571430975167;
            6'd14: xpb[147] = 1024'd93085290663434564344882887985495671581578895489548661512193564060189065272647550133111626556562368980540802495940236888597532374279007735203208043936276939899739130123419870120641114405165800353084674197750263064594092858478855264891571648688977704993421227542714606606335202265313673544817336319625231236461;
            6'd15: xpb[147] = 1024'd19977078485313985184575212367078941358671256300829197537836911808431708646709357271895625529751176137365978055141865172696529360472438072646548538135512480720919348623225506840781754525273725271748452463626341953688010373228197001192054828798971466535709948743833255487433520093881957572727988311053437013424;
            6'd16: xpb[147] = 1024'd70935561991318147423066464153476643880462044237845417691612114621651247358080303320694695717597657603634303021800986891374590187507088744645049157351079062475790241692602360898552633836898855911722428337889660689146288738198435510457516578592194677344818573359068962398638365996378874617757330129107237274718;
            6'd17: xpb[147] = 1024'd121894045497322309661557715939874346402252832174861637845387317434870786069451249369493765905444139069902627988460108610052651014541739416643549776566645644230661134761979214956323513148523986551696404212152979424604567103168674019722978328385417888153927197974304669309843211898875791662786671947161037536012;
            6'd18: xpb[147] = 1024'd48785833319201730501250040321457616179345192986142173871030665183113429443513056508277764878632946226727803547661736894151648000735169754086890270765881185051841353261784851676464153268631911470360182478029058313698484617918015756023461508495411649696215919175423318190941529727444075690697323938589243312975;
            6'd19: xpb[147] = 1024'd99744316825205892739741292107855318701135980923158394024805867996332968154884002557076835066479427692996128514320858612829708827769820426085390889981447766806712246331161705734235032580257042110334158352292377049156762982888254265288923258288634860505324543790659025102146375629940992735726665756643043574269;
            6'd20: xpb[147] = 1024'd26636104647085313579433616489438588478228341734438930050449215744575611528945809695860834039668234849821304073522486896928705813963250763528731384180683307627892464830967342454375672700364967028997936618168455938250680497637596001589406438398628622047613264991777673983244693458509276763637317748071249351232;
            6'd21: xpb[147] = 1024'd77594588153089475817924868275836291000019129671455150204224418557795150240316755744659904227514716316089629040181608615606766640997901435527232003396249889382763357900344196512146552011990097668971912492431774673708958862607834510854868188191851832856721889607013380894449539361006193808666659566125049612526;
            6'd22: xpb[147] = 1024'd4486375974968896657617192657419560777111490482735686229867766306037793614378562883443903200703523472914804599383236899705763627191331772970572497595485430203943576400149833232287192132098022587635690758307853562802876377357176247155351368301845594399010610808132029775547857189574477836577311557553255389489;
            6'd23: xpb[147] = 1024'd55444859480973058896108444443817263298902278419751906383642969119257332325749508932242973388550004939183129566042358618383824454225982444969073116811052011958814469469526687290058071443723153227609666632571172298261154742327414756420813118095068805208119235423367736686752703092071394881606653375607055650783;
            6'd24: xpb[147] = 1024'd106403342986977221134599696230214965820693066356768126537418171932476871037120454981042043576396486405451454532701480337061885281260633116967573736026618593713685362538903541347828950755348283867583642506834491033719433107297653265686274867888292016017227860038603443597957548994568311926635995193660855912077;
            6'd25: xpb[147] = 1024'd33295130808856641974292020611798235597785427168048662563061519680719514411182262119826042549585293562276630091903108621160882267454063454410914230225854134534865581038709178067969590875456208786247420772710569922813350622046995001986758047998285777559516581239722092479055866823136595954546647185089061689040;
            6'd26: xpb[147] = 1024'd84253614314860804212783272398195938119576215105064882716836722493939053122553208168625112737431775028544955058562230339838943094488714126409414849441420716289736474108086032125740470187081339426221396646973888658271628987017233511252219797791508988368625205854957799390260712725633512999575989003142861950334;
            6'd27: xpb[147] = 1024'd11145402136740225052475596779779207896668575916345418742480070242181696496615015307409111710620582185370130617763858623937940080682144463852755343640656257110916692607891668845881110307189264344885174912849967547365546501766575247552702977901502749910913927056076448271359030554201797027486640994571067727297;
            6'd28: xpb[147] = 1024'd62103885642744387290966848566176910418459363853361638896255273055401235207985961356208181898467063651638455584422980342616000907716795135851255962856222838865787585677268522903651989618814394984859150787113286282823824866736813756818164727694725960720022551671312155182563876456698714072515982812624867988591;
            6'd29: xpb[147] = 1024'd113062369148748549529458100352574612940250151790377859050030475868620773919356907405007252086313545117906780551082102061294061734751445807849756582071789420620658478746645376961422868930439525624833126661376605018282103231707052266083626477487949171529131176286547862093768722359195631117545324630678668249885;
            6'd30: xpb[147] = 1024'd39954156970627970369150424734157882717342512601658395075673823616863417293418714543791251059502352274731956110283730345393058720944876145293097076271024961441838697246451013681563509050547450543496904927252683907376020746456394002384109657597942933071419897487666510974867040187763915145455976622106874026848;
            6'd31: xpb[147] = 1024'd90912640476632132607641676520555585239133300538674615229449026430082956004789660592590321247348833741000281076942852064071119547979526817291597695486591543196709590315827867739334388362172581183470880801516002642834299111426632511649571407391166143880528522102902217886071886090260832190485318440160674288142;
            6'd32: xpb[147] = 1024'd17804428298511553447334000902138855016225661349955151255092374178325599378851467731374320220537640897825456636144480348170116534172957154734938189685827084017889808815633504459475028482280506102134659067392081531928216626175974247950054587501159905422817243304020866767170203918829116218395970431588880065105;
            6'd33: xpb[147] = 1024'd68762911804515715685825252688536557538016449286971371408867576991545138090222413780173390408384122364093781602803602066848177361207607826733438808901393665772760701885010358517245907793905636742108634941655400267386494991146212757215516337294383116231925867919256573678375049821326033263425312249642680326399;
            6'd34: xpb[147] = 1024'd119721395310519877924316504474934260059807237223987591562642779804764676801593359828972460596230603830362106569462723785526238188242258498731939428116960247527631594954387212575016787105530767382082610815918719002844773356116451266480978087087606327041034492534492280589579895723822950308454654067696480587693;
            6'd35: xpb[147] = 1024'd46613183132399298764008828856517529836899598035268127588286127553007320175655166967756459569419410987187282128664352069625235174435688836175279922316195788348811813454192849295157427225638692300746389081794797891938690870865793002781461267197600088583323213735610929470678213552391234336365306059124686364656;
            6'd36: xpb[147] = 1024'd97571666638403461002500080642915232358690385972284347742061330366226858887026113016555529757265892453455607095323473788303296001470339508173780541531762370103682706523569703352928306537263822940720364956058116627396969235836031512046923016990823299392431838350846636381883059454888151381394647877178486625950;
            6'd37: xpb[147] = 1024'd24463454460282881842192405024498502135782746783564883767704678114469502261087920155339528730454699610280782654525102072402292987663769845617121035730997910924862925023375340073068946657371747859384143221934195516490886750585373248347406197100817060934720559551965285262981377283456435409305299868606692402913;
            6'd38: xpb[147] = 1024'd75421937966287044080683656810896204657573534720581103921479880927689040972458866204138598918301181076549107621184223791080353814698420517615621654946564492679733818092752194130839825968996878499358119096197514251949165115555611757612867946894040271743829184167200992174186223185953352454334641686660492664207;
            6'd39: xpb[147] = 1024'd2313725788166464920375981192479474434665895531861639947123228675931684346520673342922597891489988233374283180385852075179350800891850855058962149145800033500914036592557830850980466089104803418021897362073593141043082630304953493913351127004034033286117905368319641055284541014521636482245293678088698441170;
            6'd40: xpb[147] = 1024'd53272209294170627158867232978877176956456683468877860100898431489151223057891619391721668079336469699642608147044973793857411627926501527057462768361366615255784929661934684908751345400729934057995873236336911876501360995275192003178812876797257244095226529983555347966489386917018553527274635496142498702464;
            6'd41: xpb[147] = 1024'd104230692800174789397358484765274879478247471405894080254673634302370761769262565440520738267182951165910933113704095512535472454961152199055963387576933197010655822731311538966522224712355064697969849110600230611959639360245430512444274626590480454904335154598791054877694232819515470572303977314196298963758;
            6'd42: xpb[147] = 1024'd31122480622054210237050809146858149255339832217174616280316982050613405143324372579304737240371758322736108672905723796634469441154582536499303881776168737831836041231117175686662864832462989616633627376476309501053556874994772248744757806700474216446623875799909703758792550648083754600214629305624504740721;
            6'd43: xpb[147] = 1024'd82080964128058372475542060933255851777130620154190836434092184863832943854695318628103807428218239789004433639564845515312530268189233208497804500991735319586706934300494029744433744144088120256607603250739628236511835239965010758010219556493697427255732500415145410669997396550580671645243971123678305002015;
            6'd44: xpb[147] = 1024'd8972751949937793315234385314839121554222980965471372459735532612075587228757125766887806401407046945829609198766473799411527254382663545941144995190970860407887152800299666464574384264196045175271381516615707125605752754714352494310702736603691188798021221616264059551095714379148955673154623115106510778978;
            6'd45: xpb[147] = 1024'd59931235455941955553725637101236824076013768902487592613510735425295125940128071815686876589253528412097934165425595518089588081417314217939645614406537442162758045869676520522345263575821175815245357390879025861064031119684591003576164486396914399607129846231499766462300560281645872718183964933160311040272;
            6'd46: xpb[147] = 1024'd110889718961946117792216888887634526597804556839503812767285938238514664651499017864485946777100009878366259132084717236767648908451964889938146233622104023917628938939053374580116142887446306455219333265142344596522309484654829512841626236190137610416238470846735473373505406184142789763213306751214111301566;
            6'd47: xpb[147] = 1024'd37781506783825538631909213269217796374896917650784348792929285986757308025560825003269945750288817035191434691286345520866645894645395227381486727821339564738809157438859011300256783007554231373883111531018423485616226999404171249142109416300131371958527192047854122254603724012711073791123958742642317078529;
            6'd48: xpb[147] = 1024'd88739990289829700870400465055615498896687705587800568946704488799976846736931771052069015938135298501459759657945467239544706721680045899379987347036906146493680050508235865358027662319179362013857087405281742221074505364374409758407571166093354582767635816663089829165808569915207990836153300560696117339823;
            6'd49: xpb[147] = 1024'd15631778111709121710092789437198768673780066399081104972347836548219490110993578190853014911324105658284935217147095523643703707873476236823327841236141687314860269008041502078168302439287286932520865671157821110168422879123751494708054346203348344309924537864208478046906887743776274864063952552124323116786;
            6'd50: xpb[147] = 1024'd66590261617713283948584041223596471195570854336097325126123039361439028822364524239652085099170587124553260183806217242321764534908126908821828460451708269069731162077418356135939181750912417572494841545421139845626701244093990003973516095996571555119033162479444184958111733646273191909093294370178123378080;
            6'd51: xpb[147] = 1024'd117548745123717446187075293009994173717361642273113545279898242174658567533735470288451155287017068590821585150465338960999825361942777580820329079667274850824602055146795210193710061062537548212468817419684458581084979609064228513238977845789794765928141787094679891869316579548770108954122636188231923639374;
            6'd52: xpb[147] = 1024'd44440532945596867026767617391577443494454003084394081305541589922901210907797277427235154260205875747646760709666967245098822348136207918263669573866510391645782273646600846913850701182645473131132595685560537470178897123813570249539461025899788527470430508295798540750414897377338392982033288179660129416337;
            6'd53: xpb[147] = 1024'd95399016451601029265258869177975146016244791021410301459316792736120749619168223476034224448052357213915085676326088963776883175170858590262170193082076973400653166715977700971621580494270603771106571559823856205637175488783808758804922775693011738279539132911034247661619743279835310027062629997713929677631;
            6'd54: xpb[147] = 1024'd22290804273480450104951193559558415793337151832690837484960140484363392993230030614818223421241164370740261235527717247875880161364288927705510687281312514221833385215783337691762220614378528689770349825699935094731093003533150495105405955803005499821827854112152896542718061108403594054973281989142135454594;
            6'd55: xpb[147] = 1024'd73249287779484612343442445345956118315127939769707057638735343297582931704600976663617293609087645837008586202186838966553940988398939599704011306496879095976704278285160191749533099926003659329744325699963253830189371368503389004370867705596228710630936478727388603453922907010900511100002623807195935715888;
            6'd56: xpb[147] = 1024'd141075601364033183134769727539388092220300580987593664378691045825575078662783802401292582276452993833761761388467250652937974592369937147351800696114636797884496784965828469673740046111584248408103965839332719283288883252730740671350885706222472173225199928507252335021224839468795127913275798624141492851;
            6'd57: xpb[147] = 1024'd51099559107368195421626021513937090614011088518003813818153893859045113790033729851200362770122934460102086728047588969330998801627020609145852419911681218552755389854342682527444619357736714888382079840102651454741567248222969249936812635499445682982333824543742959246226070741965712172942617616677941754145;
            6'd58: xpb[147] = 1024'd102058042613372357660117273300334793135801876455020033971929096672264652501404675899999432957969415926370411694706710688009059628661671281144353039127247800307626282923719536585215498669361845528356055714365970190199845613193207759202274385292668893791442449158978666157430916644462629217971959434731742015439;
            6'd59: xpb[147] = 1024'd28949830435251778499809597681918062912894237266300569997572444420507295875466483038783431931158223083195587253908338972108056614855101618587693533326483341128806501423525173305356138789469770447019833980242049079293763127942549495502757565402662655333731170360097315038529234473030913245882611426159947792402;
            6'd60: xpb[147] = 1024'd79908313941255940738300849468315765434685025203316790151347647233726834586837429087582502119004704549463912220567460690786117441889752290586194152542049922883677394492902027363127018101094901086993809854505367814752041492912788004768219315195885866142839794975333021949734080375527830290911953244213748053696;
            6'd61: xpb[147] = 1024'd6800101763135361577993173849899035211777386014597326176990994981969477960899236226366501092193511706289087779769088974885114428083182628029534646741285463704857612992707664083267658221202826005657588120381446703845959007662129741068702495305879627685128516176451670830832398204096114318822605235641953830659;
            6'd62: xpb[147] = 1024'd57758585269139523816484425636296737733568173951613546330766197795189016672270182275165571280039993172557412746428210693563175255117833300028035265956852045459728506062084518141038537532827956645631563994644765439304237372632368250334164245099102838494237140791687377742037244106593031363851947053695754091953;
            6'd63: xpb[147] = 1024'd108717068775143686054975677422694440255358961888629766484541400608408555383641128323964641467886474638825737713087332412241236082152483972026535885172418627214599399131461372198809416844453087285605539868908084174762515737602606759599625994892326049303345765406923084653242090009089948408881288871749554353247;
        endcase
    end

    always_comb begin
        case(flag[49][11:6])
            6'd0: xpb[148] = 1024'd0;
            6'd1: xpb[148] = 1024'd35608856597023106894668001804277710032451322699910302510184748356651198757702935462748640441075281795650913272288960696340233068345914309469876379371654168035779617631267008918950056964561012204269318134784163063856433252351948495900109175002319810845634486608041733534340407837658232436791940863177760130210;
            6'd2: xpb[148] = 1024'd71217713194046213789336003608555420064902645399820605020369496713302397515405870925497280882150563591301826544577921392680466136691828618939752758743308336071559235262534017837900113929122024408538636269568326127712866504703896991800218350004639621691268973216083467068680815675316464873583881726355520260420;
            6'd3: xpb[148] = 1024'd106826569791069320684004005412833130097353968099730907530554245069953596273108806388245921323225845386952739816866882089020699205037742928409629138114962504107338852893801026756850170893683036612807954404352489191569299757055845487700327525006959432536903459824125200603021223512974697310375822589533280390630;
            6'd4: xpb[148] = 1024'd18368730703967686179873079812296407385106863673905525912607138361627899693502602940979490549643452873160503681698349350781868432542436903324345392470285631209427795955496818338169988666726843095767074930749412409061372159186897210635458130326049794115718043018049876107255103276704296730049073626085446036509;
            6'd5: xpb[148] = 1024'd53977587300990793074541081616574117417558186373815828422791886718279098451205538403728130990718734668811416953987310047122101500888351212794221771841939799245207413586763827257120045631287855300036393065533575472917805411538845706535567305328369604961352529626091609641595511114362529166841014489263206166719;
            6'd6: xpb[148] = 1024'd89586443898013899969209083420851827450009509073726130932976635074930297208908473866476771431794016464462330226276270743462334569234265522264098151213593967280987031218030836176070102595848867504305711200317738536774238663890794202435676480330689415806987016234133343175935918952020761603632955352440966296929;
            6'd7: xpb[148] = 1024'd1128604810912265465078157820315104737762404647900749315029528366604600629302270419210340658211623950670094091107738005223503796738959497178814405568917094383075974279726627757389920368892673987264831726714661754266311066021845925370807085649779777385801599428058018680169798715750361023306206388993131942808;
            6'd8: xpb[148] = 1024'd36737461407935372359746159624592814770213727347811051825214276723255799387005205881958981099286905746321007363396698701563736865084873806648690784940571262418855591910993636676339977333453686191534149861498824818122744318373794421270916260652099588231436086036099752214510206553408593460098147252170892073018;
            6'd9: xpb[148] = 1024'd72346318004958479254414161428870524802665050047721354335399025079906998144708141344707621540362187541971920635685659397903969933430788116118567164312225430454635209542260645595290034298014698395803467996282987881979177570725742917171025435654419399077070572644141485748850614391066825896890088115348652203228;
            6'd10: xpb[148] = 1024'd107955174601981586149082163233148234835116372747631656845583773436558196902411076807456261981437469337622833907974620094244203001776702425588443543683879598490414827173527654514240091262575710600072786131067150945835610823077691413071134610656739209922705059252183219283191022228725058333682028978526412333438;
            6'd11: xpb[148] = 1024'd19497335514879951644951237632611512122869268321806275227636666728232500322804873360189831207855076823830597772806087356005372229281396400503159798039202725592503770235223446095559909035619517083031906657464074163327683225208743136006265215975829571501519642446107894787424901992454657753355280015078577979317;
            6'd12: xpb[148] = 1024'd55106192111903058539619239436889222155320591021716577737821415084883699080507808822938471648930358619481511045095048052345605297627310709973036177410856893628283387866490455014509966000180529287301224792248237227184116477560691631906374390978149382347154129054149628321765309830112890190147220878256338109527;
            6'd13: xpb[148] = 1024'd90715048708926165434287241241166932187771913721626880248006163441534897838210744285687112090005640415132424317384008748685838365973225019442912556782511061664063005497757463933460022964741541491570542927032400291040549729912640127806483565980469193192788615662191361856105717667771122626939161741434098239737;
            6'd14: xpb[148] = 1024'd2257209621824530930156315640630209475524809295801498630059056733209201258604540838420681316423247901340188182215476010447007593477918994357628811137834188766151948559453255514779840737785347974529663453429323508532622132043691850741614171299559554771603198856116037360339597431500722046612412777986263885616;
            6'd15: xpb[148] = 1024'd37866066218847637824824317444907919507976131995711801140243805089860400016307476301169321757498529696991101454504436706787240661823833303827505190509488356801931566190720264433729897702346360178798981588213486572389055384395640346641723346301879365617237685464157770894680005269158954483404353641164024015826;
            6'd16: xpb[148] = 1024'd73474922815870744719492319249185629540427454695622103650428553446511598774010411763917962198573811492642014726793397403127473730169747613297381569881142524837711183821987273352679954666907372383068299722997649636245488636747588842541832521304199176462872172072199504429020413106817186920196294504341784146036;
            6'd17: xpb[148] = 1024'd109083779412893851614160321053463339572878777395532406160613301803162797531713347226666602639649093288292927999082358099467706798515661922767257949252796692873490801453254282271630011631468384587337617857781812700101921889099537338441941696306518987308506658680241237963360820944475419356988235367519544276246;
            6'd18: xpb[148] = 1024'd20625940325792217110029395452926616860631672969707024542666195094837100952107143779400171866066700774500691863913825361228876026020355897681974203608119819975579744514950073852949829404512191070296738384178735917593994291230589061377072301625609348887321241874165913467594700708205018776661486404071709922125;
            6'd19: xpb[148] = 1024'd56234796922815324004697397257204326893082995669617327052850943451488299709810079242148812307141982570151605136202786057569109094366270207151850582979773988011359362146217082771899886369073203274566056518962898981450427543582537557277181476627929159732955728482207647001935108545863251213453427267249470052335;
            6'd20: xpb[148] = 1024'd91843653519838430899365399061482036925534318369527629563035691808139498467513014704897452748217264365802518408491746753909342162712184516621726962351428156047138979777484091690849943333634215478835374653747062045306860795934486053177290651630248970578590215090249380536275516383521483650245368130427230182545;
            6'd21: xpb[148] = 1024'd3385814432736796395234473460945314213287213943702247945088585099813801887906811257631021974634871852010282273323214015670511390216878491536443216706751283149227922839179883272169761106678021961794495180143985262798933198065537776112421256949339332157404798284174056040509396147251083069918619166979395828424;
            6'd22: xpb[148] = 1024'd38994671029759903289902475265223024245738536643612550455273333456465000645609746720379662415710153647661195545612174712010744458562792801006319596078405451185007540470446892191119818071239034166063813314928148326655366450417486272012530431951659143003039284892215789574849803984909315506710560030157155958634;
            6'd23: xpb[148] = 1024'd74603527626783010184570477069500734278189859343522852965458081813116199403312682183128302856785435443312108817901135408350977526908707110476195975450059619220787158101713901110069875035800046370333131449712311390511799702769434767912639606953978953848673771500257523109190211822567547943502500893334916088844;
            6'd24: xpb[148] = 1024'd110212384223806117079238478873778444310641182043433155475642830169767398161015617645876943297860717238963022090190096104691210595254621419946072354821713787256566775732980910029019932000361058574602449584496474454368232955121383263812748781956298764694308258108299256643530619660225780380294441756512676219054;
            6'd25: xpb[148] = 1024'd21754545136704482575107553273241721598394077617607773857695723461441701581409414198610512524278324725170785955021563366452379822759315394860788609177036914358655718794676701610339749773404865057561570110893397671860305357252434986747879387275389126273122841302223932147764499423955379799967692793064841864933;
            6'd26: xpb[148] = 1024'd57363401733727589469775555077519431630845400317518076367880471818092900339112349661359152965353606520821699227310524062792612891105229704330664988548691082394435336425943710529289806737965877261830888245677560735716738609604383482647988562277708937118757327910265665682104907261613612236759633656242601995143;
            6'd27: xpb[148] = 1024'd92972258330750696364443556881797141663296723017428378878065220174744099096815285124107793406428888316472612499599484759132845959451144013800541367920345250430214954057210719448239863702526889466100206380461723799573171861956331978548097737280028747964391814518307399216445315099271844673551574519420362125353;
            6'd28: xpb[148] = 1024'd4514419243649061860312631281260418951049618591602997260118113466418402517209081676841362632846495802680376364430952020894015186955837988715257622275668377532303897118906511029559681475570695949059326906858647017065244264087383701483228342599119109543206397712232074720679194863001444093224825555972527771232;
            6'd29: xpb[148] = 1024'd40123275840672168754980633085538128983500941291513299770302861823069601274912017139590003073921777598331289636719912717234248255301752298185134001647322545568083514750173519948509738440131708153328645041642810080921677516439332197383337517601438920388840884320273808255019602700659676530016766419150287901442;
            6'd30: xpb[148] = 1024'd75732132437695275649648634889815839015952263991423602280487610179720800032614952602338643514997059393982202909008873413574481323647666607655010381018976713603863132381440528867459795404692720357597963176426973144778110768791280693283446692603758731234475370928315541789360010538317908966808707282328048031652;
            6'd31: xpb[148] = 1024'd111340989034718382544316636694093549048403586691333904790672358536371998790317888065087283956072341189633116181297834109914714391993580917124886760390630881639642750012707537786409852369253732561867281311211136208634544021143229189183555867606078542080109857536357275323700418375976141403600648145505808161862;
            6'd32: xpb[148] = 1024'd22883149947616748040185711093556826336156482265508523172725251828046302210711684617820853182489948675840880046129301371675883619498274892039603014745954008741731693074403329367729670142297539044826401837608059426126616423274280912118686472925168903658924440730281950827934298139705740823273899182057973807741;
            6'd33: xpb[148] = 1024'd58492006544639854934853712897834536368607804965418825682910000184697500968414620080569493623565230471491793318418262068016116687844189201509479394117608176777511310705670338286679727106858551249095719972392222489983049675626229408018795647927488714504558927338323684362274705977363973260065840045235733937951;
            6'd34: xpb[148] = 1024'd94100863141662961829521714702112246401059127665329128193094748541348699726117555543318134064640512267142706590707222764356349756190103510979355773489262344813290928336937347205629784071419563453365038107176385553839482927978177903918904822929808525350193413946365417896615113815022205696857780908413494068161;
            6'd35: xpb[148] = 1024'd5643024054561327325390789101575523688812023239503746575147641833023003146511352096051703291058119753350470455538690026117518983694797485894072027844585471915379871398633138786949601844463369936324158633573308771331555330109229626854035428248898886929007997140290093400848993578751805116531031944965659714040;
            6'd36: xpb[148] = 1024'd41251880651584434220058790905853233721263345939414049085332390189674201904214287558800343732133401549001383727827650722457752052040711795363948407216239639951159489029900147705899658809024382140593476768357471835187988582461178122754144603251218697774642483748331826935189401416410037553322972808143419844250;
            6'd37: xpb[148] = 1024'd76860737248607541114726792710130943753714668639324351595517138546325400661917223021548984173208683344652297000116611418797985120386626104833824786587893807986939106661167156624849715773585394344862794903141634899044421834813126618654253778253538508620276970356373560469529809254068269990114913671321179974460;
            6'd38: xpb[148] = 1024'd112469593845630648009394794514408653786165991339234654105701886902976599419620158484297624614283965140303210272405572115138218188732540414303701165959547976022718724292434165543799772738146406549132113037925797962900855087165075114554362953255858319465911456964415294003870217091726502426906854534498940104670;
            6'd39: xpb[148] = 1024'd24011754758529013505263868913871931073918886913409272487754780194650902840013955037031193840701572626510974137237039376899387416237234389218417420314871103124807667354129957125119590511190213032091233564322721180392927489296126837489493558574948681044726040158339969508104096855456101846580105571051105750549;
            6'd40: xpb[148] = 1024'd59620611355552120399931870718149641106370209613319574997939528551302101597716890499779834281776854422161887409526000073239620484583148698688293799686525271160587284985396966044069647475751225236360551699106884244249360741648075333389602733577268491890360526766381703042444504693114334283372046434228865880759;
            6'd41: xpb[148] = 1024'd95229467952575227294599872522427351138821532313229877508124276907953300355419825962528474722852136217812800681814960769579853552929063008158170179058179439196366902616663974963019704440312237440629869833891047308105793994000023829289711908579588302735995013374423436576784912530772566720163987297406626010969;
            6'd42: xpb[148] = 1024'd6771628865473592790468946921890628426574427887404495890177170199627603775813622515262043949269743704020564546646428031341022780433756983072886433413502566298455845678359766544339522213356043923588990360287970525597866396131075552224842513898678664314809596568348112081018792294502166139837238333958791656848;
            6'd43: xpb[148] = 1024'd42380485462496699685136948726168338459025750587314798400361918556278802533516557978010684390345025499671477818935388727681255848779671292542762812785156734334235463309626775463289579177917056127858308495072133589454299648483024048124951688900998475160444083176389845615359200132160398576629179197136551787058;
            6'd44: xpb[148] = 1024'd77989342059519806579804950530446048491477073287225100910546666912930001291219493440759324831420307295322391091224349424021488917125585602012639192156810902370015080940893784382239636142478068332127626629856296653310732900834972544025060863903318286006078569784431579149699607969818631013421120060314311917268;
            6'd45: xpb[148] = 1024'd113598198656542913474472952334723758523928395987135403420731415269581200048922428903507965272495589090973304363513310120361721985471499911482515571528465070405794698572160793301189693107039080536396944764640459717167166153186921039925170038905638096851713056392473312684040015807476863450213060923492072047478;
            6'd46: xpb[148] = 1024'd25140359569441278970342026734187035811681291561310021802784308561255503469316225456241534498913196577181068228344777382122891212976193886397231825883788197507883641633856584882509510880082887019356065291037382934659238555317972762860300644224728458430527639586397988188273895571206462869886311960044237693357;
            6'd47: xpb[148] = 1024'd60749216166464385865010028538464745844132614261220324312969056917906702227019160918990174939988478372831981500633738078463124281322108195867108205255442365543663259265123593801459567844643899223625383425821545998515671807669921258760409819227048269276162126194439721722614303408864695306678252823221997823567;
            6'd48: xpb[148] = 1024'd96358072763487492759678030342742455876583936961130626823153805274557900984722096381738815381063760168482894772922698774803357349668022505336984584627096533579442876896390602720409624809204911427894701560605709062372105060021869754660518994229368080121796612802481455256954711246522927743470193686399757953777;
            6'd49: xpb[148] = 1024'd7900233676385858255547104742205733164336832535305245205206698566232204405115892934472384607481367654690658637754166036564526577172716480251700838982419660681531819958086394301729442582248717910853822087002632279864177462152921477595649599548458441700611195996406130761188591010252527163143444722951923599656;
            6'd50: xpb[148] = 1024'd43509090273408965150215106546483443196788155235215547715391446922883403162818828397221025048556649450341571910043126732904759645518630789721577218354073828717311437589353403220679499546809730115123140221786795343720610714504869973495758774550778252546245682604447864295528998847910759599935385586129683729866;
            6'd51: xpb[148] = 1024'd79117946870432072044883108350761153229239477935125850225576195279534601920521763859969665489631931245992485182332087429244992713864545099191453597725727996753091055220620412139629556511370742319392458356570958407577043966856818469395867949553098063391880169212489597829869406685568992036727326449307443860076;
            6'd52: xpb[148] = 1024'd114726803467455178939551110155038863261690800635036152735760943636185800678224699322718305930707213041643398454621048125585225782210459408661329977097382164788870672851887421058579613475931754523661776491355121471433477219208766965295977124555417874237514655820531331364209814523227224473519267312485203990286;
            6'd53: xpb[148] = 1024'd26268964380353544435420184554502140549443696209210771117813836927860104098618495875451875157124820527851162319452515387346395009715153383576046231452705291890959615913583212639899431248975561006620897017752044688925549621339818688231107729874508235816329239014456006868443694286956823893192518349037369636165;
            6'd54: xpb[148] = 1024'd61877820977376651330088186358779850581895018909121073627998585284511302856321431338200515598200102323502075591741476083686628078061067693045922610824359459926739233544850221558849488213536573210890215152536207752781982873691767184131216904876828046661963725622497740402784102124615056329984459212215129766375;
            6'd55: xpb[148] = 1024'd97486677574399758224756188163057560614346341609031376138183333641162501614024366800949156039275384119152988864030436780026861146406982002515798990196013627962518851176117230477799545178097585415159533287320370816638416126043715680031326079879147857507598212230539473937124509962273288766776400075392889896585;
            6'd56: xpb[148] = 1024'd9028838487298123720625262562520837902099237183205994520236226932836805034418163353682725265692991605360752728861904041788030373911675977430515244551336755064607794237813022059119362951141391898118653813717294034130488528174767402966456685198238219086412795424464149441358389726002888186449651111945055542464;
            6'd57: xpb[148] = 1024'd44637695084321230615293264366798547934550559883116297030420975289488003792121098816431365706768273401011666001150864738128263442257590286900391623922990923100387411869080030978069419915702404102387971948501457097986921780526715898866565860200558029932047282032505882975698797563661120623241591975122815672674;
            6'd58: xpb[148] = 1024'd80246551681344337509961266171076257967001882583026599540605723646139202549824034279180006147843555196662579273439825434468496510603504596370268003294645091136167029500347039897019476880263416306657290083285620161843355032878664394766675035202877840777681768640547616510039205401319353060033532838300575802884;
            6'd59: xpb[148] = 1024'd115855408278367444404629267975353967999453205282936902050790472002790401307526969741928646588918836992313492545728786130808729578949418905840144382666299259171946647131614048815969533844824428510926608218069783225699788285230612890666784210205197651623316255248589350044379613238977585496825473701478335933094;
            6'd60: xpb[148] = 1024'd27397569191265809900498342374817245287206100857111520432843365294464704727920766294662215815336444478521256410560253392569898806454112880754860637021622386274035590193309840397289351617868234993885728744466706443191860687361664613601914815524288013202130838442514025548613493002707184916498724738030501578973;
            6'd61: xpb[148] = 1024'd63006425788288916795166344179094955319657423557021822943028113651115903485623701757410856256411726274172169682849214088910131874800027190224737016393276554309815207824576849316239408582429247198155046879250869507048293939713613109502023990526607824047765325050555759082953900840365417353290665601208261709183;
            6'd62: xpb[148] = 1024'd98615282385312023689834345983372665352108746256932125453212862007767102243326637220159496697487008069823082955138174785250364943145941499694613395764930722345594825455843858235189465546990259402424365014035032570904727192065561605402133165528927634893399811658597492617294308678023649790082606464386021839393;
            6'd63: xpb[148] = 1024'd10157443298210389185703420382835942639861641831106743835265755299441405663720433772893065923904615556030846819969642047011534170650635474609329650120253849447683768517539649816509283320034065885383485540431955788396799594196613328337263770848017996472214394852522168121528188441753249209755857500938187485272;
        endcase
    end

    always_comb begin
        case(flag[49][16:12])
            5'd0: xpb[149] = 1024'd0;
            5'd1: xpb[149] = 1024'd45766299895233496080371422187113652672312964531017046345450503656092604421423369235641706364979897351681760092258602743351767238996549784079206029491908017483463386148806658735459340284595078089652803675216118852253232846548561824237372945850337807317848881460563901655868596279411481646547798364115947615482;
            5'd2: xpb[149] = 1024'd91532599790466992160742844374227305344625929062034092690901007312185208842846738471283412729959794703363520184517205486703534477993099568158412058983816034966926772297613317470918680569190156179305607350432237704506465693097123648474745891700675614635697762921127803311737192558822963293095596728231895230964;
            5'd3: xpb[149] = 1024'd13232204001575746842315339156526525272240466467315454908219655903300917926960968796910047880282017745602130869318314795476237876148429017682457963459393011516699483876848758868747781662268028547648213417261116710395337689424788699747140267867783972686726740967574646937499260764305811922524705265722248362115;
            5'd4: xpb[149] = 1024'd58998503896809242922686761343640177944553430998332501253670159559393522348384338032551754245261915097283890961576917538828005115144978801761663992951301029000162870025655417604207121946863106637301017092477235562648570535973350523984513213718121780004575622428138548593367857043717293569072503629838195977597;
            5'd5: xpb[149] = 1024'd104764803792042739003058183530753830616866395529349547599120663215486126769807707268193460610241812448965651053835520282179772354141528585840870022443209046483626256174462076339666462231458184726953820767693354414901803382521912348221886159568459587322424503888702450249236453323128775215620301993954143593079;
            5'd6: xpb[149] = 1024'd26464408003151493684630678313053050544480932934630909816439311806601835853921937593820095760564035491204261738636629590952475752296858035364915926918786023033398967753697517737495563324536057095296426834522233420790675378849577399494280535735567945373453481935149293874998521528611623845049410531444496724230;
            5'd7: xpb[149] = 1024'd72230707898384989765002100500166703216793897465647956161889815462694440275345306829461802125543932842886021830895232334304242991293407819444121956410694040516862353902504176472954903609131135184949230509738352273043908225398139223731653481585905752691302363395713195530867117808023105491597208895560444339712;
            5'd8: xpb[149] = 1024'd117997007793618485845373522687280355889106861996665002507340319118787044696768676065103508490523830194567781923153835077656010230289957603523327985902602058000325740051310835208414243893726213274602034184954471125297141071946701047969026427436243560009151244856277097186735714087434587138145007259676391955194;
            5'd9: xpb[149] = 1024'd39696612004727240526946017469579575816721399401946364724658967709902753780882906390730143640846053236806392607954944386428713628445287053047373890378179034550098451630546276606243344986804085642944640251783350131186013068274366099241420803603351918060180222902723940812497782292917435767574115797166745086345;
            5'd10: xpb[149] = 1024'd85462911899960736607317439656693228489034363932963411070109471365995358202306275626371850005825950588488152700213547129780480867441836837126579919870087052033561837779352935341702685271399163732597443926999468983439245914822927923478793749453689725378029104363287842468366378572328917414121914161282692701827;
            5'd11: xpb[149] = 1024'd7162516111069491288889934438992448416648901338244773287428119957111067286420505951998485156148173630726763385014656438553184265597166286650625824345664028583334549358588376739531786364477036100940049993828347989328117911150592974751188125620798083429058082409734686094128446777811766043551022698773045832978;
            5'd12: xpb[149] = 1024'd52928816006302987369261356626106101088961865869261819632878623613203671707843875187640191521128070982408523477273259181904951504593716070729831853837572046066797935507395035474991126649072114190592853669044466841581350757699154798988561071471135890746906963870298587749997043057223247690098821062888993448460;
            5'd13: xpb[149] = 1024'd98695115901536483449632778813219753761274830400278865978329127269296276129267244423281897886107968334090283569531861925256718743590265854809037883329480063550261321656201694210450466933667192280245657344260585693834583604247716623225934017321473698064755845330862489405865639336634729336646619427004941063942;
            5'd14: xpb[149] = 1024'd20394720112645238131205273595518973688889367805560228195647775860411985213381474748908533036430191376328894254332971234029422141745595304333083787805057040100034033235437135608279568026745064648588263411089464699723455600575381674498328393488582056115784823377309333031627707542117577966075727964495294195093;
            5'd15: xpb[149] = 1024'd66161020007878734211576695782632626361202332336577274541098279516504589634804843984550239401410088728010654346591573977381189380742145088412289817296965057583497419384243794343738908311340142738241067086305583551976688447123943498735701339338919863433633704837873234687496303821529059612623526328611241810575;
            5'd16: xpb[149] = 1024'd111927319903112230291948117969746279033515296867594320886548783172597194056228213220191945766389986079692414438850176720732956619738694872491495846788873075066960805533050453079198248595935220827893870761521702404229921293672505322973074285189257670751482586298437136343364900100940541259171324692727189426057;
            5'd17: xpb[149] = 1024'd33626924114220984973520612752045498961129834272875683103867431763712903140342443545818580916712209121931025123651286029505660017894024322015541751264450051616733517112285894477027349689013093196236476828350581410118793290000170374245468661356366028802511564344883979969126968306423389888600433230217542557208;
            5'd18: xpb[149] = 1024'd79393224009454481053892034939159151633442798803892729449317935419805507561765812781460287281692106473612785215909888772857427256890574106094747780756358069100196903261092553212486689973608171285889280503566700262372026136548732198482841607206703836120360445805447881624995564585834871535148231594333490172690;
            5'd19: xpb[149] = 1024'd1092828220563235735464529721458371561057336209174091666636584010921216645880043107086922432014329515851395900710998081630130655045903555618793685231935045649969614840327994610315791066686043654231886570395579268260898132876397249755235983373812194171389423851894725250757632791317720164577340131823843303841;
            5'd20: xpb[149] = 1024'd46859128115796731815835951908572024233370300740191138012087087667013821067303412342728628796994226867533155992969600824981897894042453339697999714723843063133433000989134653345775131351281121743884690245611698120514130979424959073992608929224150001489238305312458626906626229070729201811125138495939790919323;
            5'd21: xpb[149] = 1024'd92625428011030227896207374095685676905683265271208184357537591323106425488726781578370335161974124219214916085228203568333665133039003123777205744215751080616896387137941312081234471635876199833537493920827816972767363825973520898229981875074487808807087186773022528562494825350140683457672936860055738534805;
            5'd22: xpb[149] = 1024'd14325032222138982577779868877984896833297802676489546574856239914222134572841011903996970312296347261453526770029312877106368531194332573301251648691328057166669098717176753479063572728954072201880099987656695978656235822301185949502376251241596166858116164819469372188256893555623532087102045397546091665956;
            5'd23: xpb[149] = 1024'd60091332117372478658151291065098549505610767207506592920306743570314738994264381139638676677276244613135286862287915620458135770190882357380457678183236074650132484865983412214522913013549150291532903662872814830909468668849747773739749197091933974175965046280033273844125489835035013733649843761662039281438;
            5'd24: xpb[149] = 1024'd105857632012605974738522713252212202177923731738523639265757247226407343415687750375280383042256141964817046954546518363809903009187432141459663707675144092133595871014790070949982253298144228381185707338088933683162701515398309597977122142942271781493813927740597175499994086114446495380197642125777986896920;
            5'd25: xpb[149] = 1024'd27557236223714729420095208034511422105538269143805001483075895817523052499801980700907018192578365007055657639347627672582606407342761590983709612150721068683368582594025512347811354391222100749528313404917812689051573511725974649249516519109380139544842905787044019125756154319929344009626750663268340028071;
            5'd26: xpb[149] = 1024'd73323536118948225500466630221625074777851233674822047828526399473615656921225349936548724557558262358737417731606230415934373646339311375062915641642629086166831968742832171083270694675817178839181117080133931541304806358274536473486889464959717946862691787247607920781624750599340825656174549027384287643553;
            5'd27: xpb[149] = 1024'd119089836014181721580838052408738727450164198205839094173976903129708261342648719172190430922538159710419177823864833159286140885335861159142121671134537103650295354891638829818730034960412256928833920755350050393558039204823098297724262410810055754180540668708171822437493346878752307302722347391500235259035;
            5'd28: xpb[149] = 1024'd40789440225290476262410547191037947377778735611120456391295551720823970426762949497817066072860382752657788508665942468058844283491190608666167575610114080200068066470874271216559136053490129297176526822178929399446911201150763348996656786977164112231569646754618666063255415084235155932151455928990588390186;
            5'd29: xpb[149] = 1024'd86555740120523972342781969378151600050091700142137502736746055376916574848186318733458772437840280104339548600924545211410611522487740392745373605102022097683531452619680929952018476338085207386829330497395048251700144047699325173234029732827501919549418528215182567719124011363646637578699254293106536005668;
            5'd30: xpb[149] = 1024'd8255344331632727024354464160450819977706237547418864954064703968032283932300549059085407588162503146578159285725654520183314920643069842269419509577599074233304164198916371349847577431163079755171936564223927257589016044026990224506424108994610277600447506261629411344886079569129486208128362830596889136819;
            5'd31: xpb[149] = 1024'd54021644226866223104725886347564472650019202078435911299515207624124888353723918294727113953142400498259919377984257263535082159639619626348625539069507091716767550347723030085306917715758157844824740239440046109842248890575552048743797054844948084918296387722193313000754675848540967854676161194712836752301;
        endcase
    end

    always_comb begin
        case(flag[50][5:0])
            6'd0: xpb[150] = 1024'd0;
            6'd1: xpb[150] = 1024'd111927319903112230291948117969746279033515296867594320886548783172597194056228213220191945766389986079692414438850176720732956619738694872491495846788873075066960805533050453079198248595935220827893870761521702404229921293672505322973074285189257670751482586298437136343364900100940541259171324692727189426057;
            6'd2: xpb[150] = 1024'd99787944122099719185097308534678125322332166609452957644965711280217492775147287530368820318122297849941679470242860006886849398636169410427831568561415109200230936496529688820766258000353235934477543914656164962095481737124113872981170000695285892236145269182757214656623272127952449501223959558828784367783;
            6'd3: xpb[150] = 1024'd87648568341087208078246499099609971611149036351311594403382639387837791494066361840545694869854609620190944501635543293040742177533643948364167290333957143333501067460008924562334267404771251041061217067790627519961042180575722422989265716201314113720807952067077292969881644154964357743276594424930379309509;
            6'd4: xpb[150] = 1024'd75509192560074696971395689664541817899965906093170231161799567495458090212985436150722569421586921390440209533028226579194634956431118486300503012106499177466771198423488160303902276809189266147644890220925090077826602624027330972997361431707342335205470634951397371283140016181976265985329229291031974251235;
            6'd5: xpb[150] = 1024'd63369816779062185864544880229473664188782775835028867920216495603078388931904510460899443973319233160689474564420909865348527735328593024236838733879041211600041329386967396045470286213607281254228563374059552635692163067478939523005457147213370556690133317835717449596398388208988174227381864157133569192961;
            6'd6: xpb[150] = 1024'd51230440998049674757694070794405510477599645576887504678633423710698687650823584771076318525051544930938739595813593151502420514226067562173174455651583245733311460350446631787038295618025296360812236527194015193557723510930548073013552862719398778174796000720037527909656760236000082469434499023235164134687;
            6'd7: xpb[150] = 1024'd39091065217037163650843261359337356766416515318746141437050351818318986369742659081253193076783856701188004627206276437656313293123542100109510177424125279866581591313925867528606305022443311467395909680328477751423283954382156623021648578225426999659458683604357606222915132263011990711487133889336759076413;
            6'd8: xpb[150] = 1024'd26951689436024652543992451924269203055233385060604778195467279925939285088661733391430067628516168471437269658598959723810206072021016638045845899196667313999851722277405103270174314426861326573979582833462940309288844397833765173029744293731455221144121366488677684536173504290023898953539768755438354018139;
            6'd9: xpb[150] = 1024'd14812313655012141437141642489201049344050254802463414953884208033559583807580807701606942180248480241686534689991643009964098850918491175982181620969209348133121853240884339011742323831279341680563255986597402867154404841285373723037840009237483442628784049372997762849431876317035807195592403621539948959865;
            6'd10: xpb[150] = 1024'd2672937873999630330290833054132895632867124544322051712301136141179882526499882011783816731980792011935799721384326296117991629815965713918517342741751382266391984204363574753310333235697356787146929139731865425019965284736982273045935724743511664113446732257317841162690248344047715437645038487641543901591;
            6'd11: xpb[150] = 1024'd114600257777111860622238951023879174666382421411916372598849919313777076582728095231975762498370778091628214160234503016850948249554660586410013189530624457333352789737414027832508581831632577615040799901253567829249886578409487596019010009932769334864929318555754977506055148444988256696816363180368733327648;
            6'd12: xpb[150] = 1024'd102460881996099349515388141588811020955199291153775009357266847421397375301647169542152637050103089861877479191627186303004841028452135124346348911303166491466622920700893263574076591236050592721624473054388030387115447021861096146027105725438797556349592001440075055819313520472000164938868998046470328269374;
            6'd13: xpb[150] = 1024'd90321506215086838408537332153742867244016160895633646115683775529017674020566243852329511601835401632126744223019869589158733807349609662282684633075708525599893051664372499315644600640468607828208146207522492944981007465312704696035201440944825777834254684324395134132571892499012073180921632912571923211100;
            6'd14: xpb[150] = 1024'd78182130434074327301686522718674713532833030637492282874100703636637972739485318162506386153567713402376009254412552875312626586247084200219020354848250559733163182627851735057212610044886622934791819360656955502846567908764313246043297156450853999318917367208715212445830264526023981422974267778673518152826;
            6'd15: xpb[150] = 1024'd66042754653061816194835713283606559821649900379350919632517631744258271458404392472683260705300025172625274285805236161466519365144558738155356076620792593866433313591330970798780619449304638041375492513791418060712128352215921796051392871956882220803580050093035290759088636553035889665026902644775113094552;
            6'd16: xpb[150] = 1024'd53903378872049305087984903848538406110466770121209556390934559851878570177323466782860135257032336942874539317197919447620412144042033276091691798393334627999703444554810206540348628853722653147959165666925880618577688795667530346059488587462910442288242732977355369072347008580047797907079537510876708036278;
            6'd17: xpb[150] = 1024'd41764003091036793981134094413470252399283639863068193149351487959498868896242541093037009808764648713123804348590602733774304922939507814028027520165876662132973575518289442281916638258140668254542838820060343176443249239119138896067584302968938663772905415861675447385605380607059706149132172376978302978004;
            6'd18: xpb[150] = 1024'd29624627310024282874283284978402098688100509604926829907768416067119167615161615403213884360496960483373069379983286019928197701836982351964363241938418696266243706481768678023484647662558683361126511973194805734308809682570747446075680018474966885257568098745995525698863752634071614391184807243079897919730;
            6'd19: xpb[150] = 1024'd17485251529011771767432475543333944976917379346785466666185344174739466334080689713390758912229272253622334411375969306082090480734456889900698963710960730399513837445247913765052657066976698467710185126329268292174370126022355996083775733980995106742230781630315604012122124661083522633237442109181492861456;
            6'd20: xpb[150] = 1024'd5345875747999260660581666108265791265734249088644103424602272282359765052999764023567633463961584023871599442768652592235983259631931427837034685483502764532783968408727149506620666471394713574293858279463730850039930569473964546091871449487023328226893464514635682325380496688095430875290076975283087803182;
            6'd21: xpb[150] = 1024'd117273195651111490952529784078012070299249545956238424311151055454956959109227977243759579230351570103564013881618829312968939879370626300328530532272375839599744773941777602585818915067329934402187729040985433254269851863146469869064945734676280998978376050813072818668745396789035972134461401668010277229239;
            6'd22: xpb[150] = 1024'd105133819870098979845678974642943916588066415698097061069567983562577257828147051553936453782083881873813278913011512599122832658268100838264866254044917873733014904905256838327386924471747949508771402194119895812135412306598078419073041450182309220463038733697392896982003768816047880376514036534111872170965;
            6'd23: xpb[150] = 1024'd92994444089086468738828165207875762876883285439955697827984911670197556547066125864113328333816193644062543944404195885276725437165575376201201975817459907866285035868736074068954933876165964615355075347254358370000972750049686969081137165688337441947701416581712975295262140843059788618566671400213467112691;
            6'd24: xpb[150] = 1024'd80855068308073957631977355772807609165700155181814334586401839777817855265985200174290202885548505414311808975796879171430618216063049914137537697590001941999555166832215309810522943280583979721938748500388820927866533193501295519089232881194365663432364099466033053608520512870071696860619306266315062054417;
            6'd25: xpb[150] = 1024'd68715692527061446525126546337739455454517024923672971344818767885438153984904274484467077437280817184561074007189562457584510994960524452073873419362543976132825297795694545552090952685001994828522421653523283485732093636952904069097328596700393884917026782350353131921778884897083605102671941132416656996143;
            6'd26: xpb[150] = 1024'd56576316746048935418275736902671301743333894665531608103235695993058452703823348794643951989013128954810339038582245743738403773857998990010209141135086010266095428759173781293658962089420009935106094806657746043597654080404512619105424312206422106401689465234673210235037256924095513344724575998518251937869;
            6'd27: xpb[150] = 1024'd44436940965036424311424927467603148032150764407390244861652624100678751422742423104820826540745440725059604069974929029892296552755473527946544862907628044399365559722653017035226971493838025041689767959792208601463214523856121169113520027712450327886352148118993288548295628951107421586777210864619846879595;
            6'd28: xpb[150] = 1024'd32297565184023913204574118032534994320967634149248881620069552208299050141661497414997701092477752495308869101367612316046189331652948065882880584680170078532635690686132252776794980898256040148273441112926671159328774967307729719121615743218478549371014831003313366861554000978119329828829845730721441821321;
            6'd29: xpb[150] = 1024'd20158189403011402097723308597466840609784503891107518378486480315919348860580571725174575644210064265558134132760295602200082110550422603819216306452712112665905821649611488518362990302674055254857114266061133717194335410759338269129711458724506770855677513887633445174812373005131238070882480596823036763047;
            6'd30: xpb[150] = 1024'd8018813621998890990872499162398686898601373632966155136903408423539647579499646035351450195942376035807399164152978888353974889447897141755552028225254146799175952613090724259930999707092070361440787419195596275059895854210946819137807174230534992340340196771953523488070745032143146312935115462924631704773;
            6'd31: xpb[150] = 1024'd119946133525111121282820617132144965932116670500560476023452191596136841635727859255543395962332362115499813603003155609086931509186592014247047875014127221866136758146141177339129248303027291189334658180717298679289817147883452142110881459419792663091822783070390659831435645133083687572106440155651821130830;
            6'd32: xpb[150] = 1024'd107806757744098610175969807697076812220933540242419112781869119703757140354646933565720270514064673885749078634395838895240824288084066552183383596786669255999406889109620413080697257707445306295918331333851761237155377591335060692118977174925820884576485465954710738144694017160095595814159075021753416072556;
            6'd33: xpb[150] = 1024'd95667381963086099069118998262008658509750409984277749540286047811377439073566007875897145065796985655998343665788522181394717066981541090119719318559211290132677020073099648822265267111863321402502004486986223795020938034786669242127072890431849106061148148839030816457952389187107504056211709887855011014282;
            6'd34: xpb[150] = 1024'd83528006182073587962268188826940504798567279726136386298702975918997737792485082186074019617529297426247608697181205467548609845879015628056055040331753324265947151036578884563833276516281336509085677640120686352886498478238277792135168605937877327545810831723350894771210761214119412298264344753956605956008;
            6'd35: xpb[150] = 1024'd71388630401061076855417379391872351087384149467995023057119904026618036511404156496250894169261609196496873728573888753702502624776490165992390762104295358399217282000058120305401285920699351615669350793255148910752058921689886342143264321443905549030473514607670973084469133241131320540316979620058200897734;
            6'd36: xpb[150] = 1024'd59249254620048565748566569956804197376201019209853659815536832134238335230323230806427768720993920966746138759966572039856395403673964703928726483876837392532487412963537356046969295325117366722253023946389611468617619365141494892151360036949933770515136197491991051397727505268143228782369614486159795839460;
            6'd37: xpb[150] = 1024'd47109878839036054641715760521736043665017888951712296573953760241858633949242305116604643272726232736995403791359255326010288182571439241865062205649379426665757543927016591788537304729535381828836697099524074026483179808593103442159455752455961991999798880376311129710985877295155137024422249352261390781186;
            6'd38: xpb[150] = 1024'd34970503058023543534864951086667889953834758693570933332370688349478932668161379426781517824458544507244668822751938612164180961468913779801397927421921460799027674890495827530105314133953396935420370252658536584348740252044711992167551467961990213484461563260631208024244249322167045266474884218362985722912;
            6'd39: xpb[150] = 1024'd22831127277011032428014141651599736242651628435429570090787616457099231387080453736958392376190856277493933854144621898318073740366388317737733649194463494932297805853975063271673323538371412042004043405792999142214300695496320542175647183468018434969124246144951286337502621349178953508527519084464580664638;
            6'd40: xpb[150] = 1024'd10691751495998521321163332216531582531468498177288206849204544564719530105999528047135266927923168047743198885537305184471966519263862855674069370967005529065567936817454299013241332942789427148587716558927461700079861138947929092183742898974046656453786929029271364650760993376190861750580153950566175606364;
            6'd41: xpb[150] = 1024'd122619071399110751613111450186277861564983795044882527735753327737316724162227741267327212694313154127435613324387481905204923139002557728165565217755878604132528742350504752092439581538724647976481587320449164104309782432620434415156817184163304327205269515327708500994125893477131403009751478643293365032421;
            6'd42: xpb[150] = 1024'd110479695618098240506260640751209707853800664786741164494170255844937022881146815577504087246045465897684878355780165191358815917900032266101900939528420638265798873313983987834007590943142663083065260473583626662175342876072042965164912899669332548689932198212028579307384265504143311251804113509394959974147;
            6'd43: xpb[150] = 1024'd98340319837085729399409831316141554142617534528599801252587183952557321600065889887680961797777777667934143387172848477512708696797506804038236661300962672399069004277463223575575600347560678189648933626718089220040903319523651515173008615175360770174594881096348657620642637531155219493856748375496554915873;
            6'd44: xpb[150] = 1024'd86200944056073218292559021881073400431434404270458438011004112060177620318984964197857836349510089438183408418565531763666601475694981341974572383073504706532339135240942459317143609751978693296232606779852551777906463762975260065181104330681388991659257563980668735933901009558167127735909383241598149857599;
            6'd45: xpb[150] = 1024'd74061568275060707185708212446005246720251274012317074769421040167797919037904038508034710901242401208432673449958215049820494254592455879910908104846046740665609266204421695058711619156396708402816279932987014335772024206426868615189200046187417213143920246864988814247159381585179035977962018107699744799325;
            6'd46: xpb[150] = 1024'd61922192494048196078857403010937093009068143754175711527837968275418217756823112818211585452974712978681938481350898335974387033489930417847243826618588774798879397167900930800279628560814723509399953086121476893637584649878477165197295761693445434628582929749308892560417753612190944220014652973801339741051;
            6'd47: xpb[150] = 1024'd49782816713035684972006593575868939297885013496034348286254896383038516475742187128388460004707024748931203512743581622128279812387404955783579548391130808932149528131380166541847637965232738615983626239255939451503145093330085715205391477199473656113245612633628970873676125639202852462067287839902934682777;
            6'd48: xpb[150] = 1024'd37643440932023173865155784140800785586701883237892985044671824490658815194661261438565334556439336519180468544136264908282172591284879493719915270163672843065419659094859402283415647369650753722567299392390402009368705536781694265213487192705501877597908295517949049186934497666214760704119922706004529624503;
            6'd49: xpb[150] = 1024'd25504065151010662758304974705732631875518752979751621803088752598279113913580335748742209108171648289429733575528948194436065370182354031656250991936214877198689790058338638024983656774068768829150972545524864567234265980233302815221582908211530099082570978402269127500192869693226668946172557572106124566229;
            6'd50: xpb[150] = 1024'd13364689369998151651454165270664478164335622721610258561505680705899412632499410058919083659903960059678998606921631480589958149079828569592586713708756911331959921021817873766551666178486783935734645698659327125099826423684911365229678623717558320567233661286589205813451241720238577188225192438207719507955;
            6'd51: xpb[150] = 1024'd1225313588985640544603355835596324453152492463468895319922608813519711351418484369095958211636271829928263638314314766743850927977303107528922435481298945465230051985297109508119675582904799042318318851793789682965386867136519915237774339223586542051896344170909284126709613747250485430277827304309314449681;
            6'd52: xpb[150] = 1024'd113152633492097870836551473805342603486667789331063216206471391986116905407646697589287903978026257909620678077164491487476807547715997980020418282270172020532190857518347562587317924178840019870212189613315492087195308160809025238210848624412844212803378930469346420470074513848191026689449151997036503875738;
            6'd53: xpb[150] = 1024'd101013257711085359729700664370274449775484659072921852964888320093737204126565771899464778529758569679869943108557174773630700326613472517956754004042714054665460988481826798328885933583258034976795862766449954645060868604260633788218944339918872434288041613353666498783332885875202934931501786863138098817464;
            6'd54: xpb[150] = 1024'd88873881930072848622849854935206296064301528814780489723305248201357502845484846209641653081490881450119208139949858059784593105510947055893089725815256088798731119445306034070453942987676050083379535919584417202926429047712242338227040055424900655772704296237986577096591257902214843173554421729239693759190;
            6'd55: xpb[150] = 1024'd76734506149060337515999045500138142353118398556639126481722176308977801564403920519818527633223193220368473171342541345938485884408421593829425447587798122932001250408785269812021952392094065189963209072718879760791989491163850888235135770930928877257366979122306655409849629929226751415607056595341288700916;
            6'd56: xpb[150] = 1024'd64595130368047826409148236065069988641935268298497763240139104416598100283322994829995402184955504990617738202735224632092378663305896131765761169360340157065271381372264505553589961796512080296546882225853342318657549934615459438243231486436957098742029662006626733723108001956238659657659691461442883642642;
            6'd57: xpb[150] = 1024'd52455754587035315302297426630001834930752138040356399998556032524218399002242069140172276736687816760867003234127907918246271442203370669702096891132882191198541512335743741295157971200930095403130555378987804876523110378067067988251327201942985320226692344890946812036366373983250567899712326327544478584368;
            6'd58: xpb[150] = 1024'd40316378806022804195446617194933681219569007782215036756972960631838697721161143450349151288420128531116268265520591204400164221100845207638432612905424225331811643299222977036725980605348110509714228532122267434388670821518676538259422917449013541711355027775266890349624746010262476141764961193646073526094;
            6'd59: xpb[150] = 1024'd28177003025010293088595807759865527508385877524073673515389888739458996440080217760526025840152440301365533296913274490554056999998319745574768334677966259465081774262702212778293990009766125616297901685256729992254231264970285088267518632955041763196017710659586968662883118037274384383817596059747668467820;
            6'd60: xpb[150] = 1024'd16037627243997781981744998324797373797202747265932310273806816847079295158999292070702900391884752071614798328305957776707949778895794283511104056450508293598351905226181448519861999414184140722881574838391192550119791708421893638275614348461069984680680393543907046976141490064286292625870230925849263409546;
            6'd61: xpb[150] = 1024'd3898251462985270874894188889729220086019617007790947032223744954699593877918366380879774943617063841864063359698641062861842557793268821447439778223050327731622036189660684261430008818602155829465247991525655107985352151873502188283710063967098206165343076428227125289399862091298200867922865791950858351272;
            6'd62: xpb[150] = 1024'd115825571366097501166842306859475499119534913875385267918772528127296787934146579601071720710007049921556477798548817783594799177531963693938935625011923402798582841722711137340628257414537376657359118753047357512215273445546007511256784349156355876916825662726664261632764762192238742127094190484678047777329;
            6'd63: xpb[150] = 1024'd103686195585084990059991497424407345408351783617243904677189456234917086653065653911248595261739361691805742829941501069748691956429438231875271346784465436931852972686190373082196266818955391763942791906181820070080833888997616061264880064662384098401488345610984339946023134219250650369146825350779642719055;
        endcase
    end

    always_comb begin
        case(flag[50][11:6])
            6'd0: xpb[151] = 1024'd0;
            6'd1: xpb[151] = 1024'd91546819804072478953140687989339191697168653359102541435606384342537385371984728221425469813471673462055007861334184355902584735326912769811607068557007471065123103649669608823764276223373406870526465059316282627946394332449224611272975780168412319886151028495304418259281506246262558611199460216881237660781;
            6'd2: xpb[151] = 1024'd59026943924020216507482448573863950649638879592469398743080913620097875406660317532835868412285672614666866315210875277226105629812605205068054012097683901196555532729768000309898313255229608019742732510245325409528427814677552449580972990653595190505482153576491778488456484418596484205280230607136880837231;
            6'd3: xpb[151] = 1024'd26507068043967954061824209158388709602109105825836256050555442897658365441335906844246267011099671767278724769087566198549626524298297640324500955638360331327987961809866391796032350287085809168958999961174368191110461296905880287888970201138778061124813278657679138717631462590930409799361000997392524013681;
            6'd4: xpb[151] = 1024'd118053887848040433014964897147727901299277759184938797486161827240195750813320635065671736824571345229333732630421750554452211259625210410136108024195367802393111065459536000619796626510459216039485465020490650819056855629355104899161945981307190381010964307152983556976912968837192968410560461214273761674462;
            6'd5: xpb[151] = 1024'd85534011967988170569306657732252660251747985418305654793636356517756240847996224377082135423385344381945591084298441475775732154110902845392554967736044232524543494539634392105930663542315417188701732471419693600638889111583432737469943191792373251630295432234170917206087947009526894004641231604529404850912;
            6'd6: xpb[151] = 1024'd53014136087935908123648418316777419204218211651672512101110885795316730882671813688492534022199343534557449538175132397099253048596595280649001911276720662655975923619732783592064700574171618337917999922348736382220922593811760575777940402277556122249626557315358277435262925181860819598722001994785048027362;
            6'd7: xpb[151] = 1024'd20494260207883645677990178901302178156688437885039369408585415072877220917347402999902932621013342687169307992051823318422773943082287715905448854817397092787408352699831175078198737606027819487134267373277779163802956076040088414085937612762738992868957682396545637664437903354194745192802772385040691203812;
            6'd8: xpb[151] = 1024'd112041080011956124631130866890641369853857091244141910844191799415414606289332131221328402434485016149224315853386007674325358678409200485717055923374404563852531456349500783901963013829401226357660732432594061791749350408489313025358913392931151312755108710891850055923719409600457303804002232601921928864593;
            6'd9: xpb[151] = 1024'd79521204131903862185472627475166128806327317477508768151666328692975096324007720532738801033299015301836174307262698595648879572894892920973502866915080993983963885429599175388097050861257427506876999883523104573331383890717640863666910603416334183374439835973037416152894387772791229398083002992177572041043;
            6'd10: xpb[151] = 1024'd47001328251851599739814388059690887758797543710875625459140857970535586358683309844149199632113014454448032761139389516972400467380585356229949810455757424115396314509697566874231087893113628656093267334452147354913417372945968701974907813901517053993770961054224776382069365945125154992163773382433215217493;
            6'd11: xpb[151] = 1024'd14481452371799337294156148644215646711267769944242482766615387248096076393358899155559598230927013607059891215016080438295921361866277791486396753996433854246828743589795958360365124924969829805309534785381190136495450855174296540282905024386699924613102086135412136611244344117459080586244543772688858393943;
            6'd12: xpb[151] = 1024'd106028272175871816247296836633554838408436423303345024202221771590633461765343627376985068044398687069114899076350264794198506097193190561298003822553441325311951847239465567184129401148343236675835999844697472764441845187623521151555880804555112244499253114630716554870525850363721639197444003989570096054724;
            6'd13: xpb[151] = 1024'd73508396295819553801638597218079597360906649536711881509696300868193951800019216688395466643212686221726757530226955715522026991678882996554450766094117755443384276319563958670263438180199437825052267295626515546023878669851848989863878015040295115118584239711903915099700828536055564791524774379825739231174;
            6'd14: xpb[151] = 1024'd40988520415767291355980357802604356313376875770078738817170830145754441834694805999805865242026685374338615984103646636845547886164575431810897709634794185574816705399662350156397475212055638974268534746555558327605912152080176828171875225525477985737915364793091275328875806708389490385605544770081382407624;
            6'd15: xpb[151] = 1024'd8468644535715028910322118387129115265847102003445596124645359423314931869370395311216263840840684526950474437980337558169068780650267867067344653175470615706249134479760741642531512243911840123484802197484601109187945634308504666479872436010660856357246489874278635558050784880723415979686315160337025584074;
            6'd16: xpb[151] = 1024'd100015464339787507863462806376468306963015755362548137560251743765852317241355123532641733654312357989005482299314521914071653515977180636878951721732478086771372238129430350466295788467285246994011267256800883737134339966757729277752848216179073176243397518369583053817332291126985974590885775377218263244855;
            6'd17: xpb[151] = 1024'd67495588459735245417804566960993065915485981595914994867726273043412807276030712844052132253126357141617340753191212835395174410462873072135398665273154516902804667209528741952429825499141448143227534707729926518716373448986057116060845426664256046862728643450770414046507269299319900184966545767473906421305;
            6'd18: xpb[151] = 1024'd34975712579682982972146327545517824867956207829281852175200802320973297310706302155462530851940356294229199207067903756718695304948565507391845608813830947034237096289627133438563862530997649292443802158658969300298406931214384954368842637149438917482059768531957774275682247471653825779047316157729549597755;
            6'd19: xpb[151] = 1024'd2455836699630720526488088130042583820426434062648709482675331598533787345381891466872929450754355446841057660944594678042216199434257942648292552354507377165669525369725524924697899562853850441660069609588012081880440413442712792676839847634621788101390893613145134504857225643987751373128086547985192774205;
            6'd20: xpb[151] = 1024'd94002656503703199479628776119381775517595087421751250918281715941071172717366619688298399264226028908896065522278779033944800934761170712459899620911514848230792629019395133748462175786227257312186534668904294709826834745891937403949815627803034107987541922108449552764138731890250309984327546764866430434986;
            6'd21: xpb[151] = 1024'd61482780623650937033970536703906534470065313655118108225756245218631662752042208999708797863040028061507923976155469955268321829246863147716346564452191278362225058099493525234596212818083458461402802119833337491408868228120265242257812838288216978606873047189636912993313710062584235578408317155122073611436;
            6'd22: xpb[151] = 1024'd28962904743598674588312297288431293422535539888484965533230774496192152786717798311119196461854027214119782430032160876591842723732555582972793507992867708493657487179591916720730249849939659610619069570762380272990901710348593080565810048773399849226204172270824273222488688234918161172489087545377716787886;
            6'd23: xpb[151] = 1024'd120509724547671153541452985277770485119704193247587506968837158838729538158702526532544666275325700676174790291366345232494427459059468352784400576549875179558780590829261525544494526073313066481145534630078662900937296042797817691838785828941812169112355200766128691481770194481180719783688547762258954448667;
            6'd24: xpb[151] = 1024'd87989848667618891095794745862295244072174419480954364276311688116290028193378115843955064874139699828786648745243036153817948353545160788040847520090551609690213019909359917030628563105169267630361802081007705682519329525026145530146783039426995039731686325847316051710945172653514645377769318152514597625117;
            6'd25: xpb[151] = 1024'd55469972787566628650136506446820003024644645714321221583786217393850518228053705155365463472953698981398507199119727075141469248030853223297294463631228039821645448989458308516762600137025468779578069531936748464101363007254473368454780249912177910351017450928503411940120150825848570971850088542770240801567;
            6'd26: xpb[151] = 1024'd22950096907514366204478267031344761977114871947688078891260746671411008262729294466775862071767698134010365652996417996464990142516545658553741407171904469953077878069556700002896637168881669928794336982865791245683396489482801206762777460397360780970348576009690772169295128998182496565930858933025883978017;
            6'd27: xpb[151] = 1024'd114496916711586845157618955020683953674283525306790620326867131013948393634714022688201331885239371596065373514330602352367574877843458428365348475728911941018200981719226308826660913392255076799320802042182073873629790821932025818035753240565773100856499604504995190428576635244445055177130319149907121638798;
            6'd28: xpb[151] = 1024'd81977040831534582711960715605208712626753751540157477634341660291508883669389611999611730484053370748677231968207293273691095772329150863621795419269588371149633410799324700312794950424111277948537069493111116655211824304160353656343750451050955971475830729586182550657751613416778980771211089540162764815248;
            6'd29: xpb[151] = 1024'd49457164951482320266302476189733471579223977773524334941816189569069373704065201311022129082867369901289090422083984195014616666814843298878242362810264801281065839879423091798928987455967479097753336944040159436793857786388681494651747661536138842095161854667369910886926591589112906365291859930418407991698;
            6'd30: xpb[151] = 1024'd16937289071430057820644236774258230531694204006891192249290718846629863738740790622432527681681369053900948875960675116338137561300535734134689306350941231412498268959521483285063024487823680246969604394969202218375891268617009332959744872021321712714492979748557271116101569761446831959372630320674051168148;
            6'd31: xpb[151] = 1024'd108484108875502536773784924763597422228862857365993733684897103189167249110725518843857997495153042515955956737294859472240722296627448503946296374907948702477621372609191092108827300711197087117496069454285484846322285601066233944232720652189734032600644008243861689375383076007709390570572090537555288828929;
            6'd32: xpb[151] = 1024'd75964232995450274328126685348122181181333083599360590992371632466727739145401108155268396093967041668567815191171550393564243191113140939202743318448625132609053801689289483594961337743053288266712336905214527627904319083294561782540717862674916903219975133325049049604558054180043316164652860927810932005379;
            6'd33: xpb[151] = 1024'd43444357115398011882468445932646940133803309832727448299846161744288229180076697466678794692781040821179673645048241314887764085598833374459190261989301562740486230769387875081095374774909489415928604356143570409486352565522889620848715073160099773839306258406236409833733032352377241758733631318066575181829;
            6'd34: xpb[151] = 1024'd10924481235345749436810206517171699086273536066094305607320691021848719214752286778089193291595039973791532098924932236211284980084525809715637205529977992871918659849486266567229411806765690565144871807072613191068386047751217459156712283645282644458637383487423770062908010524711167352814401708322218358279;
            6'd35: xpb[151] = 1024'd102471301039418228389950894506510890783442189425196847042927075364386104586737014999514663105066713435846539960259116592113869715411438579527244274086985463937041763499155875390993688030139097435671336866388895819014780380200442070429688063813694964344788411982728188322189516770973725964013861925203456019060;
            6'd36: xpb[151] = 1024'd69951425159365965944292655091035649735912415658563704350401604641946594621412604310925061703880712588458398414135807513437390609897131014783691217627661894068474192579254266877127725061995298584887604317317938600596813862428769908737685274298877834964119537063915548551364494943307651558094632315459099195510;
            6'd37: xpb[151] = 1024'd37431549279313703498634415675560408688382641891930561657876133919507084656088193622335460302694711741070256868012498434760911504382823450040138161168338324199906621659352658363261762093851499734103871768246981382178847344657097747045682484784060705583450662145102908780539473115641577152175402705714742371960;
            6'd38: xpb[151] = 1024'd4911673399261441052976176260085167640852868125297418965350663197067574690763782933745858901508710893682115321889189356084432398868515885296585104709014754331339050739451049849395799125707700883320139219176024163760880826885425585353679695269243576202781787226290269009714451287975502746256173095970385548410;
            6'd39: xpb[151] = 1024'd96458493203333920006116864249424359338021521484399960400957047539604960062748511155171328714980384355737123183223373711987017134195428655108192173266022225396462154389120658673160075349081107753846604278492306791707275159334650196626655475437655896088932815721594687268995957534238061357455633312851623209191;
            6'd40: xpb[151] = 1024'd63938617323281657560458624833949118290491747717766817708431576817165450097424100466581727313794383508348981637100064633310538028681121090364639116806698655527894583469219050159294112380937308903062871729421349573289308641562978034934652685922838766708263940802782047498170935706571986951536403703107266385641;
            6'd41: xpb[151] = 1024'd31418741443229395114800385418473877242961973951133675015906106094725940132099689777992125912608382660960840090976755554634058923166813525621086060347375085659327012549317441645428149412793510052279139180350392354871342123791305873242649896408021637327595065883969407727345913878905912545617174093362909562091;
            6'd42: xpb[151] = 1024'd122965561247301874067941073407813068940130627310236216451512490437263325504084417999417595726080056123015847952310939910536643658493726295432693128904382556724450116198987050469192425636166916922805604239666674982817736456240530484515625676576433957213746094379273825986627420125168471156816634310244147222872;
            6'd43: xpb[151] = 1024'd90445685367249611622282833992337827892600853543603073758987019714823815538760007310827994324894055275627706406187630831860164552979418730689140072445058986855882545279085441955326462668023118072021871690595717764399769938468858322823622887061616827833077219460461186215802398297502396750897404700499790399322;
            6'd44: xpb[151] = 1024'd57925809487197349176624594576862586845071079776969931066461548992384305573435596622238392923708054428239564860064321753183685447465111165945587015985735416987314974359183833441460499699879319221238139141524760545981803420697186161131620097546799698452408344541648546444977376469836322344978175090755433575772;
            6'd45: xpb[151] = 1024'd25405933607145086730966355161387345797541306010336788373936078269944795608111185933648791522522053580851423313941012674507206341950803601202033959526411847118747403439282224927594536731735520370454406592453803327563836902925513999439617308031982569071739469622835906674152354642170247939058945481011076752222;
            6'd46: xpb[151] = 1024'd116952753411217565684107043150726537494709959369439329809542462612482180980095914155074261335993727042906431175275197030409791077277716371013641028083419318183870507088951833751358812955108927240980871651770085955510231235374738610712593088200394888957890498118140324933433860888432806550258405697892314413003;
            6'd47: xpb[151] = 1024'd84432877531165303238448803735251296447180185602806187117016991890042671014771503466484659934807726195518289629151887951733311971763408806270087971624095748315302936169050225237492849986965128390197139102699128737092264717603066449020590298685577759577221623199327685162608839060766732144339176088147957589453;
            6'd48: xpb[151] = 1024'd51913001651113040792790564319776055399650411836173044424491521167603161049447092777895058533621725348130148083028578873056832866249101241526534915164772178446735365249148616723626887018821329539413406553628171518674298199831394287328587509170760630196552748280515045391783817233100657738419946478403600765903;
            6'd49: xpb[151] = 1024'd19393125771060778347132324904300814352120638069539901731966050445163651084122682089305457132435724500742006536905269794380353760734793676782981858705448608578167794329247008209760924050677530688629674004557214300256331682059722125636584719655943500815883873361702405620958795405434583332500716868659243942353;
            6'd50: xpb[151] = 1024'd110939945575133257300273012893640006049289291428642443167572434787701036456107410310730926945907397962797014398239454150282938496061706446594588927262456079643290897978916617033525200274050937559156139063873496928202726014508946736909560499824355820702034901857006823880240301651697141943700177085540481603134;
            6'd51: xpb[151] = 1024'd78420069695080994854614773478164765001759517662009300475046964065261526490782999622141325544721397115408872852116145071606459390547398881851035870803132509774723327059015008519659237305907138708372406514802539709784759496737274575217557710309538691321366026938194184109415279824031067537780947475796124779584;
            6'd52: xpb[151] = 1024'd45900193815028732408956534062689523954229743895376157782521493342822016525458588933551724143535396268020731305992835992929980285033091317107482814343808939906155756139113400005793274337763339857588673965731582491366792978965602413525554920794721561940697152019381544338590257996364993131861717866051767956034;
            6'd53: xpb[151] = 1024'd13380317934976469963298294647214282906699970128743015089996022620382506560134178244962122742349395420632589759869526914253501179518783752363929757884485370037588185219211791491927311369619541006804941416660625272948826461193930251833552131279904432560028277100568904567765236168698918725942488256307411132484;
            6'd54: xpb[151] = 1024'd104927137739048948916438982636553474603868623487845556525602406962919891932118906466387592555821068882687597621203711270156085914845696522175536826441492841102711288868881400315691587592992947877331406475976907900895220793643154863106527911448316752446179305595873322827046742414961477337141948473188648793265;
            6'd55: xpb[151] = 1024'd72407261858996686470780743221078233556338849721212413833076936240480381966794495777797991154635068035299456075080402191479606809331388957431983769982169271234143717948979791801825624624849149026547673926905950682477254275871482701414525121933499623065510430677060683056221720587295402931222718863444291969715;
            6'd56: xpb[151] = 1024'd39887385978944424025122503805602992508809075954579271140551465518040872001470085089208389753449067187911314528957093112803127703817081392688430713522845701365576147029078183287959661656705350175763941377834993464059287758099810539722522332418682493684841555758248043285396698759629328525303489253699935146165;
            6'd57: xpb[151] = 1024'd7367510098892161579464264390127751461279302187946128448025994795601362036145674400618788352263066340523172982833784034126648598302773827944877657063522131497008576109176574774093698688561551324980208828764036245641321240328138378030519542903865364304172680839435403514571676931963254119384259643955578322615;
            6'd58: xpb[151] = 1024'd98914329902964640532604952379466943158447955547048669883632379138138747408130402622044258165734739802578180844167968390029233333629686597756484725620529602562131679758846183597857974911934958195506673888080318873587715572777362989303495323072277684190323709334739821773853183178225812730583719860836815983396;
            6'd59: xpb[151] = 1024'd66394454022912378086946712963991702110918181780415527191106908415699237442805991933454656764548738955190039298044659311352754228115379033012931669161206032693564108838944575083992011943791159344722941339009361655169749055005690827611492533557460554809654834415927182003028161350559738324664490251092459159846;
            6'd60: xpb[151] = 1024'd33874578142860115641288473548516461063388408013782384498581437693259727477481581244865055363362738107801897751921350232676275122601071468269378612701882462824996537919042966570126048975647360493939208789938404436751782537234018665919489744042643425428985959497114542232203139522893663918745260641348102336296;
            6'd61: xpb[151] = 1024'd1354702262807853195630234133041220015858634247149241806055966970820217512157170556275453962176737260413756205798041153999796017086763903525825556242558892956428966999141358056260086007503561643155476240867447218333816019462346504227486954527826296048317084578301902461378117695227589512826031031603745512746;
            6'd62: xpb[151] = 1024'd92901522066880332148770922122380411713027287606251783241662351313357602884141898777700923775648410722468764067132225509902380752413676673337432624799566364021552070648810966880024362230876968513681941300183729846280210351911571115500462734696238615934468113073606320720659623941490148124025491248484983173527;
            6'd63: xpb[151] = 1024'd60381646186828069703112682706905170665497513839618640549136880590918092918817488089111322374462409875080622521008916431225901646899369108593879568340242794152984499728909358366158399262733169662898208751112772627862243834139898953808459945181421486553799238154793680949834602113824073718106261638740626349977;
        endcase
    end

    always_comb begin
        case(flag[50][16:12])
            5'd0: xpb[152] = 1024'd0;
            5'd1: xpb[152] = 1024'd27861770306775807257454443291429929617967740072985497856611409868478582953493077400521720973276409027692480974885607352549422541385061543850326511880919224284416928809007749852292436294589370812114476202041815409444277316368226792116457155666604357173130363235981041179009580286157999312187032028996269526427;
            5'd2: xpb[152] = 1024'd55723540613551614514908886582859859235935480145970995713222819736957165906986154801043441946552818055384961949771214705098845082770123087700653023761838448568833857618015499704584872589178741624228952404083630818888554632736453584232914311333208714346260726471962082358019160572315998624374064057992539052854;
            5'd3: xpb[152] = 1024'd83585310920327421772363329874289788853903220218956493569834229605435748860479232201565162919829227083077442924656822057648267624155184631550979535642757672853250786427023249556877308883768112436343428606125446228332831949104680376349371466999813071519391089707943123537028740858473997936561096086988808579281;
            5'd4: xpb[152] = 1024'd111447081227103229029817773165719718471870960291941991426445639473914331813972309602086883893105636110769923899542429410197690165540246175401306047523676897137667715236030999409169745178357483248457904808167261637777109265472907168465828622666417428692521452943924164716038321144631997248748128115985078105708;
            5'd5: xpb[152] = 1024'd15242155849754294888473289052335215345140273239191805154925194277416019430156248092593533651724370829019255466970543328168048866084087384696472434388265080488393969475467531923831942281429648339262183401821837200857025731620237187617307208649792336598831912765788147864941373356861363543816470318355753147804;
            5'd6: xpb[152] = 1024'd43103926156530102145927732343765144963108013312177303011536604145894602383649325493115254625000779856711736441856150680717471407469148928546798946269184304772810898284475281776124378576019019151376659603863652610301303047988463979733764364316396693771962276001769189043950953643019362856003502347352022674231;
            5'd7: xpb[152] = 1024'd70965696463305909403382175635195074581075753385162800868148014014373185337142402893636975598277188884404217416741758033266893948854210472397125458150103529057227827093483031628416814870608389963491135805905468019745580364356690771850221519983001050945092639237750230222960533929177362168190534376348292200658;
            5'd8: xpb[152] = 1024'd98827466770081716660836618926625004199043493458148298724759423882851768290635480294158696571553597912096698391627365385816316490239272016247451970031022753341644755902490781480709251165197760775605612007947283429189857680724917563966678675649605408118223002473731271401970114215335361480377566405344561727085;
            5'd9: xpb[152] = 1024'd2622541392732782519492134813240501072312806405398112453238978686353455906819418784665346330172332630346029959055479303786675190783113225542618356895610936692371010141927313995371448268269925866409890601601858992269774146872247583118157261632980316024533462295595254550873166427564727775445908607715236769181;
            5'd10: xpb[152] = 1024'd30484311699508589776946578104670430690280546478383610309850388554832038860312496185187067303448741658038510933941086656336097732168174769392944868776530160976787938950935063847663884562859296678524366803643674401714051463240474375234614417299584673197663825531576295729882746713722727087632940636711506295608;
            5'd11: xpb[152] = 1024'd58346082006284397034401021396100360308248286551369108166461798423310621813805573585708788276725150685730991908826694008885520273553236313243271380657449385261204867759942813699956320857448667490638843005685489811158328779608701167351071572966189030370794188767557336908892326999880726399819972665707775822035;
            5'd12: xpb[152] = 1024'd86207852313060204291855464687530289926216026624354606023073208291789204767298650986230509250001559713423472883712301361434942814938297857093597892538368609545621796568950563552248757152038038302753319207727305220602606095976927959467528728632793387543924552003538378087901907286038725712007004694704045348462;
            5'd13: xpb[152] = 1024'd114069622619836011549309907978960219544183766697340103879684618160267787720791728386752230223277968741115953858597908713984365356323359400943924404419287833830038725377958313404541193446627409114867795409769120630046883412345154751583985884299397744717054915239519419266911487572196725024194036723700314874889;
            5'd14: xpb[152] = 1024'd17864697242487077407965423865575716417453079644589917608164172963769475336975666877258879981896703459365285426026022631954724056867200610239090791283876017180764979617394845919203390549699574205672074003423696193126799878492484770735464470282772652623365375061383402415814539784426091319262378926070989916985;
            5'd15: xpb[152] = 1024'd45726467549262884665419867157005646035420819717575415464775582832248058290468744277780600955173112487057766400911629984504146598252262154089417303164795241465181908426402595771495826844288945017786550205465511602571077194860711562851921625949377009796495738297364443594824120070584090631449410955067259443412;
            5'd16: xpb[152] = 1024'd73588237856038691922874310448435575653388559790560913321386992700726641243961821678302321928449521514750247375797237337053569139637323697939743815045714465749598837235410345623788263138878315829901026407507327012015354511228938354968378781615981366969626101533345484773833700356742089943636442984063528969839;
            5'd17: xpb[152] = 1024'd101450008162814499180328753739865505271356299863546411177998402569205224197454899078824042901725930542442728350682844689602991681022385241790070326926633690034015766044418095476080699433467686642015502609549142421459631827597165147084835937282585724142756464769326525952843280642900089255823475013059798496266;
            5'd18: xpb[152] = 1024'd5245082785465565038984269626481002144625612810796224906477957372706911813638837569330692660344665260692059918110958607573350381566226451085236713791221873384742020283854627990742896536539851732819781203203717984539548293744495166236314523265960632049066924591190509101746332855129455550891817215430473538362;
            5'd19: xpb[152] = 1024'd33106853092241372296438712917910931762593352883781722763089367241185494767131914969852413633621074288384540892996565960122772922951287994935563225672141097669158949092862377843035332831129222544934257405245533393983825610112721958352771678932564989222197287827171550280755913141287454863078849244426743064789;
            5'd20: xpb[152] = 1024'd60968623399017179553893156209340861380561092956767220619700777109664077720624992370374134606897483316077021867882173312672195464336349538785889737553060321953575877901870127695327769125718593357048733607287348803428102926480948750469228834599169346395327651063152591459765493427445454175265881273423012591216;
            5'd21: xpb[152] = 1024'd88830393705792986811347599500770790998528833029752718476312186978142660674118069770895855580173892343769502842767780665221618005721411082636216249433979546237992806710877877547620205420307964169163209809329164212872380242849175542585685990265773703568458014299133632638775073713603453487452913302419282117643;
            5'd22: xpb[152] = 1024'd116692164012568794068802042792200720616496573102738216332923596846621243627611147171417576553450301371461983817653388017771040547106472626486542761314898770522409735519885627399912641714897334981277686011370979622316657559217402334702143145932378060741588377535114673817784653999761452799639945331415551644070;
            5'd23: xpb[152] = 1024'd20487238635219859927457558678816217489765886049988030061403151650122931243795085661924226312069036089711315385081501935741399247650313835781709148179486953873135989759322159914574838817969500072081964605025555185396574025364732353853621731915752968647898837356978656966687706211990819094708287533786226686166;
            5'd24: xpb[152] = 1024'd48349008941995667184912001970246147107733626122973527918014561518601514197288163062445947285345445117403796359967109288290821789035375379632035660060406178157552918568329909766867275112558870884196440807067370594840851341732959145970078887582357325821029200592959698145697286498148818406895319562782496212593;
            5'd25: xpb[152] = 1024'd76210779248771474442366445261676076725701366195959025774625971387080097150781240462967668258621854145096277334852716640840244330420436923482362171941325402441969847377337659619159711407148241696310917009109186004285128658101185938086536043248961682994159563828940739324706866784306817719082351591778765739020;
            5'd26: xpb[152] = 1024'd104072549555547281699820888553106006343669106268944523631237381255558680104274317863489389231898263172788758309738323993389666871805498467332688683822244626726386776186345409471452147701737612508425393211151001413729405974469412730202993198915566040167289927064921780503716447070464817031269383620775035265447;
            5'd27: xpb[152] = 1024'd7867624178198347558476404439721503216938419216194337359716936059060367720458256353996038990516997891038089877166437911360025572349339676627855070686832810077113030425781941986114344804809777599229671804805576976809322440616742749354471784898940948073600386886785763652619499282694183326337725823145710307543;
            5'd28: xpb[152] = 1024'd35729394484974154815930847731151432834906159289179835216328345927538950673951333754517759963793406918730570852052045263909448113734401220478181582567752034361529959234789691838406781099399148411344148006847392386253599756984969541470928940565545305246730750122766804831629079568852182638524757852141979833970;
            5'd29: xpb[152] = 1024'd63591164791749962073385291022581362452873899362165333072939755796017533627444411155039480937069815946423051826937652616458870655119462764328508094448671258645946888043797441690699217393988519223458624208889207795697877073353196333587386096232149662419861113358747846010638659855010181950711789881138249360397;
            5'd30: xpb[152] = 1024'd91452935098525769330839734314011292070841639435150830929551165664496116580937488555561201910346224974115532801823259969008293196504524308178834606329590482930363816852805191542991653688577890035573100410931023205142154389721423125703843251898754019592991476594728887189648240141168181262898821910134518886824;
            5'd31: xpb[152] = 1024'd119314705405301576588294177605441221688809379508136328786162575532974699534430565956082922883622634001808013776708867321557715737889585852029161118210509707214780745661812941395284089983167260847687576612972838614586431706089649917820300407565358376766121839830709928368657820427326180575085853939130788413251;
        endcase
    end

    always_comb begin
        case(flag[51][5:0])
            6'd0: xpb[153] = 1024'd0;
            6'd1: xpb[153] = 1024'd73588237856038691922874310448435575653388559790560913321386992700726641243961821678302321928449521514750247375797237337053569139637323697939743815045714465749598837235410345623788263138878315829901026407507327012015354511228938354968378781615981366969626101533345484773833700356742089943636442984063528969839;
            6'd2: xpb[153] = 1024'd23109780027952642446949693492056718562078692455386142514642130336476387150614504446589572642241368720057345344136981239528074438433427061324327505075097890565506999901249473909946287086239425938491855206627414177666348172236979936971778993548733284672432299652573911517560872639555546870154196141501463455347;
            6'd3: xpb[153] = 1024'd96698017883991334369824003940492294215467252245947055836029123037203028394576326124891894570690890234807592719934218576581643578070750759264071320120812356315105837136659819533734550225117741768392881614134741189681702683465918291940157775164714651642058401185919396291394572996297636813790639125564992425186;
            6'd4: xpb[153] = 1024'd46219560055905284893899386984113437124157384910772285029284260672952774301229008893179145284482737440114690688273962479056148876866854122648655010150195781131013999802498947819892574172478851876983710413254828355332696344473959873943557987097466569344864599305147823035121745279111093740308392283002926910694;
            6'd5: xpb[153] = 1024'd119807797911943976816773697432549012777545944701333198350671253373679415545190830571481467212932258954864938064071199816109718016504177820588398825195910246880612837037909293443680837311357167706884736820762155367348050855702898228911936768713447936314490700838493307808955445635853183683944835267066455880533;
            6'd6: xpb[153] = 1024'd69329340083857927340849080476170155686236077366158427543926391009429161451843513339768717926724106160172036032410943718584223315300281183972982515225293671696520999703748421729838861258718277815475565619882242532999044516710939810915336980646199854017296898957721734552682617918666640610462588424504390366041;
            6'd7: xpb[153] = 1024'd18850882255771877864924463519791298594926210030983656737181528645178907358496196108055968640515953365479134000750687621058728614096384547357566205254677096512429162369587550015996885206079387924066394419002329698650038177718981392918737192578951771720103097076950161296409790201480097536980341581942324851549;
            6'd8: xpb[153] = 1024'd92439120111810569787798773968226874248314769821544570058568521345905548602458017786358290568965474880229381376547924958112297753733708245297310020300391562262027999604997895639785148344957703753967420826509656710665392688947919747887115974194933138689729198610295646070243490558222187480616784566005853821388;
            6'd9: xpb[153] = 1024'd41960662283724520311874157011848017157004902486369799251823658981655294509110700554645541282757322085536479344887668860586803052529811608681893710329774987077936162270837023925943172292318813862558249625629743876316386349955961329890516186127685056392535396729524072813970662841035644407134537723443788306896;
            6'd10: xpb[153] = 1024'd115548900139763212234748467460283592810393462276930712573210651682381935753072522232947863211206843600286726720684906197640372192167135306621637525375489452827534999506247369549731435431197129692459276033137070888331740861184899684858894967743666423362161498262869557587804363197777734350770980707507317276735;
            6'd11: xpb[153] = 1024'd65070442311677162758823850503904735719083594941755941766465789318131681659725205001235113924998690805593824689024650100114877490963238670006221215404872877643443162172086497835889459378558239801050104832257158053982734522192941266862295179676418341064967696382097984331531535480591191277288733864945251762243;
            6'd12: xpb[153] = 1024'd14591984483591113282899233547525878627773727606581170959720926953881427566377887769522364638790538010900922657364394002589382789759342033390804905434256302459351324837925626122047483325919349909640933631377245219633728183200982848865695391609170258767773894501326411075258707763404648203806487022383186247751;
            6'd13: xpb[153] = 1024'd88180222339629805205773543995961454281162287397142084281107919654608068810339709447824686567240059525651170033161631339642951929396665731330548720479970768208950162073335971745835746464797665739541960038884572231649082694429921203834074173225151625737399996034671895849092408120146738147442930006446715217590;
            6'd14: xpb[153] = 1024'd37701764511543755729848927039582597189852420061967313474363057290357814716992392216111937281031906730958268001501375242117457228192769094715132410509354193024858324739175100031993770412158775848132788838004659397300076355437962785837474385157903543440206194153900322592819580402960195073960683163884649703098;
            6'd15: xpb[153] = 1024'd111290002367582447652723237488018172843240979852528226795750049991084455960954213894414259209481428245708515377298612579171026367830092792654876225555068658774457161974585445655782033551037091678033815245511986409315430866666901140805853166773884910409832295687245807366653280759702285017597126147948178672937;
            6'd16: xpb[153] = 1024'd60811544539496398176798620531639315751931112517353455989005187626834201867606896662701509923273275451015613345638356481645531666626196156039459915584452083590365324640424573941940057498398201786624644044632073574966424527674942722809253378706636828112638493806474234110380453042515741944114879305386113158445;
            6'd17: xpb[153] = 1024'd10333086711410348700874003575260458660621245182178685182260325262583947774259579430988760637065122656322711313978100384120036965422299519424043605613835508406273487306263702228098081445759311895215472843752160740617418188682984304812653590639388745815444691925702660854107625325329198870632632462824047643953;
            6'd18: xpb[153] = 1024'd83921324567449040623748314023696034314009804972739598503647317963310589018221401109291082565514644171072958689775337721173606105059623217363787420659549974155872324541674047851886344584637627725116499251259487752632772699911922659781032372255370112785070793459048145627941325682071288814269075446887576613792;
            6'd19: xpb[153] = 1024'd33442866739362991147823697067317177222699937637564827696902455599060334924874083877578333279306491376380056658115081623648111403855726580748371110688933398971780487207513176138044368531998737833707328050379574918283766360919964241784432584188122030487876991578276572371668497964884745740786828604325511099300;
            6'd20: xpb[153] = 1024'd107031104595401683070698007515752752876088497428125741018289448299786976168835905555880655207756012891130304033912318960701680543493050278688114925734647864721379324442923521761832631670877053663608354457886901930299120872148902596752811365804103397457503093111622057145502198321626835684423271588389040069139;
            6'd21: xpb[153] = 1024'd56552646767315633594773390559373895784778630092950970211544585935536722075488588324167905921547860096437402002252062863176185842289153642072698615764031289537287487108762650047990655618238163772199183257006989095950114533156944178756211577736855315160309291230850483889229370604440292610941024745826974554647;
            6'd22: xpb[153] = 1024'd6074188939229584118848773602995038693468762757776199404799723571286467982141271092455156635339707301744499970591806765650691141085257005457282305793414714353195649774601778334148679565599273880790012056127076261601108194164985760759611789669607232863115489350078910632956542887253749537458777903264909040155;
            6'd23: xpb[153] = 1024'd79662426795268276041723084051430614346857322548337112726186716272013109226103092770757478563789228816494747346389044102704260280722580703397026120839129180102794487010012123957936942704477589710691038463634403273616462705393924115727990571285588599832741590883424395406790243243995839481095220887328438009994;
            6'd24: xpb[153] = 1024'd29183968967182226565798467095051757255547455213162341919441853907762855132755775539044729277581076021801845314728788005178765579518684066781609810868512604918702649675851252244094966651838699819281867262754490439267456366401965697731390783218340517535547789002652822150517415526809296407612974044766372495502;
            6'd25: xpb[153] = 1024'd102772206823220918488672777543487332908936015003723255240828846608489496376717597217347051206030597536552092690526025342232334719156007764721353625914227070668301486911261597867883229790717015649182893670261817451282810877630904052699769564834321884505173890535998306924351115883551386351249417028829901465341;
            6'd26: xpb[153] = 1024'd52293748995134869012748160587108475817626147668548484434083984244239242283370279985634301919822444741859190658865769244706840017952111128105937315943610495484209649577100726154041253738078125757773722469381904616933804538638945634703169776767073802207980088655226733668078288166364843277767170186267835950849;
            6'd27: xpb[153] = 1024'd1815291167048819536823543630729618726316280333373713627339121879988988190022962753921552633614291947166288627205513147181345316748214491490521005972993920300117812242939854440199277685439235866364551268501991782584798199646987216706569988699825719910786286774455160411805460449178300204284923343705770436357;
            6'd28: xpb[153] = 1024'd75403529023087511459697854079165194379704840123934626948726114580715629433984784432223874562063813461916536003002750484234914456385538189430264821018708386049716649478350200063987540824317551696265577676009318794600152710875925571674948770315807086880412388307800645185639160805920390147921366327769299406196;
            6'd29: xpb[153] = 1024'd24925071195001461983773237122786337288394972788759856141981252216465375340637467200511125275855660667223633971342494386709419755181641552814848511048091810865624812144189328350145564771678661804856406475129405960251146371883967153678348982248559004583218586427029071929366333088733847074439119485207233891704;
            6'd30: xpb[153] = 1024'd98513309051040153906647547571221912941783532579320769463368244917192016584599288878813447204305182181973881347139731723762988894818965250754592326093806276615223649379599673973933827910556977634757432882636732972266500883112905508646727763864540371552844687960374556703200033445475937018075562469270762861543;
            6'd31: xpb[153] = 1024'd48034851222954104430722930614843055850473665244145998656623382552941762491251971647100697918097029387280979315479475626237494193615068614139176016123189701431131812045438802260091851857918087743348261681756820137917494544120947090650127975797292289255650886079602983446927205728289393944593315626708697347051;
            6'd32: xpb[153] = 1024'd121623089078992796353597241063278631503862225034706911978010375253668403735213793325403019846546550902031226691276712963291063333252392312078919831168904167180730649280849147883880114996796403573249288089264147149932849055349885445618506757413273656225276987612948468220760906085031483888229758610772226316890;
            6'd33: xpb[153] = 1024'd71144631250906746877672624106899774412552357699532141171265512889418149641866476093690270560338398107338324659616456865765568632048495675463503521198287591996638811946688276170038138944157513681840116888384234315583842716357927027621906969346025573928083185732176894964488078367844940814747511768210160802398;
            6'd34: xpb[153] = 1024'd20666173422820697401748007150520917321242490364357370364520650525167895548519158861977521274130245312645422627956200768240073930844599038848087211227671016812546974612527404456196162891518623790430945687504321481234836377365968609625307181278777491630889383851405321708215250650658397741265264925648095287906;
            6'd35: xpb[153] = 1024'd94254411278859389324622317598956492974631050154918283685907643225894536792480980540279843202579766827395670003753438105293643070481922736787831026273385482562145811847937750079984426030396939620331972095011648493250190888594906964593685962894758858600515485384750806482048951007400487684901707909711624257745;
            6'd36: xpb[153] = 1024'd43775953450773339848697700642577635883321182819743512879162780861644282699133663308567093916371614032702767972093182007768148369278026100172414716302768907378053974513776878366142449977758049728922800894131735658901184549602948546597086174827510776303321683503979233225776123290213944611419461067149558743253;
            6'd37: xpb[153] = 1024'd117364191306812031771572011091013211536709742610304426200549773562370923943095484986869415844821135547453015347890419344821717508915349798112158531348483373127652811749187223989930713116636365558823827301639062670916539060831886901565464956443492143272947785037324717999609823646956034555055904051213087713092;
            6'd38: xpb[153] = 1024'd66885733478725982295647394134634354445399875275129655393804911198120669849748167755156666558612982752760113316230163247296222807711453161496742221377866797943560974415026352276088737063997475667414656100759149836567532721839928483568865168376244060975753983156553144743336995929769491481573657208651022198600;
            6'd39: xpb[153] = 1024'd16407275650639932819722777178255497354090007939954884587060048833870415756400850523443917272404829958067211284569907149770728106507556524881325911407250222759469137080865480562246761011358585776005484899879237002218526382847970065572265380308995978678560181275781571487064168212582948408091410366088956684108;
            6'd40: xpb[153] = 1024'd89995513506678624742597087626691073007478567730515797908447041534597057000362672201746239200854351472817458660367144486824297246144880222821069726452964688509067974316275826186035024150236901605906511307386564014233880894076908420540644161924977345648186282809127056260897868569325038351727853350152485653947;
            6'd41: xpb[153] = 1024'd39517055678592575266672470670312215916168700395341027101702179170346802907015354970033489914646198678124556628706888389298802544940983586205653416482348113324976136982114954472193048097598011714497340106506651179884874555084950002544044373857729263350992480928355483004625040852138495278245606507590420139455;
            6'd42: xpb[153] = 1024'd113105293534631267189546781118747791569557260185901940423089171871073444150977176648335811843095720192874804004504125726352371684578307284145397231528062579074574974217525300095981311236476327544398366514013978191900229066313888357512423155473710630320618582461700967778458741208880585221882049491653949109294;
            6'd43: xpb[153] = 1024'd62626835706545217713622164162368934478247392850727169616344309506823190057629859416623062556887567398181901972843869628826876983374410647529980921557446003890483136883364428382139335183837437652989195313134065357551222727321929939515823367406462548023424780580929394522185913491694042148399802649091883594802;
            6'd44: xpb[153] = 1024'd12148377878459168237697547205990077386937525515552398809599447142572935964282542184910313270679414603488999941183613531301382282170514010914564611586829428706391299549203556668297359131198547761580024112254152523202216388329971521519223579339214465726230978700157821265913085774507499074917555806529818080310;
            6'd45: xpb[153] = 1024'd85736615734497860160571857654425653040326085306113312130986439843299577208244363863212635199128936118239247316980850868354951421807837708854308426632543894455990136784613902292085622270076863591481050519761479535217570899558909876487602360955195832695857080233503306039746786131249589018553998790593347050149;
            6'd46: xpb[153] = 1024'd35258157906411810684647240698046795949016217970938541324241577479049323114897046631499885912920783323546345285320594770829456720603941072238892116661927319271898299450453030578243646217437973700071879318881566700868564560566951458491002572887947750398663278352731732783473958414063045945071751948031281535657;
            6'd47: xpb[153] = 1024'd108846395762450502607521551146482371602404777761499454645628570179775964358858868309802207841370304838296592661117832107883025860241264770178635931707641785021497136685863376202031909356316289529972905726388893712883919071795889813459381354503929117368289379886077217557307658770805135888708194932094810505496;
            6'd48: xpb[153] = 1024'd58367937934364453131596934190103514511094910426324683838883707815525710265511551078089458555162152043603690629457576010357531159037368133563219621737025209837405299351702504488189933303677399638563734525508980878534912732803931395462781566436681035071095578005305644301034831053618592815225948089532744991004;
            6'd49: xpb[153] = 1024'd7889480106278403655672317233724657419785043091149913032138845451275456172164233846376709268953999248910788597797319912832036457833471496947803311766408634653313462017541632774347957251038509747154563324629068044185906393811972977466181778369432952773901776124534071044762003336432049741743701246970679476512;
            6'd50: xpb[153] = 1024'd81477717962317095578546627682160233073173602881710826353525838152002097416126055524679031197403520763661035973594557249885605597470795194887547126812123100402912299252951978398136220389916825577055589732136395056201260905040911332434560559985414319743527877657879555818595703693174139685380144231034208446351;
            6'd51: xpb[153] = 1024'd30999260134231046102622010725781375981863735546536055546780975787751843322778738292966281911195367968968133941934301152360110896266898558272130816841506525218820461918791106684294244337277935685646418531256482221852254566048952914437960771918166237446334075777107982562322875975987596611897897388472142931859;
            6'd52: xpb[153] = 1024'd104587497990269738025496321174216951635252295337096968868167968488478484566740559971268603839644889483718381317731538489413680035904222256211874631887220990968419299154201452308082507476156251515547444938763809233867609077277891269406339553534147604415960177310453467336156576332729686555534340372535671901698;
            6'd53: xpb[153] = 1024'd54109040162183688549571704217838094543942428001922198061423106124228230473393242739555854553436736689025479286071282391888185334700325619596458321916604415784327461820040580594240531423517361624138273737883896399518602738285932851409739765466899522118766375429681894079883748615543143482052093529973606387206;
            6'd54: xpb[153] = 1024'd3630582334097639073647087261459237452632560666747427254678243759977976380045925507843105267228583894332577254411026294362690633496428982981042011945987840600235624485879708880398555370878471732729102537003983565169596399293974433413139977399651439821572573548910320823610920898356600408569846687411540872714;
            6'd55: xpb[153] = 1024'd77218820190136330996521397709894813106021120457308340576065236460704617624007747186145427195678105409082824630208263631416259773133752680920785826991702306349834461721290054504186818509756787562630128944511310577184950910522912788381518759015632806791198675082255805597444621255098690352206289671475069842553;
            6'd56: xpb[153] = 1024'd26740362362050281520596780753515956014711253122133569769320374096454363530660429954432677909469952614389922598548007533890765071929856044305369517021085731165742624387129182790344842457117897671220957743631397742835944571530954370384918970948384724494004873201484232341171793537912147278724042828913004328061;
            6'd57: xpb[153] = 1024'd100328600218088973443471091201951531668099812912694483090707366797181004774622251632734999837919474129140169974345244870944334211567179742245113332066800196915341461622539528414133105595996213501121984151138724754851299082759892725353297752564366091463630974734829717115005493894654237222360485812976533297900;
            6'd58: xpb[153] = 1024'd49850142390002923967546474245572674576789945577519712283962504432930750681274934401022250551711321334447267942684988773418839510363283105629697022096183621731249624288378656700291129543357323609712812950258811920502292743767934307356697964497118009166437172854058143858732666177467694148878238970414467783408;
            6'd59: xpb[153] = 1024'd123438380246041615890420784694008250230178505368080625605349497133657391925236756079324572480160842849197515318482226110472408650000606803569440837141898087480848461523789002324079392682235639439613839357766138932517647254996872662325076746113099376136063274387403628632566366534209784092514681954477996753247;
            6'd60: xpb[153] = 1024'd72959922417955566414496167737629393138868638032905854798604634769407137831889438847611823193952690054504613286821970012946913948796710166954024527171281512296756624189628130610237416629596749548204668156886226098168640916004914244328476958045851293838869472506632055376293538817023241019032435111915931238755;
            6'd61: xpb[153] = 1024'd22481464589869516938571550781250536047558770697731083991859772405156883738542121615899073907744537259811711255161713915421419247592813530338608217200664937112664786855467258896395440576957859656795496956006313263819634577012955826331877169978603211541675670625860482120020711099836697945550188269353865724263;
            6'd62: xpb[153] = 1024'd96069702445908208861445861229686111700947330488291997313246765105883524982503943294201395836194058774561958630958951252474988387230137228278352032246379402862263624090877604520183703715836175486696523363513640275834989088241894181300255951594584578511301772159205966893854411456578787889186631253417394694102;
            6'd63: xpb[153] = 1024'd45591244617822159385521244273307254609637463153117226506501902741633270889156626062488646549985905979869056599298695154949493686026240591662935722275762827678171786756716732806341727663197285595287352162633727441485982749249935763303656163527336496214107970278434393637581583739392244815704384410855329179610;
        endcase
    end

    always_comb begin
        case(flag[51][11:6])
            6'd0: xpb[154] = 1024'd0;
            6'd1: xpb[154] = 1024'd119179482473860851308395554721742830263026022943678139827888895442359912133118447740790968478435427494619303975095932492003062825663564289602679537321477293427770623992127078430129990802075601425188378570141054453501337260478874118272034945143317863183734071811779878411415284096134334759340827394918858149449;
            6'd2: xpb[154] = 1024'd114292269263596961217992182038671227781353618761620595527645935819742928928927756571566865742213180679795458542734371549427061810485908244650198949626623545921850573414682939522629742412633997129066559531894869060638313670736851463579091320603406277100648240209442698792724040118340036501562964963212121814567;
            6'd3: xpb[154] = 1024'd109405056053333071127588809355599625299681214579563051227402976197125945724737065402342763005990933864971613110372810606851060795308252199697718361931769798415930522837238800615129494023192392832944740493648683667775290080994828808886147696063494691017562408607105519174032796140545738243785102531505385479685;
            6'd4: xpb[154] = 1024'd104517842843069181037185436672528022818008810397505506927160016574508962520546374233118660269768687050147767678011249664275059780130596154745237774236916050910010472259794661707629245633750788536822921455402498274912266491252806154193204071523583104934476577004768339555341552162751439986007240099798649144803;
            6'd5: xpb[154] = 1024'd99630629632805290946782063989456420336336406215447962626917056951891979316355683063894557533546440235323922245649688721699058764952940109792757186542062303404090421682350522800128997244309184240701102417156312882049242901510783499500260446983671518851390745402431159936650308184957141728229377668091912809921;
            6'd6: xpb[154] = 1024'd94743416422541400856378691306384817854664002033390418326674097329274996112164991894670454797324193420500076813288127779123057749775284064840276598847208555898170371104906383892628748854867579944579283378910127489186219311768760844807316822443759932768304913800093980317959064207162843470451515236385176475039;
            6'd7: xpb[154] = 1024'd89856203212277510765975318623313215372991597851332874026431137706658012907974300725446352061101946605676231380926566836547056734597628019887796011152354808392250320527462244985128500465425975648457464340663942096323195722026738190114373197903848346685219082197756800699267820229368545212673652804678440140157;
            6'd8: xpb[154] = 1024'd84968990002013620675571945940241612891319193669275329726188178084041029703783609556222249324879699790852385948565005893971055719419971974935315423457501060886330269950018106077628252075984371352335645302417756703460172132284715535421429573363936760602133250595419621080576576251574246954895790372971703805275;
            6'd9: xpb[154] = 1024'd80081776791749730585168573257170010409646789487217785425945218461424046499592918386998146588657452976028540516203444951395054704242315929982834835762647313380410219372573967170128003686542767056213826264171571310597148542542692880728485948824025174519047418993082441461885332273779948697117927941264967470393;
            6'd10: xpb[154] = 1024'd75194563581485840494765200574098407927974385305160241125702258838807063295402227217774043852435206161204695083841884008819053689064659885030354248067793565874490168795129828262627755297101162760092007225925385917734124952800670226035542324284113588435961587390745261843194088295985650439340065509558231135511;
            6'd11: xpb[154] = 1024'd70307350371221950404361827891026805446301981123102696825459299216190080091211536048549941116212959346380849651480323066243052673887003840077873660372939818368570118217685689355127506907659558463970188187679200524871101363058647571342598699744202002352875755788408082224502844318191352181562203077851494800629;
            6'd12: xpb[154] = 1024'd65420137160958060313958455207955202964629576941045152525216339593573096887020844879325838379990712531557004219118762123667051658709347795125393072678086070862650067640241550447627258518217954167848369149433015132008077773316624916649655075204290416269789924186070902605811600340397053923784340646144758465747;
            6'd13: xpb[154] = 1024'd60532923950694170223555082524883600482957172758987608224973379970956113682830153710101735643768465716733158786757201181091050643531691750172912484983232323356730017062797411540127010128776349871726550111186829739145054183574602261956711450664378830186704092583733722987120356362602755666006478214438022130865;
            6'd14: xpb[154] = 1024'd55645710740430280133151709841811998001284768576930063924730420348339130478639462540877632907546218901909313354395640238515049628354035705220431897288378575850809966485353272632626761739334745575604731072940644346282030593832579607263767826124467244103618260981396543368429112384808457408228615782731285795983;
            6'd15: xpb[154] = 1024'd50758497530166390042748337158740395519612364394872519624487460725722147274448771371653530171323972087085467922034079295939048613176379660267951309593524828344889915907909133725126513349893141279482912034694458953419007004090556952570824201584555658020532429379059363749737868407014159150450753351024549461101;
            6'd16: xpb[154] = 1024'd45871284319902499952344964475668793037939960212814975324244501103105164070258080202429427435101725272261622489672518353363047597998723615315470721898671080838969865330464994817626264960451536983361092996448273560555983414348534297877880577044644071937446597776722184131046624429219860892672890919317813126219;
            6'd17: xpb[154] = 1024'd40984071109638609861941591792597190556267556030757431024001541480488180866067389033205324698879478457437777057310957410787046582821067570362990134203817333333049814753020855910126016571009932687239273958202088167692959824606511643184936952504732485854360766174385004512355380451425562634895028487611076791337;
            6'd18: xpb[154] = 1024'd36096857899374719771538219109525588074595151848699886723758581857871197661876697863981221962657231642613931624949396468211045567643411525410509546508963585827129764175576717002625768181568328391117454919955902774829936234864488988491993327964820899771274934572047824893664136473631264377117166055904340456455;
            6'd19: xpb[154] = 1024'd31209644689110829681134846426453985592922747666642342423515622235254214457686006694757119226434984827790086192587835525635044552465755480458028958814109838321209713598132578095125519792126724094995635881709717381966912645122466333799049703424909313688189102969710645274972892495836966119339303624197604121573;
            6'd20: xpb[154] = 1024'd26322431478846939590731473743382383111250343484584798123272662612637231253495315525533016490212738012966240760226274583059043537288099435505548371119256090815289663020688439187625271402685119798873816843463531989103889055380443679106106078884997727605103271367373465656281648518042667861561441192490867786691;
            6'd21: xpb[154] = 1024'd21435218268583049500328101060310780629577939302527253823029702990020248049304624356308913753990491198142395327864713640483042522110443390553067783424402343309369612443244300280125023013243515502751997805217346596240865465638421024413162454345086141522017439765036286037590404540248369603783578760784131451809;
            6'd22: xpb[154] = 1024'd16548005058319159409924728377239178147905535120469709522786743367403264845113933187084811017768244383318549895503152697907041506932787345600587195729548595803449561865800161372624774623801911206630178766971161203377841875896398369720218829805174555438931608162699106418899160562454071346005716329077395116927;
            6'd23: xpb[154] = 1024'd11660791848055269319521355694167575666233130938412165222543783744786281640923242017860708281545997568494704463141591755331040491755131300648106608034694848297529511288356022465124526234360306910508359728724975810514818286154375715027275205265262969355845776560361926800207916584659773088227853897370658782045;
            6'd24: xpb[154] = 1024'd6773578637791379229117983011095973184560726756354620922300824122169298436732550848636605545323750753670859030780030812755039476577475255695626020339841100791609460710911883557624277844918702614386540690478790417651794696412353060334331580725351383272759944958024747181516672606865474830449991465663922447163;
            6'd25: xpb[154] = 1024'd1886365427527489138714610328024370702888322574297076622057864499552315232541859679412502809101503938847013598418469870179038461399819210743145432644987353285689410133467744650124029455477098318264721652232605024788771106670330405641387956185439797189674113355687567562825428629071176572672129033957186112281;
            6'd26: xpb[154] = 1024'd121065847901388340447110165049767200965914345517975216449946759941912227365660307420203471287536931433466317573514402362182101287063383500345824969966464646713460034125594823080254020257552699743453100222373659478290108367149204523913422901328757660373408185167467445974240712725205511332012956428876044261730;
            6'd27: xpb[154] = 1024'd116178634691124450356706792366695598484241941335917672149703800319295244161469616250979368551314684618642472141152841419606100271885727455393344382271610899207539983548150684172753771868111095447331281184127474085427084777407181869220479276788846074290322353565130266355549468747411213074235093997169307926848;
            6'd28: xpb[154] = 1024'd111291421480860560266303419683623996002569537153860127849460840696678260957278925081755265815092437803818626708791280477030099256708071410440863794576757151701619932970706545265253523478669491151209462145881288692564061187665159214527535652248934488207236521962793086736858224769616914816457231565462571591966;
            6'd29: xpb[154] = 1024'd106404208270596670175900047000552393520897132971802583549217881074061277753088233912531163078870190988994781276429719534454098241530415365488383206881903404195699882393262406357753275089227886855087643107635103299701037597923136559834592027709022902124150690360455907118166980791822616558679369133755835257084;
            6'd30: xpb[154] = 1024'd101516995060332780085496674317480791039224728789745039248974921451444294548897542743307060342647944174170935844068158591878097226352759320535902619187049656689779831815818267450253026699786282558965824069388917906838014008181113905141648403169111316041064858758118727499475736814028318300901506702049098922202;
            6'd31: xpb[154] = 1024'd96629781850068889995093301634409188557552324607687494948731961828827311344706851574082957606425697359347090411706597649302096211175103275583422031492195909183859781238374128542752778310344678262844005031142732513974990418439091250448704778629199729957979027155781547880784492836234020043123644270342362587320;
            6'd32: xpb[154] = 1024'd91742568639804999904689928951337586075879920425629950648489002206210328140516160404858854870203450544523244979345036706726095195997447230630941443797342161677939730660929989635252529920903073966722185992896547121111966828697068595755761154089288143874893195553444368262093248858439721785345781838635626252438;
            6'd33: xpb[154] = 1024'd86855355429541109814286556268265983594207516243572406348246042583593344936325469235634752133981203729699399546983475764150094180819791185678460856102488414172019680083485850727752281531461469670600366954650361728248943238955045941062817529549376557791807363951107188643402004880645423527567919406928889917556;
            6'd34: xpb[154] = 1024'd81968142219277219723883183585194381112535112061514862048003082960976361732134778066410649397758956914875554114621914821574093165642135140725980268407634666666099629506041711820252033142019865374478547916404176335385919649213023286369873905009464971708721532348770009024710760902851125269790056975222153582674;
            6'd35: xpb[154] = 1024'd77080929009013329633479810902122778630862707879457317747760123338359378527944086897186546661536710100051708682260353878998092150464479095773499680712780919160179578928597572912751784752578261078356728878157990942522896059471000631676930280469553385625635700746432829406019516925056827012012194543515417247792;
            6'd36: xpb[154] = 1024'd72193715798749439543076438219051176149190303697399773447517163715742395323753395727962443925314463285227863249898792936422091135286823050821019093017927171654259528351153434005251536363136656782234909839911805549659872469728977976983986655929641799542549869144095649787328272947262528754234332111808680912910;
            6'd37: xpb[154] = 1024'd67306502588485549452673065535979573667517899515342229147274204093125412119562704558738341189092216470404017817537231993846090120109167005868538505323073424148339477773709295097751287973695052486113090801665620156796848879986955322291043031389730213459464037541758470168637028969468230496456469680101944578028;
            6'd38: xpb[154] = 1024'd62419289378221659362269692852907971185845495333284684847031244470508428915372013389514238452869969655580172385175671051270089104931510960916057917628219676642419427196265156190251039584253448189991271763419434763933825290244932667598099406849818627376378205939421290549945784991673932238678607248395208243146;
            6'd39: xpb[154] = 1024'd57532076167957769271866320169836368704173091151227140546788284847891445711181322220290135716647722840756326952814110108694088089753854915963577329933365929136499376618821017282750791194811843893869452725173249371070801700502910012905155782309907041293292374337084110931254541013879633980900744816688471908264;
            6'd40: xpb[154] = 1024'd52644862957693879181462947486764766222500686969169596246545325225274462506990631051066032980425476025932481520452549166118087074576198871011096742238512181630579326041376878375250542805370239597747633686927063978207778110760887358212212157769995455210206542734746931312563297036085335723122882384981735573382;
            6'd41: xpb[154] = 1024'd47757649747429989091059574803693163740828282787112051946302365602657479302799939881841930244203229211108636088090988223542086059398542826058616154543658434124659275463932739467750294415928635301625814648680878585344754521018864703519268533230083869127120711132409751693872053058291037465345019953274999238500;
            6'd42: xpb[154] = 1024'd42870436537166099000656202120621561259155878605054507646059405980040496098609248712617827507980982396284790655729427280966085044220886781106135566848804686618739224886488600560250046026487031005503995610434693192481730931276842048826324908690172283044034879530072572075180809080496739207567157521568262903618;
            6'd43: xpb[154] = 1024'd37983223326902208910252829437549958777483474422996963345816446357423512894418557543393724771758735581460945223367866338390084029043230736153654979153950939112819174309044461652749797637045426709382176572188507799618707341534819394133381284150260696960949047927735392456489565102702440949789295089861526568736;
            6'd44: xpb[154] = 1024'd33096010116638318819849456754478356295811070240939419045573486734806529690227866374169622035536488766637099791006305395814083013865574691201174391459097191606899123731600322745249549247603822413260357533942322406755683751792796739440437659610349110877863216325398212837798321124908142692011432658154790233854;
            6'd45: xpb[154] = 1024'd28208796906374428729446084071406753814138666058881874745330527112189546486037175204945519299314241951813254358644744453238081998687918646248693803764243444100979073154156183837749300858162218117138538495696137013892660162050774084747494035070437524794777384723061033219107077147113844434233570226448053898972;
            6'd46: xpb[154] = 1024'd23321583696110538639042711388335151332466261876824330445087567489572563281846484035721416563091995136989408926283183510662080983510262601296213216069389696595059022576712044930249052468720613821016719457449951621029636572308751430054550410530525938711691553120723853600415833169319546176455707794741317564090;
            6'd47: xpb[154] = 1024'd18434370485846648548639338705263548850793857694766786144844607866955580077655792866497313826869748322165563493921622568086079968332606556343732628374535949089138971999267906022748804079279009524894900419203766228166612982566728775361606785990614352628605721518386673981724589191525247918677845363034581229208;
            6'd48: xpb[154] = 1024'd13547157275582758458235966022191946369121453512709241844601648244338596873465101697273211090647501507341718061560061625510078953154950511391252040679682201583218921421823767115248555689837405228773081380957580835303589392824706120668663161450702766545519889916049494363033345213730949660899982931327844894326;
            6'd49: xpb[154] = 1024'd8659944065318868367832593339120343887449049330651697544358688621721613669274410528049108354425254692517872629198500682934077937977294466438771452984828454077298870844379628207748307300395800932651262342711395442440565803082683465975719536910791180462434058313712314744342101235936651403122120499621108559444;
            6'd50: xpb[154] = 1024'd3772730855054978277429220656048741405776645148594153244115728999104630465083719358825005618203007877694027196836939740358076922799638421486290865289974706571378820266935489300248058910954196636529443304465210049577542213340660811282775912370879594379348226711375135125650857258142353145344258067914372224562;
            6'd51: xpb[154] = 1024'd122952213328915829585824775377791571668802668092272293072004624441464542598202167099615974096638435372313331171932872232361139748463202711088970402611451999999149444259062567730378049713029798061717821874606264503078879473819534929554810857514197457563082298523155013537066141354276687904685085462833230374011;
            6'd52: xpb[154] = 1024'd118065000118651939495421402694719969187130263910214748771761664818847559394011475930391871360416188557489485739571311289785138733285546666136489814916598252493229393681618428822877801323588193765596002836360079110215855884077512274861867232974285871479996466920817833918374897376482389646907223031126494039129;
            6'd53: xpb[154] = 1024'd113177786908388049405018030011648366705457859728157204471518705196230576189820784761167768624193941742665640307209750347209137718107890621184009227221744504987309343104174289915377552934146589469474183798113893717352832294335489620168923608434374285396910635318480654299683653398688091389129360599419757704247;
            6'd54: xpb[154] = 1024'd108290573698124159314614657328576764223785455546099660171275745573613592985630093591943665887971694927841794874848189404633136702930234576231528639526890757481389292526730151007877304544704985173352364759867708324489808704593466965475979983894462699313824803716143474680992409420893793131351498167713021369365;
            6'd55: xpb[154] = 1024'd103403360487860269224211284645505161742113051364042115871032785950996609781439402422719563151749448113017949442486628462057135687752578531279048051832037009975469241949286012100377056155263380877230545721621522931626785114851444310783036359354551113230738972113806295062301165443099494873573635736006285034483;
            6'd56: xpb[154] = 1024'd98516147277596379133807911962433559260440647181984571570789826328379626577248711253495460415527201298194104010125067519481134672574922486326567464137183262469549191371841873192876807765821776581108726683375337538763761525109421656090092734814639527147653140511469115443609921465305196615795773304299548699601;
            6'd57: xpb[154] = 1024'd93628934067332489043404539279361956778768242999927027270546866705762643373058020084271357679304954483370258577763506576905133657397266441374086876442329514963629140794397734285376559376380172284986907645129152145900737935367399001397149110274727941064567308909131935824918677487510898358017910872592812364719;
            6'd58: xpb[154] = 1024'd88741720857068598953001166596290354297095838817869482970303907083145660168867328915047254943082707668546413145401945634329132642219610396421606288747475767457709090216953595377876310986938567988865088606882966753037714345625376346704205485734816354981481477306794756206227433509716600100240048440886076029837;
            6'd59: xpb[154] = 1024'd83854507646804708862597793913218751815423434635811938670060947460528676964676637745823152206860460853722567713040384691753131627041954351469125701052622019951789039639509456470376062597496963692743269568636781360174690755883353692011261861194904768898395645704457576587536189531922301842462186009179339694955;
            6'd60: xpb[154] = 1024'd78967294436540818772194421230147149333751030453754394369817987837911693760485946576599049470638214038898722280678823749177130611864298306516645113357768272445868989062065317562875814208055359396621450530390595967311667166141331037318318236654993182815309814102120396968844945554128003584684323577472603360073;
            6'd61: xpb[154] = 1024'd74080081226276928681791048547075546852078626271696850069575028215294710556295255407374946734415967224074876848317262806601129596686642261564164525662914524939948938484621178655375565818613755100499631492144410574448643576399308382625374612115081596732223982499783217350153701576333705326906461145765867025191;
            6'd62: xpb[154] = 1024'd69192868016013038591387675864003944370406222089639305769332068592677727352104564238150843998193720409251031415955701864025128581508986216611683937968060777434028887907177039747875317429172150804377812453898225181585619986657285727932430987575170010649138150897446037731462457598539407069128598714059130690309;
            6'd63: xpb[154] = 1024'd64305654805749148500984303180932341888733817907581761469089108970060744147913873068926741261971473594427185983594140921449127566331330171659203350273207029928108837329732900840375069039730546508255993415652039788722596396915263073239487363035258424566052319295108858112771213620745108811350736282352394355427;
        endcase
    end

    always_comb begin
        case(flag[51][16:12])
            5'd0: xpb[155] = 1024'd0;
            5'd1: xpb[155] = 1024'd59418441595485258410580930497860739407061413725524217168846149347443760943723181899702638525749226779603340551232579978873126551153674126706722762578353282422188786752288761932874820650288942212134174377405854395859572807173240418546543738495346838482966487692771678494079969642950810553572873850645658020545;
            5'd2: xpb[155] = 1024'd118836883190970516821161860995721478814122827451048434337692298694887521887446363799405277051498453559206681102465159957746253102307348253413445525156706564844377573504577523865749641300577884424268348754811708791719145614346480837093087476990693676965932975385543356988159939285901621107145747701291316041090;
            5'd3: xpb[155] = 1024'd54188629102331033832943864088767785476485814050836967378406592977354387493860406789092844362590006029366872246240246502040315812619802045565008162718728806332875685687295068460994222759349620915092325523830323341214357571298824482674652645802811066182079559664197977452133380854923798643599931725311379577304;
            5'd4: xpb[155] = 1024'd113607070697816292243524794586628524883547227776361184547252742324798148437583588688795482888339232808970212797472826480913442363773476172271730925297082088755064472439583830393869043409638563127226499901236177737073930378472064901221196384298157904665046047356969655946213350497874609197172805575957037597849;
            5'd5: xpb[155] = 1024'd48958816609176809255306797679674831545910214376149717587967036607265014043997631678483050199430785279130403941247913025207505074085929964423293562859104330243562584622301374989113624868410299618050476670254792286569142335424408546802761553110275293881192631635624276410186792066896786733626989599977101134063;
            5'd6: xpb[155] = 1024'd108377258204662067665887728177535570952971628101673934756813185954708774987720813578185688725180012058733744492480493004080631625239604091130016325437457612665751371374590136921988445518699241830184651047660646682428715142597648965349305291605622132364159119328395954904266761709847597287199863450622759154608;
            5'd7: xpb[155] = 1024'd43729004116022584677669731270581877615334614701462467797527480237175640594134856567873256036271564528893935636255579548374694335552057883281578962999479854154249483557307681517233026977470978321008627816679261231923927099549992610930870460417739521580305703607050575368240203278869774823654047474642822690822;
            5'd8: xpb[155] = 1024'd103147445711507843088250661768442617022396028426986684966373629584619401537858038467575894562020791308497276187488159527247820886705732009988301725577833136576438270309596443450107847627759920533142802194085115627783499906723233029477414198913086360063272191299822253862320172921820585377226921325288480711367;
            5'd9: xpb[155] = 1024'd38499191622868360100032664861488923684759015026775218007087923867086267144272081457263461873112343778657467331263246071541883597018185802139864363139855378064936382492313988045352429086531657023966778963103730177278711863675576675058979367725203749279418775578476874326293614490842762913681105349308544247581;
            5'd10: xpb[155] = 1024'd97917633218353618510613595359349663091820428752299435175934073214530028087995263356966100398861570558260807882495826050415010148171859928846587125718208660487125169244602749978227249736820599236100953340509584573138284670848817093605523106220550587762385263271248552820373584133793573467253979199954202268126;
            5'd11: xpb[155] = 1024'd33269379129714135522395598452395969754183415352087968216648367496996893694409306346653667709953123028420999026270912594709072858484313720998149763280230901975623281427320294573471831195592335726924930109528199122633496627801160739187088275032667976978531847549903173284347025702815751003708163223974265804340;
            5'd12: xpb[155] = 1024'd92687820725199393932976528950256709161244829077612185385494516844440654638132488246356306235702349808024339577503492573582199409637987847704872525858584184397812068179609056506346651845881277939059104486934053518493069434974401157733632013528014815461498335242674851778426995345766561557281037074619923824885;
            5'd13: xpb[155] = 1024'd28039566636559910944758532043303015823607815677400718426208811126907520244546531236043873546793902278184530721278579117876262119950441639856435163420606425886310180362326601101591233304653014429883081255952668067988281391926744803315197182340132204677644919521329472242400436914788739093735221098639987361099;
            5'd14: xpb[155] = 1024'd87458008232045169355339462541163755230669229402924935595054960474351281188269713135746512072543129057787871272511159096749388671104115766563157925998959708308498967114615363034466053954941956642017255633358522463847854199099985221861740920835479043160611407214101150736480406557739549647308094949285645381644;
            5'd15: xpb[155] = 1024'd22809754143405686367121465634210061893032216002713468635769254756818146794683756125434079383634681527948062416286245641043451381416569558714720563560981949796997079297332907629710635413713693132841232402377137013343066156052328867443306089647596432376757991492755771200453848126761727183762278973305708917858;
            5'd16: xpb[155] = 1024'd82228195738890944777702396132070801300093629728237685804615404104261907738406938025136717909383908307551402967518825619916577932570243685421443326139335232219185866049621669562585456064002635344975406779782991409202638963225569285989849828142943270859724479185527449694533817769712537737335152823951366938403;
            5'd17: xpb[155] = 1024'd17579941650251461789484399225117107962456616328026218845329698386728773344820981014824285220475460777711594111293912164210640642882697477573005963701357473707683978232339214157830037522774371835799383548801605958697850920177912931571414996955060660075871063464182070158507259338734715273789336847971430474617;
            5'd18: xpb[155] = 1024'd76998383245736720200065329722977847369518030053550436014175847734172534288544162914526923746224687557314934662526492143083767194036371604279728726279710756129872764984627976090704858173063314047933557926207460354557423727351153350117958735450407498558837551156953748652587228981685525827362210698617088495162;
            5'd19: xpb[155] = 1024'd12350129157097237211847332816024154031881016653338969054890142016639399894958205904214491057316240027475125806301578687377829904348825396431291363841732997618370877167345520685949439631835050538757534695226074904052635684303496995699523904262524887774984135435608369116560670550707703363816394722637152031376;
            5'd20: xpb[155] = 1024'd71768570752582495622428263313884893438942430378863186223736291364083160838681387803917129583065466807078466357534158666250956455502499523138014126420086280040559663919634282618824260282123992750891709072631929299912208491476737414246067642757871726257950623128380047610640640193658513917389268573282810051921;
            5'd21: xpb[155] = 1024'd7120316663943012634210266406931200101305416978651719264450585646550026445095430793604696894157019277238657501309245210545019165814953315289576763982108521529057776102351827214068841740895729241715685841650543849407420448429081059827632811569989115474097207407034668074614081762680691453843452597302873588135;
            5'd22: xpb[155] = 1024'd66538758259428271044791196904791939508366830704175936433296734993993787388818612693307335419906246056841998052541825189418145716968627441996299526560461803951246562854640589146943662391184671453849860219056398245266993255602321478374176550065335953957063695099806346568694051405631502007416326447948531608680;
            5'd23: xpb[155] = 1024'd1890504170788788056573199997838246170729817303964469474011029276460652995232655682994902730997798527002189196316911733712208427281081234147862164122484045439744675037358133742188243849956407944673836988075012794762205212554665123955741718877453343173210279378460967032667492974653679543870510471968595144894;
            5'd24: xpb[155] = 1024'd61308945766274046467154130495698985577791231029488686642857178623904413938955837582697541256747025306605529747549491712585334978434755360854584926700837327861933461789646895675063064500245350156808011365480867190621778019727905542502285457372800181656176767071232645526747462617604490097443384322614253165439;
            5'd25: xpb[155] = 1024'd120727387361759304877735060993559724984852644755012903811703327971348174882679019482400179782496252086208870298782071691458461529588429487561307689279190610284122248541935657607937885150534292368942185742886721586481350826901145961048829195868147020139143254764004324020827432260555300651016258173259911185984;
            5'd26: xpb[155] = 1024'd56079133273119821889517064086606031647215631354801436852417622253815040489093062472087747093587804556369061442557158235752524239900883279712870326841212851772620360724653202203182466609306028859766162511905336135976562783853489606630394364680264409355289839042658944484800873829577478187470442197279974722198;
            5'd27: xpb[155] = 1024'd115497574868605080300097994584466771054277045080325654021263771601258801432816244371790385619337031335972401993789738214625650791054557406419593089419566134194809147476941964136057287259594971071900336889311190531836135591026730025176938103175611247838256326735430622978880843472528288741043316047925632742743;
            5'd28: xpb[155] = 1024'd50849320779965597311879997677513077716640031680114187061978065883725667039230287361477952930428583806132593137564824758919713501367011198571155726981588375683307259659659508731301868718366707562724313658329805081331347547979073670758503271987728637054402911014085243442854285041550466277497500071945696278957;
            5'd29: xpb[155] = 1024'd110267762375450855722460928175373817123701445405638404230824215231169427982953469261180591456177810585735933688797404737792840052520685325277878489559941658105496046411948270664176689368655649774858488035735659477190920355152314089305047010483075475537369398706856921936934254684501276831070373922591354299502;
            5'd30: xpb[155] = 1024'd45619508286811372734242931268420123786064432005426937271538509513636293589367512250868158767269363055896124832572491282086902762833139117429441127121963899593994158594665815259421270827427386265682464804754274026686132312104657734886612179295192864753515982985511542400907696253523454367524557946611417835716;
            5'd31: xpb[155] = 1024'd105037949882296631144823861766280863193125845730951154440384658861080054533090694150570797293018589835499465383805071260960029313986813244136163889700317182016182945346954577192296091477716328477816639182160128422545705119277898153433155917790539703236482470678283220894987665896474264921097431797257075856261;
        endcase
    end

    always_comb begin
        case(flag[52][5:0])
            6'd0: xpb[156] = 1024'd0;
            6'd1: xpb[156] = 1024'd82228195738890944777702396132070801300093629728237685804615404104261907738406938025136717909383908307551402967518825619916577932570243685421443326139335232219185866049621669562585456064002635344975406779782991409202638963225569285989849828142943270859724479185527449694533817769712537737335152823951366938403;
            6'd2: xpb[156] = 1024'd40389695793657148156605864859327169855488832330739687481098953143546920139504737140258364604110142305659656527580157805254092024299267036287726527262339423504681057529672121787540672936488064968640615951178742972040917076230241799014721086602657092452629054956937841358961107465496442457551615821277139392475;
            6'd3: xpb[156] = 1024'd122617891532548092934308260991397971155582462058977373285714357247808827877911675165395082513494050613211059495098983425170669956869510721709169853401674655723866923579293791350126129000490700313616022730961734381243556039455811085004570914745600363312353534142465291053494925235208980194886768645228506330878;
            6'd4: xpb[156] = 1024'd80779391587314296313211729718654339710977664661479374962197906287093840279009474280516729208220284611319313055160315610508184048598534072575453054524678847009362115059344243575081345872976129937281231902357485944081834152460483598029442173205314184905258109913875682717922214930992884915103231642554278784950;
            6'd5: xpb[156] = 1024'd38940891642080499692115198445910708266372867263981376638681455326378852680107273395638375902946518609427566615221647795845698140327557423441736255647683038294857306539394695800036562745461559560946441073753237506920112265465156111054313431665028006498162685685286074382349504626776789635319694639880051239022;
            6'd6: xpb[156] = 1024'd121169087380971444469817594577981509566466496992219062443296859430640760418514211420775093812330426916978969582740473415762276072897801108863179581787018270514043172589016365362622018809464194905921847853536228916122751228690725397044163259807971277357887164870813524076883322396489327372654847463831418177425;
            6'd7: xpb[156] = 1024'd79330587435737647848721063305237878121861699594721064119780408469925772819612010535896740507056660915087223142801805601099790164626824459729462782910022461799538364069066817587577235681949624529587057024931980478961029341695397910069034518267685098950791740642223915741310612092273232092871310461157190631497;
            6'd8: xpb[156] = 1024'd37492087490503851227624532032494246677256902197223065796263957509210785220709809651018387201782894913195476702863137786437304256355847810595745984033026653085033555549117269812532452554435054153252266196327732041799307454700070423093905776727398920543696316413634307405737901788057136813087773458482963085569;
            6'd9: xpb[156] = 1024'd119720283229394796005326928164565047977350531925460751600879361613472692959116747676155105111166803220746879670381963406353882188926091496017189310172361885304219421598738939375117908618437689498227672976110723451001946417925639709083755604870342191403420795599161757100271719557769674550422926282434330023972;
            6'd10: xpb[156] = 1024'd77881783284160999384230396891821416532745734527962753277362910652757705360214546791276751805893037218855133230443295591691396280655114846883472511295366076589714613078789391600073125490923119121892882147506475013840224530930312222108626863330056012996325371370572148764699009253553579270639389279760102478044;
            6'd11: xpb[156] = 1024'd36043283338927202763133865619077785088140937130464754953846459692042717761312345906398398500619271216963386790504627777028910372384138197749755712418370267875209804558839843825028342363408548745558091318902226576678502643934984735133498121789769834589229947141982540429126298949337483990855852277085874932116;
            6'd12: xpb[156] = 1024'd118271479077818147540836261751148586388234566858702440758461863796304625499719283931535116410003179524514789758023453396945488304954381883171199038557705500094395670608461513387613798427411184090533498098685217985881141607160554021123347949932713105448954426327509990123660116719050021728191005101037241870519;
            6'd13: xpb[156] = 1024'd76432979132584350919739730478404954943629769461204442434945412835589637900817083046656763104729413522623043318084785582283002396683405234037482239680709691379890862088511965612569015299896613714198707270080969548719419720165226534148219208392426927041859002098920381788087406414833926448407468098363014324591;
            6'd14: xpb[156] = 1024'd34594479187350554298643199205661323499024972063706444111428961874874650301914882161778409799455647520731296878146117767620516488412428584903765440803713882665386053568562417837524232172382043337863916441476721111557697833169899047173090466852140748634763577870330773452514696110617831168623931095688786778663;
            6'd15: xpb[156] = 1024'd116822674926241499076345595337732124799118601791944129916044365979136558040321820186915127708839555828282699845664943387537094420982672270325208766943049114884571919618184087400109688236384678682839323221259712520760336796395468333162940294995084019494488057055858223147048513880330368905959083919640153717066;
            6'd16: xpb[156] = 1024'd74984174981007702455249064064988493354513804394446131592527915018421570441419619302036774403565789826390953405726275572874608512711695621191491968066053306170067111098234539625064905108870108306504532392655464083598614909400140846187811553454797841087392632827268614811475803576114273626175546916965926171138;
            6'd17: xpb[156] = 1024'd33145675035773905834152532792244861909909006996948133269011464057706582842517418417158421098292023824499206965787607758212122604440718972057775169189057497455562302578284991850020121981355537930169741564051215646436893022404813359212682811914511662680297208598679006475903093271898178346392009914291698625210;
            6'd18: xpb[156] = 1024'd115373870774664850611854928924315663210002636725185819073626868161968490580924356442295139007675932132050609933306433378128700537010962657479218495328392729674748168627906661412605578045358173275145148343834207055639531985630382645202532640057454933540021687784206456170436911041610716083727162738243065563613;
            6'd19: xpb[156] = 1024'd73535370829431053990758397651572031765397839327687820750110417201253502982022155557416785702402166130158863493367765563466214628739986008345501696451396920960243360107957113637560794917843602898810357515229958618477810098635055158227403898517168755132926263555616847834864200737394620803943625735568838017685;
            6'd20: xpb[156] = 1024'd31696870884197257369661866378828400320793041930189822426593966240538515383119954672538432397128400128267117053429097748803728720469009359211784897574401112245738551588007565862516011790329032522475566686625710181316088211639727671252275156976882576725830839327027239499291490433178525524160088732894610471757;
            6'd21: xpb[156] = 1024'd113925066623088202147364262510899201620886671658427508231209370344800423121526892697675150306512308435818520020947923368720306653039253044633228223713736344464924417637629235425101467854331667867450973466408701590518727174865296957242124985119825847585555318512554689193825308202891063261495241556845977410160;
            6'd22: xpb[156] = 1024'd72086566677854405526267731238155570176281874260929509907692919384085435522624691812796797001238542433926773581009255554057820744768276395499511424836740535750419609117679687650056684726817097491116182637804453153357005287869969470266996243579539669178459894283965080858252597898674967981711704554171749864232;
            6'd23: xpb[156] = 1024'd30248066732620608905171199965411938731677076863431511584176468423370447923722490927918443695964776432035027141070587739395334836497299746365794625959744727035914800597730139875011901599302527114781391809200204716195283400874641983291867502039253490771364470055375472522679887594458872701928167551497522318304;
            6'd24: xpb[156] = 1024'd112476262471511553682873596097482740031770706591669197388791872527632355662129428953055161605348684739586430108589413359311912769067543431787237952099079959255100666647351809437597357663305162459756798588983196125397922364100211269281717330182196761631088949240902922217213705364171410439263320375448889256707;
            6'd25: xpb[156] = 1024'd70637762526277757061777064824739108587165909194171199065275421566917368063227228068176808300074918737694683668650745544649426860796566782653521153222084150540595858127402261662552574535790592083422007760378947688236200477104883782306588588641910583223993525012313313881640995059955315159479783372774661710779;
            6'd26: xpb[156] = 1024'd28799262581043960440680533551995477142561111796673200741758970606202380464325027183298454994801152735802937228712077729986940952525590133519804354345088341826091049607452713887507791408276021707087216931774699251074478590109556295331459847101624404816898100783723705546068284755739219879696246370100434164851;
            6'd27: xpb[156] = 1024'd111027458319934905218382929684066278442654741524910886546374374710464288202731965208435172904185061043354340196230903349903518885095833818941247680484423574045276915657074383450093247472278657052062623711557690660277117553335125581321309675244567675676622579969251155240602102525451757617031399194051801103254;
            6'd28: xpb[156] = 1024'd69188958374701108597286398411322646998049944127412888222857923749749300603829764323556819598911295041462593756292235535241032976824857169807530881607427765330772107137124835675048464344764086675727832882953442223115395666339798094346180933704281497269527155740661546905029392221235662337247862191377573557326;
            6'd29: xpb[156] = 1024'd27350458429467311976189867138579015553445146729914889899341472789034313004927563438678466293637529039570847316353567720578547068553880520673814082730431956616267298617175287900003681217249516299393042054349193785953673779344470607371052192163995318862431731512071938569456681917019567057464325188703346011398;
            6'd30: xpb[156] = 1024'd109578654168358256753892263270649816853538776458152575703956876893296220743334501463815184203021437347122250283872393340495125001124124206095257408869767188835453164666796957462589137281252151644368448834132185195156312742570039893360902020306938589722156210697599388263990499686732104794799478012654712949801;
            6'd31: xpb[156] = 1024'd67740154223124460132795731997906185408933979060654577380440425932581233144432300578936830897747671345230503843933725525832639092853147556961540609992771380120948356146847409687544354153737581268033658005527936757994590855574712406385773278766652411315060786469009779928417789382516009515015941009980485403873;
            6'd32: xpb[156] = 1024'd25901654277890663511699200725162553964329181663156579056923974971866245545530099694058477592473905343338757403995057711170153184582170907827823811115775571406443547626897861912499571026223010891698867176923688320832868968579384919410644537226366232907965362240420171592845079078299914235232404007306257857945;
            6'd33: xpb[156] = 1024'd108129850016781608289401596857233355264422811391394264861539379076128153283937037719195195501857813650890160371513883331086731117152414593249267137255110803625629413676519531475085027090225646236674273956706679730035507931804954205400494365369309503767689841425947621287378896848012451972567556831257624796348;
            6'd34: xpb[156] = 1024'd66291350071547811668305065584489723819818013993896266538022928115413165685034836834316842196584047648998413931575215516424245208881437944115550338378114994911124605156569983700040243962711075860339483128102431292873786044809626718425365623829023325360594417197358012951806186543796356692784019828583397250420;
            6'd35: xpb[156] = 1024'd24452850126314015047208534311746092375213216596398268214506477154698178086132635949438488891310281647106667491636547701761759300610461294981833539501119186196619796636620435924995460835196505484004692299498182855712064157814299231450236882288737146953498992968768404616233476239580261413000482825909169704492;
            6'd36: xpb[156] = 1024'd106681045865204959824910930443816893675306846324635954019121881258960085824539573974575206800694189954658070459155373321678337233180704980403276865640454418415805662686242105487580916899199140828980099079281174264914703121039868517440086710431680417813223472154295854310767294009292799150335635649860536642895;
            6'd37: xpb[156] = 1024'd64842545919971163203814399171073262230702048927137955695605430298245098225637373089696853495420423952766324019216705507015851324909728331269560066763458609701300854166292557712536133771684570452645308250676925827752981234044541030464957968891394239406128047925706245975194583705076703870552098647186309096967;
            6'd38: xpb[156] = 1024'd23004045974737366582717867898329630786097251529639957372088979337530110626735172204818500190146657950874577579278037692353365416638751682135843267886462800986796045646343009937491350644170000076310517422072677390591259347049213543489829227351108060999032623697116637639621873400860608590768561644512081551039;
            6'd39: xpb[156] = 1024'd105232241713628311360420264030400432086190881257877643176704383441792018365142110229955218099530566258425980546796863312269943349208995367557286594025798033205981911695964679500076806708172635421285924201855668799793898310274782829479679055494051331858757102882644087334155691170573146328103714468463448489442;
            6'd40: xpb[156] = 1024'd63393741768394514739323732757656800641586083860379644853187932481077030766239909345076864794256800256534234106858195497607457440938018718423569795148802224491477103176015131725032023580658065044951133373251420362632176423279455342504550313953765153451661678654054478998582980866357051048320177465789220943514;
            6'd41: xpb[156] = 1024'd21555241823160718118227201484913169196981286462881646529671481520362043167337708460198511488983034254642487666919527682944971532667042069289852996271806415776972294656065583949987240453143494668616342544647171925470454536284127855529421572413478975044566254425464870663010270562140955768536640463114993397586;
            6'd42: xpb[156] = 1024'd103783437562051662895929597616983970497074916191119332334286885624623950905744646485335229398366942562193890634438353302861549465237285754711296322411141647996158160705687253512572696517146130013591749324430163334673093499509697141519271400556422245904290733610992320357544088331853493505871793287066360335989;
            6'd43: xpb[156] = 1024'd61944937616817866274833066344240339052470118793621334010770434663908963306842445600456876093093176560302144194499685488199063556966309105577579523534145839281653352185737705737527913389631559637256958495825914897511371612514369654544142659016136067497195309382402712021971378027637398226088256284392132790061;
            6'd44: xpb[156] = 1024'd20106437671584069653736535071496707607865321396123335687253983703193975707940244715578522787819410558410397754561017673536577648695332456443862724657150030567148543665788157962483130262116989260922167667221666460349649725519042167569013917475849889090099885153813103686398667723421302946304719281717905244133;
            6'd45: xpb[156] = 1024'd102334633410475014431438931203567508907958951124361021491869387807455883446347182740715240697203318865961800722079843293453155581265576141865306050796485262786334409715409827525068586326119624605897574447004657869552288688744611453558863745618793159949824364339340553380932485493133840683639872105669272182536;
            6'd46: xpb[156] = 1024'd60496133465241217810342399930823877463354153726863023168352936846740895847444981855836887391929552864070054282141175478790669672994599492731589251919489454071829601195460279750023803198605054229562783618400409432390566801749283966583735004078506981542728940110750945045359775188917745403856335102995044636608;
            6'd47: xpb[156] = 1024'd18657633520007421189245868658080246018749356329365024844836485886025908248542780970958534086655786862178307842202507664128183764723622843597872453042493645357324792675510731974979020071090483853227992789796160995228844914753956479608606262538220803135633515882161336709787064884701650124072798100320817090680;
            6'd48: xpb[156] = 1024'd100885829258898365966948264790151047318842986057602710649451889990287815986949718996095251996039695169729710809721333284044761697293866529019315779181828877576510658725132401537564476135093119198203399569579152404431483877979525765598456090681164073995357995067688786404320882654414187861407950924272184029083;
            6'd49: xpb[156] = 1024'd59047329313664569345851733517407415874238188660104712325935439029572828388047518111216898690765929167837964369782665469382275789022889879885598980304833068862005850205182853762519693007578548821868608740974903967269761990984198278623327349140877895588262570839099178068748172350198092581624413921597956483155;
            6'd50: xpb[156] = 1024'd17208829368430772724755202244663784429633391262606714002418988068857840789145317226338545385492163165946217929843997654719789880751913230751882181427837260147501041685233305987474909880063978445533817912370655530108040103988870791648198607600591717181167146610509569733175462045981997301840876918923728937227;
            6'd51: xpb[156] = 1024'd99437025107321717502457598376734585729727020990844399807034392173119748527552255251475263294876071473497620897362823274636367813322156916173325507567172492366686907734854975550060365944066613790509224692153646939310679067214440077638048435743534988040891625796037019427709279815694535039176029742875095875630;
            6'd52: xpb[156] = 1024'd57598525162087920881361067103990954285122223593346401483517941212404760928650054366596909989602305471605874457424155459973881905051180267039608708690176683652182099214905427775015582816552043414174433863549398502148957180219112590662919694203248809633796201567447411092136569511478439759392492740200868329702;
            6'd53: xpb[156] = 1024'd15760025216854124260264535831247322840517426195848403160001490251689773329747853481718556684328539469714128017485487645311395996780203617905891909813180874937677290694955879999970799689037473037839643034945150064987235293223785103687790952662962631226700777338857802756563859207262344479608955737526640783774;
            6'd54: xpb[156] = 1024'd97988220955745069037966931963318124140611055924086088964616894355951681068154791506855274593712447777265530985004313265227973929350447303327335235952516107156863156744577549562556255753040108382815049814728141474189874256449354389677640780805905902086425256524385252451097676976974882216944108561478007722177;
            6'd55: xpb[156] = 1024'd56149721010511272416870400690574492696006258526588090641100443395236693469252590621976921288438681775373784545065645450565488021079470654193618437075520298442358348224628001787511472625525538006480258986123893037028152369454026902702512039265619723679329832295795644115524966672758786937160571558803780176249;
            6'd56: xpb[156] = 1024'd14311221065277475795773869417830861251401461129090092317583992434521705870350389737098567983164915773482038105126977635903002112808494005059901638198524489727853539704678454012466689498010967630145468157519644599866430482458699415727383297725333545272234408067206035779952256368542691657377034556129552630321;
            6'd57: xpb[156] = 1024'd96539416804168420573476265549901662551495090857327778122199396538783613608757327762235285892548824081033441072645803255819580045378737690481344964337859721947039405754300123575052145562013602975120874937302636009069069445684268701717233125868276816131958887252733485474486074138255229394712187380080919568724;
            6'd58: xpb[156] = 1024'd54700916858934623952379734277158031106890293459829779798682945578068626009855126877356932587275058079141694632707135441157094137107761041347628165460863913232534597234350575800007362434499032598786084108698387571907347558688941214742104384327990637724863463024143877138913363834039134114928650377406692022796;
            6'd59: xpb[156] = 1024'd12862416913700827331283203004414399662285496062331781475166494617353638410952925992478579282001292077249948192768467626494608228836784392213911366583868104518029788714401028024962579306984462222451293280094139134745625671693613727766975642787704459317768038795554268803340653529823038835145113374732464476868;
            6'd60: xpb[156] = 1024'd95090612652591772108985599136485200962379125790569467279781898721615546149359864017615297191385200384801351160287293246411186161407028077635354692723203336737215654764022697587548035370987097567426700059877130543948264634919183013756825470930647730177492517981081718497874471299535576572480266198683831415271;
            6'd61: xpb[156] = 1024'd53252112707357975487889067863741569517774328393071468956265447760900558550457663132736943886111434382909604720348625431748700253136051428501637893846207528022710846244073149812503252243472527191091909231272882106786542747923855526781696729390361551770397093752492110162301760995319481292696729196009603869343;
            6'd62: xpb[156] = 1024'd11413612762124178866792536590997938073169530995573470632748996800185570951555462247858590580837668381017858280409957617086214344865074779367921094969211719308206037724123602037458469115957956814757118402668633669624820860928528039806567987850075373363301669523902501826729050691103386012913192193335376323415;
            6'd63: xpb[156] = 1024'd93641808501015123644494932723068739373263160723811156437364400904447478689962400272995308490221576688569261247928783237002792277435318464789364421108546951527391903773745271600043925179960592159732525182451625078827459824154097325796417815993018644223026148709429951521262868460815923750248345017286743261818;
        endcase
    end

    always_comb begin
        case(flag[52][11:6])
            6'd0: xpb[157] = 1024'd0;
            6'd1: xpb[157] = 1024'd51803308555781327023398401450325107928658363326313158113847949943732491091060199388116955184947810686677514807990115422340306369164341815655647622231551142812887095253795723824999142052446021783397734353847376641665737937158769838821289074452732465815930724480840343185690158156599828470464808014612515715890;
            6'd2: xpb[157] = 1024'd103606617111562654046796802900650215857316726652626316227695899887464982182120398776233910369895621373355029615980230844680612738328683631311295244463102285625774190507591447649998284104892043566795468707694753283331475874317539677642578148905464931631861448961680686371380316313199656940929616029225031431780;
            6'd3: xpb[157] = 1024'd31343229983219239671396276946160891041276662853203790213411994766220577935871459254335794340185757750589395016512852832441855266651805112411782741678322387504970611191815954137367186965820859628883005453154890078632852961255412743498888653674967948180972270028403971526963946395870852394275734217211952663339;
            6'd4: xpb[157] = 1024'd83146538539000566694794678396485998969935026179516948327259944709953069026931658642452749525133568437266909824502968254782161635816146928067430363909873530317857706445611677962366329018266881412280739807002266720298590898414182582320177728127700413996902994509244314712654104552470680864740542231824468379229;
            6'd5: xpb[157] = 1024'd10883151410657152319394152441996674153894962380094422312976039588708664780682719120554633495423704814501275225035590242543404164139268409167917861125093632197054127129836184449735231879195697474368276552462403515599967985352055648176488232897203430546013815575967599868237734635141876318086660419811389610788;
            6'd6: xpb[157] = 1024'd62686459966438479342792553892321782082553325706407580426823989532441155871742918508671588680371515501178790033025705664883710533303610224823565483356644775009941222383631908274734373931641719257766010906309780157265705922510825486997777307349935896361944540056807943053927892791741704788551468434423905326678;
            6'd7: xpb[157] = 1024'd114489768522219806366190955342646890011211689032720738540671939476173646962803117896788543865319326187856304841015821087224016902467952040479213105588195917822828317637427632099733515984087741041163745260157156798931443859669595325819066381802668362177875264537648286239618050948341533259016276449036421042568;
            6'd8: xpb[157] = 1024'd42226381393876391990790429388157565195171625233298212526388034354929242716554178374890427835609462565090670241548443074985259430791073521579700602803416019702024738321652138587102418845016557103251282005617293594232820946607468391675376886572171378726986085604371571395201681031012728712362394637023342274127;
            6'd9: xpb[157] = 1024'd94029689949657719014188830838482673123829988559611370640235984298661733807614377763007383020557273251768185049538558497325565799955415337235348225034967162514911833575447862412101560897462578886649016359464670235898558883766238230496665961024903844542916810085211914580891839187612557182827202651635857990017;
            6'd10: xpb[157] = 1024'd21766302821314304638788304883993348307789924760188844625952079177417329561365438241109266990847409629002550450071180485086808328278536818335835722250187264394108254259672368899470463758391394948736553104924807031199935970704111296352976465794406861092027631151935199736475469270283752636173320839622779221576;
            6'd11: xpb[157] = 1024'd73569611377095631662186706334318456236448288086502002739800029121149820652425637629226222175795220315680065258061295907427114697442878633991483344481738407206995349513468092724469605810837416732134287458772183672865673907862881135174265540247139326907958355632775542922165627426883581106638128854235294937466;
            6'd12: xpb[157] = 1024'd1306224248752217286786180379829131420408224287079476725516123999905416406176698107328106146085356692914430658593917895188357225766000115091970841696958509086191770197692599211838508671766232794221824204232320468167050994800754201030576045016642343457069176699498828077749257509554776559984247042222216169025;
            6'd13: xpb[157] = 1024'd53109532804533544310184581830154239349066587613392634839364073943637907497236897495445061331033167379591945466584033317528663594930341930747618463928509651899078865451488323036837650724212254577619558558079697109832788931959524039851865119469374809272999901180339171263439415666154605030449055056834731884915;
            6'd14: xpb[157] = 1024'd104912841360314871333582983280479347277724950939705792953212023887370398588297096883562016515980978066269460274574148739868969964094683746403266086160060794711965960705284046861836792776658276361017292911927073751498526869118293878673154193922107275088930625661179514449129573822754433500913863071447247600805;
            6'd15: xpb[157] = 1024'd32649454231971456958182457325990022461684887140283266938928118766125994342048157361663900486271114443503825675106770727630212492417805227503753583375280896591162381389508553349205695637587092423104829657387210546799903956056166944529464698691610291638041446727902799604713203905425628954259981259434168832364;
            6'd16: xpb[157] = 1024'd84452762787752783981580858776315130390343250466596425052776068709858485433108356749780855671218925130181340483096886149970518861582147043159401205606832039404049476643304277174204837690033114206502564011234587188465641893214936783350753773144342757453972171208743142790403362062025457424724789274046684548254;
            6'd17: xpb[157] = 1024'd12189375659409369606180332821825805574303186667173899038492163588614081186859417227882739641509061507415705883629508137731761389905268524259888702822052141283245897327528783661573740550961930268590100756694723983767018980152809849207064277913845774003082992275466427945986992144696652878070907462033605779813;
            6'd18: xpb[157] = 1024'd63992684215190696629578734272150913502961549993487057152340113532346572277919616615999694826456872194093220691619623560072067759069610339915536325053603284096132992581324507486572882603407952051987835110542100625432756917311579688028353352366578239819013716756306771131677150301296481348535715476646121495703;
            6'd19: xpb[157] = 1024'd115795992770972023652977135722476021431619913319800215266188063476079063368979816004116650011404682880770735499609738982412374128233952155571183947285154426909020087835120231311572024655853973835385569464389477267098494854470349526849642426819310705634944441237147114317367308457896309819000523491258637211593;
            6'd20: xpb[157] = 1024'd43532605642628609277576609767986696615579849520377689251904158354834659122730876482218533981694819258005100900142360970173616656557073636671671444500374528788216508519344737798940927516782789897473106209849614062399871941408222592705952931588813722184055262303870399472950938540567505272346641679245558443152;
            6'd21: xpb[157] = 1024'd95335914198409936300975011218311804544238212846690847365752108298567150213791075870335489166642629944682615708132476392513923025721415452327319066731925671601103603773140461623940069569228811680870840563696990704065609878566992431527242006041546187999985986784710742658641096697167333742811449693858074159042;
            6'd22: xpb[157] = 1024'd23072527070066521925574485263822479728198149047268321351468203177322745967542136348437373136932766321916981108665098380275165554044536933427806563947145773480300024457364968111308972430157627742958377309157127499366986965504865497383552510811049204549096807851434027814224726779838529196157567881844995390601;
            6'd23: xpb[157] = 1024'd74875835625847848948972886714147587656856512373581479465316153121055237058602335736554328321880577008594495916655213802615471923208878749083454186178696916293187119711160691936308114482603649526356111663004504141032724902663635336204841585263781670365027532332274370999914884936438357666622375896457511106491;
            6'd24: xpb[157] = 1024'd2612448497504434573572360759658262840816448574158953451032247999810832812353396214656212292170713385828861317187835790376714451532000230183941683393917018172383540395385198423677017343532465588443648408464640936334101989601508402061152090033284686914138353398997656155498515019109553119968494084444432338050;
            6'd25: xpb[157] = 1024'd54415757053285761596970762209983370769474811900472111564880197943543323903413595602773167477118524072506376125177951212717020820696342045839589305625468160985270635649180922248676159395978487371841382762312017577999839926760278240882441164486017152730069077879837999341188673175709381590433302099056948053940;
            6'd26: xpb[157] = 1024'd106219065609067088620369163660308478698133175226785269678728147887275814994473794990890122662066334759183890933168066635057327189860683861495236927857019303798157730902976646073675301448424509155239117116159394219665577863919048079703730238938749618545999802360678342526878831332309210060898110113669463769830;
            6'd27: xpb[157] = 1024'd33955678480723674244968637705819153882093111427362743664444242766031410748224855468992006632356471136418256333700688622818569718183805342595724425072239405677354151587201152561044204309353325217326653861619531014966954950856921145560040743708252635095110623427401627682462461414980405514244228301656385001389;
            6'd28: xpb[157] = 1024'd85758987036505001268367039156144261810751474753675901778292192709763901839285054857108961817304281823095771141690804045158876087348147158251372047303790548490241246840996876386043346361799347000724388215466907656632692888015690984381329818160985100911041347908241970868152619571580233984709036316268900717279;
            6'd29: xpb[157] = 1024'd13495599908161586892966513201654936994711410954253375764008287588519497593036115335210845787594418200330136542223426032920118615671268639351859544519010650369437667525221382873412249222728163062811924960927044451934069974953564050237640322930488117460152168974965256023736249654251429438055154504255821948838;
            6'd30: xpb[157] = 1024'd65298908463942913916364914651980044923369774280566533877856237532251988684096314723327800972542228887007651350213541455260424984835610455007507166750561793182324762779017106698411391275174184846209659314774421093599807912112333889058929397383220583276082893455805599209426407810851257908519962518868337664728;
            6'd31: xpb[157] = 1024'd117102217019724240939763316102305152852028137606879691991704187475984479775156514111444756157490039573685166158203656877600731353999952270663154788982112935995211858032812830523410533327620206629607393668621797735265545849271103727880218471835953049092013617936645942395116565967451086378984770533480853380618;
            6'd32: xpb[157] = 1024'd44838829891380826564362790147815828035988073807457165977420282354740075528907574589546640127780175950919531558736278865361973882323073751763642286197333037874408278717037337010779436188549022691694930414081934530566922936208976793736528976605456065641124439003369227550700196050122281832330888721467774612177;
            6'd33: xpb[157] = 1024'd96642138447162153587761191598140935964646437133770324091268232298472566619967773977663595312727986637597046366726394287702280251487415567419289908428884180687295373970833060835778578240995044475092664767929311172232660873367746632557818051058188531457055163484209570736390354206722110302795696736080290328067;
            6'd34: xpb[157] = 1024'd24378751318818739212360665643651611148606373334347798076984327177228162373718834455765479283018123014831411767259016275463522779810537048519777405644104282566491794655057567323147481101923860537180201513389447967534037960305619698414128555827691548006165984550932855891973984289393305756141814924067211559626;
            6'd35: xpb[157] = 1024'd76182059874600066235759067093976719077264736660660956190832277120960653464779033843882434467965933701508926575249131697803829148974878864175425027875655425379378889908853291148146623154369882320577935867236824609199775897464389537235417630280424013822096709031773199077664142445993134226606622938679727275516;
            6'd36: xpb[157] = 1024'd3918672746256651860358541139487394261224672861238430176548371999716249218530094321984318438256070078743291975781753685565071677298000345275912525090875527258575310593077797635515526015298698382665472612696961404501152984402262603091728135049927030371207530098496484233247772528664329679952741126666648507075;
            6'd37: xpb[157] = 1024'd55721981302037978883756942589812502189883036187551588290396321943448740309590293710101273623203880765420806783771869107905378046462342160931560147322426670071462405846873521460514668067744720166063206966544338046166890921561032441913017209502659496187138254579336827418937930685264158150417549141279164222965;
            6'd38: xpb[157] = 1024'd107525289857819305907155344040137610118541399513864746404244271887181231400650493098218228808151691452098321591761984530245684415626683976587207769553977812884349501100669245285513810120190741949460941320391714687832628858719802280734306283955391962003068979060177170604628088841863986620882357155891679938855;
            6'd39: xpb[157] = 1024'd35261902729475891531754818085648285302501335714442220389960366765936827154401553576320112778441827829332686992294606518006926943949805457687695266769197914763545921784893751772882712981119558011548478065851851483134005945657675346590616788724894978552179800126900455760211718924535182074228475343878601170414;
            6'd40: xpb[157] = 1024'd87065211285257218555153219535973393231159699040755378503808316709669318245461752964437067963389638516010201800284721940347233313114147273343342889000749057576433017038689475597881855033565579794946212419699228124799743882816445185411905863177627444368110524607740798945901877081135010544693283358491116886304;
            6'd41: xpb[157] = 1024'd14801824156913804179752693581484068415119635241332852489524411588424913999212813442538951933679774893244567200817343928108475841437268754443830386215969159455629437722913982085250757894494395857033749165159364920101120969754318251268216367947130460917221345674464084101485507163806205998039401546478038117863;
            6'd42: xpb[157] = 1024'd66605132712695131203151095031809176343777998567646010603372361532157405090273012830655907118627585579922082008807459350448782210601610570099478008447520302268516532976709705910249899946940417640431483519006741561766858906913088090089505442399862926733152070155304427287175665320406034468504209561090553833753;
            6'd43: xpb[157] = 1024'd118408441268476458226549496482134284272436361893959168717220311475889896181333212218772862303575396266599596816797574772789088579765952385755125630679071445081403628230505429735249041999386439423829217872854118203432596844071857928910794516852595392549082794636144770472865823477005862938969017575703069549643;
            6'd44: xpb[157] = 1024'd46145054140133043851148970527644959456396298094536642702936406354645491935084272696874746273865532643833962217330196760550331108089073866855613127894291546960600048914729936222617944860315255485916754618314254998733973931009730994767105021622098409098193615702868055628449453559677058392315135763689990781202;
            6'd45: xpb[157] = 1024'd97948362695914370874547371977970067385054661420849800816784356298377983026144472084991701458813343330511477025320312182890637477253415682511260750125842689773487144168525660047617086912761277269314488972161631640399711868168500833588394096074830874914124340183708398814139611716276886862779943778302506497092;
            6'd46: xpb[157] = 1024'd25684975567570956499146846023480742569014597621427274802500451177133578779895532563093585429103479707745842425852934170651880005576537163611748247341062791652683564852750166534985989773690093331402025717621768435701088955106373899444704600844333891463235161250431683969723241798948082316126061966289427728651;
            6'd47: xpb[157] = 1024'd77488284123352283522545247473805850497672960947740432916348401120866069870955731951210540614051290394423357233843049592992186374740878979267395869572613934465570660106545890359985131826136115114799760071469145077366826892265143738265993675297066357279165885731272027155413399955547910786590869980901943444541;
            6'd48: xpb[157] = 1024'd5224896995008869147144721519316525681632897148317906902064495999621665624706792429312424584341426771657722634375671580753428903064000460367883366787834036344767080790770396847354034687064931176887296816929281872668203979203016804122304180066569373828276706797995312310997030038219106239936988168888864676100;
            6'd49: xpb[157] = 1024'd57028205550790196170543122969641633610291260474631065015912445943354156715766991817429379769289237458335237442365787003093735272228342276023530989019385179157654176044566120672353176739510952960285031170776658514333941916361786642943593254519301839644207431278835655496687188194818934710401796183501380391990;
            6'd50: xpb[157] = 1024'd108831514106571523193941524419966741538949623800944223129760395887086647806827191205546334954237048145012752250355902425434041641392684091679178611250936321970541271298361844497352318791956974743682765524624035155999679853520556481764882328972034305460138155759675998682377346351418763180866604198113896107880;
            6'd51: xpb[157] = 1024'd36568126978228108818540998465477416722909560001521697115476490765842243560578251683648218924527184522247117650888524413195284169715805572779666108466156423849737691982586350984721221652885790805770302270084171951301056940458429547621192833741537322009248976826399283837960976434089958634212722386100817339439;
            6'd52: xpb[157] = 1024'd88371435534009435841939399915802524651567923327834855229324440709574734651638451071765174109474995208924632458878639835535590538880147388435313730697707566662624787236382074809720363705331812589168036623931548592966794877617199386442481908194269787825179701307239627023651134590689787104677530400713333055329;
            6'd53: xpb[157] = 1024'd16108048405666021466538873961313199835527859528412329215040535588330330405389511549867058079765131586158997859411261823296833067203268869535801227912927668541821207920606581297089266566260628651255573369391685388268171964555072452298792412963772804374290522373962912179234764673360982558023648588700254286888;
            6'd54: xpb[157] = 1024'd67911356961447348489937275411638307764186222854725487328888485532062821496449710937984013264712942272836512667401377245637139436367610685191448850144478811354708303174402305122088408618706650434653307723239062029933909901713842291120081487416505270190221246854803255364924922829960811028488456603312770002778;
            6'd55: xpb[157] = 1024'd119714665517228675513335676861963415692844586181038645442736435475795312587509910326100968449660752959514027475391492667977445805531952500847096472376029954167595398428198028947087550671152672218051042077086438671599647838872612129941370561869237736006151971335643598550615080986560639498953264617925285718668;
            6'd56: xpb[157] = 1024'd47451278388885261137935150907474090876804522381616119428452530354550908341260970804202852419950889336748392875924114655738688333855073981947583969591250056046791819112422535434456453532081488280138578822546575466901024925810485195797681066638740752555262792402366883706198711069231834952299382805912206950227;
            6'd57: xpb[157] = 1024'd99254586944666588161333552357799198805462885707929277542300480298283399432321170192319807604898700023425907683914230078078994703019415797603231591822801198859678914366218259259455595584527510063536313176393952108566762862969255034618970141091473218371193516883207226891888869225831663422764190820524722666117;
            6'd58: xpb[157] = 1024'd26991199816323173785933026403309873989422821908506751528016575177038995186072230670421691575188836400660273084446852065840237231342537278703719089038021300738875335050442765746824498445456326125623849921854088903868139949907128100475280645860976234920304337949930512047472499308502858876110309008511643897676;
            6'd59: xpb[157] = 1024'd78794508372104500809331427853634981918081185234819909641864525120771486277132430058538646760136647087337787892436967488180543600506879094359366711269572443551762430304238489571823640497902347909021584275701465545533877887065897939296569720313708700736235062430770855233162657465102687346575117023124159613566;
            6'd60: xpb[157] = 1024'd6531121243761086433930901899145657102041121435397383627580619999527082030883490536640530730426783464572153292969589475941786128830000575459854208484792545430958850988462996059192543358831163971109121021161602340835254974003771005152880225083211717285345883497494140388746287547773882799921235211111080845125;
            6'd61: xpb[157] = 1024'd58334429799542413457329303349470765030699484761710541741428569943259573121943689924757485915374594151249668100959704898282092497994342391115501830716343688243845946242258719884191685411277185754506855375008978982500992911162540843974169299535944183101276607978334483574436445704373711270386043225723596561015;
            6'd62: xpb[157] = 1024'd110137738355323740480727704799795872959357848088023699855276519886992064213003889312874441100322404837927182908949820320622398867158684206771149452947894831056733041496054443709190827463723207537904589728856355624166730848321310682795458373988676648917207332459174826760126603860973539740850851240336112276905;
            6'd63: xpb[157] = 1024'd37874351226980326105327178845306548143317784288601173840992614765747659966754949790976325070612541215161548309482442308383641395481805687871636950163114932935929462180278950196559730324652023599992126474316492419468107935259183748651768878758179665466318153525898111915710233943644735194196969428323033508464;
        endcase
    end

    always_comb begin
        case(flag[52][16:12])
            5'd0: xpb[158] = 1024'd0;
            5'd1: xpb[158] = 1024'd89677659782761653128725580295631656071976147614914331954840564709480151057815149179093280255560351901839063117472557730723947764646147503527284572394666075748816557434074674021558872377098045383389860828163869061133845872417953587473057953210912131282248878006738455101400392100244563664661777442935549224354;
            5'd2: xpb[158] = 1024'd55288623881398564858652233186448879399253868104092979781549274353983406778321159448171489296463029494234976827487622026868831688451074672499409019773001110563942440298578130705487505562678885045469524047940498275903330894615010401981137336738594813297677852599359852172694256126560494312204865059245503964377;
            5'd3: xpb[158] = 1024'd20899587980035476588578886077266102726531588593271627608257983998486662498827169717249698337365707086630890537502686323013715612256001841471533467151336145379068323163081587389416138748259724707549187267717127490672815916812067216489216720266277495313106827191981249243988120152876424959747952675555458704400;
            5'd4: xpb[158] = 1024'd110577247762797129717304466372897758798507736208185959563098548707966813556642318896342978592926058988469953654975244053737663376902149344998818039546002221127884880597156261410975011125357770090939048095880996551806661789230020803962274673477189626595355705198719704345388512253120988624409730118491007928754;
            5'd5: xpb[158] = 1024'd76188211861434041447231119263714982125785456697364607389807258352470069277148329165421187633828736580865867364990308349882547300707076513970942486924337255943010763461659718094903644310938609753018711315657625766576146811427077618470354057004872308610784679791341101416682376279436919271952817734800962668777;
            5'd6: xpb[158] = 1024'd41799175960070953177157772154532205453063177186543255216515967996973324997654339434499396674731414173261781075005372646027431224512003682943066934302672290758136646326163174778832277496519449415098374535434254981345631833624134432978433440532554990626213654383962498487976240305752849919495905351110917408800;
            5'd7: xpb[158] = 1024'd7410140058707864907084425045349428780340897675721903043224677641476580718160349703577605715634091765657694785020436942172315148316930851915191381681007325573262529190666631462760910682100289077178037755210884196115116855821191247486512824060237672641642628976583895559270104332068780567038992967420872148823;
            5'd8: xpb[158] = 1024'd97087799841469518035810005340981084852317045290636234998065242350956731775975498882670885971194443667496757902492994672896262912963078355442475954075673401322079086624741305484319783059198334460567898583374753257248962728239144834959570777271149803923891506983322350660670496432313344231700770410356421373177;
            5'd9: xpb[158] = 1024'd62698763940106429765736658231798308179594765779814882824773951995459987496481509151749095012097121259892671612508058969041146836768005524414600401454008436137204969489244762168248416244779174122647561803151382472018447750436201649467650160798832485939320481575943747731964360458629274879243858026666376113200;
            5'd10: xpb[158] = 1024'd28309728038743341495663311122615531506872486268993530651482661639963243216987519420827304052999798852288585322523123265186030760572932693386724848832343470952330852353748218852177049430360013784727225022928011686787932772633258463975729544326515167954749456168565144803258224484945205526786945642976330853223;
            5'd11: xpb[158] = 1024'd117987387821504994624388891418247187578848633883907862606323226349443394274802668599920584308560150754127648439995680995909978525219080196914009421227009546701147409787822892873735921807458059168117085851091880747921778645051212051448787497537427299236998334175303599904658616585189769191448723085911880077577;
            5'd12: xpb[158] = 1024'd83598351920141906354315544309064410906126354373086510433031935993946649995308678868998793349462828346523562150010745292054862449024007365886133868605344581516273292652326349557664554993038898830196749070868509962691263667248268865956866881065109981252427308767924996975952480611505699838991810702221834817600;
            5'd13: xpb[158] = 1024'd49209316018778818084242197199881634233404074862265158259740645638449905715814689138077002390365505938919475860025809588199746372828934534858258315983679616331399175516829806241593188178619738492276412290645139177460748689445325680464946264592792663267856283360546394047246344637821630486534898318531789557623;
            5'd14: xpb[158] = 1024'd14820280117415729814168850090698857560681795351443806086449355282953161436320699407155211431268183531315389570040873884344630296633861703830382763362014651146525058381333262925521821364200578154356075510421768392230233711642382494973025648120475345283285257953167791118540208664137561134077985934841744297646;
            5'd15: xpb[158] = 1024'd104497939900177382942894430386330513632657942966358138041289919992433312494135848586248491686828535433154452687513431615068578061280009207357667335756680726895341615815407936947080693741298623537745936338585637453364079584060336082446083601331387476565534135959906246219940600764382124798739763377777293522000;
            5'd16: xpb[158] = 1024'd70108903998814294672821083277147736959935663455536785867998629636936568214641858855326700727731213025550366397528495911213461985084936376329791783135015761710467498679911393631009326926879463199825599558362266668133564606257392896954162984859070158580963110552527643291234464790698055446282850994087248262023;
            5'd17: xpb[158] = 1024'd35719868097451206402747736167964960287213383944715433694707339281439823935147869124404909768633890617946280107543560207358345908889863545301916230513350796525593381544414850314937960112460302861905262778138895882903049628454449711462242368386752840596392085145149040362528328817013986093825938610397203002046;
            5'd18: xpb[158] = 1024'd1330832196088118132674389058782183614491104433894081521416048925943079655653879393483118809536568210342193817558624503503229832694790714274040677891685831340719264408918306998866593298041142523984925997915525097672534650651506525970321751914435522611821059737770437433822192843329916741369026226707157742069;
            5'd19: xpb[158] = 1024'd91008491978849771261399969354413839686467252048808413476256613635423230713469028572576399065096920112181256935031182234227177597340938217801325250286351907089535821842992981020425465675139187907374786826079394158806380523069460113443379705125347653894069937744508892535222584943574480406030803669642706966423;
            5'd20: xpb[158] = 1024'd56619456077486682991326622245231063013744972537987061302965323279926486433975038841654608105999597704577170645046246530372061521145865386773449697664686941904661704707496437704354098860720027569454450045856023373575865545266516927951459088653030335909498912337130289606516448969890411053573891285952661706446;
            5'd21: xpb[158] = 1024'd22230420176123594721253275136048286341022693027165709129674032924429742154481049110732817146902275296973084355061310826516945444950792555745574145043021976719787587571999894388282732046300867231534113265632652588345350567463573742459538472180713017924927886929751686677810312996206341701116978902262616446469;
            5'd22: xpb[158] = 1024'd111908079958885247849978855431679942412998840642080041084514597633909893212296198289826097402462627198812147472533868557240893209596940059272858717437688052468604145006074568409841604423398912614923974093796521649479196439881527329932596425391625149207176764936490141779210705096450905365778756345198165670823;
            5'd23: xpb[158] = 1024'd77519044057522159579905508322497165740276561131258688911223307278413148932802208558904306443365304791208061182548932853385777133401867228244983164816023087283730027870578025093770237608979752277003637313573150864248681462078584144440675808919307831222605739529111538850504569122766836013321843961508120410846;
            5'd24: xpb[158] = 1024'd43130008156159071309832161213314389067554281620437336737932016922916404653308218827982515484267982383603974892563997149530661057206794397217107612194358122098855910735081481777698870794560591939083300533349780079018166484275640958948755192446990513238034714121732935921798433149082766660864931577818075150869;
            5'd25: xpb[158] = 1024'd8740972254795983039758814104131612394832002109615984564640726567419660373814229097060724525170659975999888602579061445675544981011721566189232059572693156913981793599584938461627503980141431601162963753126409293787651506472697773456834575974673195253463688714354332993092297175398697308408019194128029890892;
            5'd26: xpb[158] = 1024'd98418632037557636168484394399763268466808149724530316519481291276899811431629378276154004780731011877838951720051619176399492745657869069716516631967359232662798351033659612483186376357239476984552824581290278354921497378890651360929892529185585326535712566721092788094492689275643260973069796637063579115246;
            5'd27: xpb[158] = 1024'd64029596136194547898411047290580491794085870213708964346190000921403067152135388545232213821633689470234865430066683472544376669462796238688641079345694267477924233898163069167115009542820316646632487801066907569690982401087708175437971912713268008551141541313714185165786553301959191620612884253373533855269;
            5'd28: xpb[158] = 1024'd29640560234831459628337700181397715121363590702887612172898710565906322872641398814310422862536367062630779140081747768689260593267723407660765526724029302293050116762666525851043642728401156308712151020843536784460467423284764989946051296240950690566570515906335582237080417328275122268155971869683488595292;
            5'd29: xpb[158] = 1024'd119318220017593112757063280477029371193339738317801944127739275275386473930456547993403703118096718964469842257554305499413208357913870911188050099118695378041866674196741199872602515105499201692102011849007405845594313295702718577419109249451862821848819393913074037338480809428519685932817749312619037819646;
            5'd30: xpb[158] = 1024'd84929184116230024486989933367846594520617458806980591954447984919889729650962558262481912158999396556865755967569369795558092281718798080160174546497030412856992557061244656556531148291080041354181675068784035060363798317899775391927188632979545503864248368505695434409774673454835616580360836928928992559669;
            5'd31: xpb[158] = 1024'd50540148214866936216916586258663817847895179296159239781156694564392985371468568531560121199902074149261669677584434091702976205523725249132298993875365447672118439925748113240459781476660881016261338288560664275133283340096832206435268016507228185879677343098316831481068537481151547227903924545238947299692;
        endcase
    end

    always_comb begin
        case(flag[53][5:0])
            6'd0: xpb[159] = 1024'd0;
            6'd1: xpb[159] = 1024'd70108903998814294672821083277147736959935663455536785867998629636936568214641858855326700727731213025550366397528495911213461985084936376329791783135015761710467498679911393631009326926879463199825599558362266668133564606257392896954162984859070158580963110552527643291234464790698055446282850994087248262023;
            6'd2: xpb[159] = 1024'd16151112313503847946843239149481041175172899785337887607865404208896241091974578800638330240804751741657583387599498387847860129328652418104423441253700482487244322790251569924388414662241720678341001508337293489902768362293889020943347400034910867895106317690938228552362401507467477875447012161548902039715;
            6'd3: xpb[159] = 1024'd86260016312318142619664322426628778135108563240874673475864033845832809306616437655965030968535964767207949785127994299061322114413588794434215224388716244197711821470162963555397741589121183878166601066699560158036332968551281917897510384893981026476069428243465871843596866298165533321729863155636150301738;
            6'd4: xpb[159] = 1024'd32302224627007695893686478298962082350345799570675775215730808417792482183949157601276660481609503483315166775198996775695720258657304836208846882507400964974488645580503139848776829324483441356682003016674586979805536724587778041886694800069821735790212635381876457104724803014934955750894024323097804079430;
            6'd5: xpb[159] = 1024'd102411128625821990566507561576109819310281463026212561083729438054729050398591016456603361209340716508865533172727492686909182243742241212538638665642416726684956144260414533479786156251362904556507602575036853647939101330845170938840857784928891894371175745934404100395959267805633011197176875317185052341453;
            6'd6: xpb[159] = 1024'd48453336940511543840529717448443123525518699356013662823596212626688723275923736401914990722414255224972750162798495163543580387985957254313270323761101447461732968370754709773165243986725162035023004525011880469708305086881667062830042200104732603685318953072814685657087204522402433626341036484646706119145;
            6'd7: xpb[159] = 1024'd118562240939325838513350800725590860485454362811550448691594842263625291490565595257241691450145468250523116560326991074757042373070893630643062106896117209172200467050666103404174570913604625234848604083374147137841869693139059959784205184963802762266282063625342328948321669313100489072623887478733954381168;
            6'd8: xpb[159] = 1024'd64604449254015391787372956597924164700691599141351550431461616835584964367898315202553320963219006966630333550397993551391440517314609672417693765014801929948977291161006279697553658648966882713364006033349173959611073449175556083773389600139643471580425270763752914209449606029869911501788048646195608158860;
            6'd9: xpb[159] = 1024'd10646657568704945061395112470257468915928835471152652171328391407544637245231035147864950476292545682737550540468996028025838661558325714192325423133486650725754115271346455990932746384329140191879407983324200781380277205212052207762574015315484180894568477902163499470577542746639333930952209813657261936552;
            6'd10: xpb[159] = 1024'd80755561567519239734216195747405205875864498926689438039327021044481205459872894003191651204023758708287916937997491939239300646643262090522117206268502412436221613951257849621942073311208603391705007541686467449513841811469445104716737000174554339475531588454691142761812007537337389377235060807744510198575;
            6'd11: xpb[159] = 1024'd26797769882208793008238351619738510091101735256490539779193795616440878337205613948503280717097297424395133928068494415873698790886978132296748864387187133212998438061598025915321161046570860870220409491661494271283045567505941228705921415350395048789674795593101728022939944254106811806399221975206163976267;
            6'd12: xpb[159] = 1024'd96906673881023087681059434896886247051037398712027325647192425253377446551847472803829981444828510449945500325596990327087160775971914508626540647522202894923465936741509419546330487973450324070046009050023760939416610173763334125660084400209465207370637906145629371314174409044804867252682072969293412238290;
            6'd13: xpb[159] = 1024'd42948882195712640955081590769219551266274635041828427387059199825337119429180192749141610957902049166052717315667992803721558920215630550401172305640887615700242760851849595839709575708812581548561410999998787761185813929799830249649268815385305916684781113284039956575302345761574289681846234136755066015982;
            6'd14: xpb[159] = 1024'd113057786194526935627902674046367288226210298497365213255057829462273687643822051604468311685633262191603083713196488714935020905300566926730964088775903377410710259531760989470718902635692044748387010558361054429319378536057223146603431800244376075265744223836567599866536810552272345128129085130842314278005;
            6'd15: xpb[159] = 1024'd59099994509216488901924829918700592441447534827166314994924604034233360521154771549779941198706800907710300703267491191569419049544282968505595746894588098187487083642101165764097990371054302226902412508336081251088582292093719270592616215420216784579887430974978185127664747269041767557293246298303968055697;
            6'd16: xpb[159] = 1024'd5142202823906042175946985791033896656684771156967416734791378606193033398487491495091570711780339623817517693338493668203817193787999010280227405013272818964263907752441342057477078106416559705417814458311108072857786048130215394581800630596057493894030638113388770388792683985811189986457407465765621833389;
            6'd17: xpb[159] = 1024'd75251106822720336848768069068181633616620434612504202602790008243129601613129350350418271439511552649367884090866989579417279178872935386610019188148288580674731406432352735688486405033296022905243414016673374740991350654387608291535963615455127652474993748665916413680027148776509245432740258459852870095412;
            6'd18: xpb[159] = 1024'd21293315137409890122790224940514937831857670942305304342656782815089274490462070295729900952585091365475101080937992056051677323116651428384650846266973301451508230542692911981865492768658280383758815966648401562760554410424104415525148030630968361789136955804326998941155085493278667861904419627314523873104;
            6'd19: xpb[159] = 1024'd91402219136224184795611308217662674791793334397842090210655412452025842705103929151056601680316304391025467478466487967265139308201587804714442629401989063161975729222604305612874819695537743583584415525010668230894119016681497312479311015490038520370100066356854642232389550283976723308187270621401772135127;
            6'd20: xpb[159] = 1024'd37444427450913738069633464089995979007030570727643191950522187023985515582436649096368231193389843107132684468537490443899537452445303846489074287520673783938752553332944481906253907430900001062099817474985695052663322772717993436468495430665879229684243273495265227493517487000746145737351431788863425912819;
            6'd21: xpb[159] = 1024'd107553331449728032742454547367143715966966234183179977818520816660922083797078507951694931921121056132683050866065986355112999437530240222818866070655689545649220052012855875537263234357779464261925417033347961720796887378975386333422658415524949388265206384047792870784751951791444201183634282782950674174842;
            6'd22: xpb[159] = 1024'd53595539764417586016476703239477020182203470512981079558387591232881756674411227897006561434194594848790267856136988831747397581773956264593497728774374266425996876123196051830642322093141721740440818983322988542566091135011882457411842830700790097579349591186203456045879888508213623612798443950412327952534;
            6'd23: xpb[159] = 1024'd123704443763231880689297786516624757142139133968517865426386220869818324889053086752333262161925807874340634253665484742960859566858892640923289511909390028136464374803107445461651649020021184940266418541685255210699655741269275354366005815559860256160312701738731099337114353298911679059081294944499576214557;
            6'd24: xpb[159] = 1024'd69746652077921433963319942388958061357376370298318967166252995441777997766385806697644891674999346590447851243736487219595257711102608682697921170028074748913241198913447621755030736755383442418781820491660282032468859497305771478355190230735700965474455908877141684598242290015681101488245456111961229992249;
            6'd25: xpb[159] = 1024'd15788860392610987237342098261291365572613606628120068906119770013737670643718526642956521188072885306555068233807489696229655855346324724472552828146759469690018023023787798048409824490745699897297222441635308854238063253342267602344374645911541674788599116015552269859370226732450523917409617279422883769941;
            6'd26: xpb[159] = 1024'd85897764391425281910163181538439102532549270083656854774118399650674238858360385498283221915804098332105434631335985607443117840431261100802344611281775231400485521703699191679419151417625163097122821999997575522371627859599660499298537630770611833369562226568079913150604691523148579363692468273510132031964;
            6'd27: xpb[159] = 1024'd31939972706114835184185337410772406747786506413457956513985174222633911735693105443594851428877637048212651621406988084077515984674977142576976269400459952177262345814039367972798239152987420575638223949972602344140831615636156623287722045946452542683705433706490498411732628239918001792856629440971785809656;
            6'd28: xpb[159] = 1024'd102048876704929129857006420687920143707722169868994742381983803859570479950334964298921552156608850073763018018935483995290977969759913518906768052535475713887729844493950761603807566079866883775463823508334869012274396221893549520241885030805522701264668544259018141702967093030616057239139480435059034071679;
            6'd29: xpb[159] = 1024'd48091085019618683131028576560253447922959406198795844121850578431530152827667684244233181669682388789870235009006486471925376114003629560681399710654160434664506668604290937897186653815229141253979225458309895834043599977930045644231069445981363410578811751397428726964095029747385479668303641602520687849371;
            6'd30: xpb[159] = 1024'd118199989018432977803849659837401184882895069654332629989849208068466721042309543099559882397413601815420601406534982383138838099088565937011191493789176196374974167284202331528195980742108604453804825016672162502177164584187438541185232430840433569159774861949956370255329494538083535114586492596607936111394;
            6'd31: xpb[159] = 1024'd64242197333122531077871815709734489098132305984133731729715982640426393919642263044871511910487140531527818396605984859773236243332281978785823151907860917151750991394542507821575068477470861932320226966647189323946368340223934665174416846016274278473918069088366955516457431254852957543750653764069589889086;
            6'd32: xpb[159] = 1024'd10284405647812084351893971582067793313369542313934833469582757212386066796974982990183141423560679247635035386676987336407634387575998020560454810026545637928527815504882684114954156212833119410835628916622216145715572096260430789163601261192114987788061276226777540777585367971622379972914814931531243666778;
            6'd33: xpb[159] = 1024'd80393309646626379024715054859215530273305205769471619337581386849322635011616841845509842151291892273185401784205483247621096372660934396890246593161561399638995314184794077745963483139712582610661228474984482813849136702517823686117764246051185146369024386779305184068819832762320435419197665925618491928801;
            6'd34: xpb[159] = 1024'd26435517961315932298737210731548834488542442099272721077448161421282307888949561790821471664365430989292618774276485724255494516904650438664878251280246120415772138295134254039342570875074840089176630424959509635618340458554319810106948661227025855683167593917715769329947769479089857848361827093080145706493;
            6'd35: xpb[159] = 1024'd96544421960130226971558294008696571448478105554809506945446791058218876103591420646148172392096644014842985171804981635468956501989586814994670034415261882126239636975045647670351897801954303289002229983321776303751905064811712707061111646086096014264130704470243412621182234269787913294644678087167393968516;
            6'd36: xpb[159] = 1024'd42586630274819780245580449881029875663715341884610608685313565630178548980924140591459801905170182730950202161875984112103354646233302856769301692533946602903016461085385823963730985537316560767517631933296803125521108820848208831050296061261936723578273911608653997882310170986557335723808839254629047746208;
            6'd37: xpb[159] = 1024'd112695534273634074918401533158177612623651005340147394553312195267115117195565999446786502632901395756500568559404480023316816631318239233099093475668962364613483959765297217594740312464196023967343231491659069793654673427105601728004459046121006882159237022161181641173544635777255391170091690248716296008231;
            6'd38: xpb[159] = 1024'd58737742588323628192423689030510916838888241669948496293178969839074790072898719392098132145974934472607785549475482499951214775561955274873725133787647085390260783875637393888119400199558281445858633441634096615423877183142097851993643461296847591473380229299592226434672572494024813599255851416177949785923;
            6'd39: xpb[159] = 1024'd4779950903013181466445844902844221054125477999749598033045744411034462950231439337409761659048473188715002539546484976585612919805671316648356791906331806167037607985977570181498487934920538924374035391609123437193080939178593975982827876472688300787523436438002811695800509210794236028420012583639603563615;
            6'd40: xpb[159] = 1024'd74888854901827476139266928179991958014061141455286383901044374047971031164873298192736462386779686214265368937074980887799074904890607692978148575041347567877505106665888963812507814861800002124199634949971390105326645545435986872936990861331758459368486546990530454987034974001492291474702863577726851825638;
            6'd41: xpb[159] = 1024'd20931063216517029413289084052325262229298377785087485640911148619930704042206018138048091899853224930372585927145983364433473049134323734752780233160032288654281930776229140105886902597162259602715036899946416927095849301472482996926175276507599168682629754128941040248162910718261713903867024745188505603330;
            6'd42: xpb[159] = 1024'd91039967215331324086110167329472999189234041240624271508909778256867272256847876993374792627584437955922952324674479275646935034219260111082572016295048050364749429456140533736896229524041722802540636458308683595229413907729875893880338261366669327263592864681468683539397375508959769350149875739275753865353;
            6'd43: xpb[159] = 1024'd37082175530020877360132323201806303404471277570425373248776552828826945134180596938686422140657976672030169314745481752281333178462976152857203674413732771141526253566480710030275317259403980281056038408283710416998617663766372017869522676542510036577736071819879268800525312225729191779314036906737407643045;
            6'd44: xpb[159] = 1024'd107191079528835172032953406478954040364406941025962159116775182465763513348822455794013122868389189697580535712273977663494795163547912529186995457548748532851993752246392103661284644186283443480881637966645977085132182270023764914823685661401580195158699182372406912091759777016427247225596887900824655905068;
            6'd45: xpb[159] = 1024'd53233287843524725306975562351287344579644177355763260856641957037723186226155175739324752381462728413687752702344980140129193307791628570961627115667433253628770576356732279954663731921645700959397039916621003906901386026060261038812870076577420904472842389510817497352887713733196669654761049068286309682760;
            6'd46: xpb[159] = 1024'd123342191842339019979796645628435081539579840811300046724640586674659754440797034594651453109193941439238119099873476051342655292876564947291418898802449015339238075036643673585673058848525164159222639474983270575034950632317653935767033061436491063053805500063345140644122178523894725101043900062373557944783;
            6'd47: xpb[159] = 1024'd69384400157028573253818801500768385754817077141101148464507361246619427318129754539963082622267480155345336089944478527977053437120280989066050556921133736116014899146983849879052146583887421637738041424958297396804154388354150059756217476612331772367948707201755725905250115240664147530208061229835211722475;
            6'd48: xpb[159] = 1024'd15426608471718126527840957373101689970054313470902250204374135818579100195462474485274712135341018871452553080015481004611451581363997030840682215039818456892791723257324026172431234319249679116253443374933324218573358144390646183745401891788172481682091914340166311166378051957433569959372222397296865500167;
            6'd49: xpb[159] = 1024'd85535512470532421200662040650249426929989976926439036072372765455515668410104333340601412863072231897002919477543976915824913566448933407170473998174834218603259221937235419803440561246129142316079042933295590886706922750648039080699564876647242640263055024892693954457612516748131625405655073391384113762190;
            6'd50: xpb[159] = 1024'd31577720785221974474684196522582731145227213256240137812239540027475341287437053285913042376145770613110136467614979392459311710692649448945105656293518939380036046047575596096819648981491399794594444883270617708476126506684535204688749291823083349577198232031104539718740453464901047834819234558845767539882;
            6'd51: xpb[159] = 1024'd101686624784036269147505279799730468105162876711776923680238169664411909502078912141239743103876983638660502865143475303672773695777585825274897439428534701090503544727486989727828975908370862994420044441632884376609691112941928101642912276682153508158161342583632183009974918255599103281102085552933015801905;
            6'd52: xpb[159] = 1024'd47728833098725822421527435672063772320400113041578025420104944236371582379411632086551372616950522354767719855214477780307171840021301867049529097547219421867280368837827166021208063643733120472935446391607911198378894868978424225632096691857994217472304549722042768271102854972368525710266246720394669579597;
            6'd53: xpb[159] = 1024'd117837737097540117094348518949211509280335776497114811288103573873308150594053490941878073344681735380318086252742973691520633825106238243379320880682235183577747867517738559652217390570612583672761045949970177866512459475235817122586259676717064376053267660274570411562337319763066581156549097714481917841620;
            6'd54: xpb[159] = 1024'd63879945412229670368370674821544813495573012826915913027970348445267823471386210887189702857755274096425303242813976168155031969349954285153952538800919904354524691628078735945596478305974841151276447899945204688281663231272313246575444091892905085367410867412980996823465256479836003585713258881943571619312;
            6'd55: xpb[159] = 1024'd9922153726919223642392830693878117710810249156717014767837123017227496348718930832501332370828812812532520232884978644789430113593670326928584196919604625131301515738418912238975566041337098629791849849920231510050866987308809370564628507068745794681554074551391582084593193196605426014877420049405225397004;
            6'd56: xpb[159] = 1024'd80031057725733518315213913971025854670745912612253800635835752654164064563360789687828033098560025838082886630413474556002892098678606703258375980054620386841769014418330305869984892968216561829617449408282498178184431593566202267518791491927815953262517185103919225375827657987303481461160271043492473659027;
            6'd57: xpb[159] = 1024'd26073266040423071589236069843359158885983148942054902375702527226123737440693509633139662611633564554190103620484477032637290242922322745033007638173305107618545838528670482163363980703578819308132851358257524999953635349602698391507975907103656662576660392242329810636955594704072903890324432210954127436719;
            6'd58: xpb[159] = 1024'd96182170039237366262057153120506895845918812397591688243701156863060305655335368488466363339364777579740470018012972943850752228007259121362799421308320869329013337208581875794373307630458282507958450916619791668087199955860091288462138891962726821157623502794857453928190059494770959336607283205041375698742;
            6'd59: xpb[159] = 1024'd42224378353926919536079308992840200061156048727392789983567931435019978532668088433777992852438316295847687008083975420485150372250975163137431079427005590105790161318922052087752395365820539986473852866594818489856403711896587412451323307138567530471766709933268039189317996211540381765771444372503029476434;
            6'd60: xpb[159] = 1024'd112333282352741214208900392269987937021091712182929575851566561071956546747309947289104693580169529321398053405612471331698612357335911539467222862562021351816257659998833445718761722292700003186299452424957085157989968318153980309405486291997637689052729820485795682480552461002238437212054295366590277738457;
            6'd61: xpb[159] = 1024'd58375490667430767482922548142321241236328948512730677591433335643916219624642667234416323093243068037505270395683473808333010501579627581241854520680706072593034484109173622012140810028062260664814854374932111979759172074190476433394670707173478398366873027624206267741680397719007859641218456534051931516149;
            6'd62: xpb[159] = 1024'd4417698982120320756944704014654545451566184842531779331300110215875892501975387179727952606316606753612487385754476284967408645823343623016486178799390793369811308219513798305519897763424518143330256324907138801528375830226972557383855122349319107681016234762616853002808334435777282070382617701513585293841;
            6'd63: xpb[159] = 1024'd74526602980934615429765787291802282411501848298068565199298739852812460716617246035054653334047819779162853783282972196180870630908279999346277961934406555080278806899425191936529224690303981343155855883269405469661940436484365454338018107208389266261979345315144496294042799226475337516665468695600833555864;
        endcase
    end

    always_comb begin
        case(flag[53][11:6])
            6'd0: xpb[160] = 1024'd0;
            6'd1: xpb[160] = 1024'd20568811295624168703787943164135586626739084627869666939165514424772133593949965980366282847121358495270070773353974672815268775151996041120909620053091275857055631009765368229908312425666238821671257833244432291431144192520861578327202522384229975576122552453555081555170735943244759945829629863062487333556;
            6'd2: xpb[160] = 1024'd41137622591248337407575886328271173253478169255739333878331028849544267187899931960732565694242716990540141546707949345630537550303992082241819240106182551714111262019530736459816624851332477643342515666488864582862288385041723156654405044768459951152245104907110163110341471886489519891659259726124974667112;
            6'd3: xpb[160] = 1024'd61706433886872506111363829492406759880217253883609000817496543274316400781849897941098848541364075485810212320061924018445806325455988123362728860159273827571166893029296104689724937276998716465013773499733296874293432577562584734981607567152689926728367657360665244665512207829734279837488889589187462000668;
            6'd4: xpb[160] = 1024'd82275245182496674815151772656542346506956338511478667756662057699088534375799863921465131388485433981080283093415898691261075100607984164483638480212365103428222524039061472919633249702664955286685031332977729165724576770083446313308810089536919902304490209814220326220682943772979039783318519452249949334224;
            6'd5: xpb[160] = 1024'd102844056478120843518939715820677933133695423139348334695827572123860667969749829901831414235606792476350353866769873364076343875759980205604548100265456379285278155048826841149541562128331194108356289166222161457155720962604307891636012611921149877880612762267775407775853679716223799729148149315312436667780;
            6'd6: xpb[160] = 1024'd123412867773745012222727658984813519760434507767218001634993086548632801563699795882197697082728150971620424640123848036891612650911976246725457720318547655142333786058592209379449874553997432930027546999466593748586865155125169469963215134305379853456735314721330489331024415659468559674977779178374924001336;
            6'd7: xpb[160] = 1024'd19914983385244439527716674744134673642475165269351984446026745908428039820340622952548908715191835157447346006020329275127817585222751953291207215355307890065698742498786360271727947788146466030388607224323786193653648497425134275325439087006380379766037963760768512856088623528784686603688719214811816850561;
            6'd8: xpb[160] = 1024'd40483794680868608231504617908270260269214249897221651385192260333200173414290588932915191562313193652717416779374303947943086360374747994412116835408399165922754373508551728501636260213812704852059865057568218485084792689945995853652641609390610355342160516214323594411259359472029446549518349077874304184117;
            6'd9: xpb[160] = 1024'd61052605976492776935292561072405846895953334525091318324357774757972307008240554913281474409434552147987487552728278620758355135526744035533026455461490441779810004518317096731544572639478943673731122890812650776515936882466857431979844131774840330918283068667878675966430095415274206495347978940936791517673;
            6'd10: xpb[160] = 1024'd81621417272116945639080504236541433522692419152960985263523289182744440602190520893647757256555910643257558326082253293573623910678740076653936075514581717636865635528082464961452885065145182495402380724057083067947081074987719010307046654159070306494405621121433757521600831358518966441177608803999278851229;
            6'd11: xpb[160] = 1024'd102190228567741114342868447400677020149431503780830652202688803607516574196140486874014040103677269138527629099436227966388892685830736117774845695567672993493921266537847833191361197490811421317073638557301515359378225267508580588634249176543300282070528173574988839076771567301763726387007238667061766184785;
            6'd12: xpb[160] = 1024'd122759039863365283046656390564812606776170588408700319141854318032288707790090452854380322950798627633797699872790202639204161460982732158895755315620764269350976897547613201421269509916477660138744896390545947650809369460029442166961451698927530257646650726028543920631942303245008486332836868530124253518341;
            6'd13: xpb[160] = 1024'd19261155474864710351645406324133760658211245910834301952887977392083946046731279924731534583262311819624621238686683877440366395293507865461504810657524504274341853987807352313547583150626693239105956615403140095876152802329406972323675651628530783955953375067981944157006511114324613261547808566561146367566;
            6'd14: xpb[160] = 1024'd39829966770488879055433349488269347284950330538703968892053491816856079640681245905097817430383670314894692012040658550255635170445503906582414430710615780131397484997572720543455895576292932060777214448647572387307296994850268550650878174012760759532075927521537025712177247057569373207377438429623633701122;
            6'd15: xpb[160] = 1024'd60398778066113047759221292652404933911689415166573635831219006241628213234631211885464100277505028810164762785394633223070903945597499947703324050763707055988453116007338088773364208001959170882448472281892004678738441187371130128978080696396990735108198479975092107267347983000814133153207068292686121034678;
            6'd16: xpb[160] = 1024'd80967589361737216463009235816540520538428499794443302770384520666400346828581177865830383124626387305434833558748607895886172720749495988824233670816798331845508747017103457003272520427625409704119730115136436970169585379891991707305283218781220710684321032428647188822518718944058893099036698155748608368234;
            6'd17: xpb[160] = 1024'd101536400657361385166797178980676107165167584422312969709550035091172480422531143846196665971747745800704904332102582568701441495901492029945143290869889607702564378026868825233180832853291648525790987948380869261600729572412853285632485741165450686260443584882202270377689454887303653044866328018811095701790;
            6'd18: xpb[160] = 1024'd122105211952985553870585122144811693791906669050182636648715549515944614016481109826562948818869104295974975105456557241516710271053488071066052910922980883559620009036634193463089145278957887347462245781625301553031873764933714863959688263549680661836566137335757351932860190830548412990695957881873583035346;
            6'd19: xpb[160] = 1024'd18607327564484981175574137904132847673947326552316619459749208875739852273121936896914160451332788481801896471353038479752915205364263777631802405959741118482984965476828344355367218513106920447823306006482493998098657107233679669321912216250681188145868786375195375457924398699864539919406897918310475884571;
            6'd20: xpb[160] = 1024'd39176138860109149879362081068268434300686411180186286398914723300511985867071902877280443298454146977071967244707013152568183980516259818752712026012832394340040596486593712585275530938773159269494563839726926289529801299754541247649114738634911163721991338828750457013095134643109299865236527781372963218127;
            6'd21: xpb[160] = 1024'd59744950155733318583150024232404020927425495808055953338080237725284119461021868857646726145575505472342038018060987825383452755668255859873621646065923670197096227496359080815183843364439398091165821672971358580960945492275402825976317261019141139298113891282305538568265870586354059811066157644435450551683;
            6'd22: xpb[160] = 1024'd80313761451357487286937967396539607554164580435925620277245752150056253054971834838013008992696863967612108791414962498198721530820251900994531266119014946054151858506124449045092155790105636912837079506215790872392089684796264404303519783403371114874236443735860620123436606529598819756895787507497937885239;
            6'd23: xpb[160] = 1024'd100882572746981655990725910560675194180903665063795287216411266574828386648921800818379291839818222462882179564768937171013990305972247942115440886172106221911207489515889817275000468215771875734508337339460223163823233877317125982630722305787601090450358996189415701678607342472843579702725417370560425218795;
            6'd24: xpb[160] = 1024'd121451384042605824694513853724810780807642749691664954155576780999600520242871766798745574686939580958152250338122911843829259081124243983236350506225197497768263120525655185504908780641438114556179595172704655455254378069837987560957924828171831066026481548642970783233778078416088339648555047233622912552351;
            6'd25: xpb[160] = 1024'd17953499654105251999502869484131934689683407193798936966610440359395758499512593869096786319403265143979171704019393082065464015435019689802100001261957732691628076965849336397186853875587147656540655397561847900321161412137952366320148780872831592335784197682408806758842286285404466577265987270059805401576;
            6'd26: xpb[160] = 1024'd38522310949729420703290812648267521316422491821668603905775954784167892093462559849463069166524623639249242477373367754880732790587015730923009621315049008548683707975614704627095166301253386478211913230806280191752305604658813944647351303257061567911906750135963888314013022228649226523095617133122292735132;
            6'd27: xpb[160] = 1024'd59091122245353589407078755812403107943161576449538270844941469208940025687412525829829352013645982134519313250727342427696001565739011772043919241368140284405739338985380072857003478726919625299883171064050712483183449797179675522974553825641291543488029302589518969869183758171893986468925246996184780068688;
            6'd28: xpb[160] = 1024'd79659933540977758110866698976538694569900661077407937784106983633712159281362491810195634860767340629789384024081317100511270340891007813164828861421231560262794969995145441086911791152585864121554428897295144774614593989700537101301756348025521519064151855043074051424354494115138746414754876859247267402244;
            6'd29: xpb[160] = 1024'd100228744836601926814654642140674281196639745705277604723272498058484292875312457790561917707888699125059454797435291773326539116043003854285738481474322836119850601004910809316820103578252102943225686730539577066045738182221398679628958870409751494640274407496629132979525230058383506360584506722309754735800;
            6'd30: xpb[160] = 1024'd120797556132226095518442585304809867823378830333147271662438012483256426469262423770928200555010057620329525570789266446141807891194999895406648101527414111976906232014676177546728416003918341764896944563784009357476882374742260257956161392793981470216396959950184214534695966001628266306414136585372242069356;
            6'd31: xpb[160] = 1024'd17299671743725522823431601064131021705419487835281254473471671843051664725903250841279412187473741806156446936685747684378012825505775601972397596564174346900271188454870328439006489238067374865258004788641201802543665717042225063318385345494981996525699608989622238059760173870944393235125076621809134918581;
            6'd32: xpb[160] = 1024'd37868483039349691527219544228266608332158572463150921412637186267823798319853216821645695034595100301426517710039722357193281600657771643093307216617265622757326819464635696668914801663733613686929262621885634093974809909563086641645587867879211972101822161443177319614930909814189153180954706484871622252137;
            6'd33: xpb[160] = 1024'd58437294334973860231007487392402194958897657091020588351802700692595931913803182802011977881716458796696588483393697030008550375809767684214216836670356898614382450474401064898823114089399852508600520455130066385405954102083948219972790390263441947677944713896732401170101645757433913126784336347934109585693;
            6'd34: xpb[160] = 1024'd79006105630598028934795430556537781585636741718890255290968215117368065507753148782378260728837817291966659256747671702823819150961763725335126456723448174471438081484166433128731426515066091330271778288374498676837098294604809798299992912647671923254067266350287482725272381700678673072613966210996596919249;
            6'd35: xpb[160] = 1024'd99574916926222197638583373720673368212375826346759922230133729542140199101703114762744543575959175787236730030101646375639087926113759766456036076776539450328493712493931801358639738940732330151943036121618930968268242487125671376627195435031901898830189818803842564280443117643923433018443596074059084252805;
            6'd36: xpb[160] = 1024'd120143728221846366342371316884808954839114910974629589169299243966912332695653080743110826423080534282506800803455621048454356701265755807576945696829630726185549343503697169588548051366398568973614293954863363259699386679646532954954397957416131874406312371257397645835613853587168192964273225937121571586361;
            6'd37: xpb[160] = 1024'd16645843833345793647360332644130108721155568476763571980332903326707570952293907813462038055544218468333722169352102286690561635576531514142695191866390961108914299943891320480826124600547602073975354179720555704766170021946497760316621910117132400715615020296835669360678061456484319892984165973558464435586;
            6'd38: xpb[160] = 1024'd37214655128969962351148275808265695347894653104633238919498417751479704546243873793828320902665576963603792942706076959505830410728527555263604811919482236965969930953656688710734437026213840895646612012964987996197314214467359338643824432501362376291737572750390750915848797399729079838813795836620951769142;
            6'd39: xpb[160] = 1024'd57783466424594131054936218972401281974633737732502905858663932176251838140193839774194603749786935458873863716060051632321099185880523596384514431972573512823025561963422056940642749451880079717317869846209420287628458406988220916971026954885592351867860125203945832471019533342973839784643425699683439102698;
            6'd40: xpb[160] = 1024'd78352277720218299758724162136536868601372822360372572797829446601023971734143805754560886596908293954143934489414026305136367961032519637505424052025664788680081192973187425170551061877546318538989127679453852579059602599509082495298229477269822327443982677657500914026190269286218599730473055562745926436254;
            6'd41: xpb[160] = 1024'd98921089015842468462512105300672455228111906988242239736994961025796105328093771734927169444029652449414005262768000977951636736184515678626333672078756064537136823982952793400459374303212557360660385512698284870490746792029944073625431999654052303020105230111055995581361005229463359676302685425808413769810;
            6'd42: xpb[160] = 1024'd119489900311466637166300048464808041854850991616111906676160475450568238922043737715293452291151010944684076036121975650766905511336511719747243292131847340394192454992718161630367686728878796182331643345942717161921890984550805651952634522038282278596227782564611077136531741172708119622132315288870901103366;
            6'd43: xpb[160] = 1024'd15992015922966064471289064224129195736891649118245889487194134810363477178684564785644663923614695130510997402018456889003110445647287426312992787168607575317557411432912312522645759963027829282692703570799909606988674326850770457314858474739282804905530431604049100661595949042024246550843255325307793952591;
            6'd44: xpb[160] = 1024'd36560827218590233175077007388264782363630733746115556426359649235135610772634530766010946770736053625781068175372431561818379220799283467433902407221698851174613042442677680752554072388694068104363961404044341898419818519371632035642060997123512780481652984057604182216766684985269006496672885188370281286147;
            6'd45: xpb[160] = 1024'd57129638514214401878864950552400368990369818373985223365525163659907744366584496746377229617857412121051138948726406234633647995951279508554812027274790127031668673452443048982462384814360306926035219237288774189850962711892493613969263519507742756057775536511159263771937420928513766442502515051432768619703;
            6'd46: xpb[160] = 1024'd77698449809838570582652893716535955617108903001854890304690678084679877960534462726743512464978770616321209722080380907448916771103275549675721647327881402888724304462208417212370697240026545747706477070533206481282106904413355192296466041891972731633898088964714345327108156871758526388332144914495255953259;
            6'd47: xpb[160] = 1024'd98267261105462739286440836880671542243847987629724557243856192509452011554484428707109795312100129111591280495434355580264185546255271590796631267380972678745779935471973785442279009665692784569377734903777638772713251096934216770623668564276202707210020641418269426882278892815003286334161774777557743286815;
            6'd48: xpb[160] = 1024'd118836072401086907990228780044807128870587072257594224183021706934224145148434394687476078159221487606861351268788330253079454321407267631917540887434063954602835566481739153672187322091359023391048992737022071064144395289455078348950871086660432682786143193871824508437449628758248046279991404640620230620371;
            6'd49: xpb[160] = 1024'd15338188012586335295217795804128282752627729759728206994055366294019383405075221757827289791685171792688272634684811491315659255718043338483290382470824189526200522921933304564465395325508056491410052961879263509211178631755043154313095039361433209095445842911262531962513836627564173208702344677057123469596;
            6'd50: xpb[160] = 1024'd35906999308210503999005738968263869379366814387597873933220880718791516999025187738193572638806530287958343408038786164130928030870039379604200002523915465383256153931698672794373707751174295313081310795123695800642322824275904732640297561745663184671568395364817613517684572570808933154531974540119610803152;
            6'd51: xpb[160] = 1024'd56475810603834672702793682132399456006105899015467540872386395143563650592975153718559855485927888783228414181392760836946196806022035420725109622577006741240311784941464041024282020176840534134752568628368128092073467016796766310967500084129893160247690947818372695072855308514053693100361604403182098136708;
            6'd52: xpb[160] = 1024'd77044621899458841406581625296535042632844983643337207811551909568335784186925119698926138333049247278498484954746735509761465581174031461846019242630098017097367415951229409254190332602506772956423826461612560383504611209317627889294702606514123135823813500271927776628026044457298453046191234266244585470264;
            6'd53: xpb[160] = 1024'd97613433195083010110369568460670629259584068271206874750717423993107917780875085679292421180170605773768555728100710182576734356326027502966928862683189292954423046960994777484098645028173011778095084294856992674935755401838489467621905128898353111399936052725482858183196780400543212992020864129307072803820;
            6'd54: xpb[160] = 1024'd118182244490707178814157511624806215886323152899076541689882938417880051374825051659658704027291964269038626501454684855392003131478023544087838482736280568811478677970760145714006957453839250599766342128101424966366899594359351045949107651282583086976058605179037939738367516343787972937850493992369560137376;
            6'd55: xpb[160] = 1024'd14684360102206606119146527384127369768363810401210524500916597777675289631465878730009915659755648454865547867351166093628208065788799250653587977773040803734843634410954296606285030687988283700127402352958617411433682936659315851311331603983583613285361254218475963263431724213104099866561434028806452986601;
            6'd56: xpb[160] = 1024'd35253171397830774822934470548262956395102895029080191440082112202447423225415844710376198506877006950135618640705140766443476840940795291774497597826132079591899265420719664836193343113654522521798660186203049702864827129180177429638534126367813588861483806672031044818602460156348859812391063891868940320157;
            6'd57: xpb[160] = 1024'd55821982693454943526722413712398543021841979656949858379247626627219556819365810690742481353998365445405689414059115439258745616092791332895407217879223355448954896430485033066101655539320761343469918019447481994295971321701039007965736648752043564437606359125586126373773196099593619758220693754931427653713;
            6'd58: xpb[160] = 1024'd76390793989079112230510356876534129648581064284819525318413141051991690413315776671108764201119723940675760187413090112074014391244787374016316837932314631306010527440250401296009967964987000165141175852691914285727115514221900586292939171136273540013728911579141207928943932042838379704050323617993914987269;
            6'd59: xpb[160] = 1024'd96959605284703280934298300040669716275320148912689192257578655476763824007265742651475047048241082435945830960767064784889283166396783415137226457985405907163066158450015769525918280390653238986812433685936346577158259706742762164620141693520503515589851464032696289484114667986083139649879953481056402320825;
            6'd60: xpb[160] = 1024'd117528416580327449638086243204805302902059233540558859196744169901535957601215708631841329895362440931215901734121039457704551941548779456258136078038497183020121789459781137755826592816319477808483691519180778868589403899263623742947344215904733491165974016486251371039285403929327899595709583344118889654381;
            6'd61: xpb[160] = 1024'd14030532191826876943075258964126456784099891042692842007777829261331195857856535702192541527826125117042823100017520695940756875859555162823885573075257417943486745899975288648104666050468510908844751744037971313656187241563588548309568168605734017475276665525689394564349611798644026524420523380555782503606;
            6'd62: xpb[160] = 1024'd34599343487451045646863202128262043410838975670562508946943343686103329451806501682558824374947483612312893873371495368756025651011551203944795193128348693800542376909740656878012978476134749730516009577282403605087331434084450126636770690989963993051399217979244476119520347741888786470250153243618269837162;
            6'd63: xpb[160] = 1024'd55168154783075214350651145292397630037578060298432175886108858110875463045756467662925107222068842107582964646725470041571294426163547245065704813181439969657598007919506025107921290901800988552187267410526835896518475626605311704963973213374193968627521770432799557674691083685133546416079783106680757170718;
        endcase
    end

    always_comb begin
        case(flag[53][16:12])
            5'd0: xpb[161] = 1024'd0;
            5'd1: xpb[161] = 1024'd75736966078699383054439088456533216664317144926301842825274372535647596639706433643291390069190200602853035420079444714386563201315543286186614433234531245514653638929271393337829603327467227373858525243771268187949619819126173283291175735758423944203644322886354639229861819628378306361909412969743244504274;
            5'd2: xpb[161] = 1024'd27407236473274024710079249508252000583935862726868001522416890006318297942103728376567708923722726896262921432701395994194062561789866237818068741452731450095616603288971569338028967463417249026406852879155296529534878788031449793617372901833618439140468742358592220429617111182827979706700136112860894524217;
            5'd3: xpb[161] = 1024'd103144202551973407764518337964785217248253007653169844347691262541965894581810162019859098992912927499115956852780840708580625763105409524004683174687262695610270242218242962675858570790884476400265378122926564717484498607157623076908548637592042383344113065244946859659478930811206286068609549082604139028491;
            5'd4: xpb[161] = 1024'd54814472946548049420158499016504001167871725453736003044833780012636595884207456753135417847445453792525842865402791988388125123579732475636137482905462900191233206577943138676057934926834498052813705758310593059069757576062899587234745803667236878280937484717184440859234222365655959413400272225721789048434;
            5'd5: xpb[161] = 1024'd6484743341122691075798660068222785087490443254302161741976297483307297186604751486411736701977980085935728878024743268195624484054055427267591791123663104772196170937643314676257299062784519705362033393694621400655016544968176097560942969742431373217761904189422022058989513920105632758190995368839439068377;
            5'd6: xpb[161] = 1024'd82221709419822074130237748524756001751807588180604004567250670018954893826311185129703126771168180688788764298104187982582187685369598713454206224358194350286849809866914708014086902390251747079220558637465889588604636364094349380852118705500855317421406227075776661288851333548483939120100408338582683572651;
            5'd7: xpb[161] = 1024'd33891979814396715785877909576474785671426305981170163264393187489625595128708479862979445625700706982198650310726139262389687045843921665085660532576394554867812774226614884014286266526201768731768886272849917930189895332999625891178315871576049812358230646548014242488606625102933612464891131481700333592594;
            5'd8: xpb[161] = 1024'd109628945893096098840316998033008002335743450907472006089667560025273191768414913506270835694890907585051685730805583976776250247159464951272274965810925800382466413155886277352115869853668996105627411516621186118139515152125799174469491607334473756561874969434368881718468444731311918826800544451443578096868;
            5'd9: xpb[161] = 1024'd61299216287670740495957159084726786255362168708038164786810077495943893070812208239547154549423433878461571743427535256583749607633787902903729274029126004963429377515586453352315233989619017758175739152005214459724774121031075684795688773409668251498699388906606462918223736285761592171591267594561228116811;
            5'd10: xpb[161] = 1024'd12969486682245382151597320136445570174980886508604323483952594966614594373209502972823473403955960171871457756049486536391248968108110854535183582247326209544392341875286629352514598125569039410724066787389242801310033089936352195121885939484862746435523808378844044117979027840211265516381990737678878136754;
            5'd11: xpb[161] = 1024'd88706452760944765206036408592978786839298031434906166309226967502262191012915936616114863473146160774724493176128931250777812169423654140721798015481857455059045980804558022690344201453036266784582592031160510989259652909062525478413061675243286690639168131265198683347840847468589571878291403707422122641028;
            5'd12: xpb[161] = 1024'd40376723155519406861676569644697570758916749235472325006369484972932892315313231349391182327678687068134379188750882530585311529897977092353252323700057659640008945164258198690543565588986288437130919666544539330844911877967801988739258841318481185575992550737436264547596139023039245223082126850539772660971;
            5'd13: xpb[161] = 1024'd116113689234218789916115658101230787423233894161774167831643857508580488955019664992682572396868887670987414608830327244971874731213520378539866756934588905154662584093529592028373168916453515810989444910315807518794531697093975272030434577076905129779636873623790903777457958651417551584991539820283017165245;
            5'd14: xpb[161] = 1024'd67783959628793431571755819152949571342852611962340326528786374979251190257416959725958891251401413964397300621452278524779374091687843330171321065152789109735625548453229768028572533052403537463537772545699835860379790665999251782356631743152099624716461293096028484977213250205867224929782262963400667185188;
            5'd15: xpb[161] = 1024'd19454230023368073227395980204668355262471329762906485225928892449921891559814254459235210105933940257807186634074229804586873452162166281802775373370989314316588512812929944028771897188353559116086100181083864201965049634904528292682828909227294119653285712568266066176968541760316898274572986106518317205131;
            5'd16: xpb[161] = 1024'd95191196102067456281835068661201571926788474689208328051203264985569488199520688102526600175124140860660222054153674518973436653477709567989389806605520559831242151742201337366601500515820786489944625424855132389914669454030701575974004644985718063856930035454620705406830361388695204636482399076261561709405;
            5'd17: xpb[161] = 1024'd46861466496642097937475229712920355846407192489774486748345782456240189501917982835802919029656667154070108066775625798780936013952032519620844114823720764412205116101901513366800864651770808142492953060239160731499928422935978086300201811060912558793754454926858286606585652943144877981273122219379211729348;
            5'd18: xpb[161] = 1024'd122598432575341480991914318169453572510724337416076329573620154991887786141624416479094309098846867756923143486855070513167499215267575805807458548058252009926858755031172906704630467979238035516351478304010428919449548242062151369591377546819336502997398777813212925836447472571523184343182535189122456233622;
            5'd19: xpb[161] = 1024'd74268702969916122647554479221172356430343055216642488270762672462558487444021711212370627953379394050333029499477021792974998575741898757438912856276452214507821719390873082704829832115188057168899805939394457261034807210967427879917574712894530997934223197285450507036202764125972857687973258332240106253565;
            5'd20: xpb[161] = 1024'd25938973364490764303194640272891140349961773017208646967905189933229188746419005945646946807911920343742915512098973072782497936216221709070367164494652419088784683750573258705029196251138078821448133574778485602620066179872704390243771878969725492871047616757688088235958055680422531032763981475357756273508;
            5'd21: xpb[161] = 1024'd101675939443190147357633728729424357014278917943510489793179562468876785386125439588938336877102120946595950932178417787169061137531764995256981597729183664603438322679844652042858799578605306195306658818549753790569685998998877673534947614728149437074691939644042727465819875308800837394673394445101000777782;
            5'd22: xpb[161] = 1024'd53346209837764789013273889781143140933897635744076648490322079939547486688522734322214655731634647240005836944800369066976560498006087946888435905947383869184401287039544828043058163714555327847854986453933782132154944967904154183861144780803343932011516359116280308665575166863250510739464117588218650797725;
            5'd23: xpb[161] = 1024'd5016480232339430668914050832861924853516353544642807187464597410218187990920029055490974586167173533415722957422320346784059858480410898519890214165584073765364251399245004043257527850505349500403314089317810473740203936809430694187341946878538426948340778588517889865330458417700184084254840731336300817668;
            5'd24: xpb[161] = 1024'd80753446311038813723353139289395141517833498470944650012738969945865784630626462698782364655357374136268758377501765061170623059795954184706504647400115319280017890328516397381087131177972576874261839333089078661689823755935603977478517682636962371151985101474872529095192278046078490446164253701079545321942;
            5'd25: xpb[161] = 1024'd32423716705613455378993300341113925437452216271510808709881487416536485933023757432058683509889900429678644390123716340978122420270277136337958955618315523860980854688216573381286495313922598526810166968473107003275082724840880487804714848712156866088809520947110110294947569600528163790954976844197195341885;
            5'd26: xpb[161] = 1024'd108160682784312838433432388797647142101769361197812651535155859952184082572730191075350073579080101032531679810203161055364685621585820422524573388852846769375634493617487966719116098641389825900668692212244375191224702543967053771095890584470580810292453843833464749524809389228906470152864389813940439846159;
            5'd27: xpb[161] = 1024'd59830953178887480089072549849365926021388078998378810232298377422854783875127485808626392433612627325941565822825112335172184982060143374156027697071046973956597457977188142719315462777339847553217019847628403532809961512872330281422087750545775305229278263305702330724564680783356143497655112957058089866102;
            5'd28: xpb[161] = 1024'd11501223573462121744712710901084709941006796798944968929440894893525485177524780541902711288145153619351451835447063614979684342534466325787482005289247178537560422336888318719514826913289869205765347483012431874395220481777606791748284916620969800166102682777939911924319972337805816842445836100175739886045;
            5'd29: xpb[161] = 1024'd87238189652161504799151799357617926605323941725246811754715267429173081817231214185194101357335354222204487255526508329366247543850009611974096438523778424052214061266159712057344430240757096579623872726783700062344840300903780075039460652379393744369747005664294551154181791966184123204355249069918984390319;
            5'd30: xpb[161] = 1024'd38908460046736146454791960409336710524942659525812970451857784899843783119628508918470420211867880515614373268148459609173746904324332563605550746741978628633177025625859888057543794376707118232172200362167728403930099269809056585365657818454588239306571425136532132353937083520633796549145972213036634410262;
            5'd31: xpb[161] = 1024'd114645426125435529509231048865869927189259804452114813277132157435491379759334942561761810281058081118467408688227904323560310105639875849792165179976509874147830664555131281395373397704174345606030725605938996591879719088935229868656833554213012183510215748022886771583798903149012102911055385182779878914536;
        endcase
    end

    always_comb begin
        case(flag[54][5:0])
            6'd0: xpb[162] = 1024'd0;
            6'd1: xpb[162] = 1024'd95191196102067456281835068661201571926788474689208328051203264985569488199520688102526600175124140860660222054153674518973436653477709567989389806605520559831242151742201337366601500515820786489944625424855132389914669454030701575974004644985718063856930035454620705406830361388695204636482399076261561709405;
            6'd2: xpb[162] = 1024'd66315696520010171164871209917588711108878522252680971974274674906162081061732237295038129135590607411877294700849855603367809466114198801423619488194710078728793628914831457395572761840124367258579053241323024933464978057840506378983030720288206678447040167495124352783554194703461776255846108325897528934479;
            6'd3: xpb[162] = 1024'd37440196937952886047907351173975850290968569816153615897346084826754673923943786487549658096057073963094367347546036687762182278750688034857849169783899597626345106087461577424544023164427948027213481057790917477015286661650311181992056795590695293037150299535628000160278028018228347875209817575533496159553;
            6'd4: xpb[162] = 1024'd8564697355895600930943492430362989473058617379626259820417494747347266786155335680061187056523540514311439994242217772156555091387177268292078851373089116523896583260091697453515284488731528795847908874258810020565595265460115985001082870893183907627260431576131647537001861332994919494573526825169463384627;
            6'd5: xpb[162] = 1024'd103755893457963057212778561091564561399847092068834587871620759732916754985676023782587787231647681374971662048395892291129991744864886836281468657978609676355138735002293034820116785004552315285792534299113942410480264719490817560975087515878901971484190467030752352943832222721690124131055925901431025094032;
            6'd6: xpb[162] = 1024'd74880393875905772095814702347951700581937139632307231794692169653509347847887572975099316192114147926188734695092073375524364557501376069715698339567799195252690212174923154849088046328855896054426962115581834954030573323300622363984113591181390586074300599071256000320556056036456695750419635151066992319106;
            6'd7: xpb[162] = 1024'd46004894293848486978850843604338839764027187195779875717763579574101940710099122167610845152580614477405807341788254459918737370137865303149928021156988714150241689347553274878059307653159476823061389932049727497580881927110427166993139666483879200664410731111759647697279889351223267369783344400702959544180;
            6'd8: xpb[162] = 1024'd17129394711791201861886984860725978946117234759252519640834989494694533572310671360122374113047081028622879988484435544313110182774354536584157702746178233047793166520183394907030568977463057591695817748517620041131190530920231970002165741786367815254520863152263295074003722665989838989147053650338926769254;
            6'd9: xpb[162] = 1024'd112320590813858658143722053521927550872905709448460847692038254480264021771831359462648974288171221889283102042638110063286546836252064104573547509351698792879035318262384732273632069493283844081640443173372752431045859984950933545976170386772085879111450898606884000480834084054685043625629452726600488478659;
            6'd10: xpb[162] = 1024'd83445091231801373026758194778314690054995757011933491615109664400856614634042908655160503248637688440500174689334291147680919648888553338007777190940888311776586795435014852302603330817587424850274870989840644974596168588760738348985196462074574493701561030647387647857557917369451615244993161976236455703733;
            6'd11: xpb[162] = 1024'd54569591649744087909794336034701829237085804575406135538181074321449207496254457847672032209104154991717247336030472232075292461525042571442006872530077830674138272607644972331574592141891005618909298806308537518146477192570543151994222537377063108291671162687891295234281750684218186864356871225872422928807;
            6'd12: xpb[162] = 1024'd25694092067686802792830477291088968419175852138878779461252484242041800358466007040183561169570621542934319982726653316469665274161531804876236554119267349571689749780275092360545853466194586387543726622776430061696785796380347955003248612679551722881781294728394942611005583998984758483720580475508390153881;
            6'd13: xpb[162] = 1024'd120885288169754259074665545952290540345964326828087107512455749227611288557986695142710161344694762403594542036880327835443101927639241372865626360724787909402931901522476429727147353982015372877488352047631562451611455250411049530977253257665269786738711330183015648017835945387679963120202979551769951863286;
            6'd14: xpb[162] = 1024'd92009788587696973957701687208677679528054374391559751435527159148203881420198244335221690305161228954811614683576508919837474740275730606299856042313977428300483378695106549756118615306318953646122779864099454995161763854220854333986279332967758401328821462223519295394559778702446534739566688801405919088360;
            6'd15: xpb[162] = 1024'd63134289005639688840737828465064818710144421955032395358598569068796474282409793527733219265627695506028687330272690004231847552912219839734085723903166947198034855867736669785089876630622534414757207680567347538712072458030659136995305408270247015918931594264022942771283612017213106358930398051041886313434;
            6'd16: xpb[162] = 1024'd34258789423582403723773969721451957892234469518505039281669978989389067144621342720244748226094162057245759976968871088626220365548709073168315405492356466095586333040366789814061137954926115183391635497035240082262381061840463940004331483572735630509041726304526590148007445331979677978294107300677853538508;
            6'd17: xpb[162] = 1024'd5383289841525118606810110977839097074324517081977683204741388909981660006832891912756277186560628608462832623665052173020593178185198306602545087081545984993137810212996909843032399279229695952026063313503132625812689665650268743013357558875224245099151858345030237524731278646746249597657816550313820763582;
            6'd18: xpb[162] = 1024'd100574485943592574888645179639040669001112991771186011255944653895551148206353580015282877361684769469123054677818726691994029831662907874591934893687066544824379961955198247209633899795050482441970688738358265015727359119680970318987362203860942308956081893799650942931561640035441454234140215626575382472987;
            6'd19: xpb[162] = 1024'd71698986361535289771681320895427808183203039334658655179016063816143741068565129207794406322151236020340127324514907776388402644299397108026164575276256063721931439127828367238605161119354063210605116554826157559277667723490775121996388279163430923546192025840154590308285473350208025853503924876211349698061;
            6'd20: xpb[162] = 1024'd42823486779478004654717462151814947365293086898131299102087473736736333930776678400305935282617702571557199971211088860782775456935886341460394256865445582619482916300458487267576422443657643979239544371294050102827976327300579925005414354465919538136302157880658237685009306664974597472867634125847316923135;
            6'd21: xpb[162] = 1024'd13947987197420719537753603408202086547383134461603943025158883657328926792988227592817464243084169122774272617907269945177148269572375574894623938454635101517034393473088607296547683767961224747873972187761942646378284931110384728014440429768408152726412289921161885061733139979741169092231343375483284148209;
            6'd22: xpb[162] = 1024'd109139183299488175819588672069403658474171609150812271076362148642898414992508915695344064418208309983434494672060944464150584923050085142884013745060155661348276545215289944663149184283782011237818597612617075036292954385141086303988445074754126216583342325375782590468563501368436373728713742451744845857614;
            6'd23: xpb[162] = 1024'd80263683717430890702624813325790797656261656714284914999433558563491007854720464887855593378674776534651567318757125548544957735686574376318243426649345180245828022387920064692120445608085592006453025429084967579843262988950891106997471150056614831173452457416286237845287334683202945348077451701380813082688;
            6'd24: xpb[162] = 1024'd51388184135373605585660954582177936838351704277757558922504968484083600716932014080367122339141243085868639965453306632939330548323063609752473108238534699143379499560550184721091706932389172775087453245552860123393571592760695910006497225359103445763562589456789885222011167997969516967441160951016780307762;
            6'd25: xpb[162] = 1024'd22512684553316320468697095838565076020441751841230202845576378404676193579143563272878651299607709637085712612149487717333703360959552843186702789827724218040930976733180304750062968256692753543721881062020752666943880196570500713015523300661592060353672721497293532598735001312736088586804870200652747532836;
            6'd26: xpb[162] = 1024'd117703880655383776750532164499766647947230226530438530896779643390245681778664251375405251474731850497745934666303162236307140014437262411176092596433244777872173128475381642116664468772513540033666506486875885056858549650601202288989527945647310124210602756951914238005565362701431293223287269276914309242241;
            6'd27: xpb[162] = 1024'd88828381073326491633568305756153787129320274093911174819851053310838274640875800567916780435198317048963007312999343320701512827073751644610322278022434296769724605648011762145635730096817120802300934303343777600408858254411007091998554020949798738800712888992417885382289196016197864842650978526550276467315;
            6'd28: xpb[162] = 1024'd59952881491269206516604447012540926311410321657383818742922463231430867503087349760428309395664783600180079959695524405095885639710240878044551959611623815667276082820641882174606991421120701570935362119811670143959166858220811895007580096252287353390823021032921532759013029330964436462014687776186243692389;
            6'd29: xpb[162] = 1024'd31077381909211921399640588268928065493500369220856462665993873152023460365298898952939838356131250151397152606391705489490258452346730111478781641200813334564827559993272002203578252745424282339569789936279562687509475462030616698016606171554775967980933153073425180135736862645731008081378397025822210917463;
            6'd30: xpb[162] = 1024'd2201882327154636282676729525315204675590416784329106589065283072616053227510448145451367316597716702614225253087886573884631264983219344913011322790002853462379037165902122232549514069727863108204217752747455231059784065840421501025632246857264582571043285113928827512460695960497579700742106275458178142537;
            6'd31: xpb[162] = 1024'd97393078429222092564511798186516776602378891473537434640268548058185541427031136247977967491721857563274447307241561092858067918460928912902401129395523413293621188908103459599151014585548649598148843177602587620974453519871123076999636891842982646427973320568549532919291057349192784337224505351719739851942;
            6'd32: xpb[162] = 1024'd68517578847164807447547939442903915784468939037010078563339957978778134289242685440489496452188324114491519953937742177252440731097418146336630810984712932191172666080733579628122275909852230366783270994070480164524762123680927880008662967145471261018083452609053180296014890663959355956588214601355707077016;
            6'd33: xpb[162] = 1024'd39642079265107522330584080699291054966558986600482722486411367899370727151454234633001025412654790665708592600633923261646813543733907379770860492573902451088724143253363699657093537234155811135417698810538372708075070727490732683017689042447959875608193584649556827672738723978725927575951923850991674302090;
            6'd34: xpb[162] = 1024'd10766579683050237213620221955678194148649034163955366409482777819963320013665783825512554373121257216925665247330104346041186356370396613205090174163091969986275620425993819686064798558459391904052126627006265251625379331300537486026715117750448490198303716690060475049462557293492499195315633100627641527164;
            6'd35: xpb[162] = 1024'd105957775785117693495455290616879766075437508853163694460686042805532808213186471928039154548245398077585887301483778865014623009848106181194479980768612529817517772168195157052666299074280178393996752051861397641540048785331239062000719762736166554055233752144681180456292918682187703831798032176889203236569;
            6'd36: xpb[162] = 1024'd77082276203060408378491431873266905257527556416636338383757452726125401075398021120550683508711864628802959948179959949408995822484595414628709662357802048715069249340825277081637560398583759162631179868329290185090357389141043865009745838038655168645343884185184827833016751996954275451161741426525170461643;
            6'd37: xpb[162] = 1024'd48206776621003123261527573129654044439617603980108982306828862646717993937609570313062212469178331180020032594876141033803368635121084648062939343946991567612620726513455397110608821722887339931265607684797182728640665992950848668018771913341143783235454016225688475209740585311720847070525450676161137686717;
            6'd38: xpb[162] = 1024'd19331277038945838144563714386041183621707651543581626229900272567310586799821119505573741429644797731237105241572322118197741447757573881497169025536181086510172203686085517139580083047190920699900035501265075272190974596760653471027797988643632397825564148266192122586464418626487418689889159925797104911791;
            6'd39: xpb[162] = 1024'd114522473141013294426398783047242755548496126232789954281103537552880074999341807608100341604768938591897327295725996637171178101235283449486558832141701646341414355428286854506181583563011707189844660926120207662105644050791355047001802633629350461682494183720812827993294780015182623326371559002058666621196;
            6'd40: xpb[162] = 1024'd85646973558956009309434924303629894730586173796262598204174947473472667861553356800611870565235405143114399942422177721565550913871772682920788513730891165238965832600916974535152844887315287958479088742588100205655952654601159850010828708931839076272604315761316475370018613329949194945735268251694633846270;
            6'd41: xpb[162] = 1024'd56771473976898724192471065560017033912676221359735242127246357394065260723764905993123399525701871694331472589118358805959923726508261916355018195320080684136517309773547094564124106211618868727113516559055992749206261258410964653019854784234327690862714447801820122746742446644715766565098977501330601071344;
            6'd42: xpb[162] = 1024'd27895974394841439075507206816404173094766268923207886050317767314657853585976455185634928486168338245548545235814539890354296539144751149789247876909270203034068786946177214593095367535922449495747944375523885292756569862220769456028880859536816305452824579842323770123466279959482338184462686750966568296418;
            6'd43: xpb[162] = 1024'd123087170496908895357342275477605745021554743612416214101521032300227341785497143288161528661292479106208767289968214409327733192622460717778637683514790762865310938688378551959696868051743235985692569800379017682671239316251471032002885504522534369309754615296944475530296641348177542820945085827228130005823;
            6'd44: xpb[162] = 1024'd94211670914851610240378416733992884203644791175888858024592442220819934647708692480673057621758945657425839936664395493722106005258949951212867365103980281762862415861008671988668129376046816754326997616846910226221547920061275835011911579825022983899864747337448122907020474662944114440308795076864097230897;
            6'd45: xpb[162] = 1024'd65336171332794325123414557990380023385734838739361501947663852141412527509920241673184586582225412208642912583360576578116478817895439184647097046693169800660413893033638792017639390700350397522961425433314802769771856523871080638020937655127511598489974879377951770283744307977710686059672504326500064455971;
            6'd46: xpb[162] = 1024'd36460671750737040006450699246767162567824886302834145870735262062005120372131790865696115542691878759859985230056757662510851630531928418081326728282359319557965370206268912046610652024653978291595853249782695313322165127680885441029963730430000213080085011418455417660468141292477257679036213576136031681045;
            6'd47: xpb[162] = 1024'd7585172168679754889486840503154301749914933866306789793806671982597713234343340058207644503158345311077057876752938746905224443168417651515556409871548838455516847378899032075581913348957559060230281066250587856872473731490690244038989805732488827670195143458959065037191974607243829298399922825771998906119;
            6'd48: xpb[162] = 1024'd102776368270747211171321909164355873676703408555515117845009936968167201433864028160734244678282486171737279930906613265878661096646127219504946216477069398286758999121100369442183413864778345550174906491105720246787143185521391820012994450718206891527125178913579770444022335995939033934882321902033560615524;
            6'd49: xpb[162] = 1024'd73900868688689926054358050420743012858793456118987761768081346888759794296075577353245773638748952722954352577602794350273033909282616452939175898066258917184310476293730489471154675189081926318809334307573612790337451789331196623022020526020695506117235310954083417820746169310705605554246031151669527840598;
            6'd50: xpb[162] = 1024'd45025369106632640937394191677130152040883503682460405691152756809352387158287126545757302599215419274171425224298975434667406721919105686373405579655448436081861953466360609500125936513385507087443762124041505333887760393141001426031046601323184120707345442994587065197470002625472177173609740401305495065672;
            6'd51: xpb[162] = 1024'd16149869524575355820430332933517291222973551245933049614224166729944980020498675738268831559681885825388497870995156519061779534555594919807635261244637954979413430638990729529097197837689087856078189940509397877438068996950806229040072676625672735297455575035090712574193835940238748792973449650941462290746;
            6'd52: xpb[162] = 1024'd111341065626642812102265401594718863149762025935141377665427431715514468220019363840795431734806026686048719925148831038035216188033304487797025067850158514810655582381192066895698698353509874346022815365364530267352738450981507805014077321611390799154385610489711417981024197328933953429455848727203024000151;
            6'd53: xpb[162] = 1024'd82465566044585526985301542851106002331852073498614021588498841636107061082230913033306960695272493237265792571845012122429589000669793721231254749439348033708207059553822186924669959677813455114657243181832422810903047054791312608023103396913879413744495742530215065357748030643700525048819557976838991225225;
            6'd54: xpb[162] = 1024'd53590066462528241868337684107493141513942121062086665511570251556699653944442462225818489655738959788482865218541193206823961813306282954665484431028537552605758536726452306953641221002117035883291670998300315354453355658601117411032129472216368028334605874570718712734471863958467096668183267226474958450299;
            6'd55: xpb[162] = 1024'd24714566880470956751373825363880280696032168625559309434641661477292246806654011418330018616205426339699937865237374291218334625942772188099714112617727071503310013899082426982612482326420616651926098814768207898003664262410922214041155547518856642924716006611222360111195697273233668287546976476110925675373;
            6'd56: xpb[162] = 1024'd119905762982538413033208894025081852622820643314767637485844926462861735006174699520856618791329567200360159919391048810191771279420481756089103919223247631334552165641283764349213982842241403141870724239623340287918333716441623790015160192504574706781646042065843065518026058661928872924029375552372487384778;
            6'd57: xpb[162] = 1024'd91030263400481127916245035281468991804910690878240281408916336383454327868386248713368147751796033751577232566087229894586144092056970989523333600812437150232103642813913884378185244166544983910505152056091232831468642320251428593024186267807063321371756174106346712894749891976695444543393084802008454609852;
            6'd58: xpb[162] = 1024'd62154763818423842799281176537856130987000738441712925331987746304046920730597797905879676712262500302794305212783410978980516904693460222957563282401626669129655119986544004407156505490848564679139579872559125375018950924061233396033212343109551935961866306146850360271473725291462016162756794051644421834926;
            6'd59: xpb[162] = 1024'd33279264236366557682317317794243270169090786005185569255059156224639513592809347098391205672728966854011377859479592063374889717329949456391792963990816188027206597159174124436127766815152145447774007689027017918569259527871038199042238418412040550551976438187354007648197558606228587782120503301280389060000;
            6'd60: xpb[162] = 1024'd4403764654309272565353459050630409351180833568658213178130566145232106455020896290902734633195433405228450506175773147769262529966438689826022645580005706924758074331804244465099028139455726216408435505494910462119568131680843002051264493714529165142086570227857655024921391920995159401484212550916356285074;
            6'd61: xpb[162] = 1024'd99594960756376728847188527711831981277969308257866541229333831130801594654541584393429334808319574265888672560329447666742699183444148257815412452185526266756000226074005581831700528655276512706353060930350042852034237585711544578025269138700247228999016605682478360431751753309690364037966611627177917994479;
            6'd62: xpb[162] = 1024'd70719461174319443730224668968219120460059355821339185152405241051394187516753133585940863768786040817105745207025628751137071996080637491249642133774715785653551703246635701860671789979580093474987488746817935395584546189521349381034295214002735843589126737722982007808475586624456935657330320876813885219553;
            6'd63: xpb[162] = 1024'd41843961592262158613260810224606259642149403384811829075476650971986780378964682778452392729252507368322817853721809835531444808717126724683871815363905304551103180419265821889643051303883674243621916563285827939134854793331154184043321289305224458179236869763485655185199419939223507276694030126449852444627;
        endcase
    end

    always_comb begin
        case(flag[54][11:6])
            6'd0: xpb[163] = 1024'd0;
            6'd1: xpb[163] = 1024'd12968462010204873496296951480993398824239450948284472998548060892579373241176231970963921689718973919539890500417990919925817621353615958118101496953094823448654657591895941918614312628187255012256344379753720482685163397140958987052347364607713072769347001803989302561923253253990078896057739376085819669701;
            6'd2: xpb[163] = 1024'd25936924020409746992593902961986797648478901896568945997096121785158746482352463941927843379437947839079781000835981839851635242707231916236202993906189646897309315183791883837228625256374510024512688759507440965370326794281917974104694729215426145538694003607978605123846506507980157792115478752171639339402;
            6'd3: xpb[163] = 1024'd38905386030614620488890854442980196472718352844853418995644182677738119723528695912891765069156921758619671501253972759777452864060847874354304490859284470345963972775687825755842937884561765036769033139261161448055490191422876961157042093823139218308041005411967907685769759761970236688173218128257459009103;
            6'd4: xpb[163] = 1024'd51873848040819493985187805923973595296957803793137891994192243570317492964704927883855686758875895678159562001671963679703270485414463832472405987812379293794618630367583767674457250512749020049025377519014881930740653588563835948209389458430852291077388007215957210247693013015960315584230957504343278678804;
            6'd5: xpb[163] = 1024'd64842310051024367481484757404966994121197254741422364992740304462896866205881159854819608448594869597699452502089954599629088106768079790590507484765474117243273287959479709593071563140936275061281721898768602413425816985704794935261736823038565363846735009019946512809616266269950394480288696880429098348505;
            6'd6: xpb[163] = 1024'd77810772061229240977781708885960392945436705689706837991288365355476239447057391825783530138313843517239343002507945519554905728121695748708608981718568940691927945551375651511685875769123530073538066278522322896110980382845753922314084187646278436616082010823935815371539519523940473376346436256514918018206;
            6'd7: xpb[163] = 1024'd90779234071434114474078660366953791769676156637991310989836426248055612688233623796747451828032817436779233502925936439480723349475311706826710478671663764140582603143271593430300188397310785085794410658276043378796143779986712909366431552253991509385429012627925117933462772777930552272404175632600737687907;
            6'd8: xpb[163] = 1024'd103747696081638987970375611847947190593915607586275783988384487140634985929409855767711373517751791356319124003343927359406540970828927664944811975624758587589237260735167535348914501025498040098050755038029763861481307177127671896418778916861704582154776014431914420495386026031920631168461915008686557357608;
            6'd9: xpb[163] = 1024'd116716158091843861466672563328940589418155058534560256986932548033214359170586087738675295207470765275859014503761918279332358592182543623062913472577853411037891918327063477267528813653685295110307099417783484344166470574268630883471126281469417654924123016235903723057309279285910710064519654384772377027309;
            6'd10: xpb[163] = 1024'd5617924417923993564170587405119555497696082357109045857348753860816837074453180799624145682532064885955755596722415764679112372694939246625854844514617193552855901349388201848512887090355344401253246189149964980487273121188693097558495076393901278426650114625775967589126004465972155943458703934232602212679;
            6'd11: xpb[163] = 1024'd18586386428128867060467538886112954321935533305393518855896814753396210315629412770588067372251038805495646097140406684604929994048555204743956341467712017001510558941284143767127199718542599413509590568903685463172436518329652084610842441001614351195997116429765270151049257719962234839516443310318421882380;
            6'd12: xpb[163] = 1024'd31554848438333740556764490367106353146174984253677991854444875645975583556805644741551989061970012725035536597558397604530747615402171162862057838420806840450165216533180085685741512346729854425765934948657405945857599915470611071663189805609327423965344118233754572712972510973952313735574182686404241552081;
            6'd13: xpb[163] = 1024'd44523310448538614053061441848099751970414435201962464852992936538554956797981876712515910751688986644575427097976388524456565236755787120980159335373901663898819874125076027604355824974917109438022279328411126428542763312611570058715537170217040496734691120037743875274895764227942392631631922062490061221782;
            6'd14: xpb[163] = 1024'd57491772458743487549358393329093150794653886150246937851540997431134330039158108683479832441407960564115317598394379444382382858109403079098260832326996487347474531716971969522970137603104364450278623708164846911227926709752529045767884534824753569504038121841733177836819017481932471527689661438575880891483;
            6'd15: xpb[163] = 1024'd70460234468948361045655344810086549618893337098531410850089058323713703280334340654443754131126934483655208098812370364308200479463019037216362329280091310796129189308867911441584450231291619462534968087918567393913090106893488032820231899432466642273385123645722480398742270735922550423747400814661700561184;
            6'd16: xpb[163] = 1024'd83428696479153234541952296291079948443132788046815883848637119216293076521510572625407675820845908403195098599230361284234018100816634995334463826233186134244783846900763853360198762859478874474791312467672287876598253504034447019872579264040179715042732125449711782960665523989912629319805140190747520230885;
            6'd17: xpb[163] = 1024'd96397158489358108038249247772073347267372238995100356847185180108872449762686804596371597510564882322734989099648352204159835722170250953452565323186280957693438504492659795278813075487666129487047656847426008359283416901175406006924926628647892787812079127253701085522588777243902708215862879566833339900586;
            6'd18: xpb[163] = 1024'd109365620499562981534546199253066746091611689943384829845733241001451823003863036567335519200283856242274879600066343124085653343523866911570666820139375781142093162084555737197427388115853384499304001227179728841968580298316364993977273993255605860581426129057690388084512030497892787111920618942919159570287;
            6'd19: xpb[163] = 1024'd122334082509767855030843150734060144915851140891669302844281301894031196245039268538299440890002830161814770100484334044011470964877482869688768317092470604590747819676451679116041700744040639511560345606933449324653743695457323981029621357863318933350773130861679690646435283751882866007978358319004979239988;
            6'd20: xpb[163] = 1024'd11235848835847987128341174810239110995392164714218091714697507721633674148906361599248291365064129771911511193444831529358224745389878493251709689029234387105711802698776403697025774180710688802506492378299929960974546242377386195116990152787802556853300229251551935178252008931944311886917407868465204425358;
            6'd21: xpb[163] = 1024'd24204310846052860624638126291232509819631615662502564713245568614213047390082593570212213054783103691451401693862822449284042366743494451369811185982329210554366460290672345615640086808897943814762836758053650443659709639518345182169337517395515629622647231055541237740175262185934390782975147244551024095059;
            6'd22: xpb[163] = 1024'd37172772856257734120935077772225908643871066610787037711793629506792420631258825541176134744502077610991292194280813369209859988097110409487912682935424034003021117882568287534254399437085198827019181137807370926344873036659304169221684882003228702391994232859530540302098515439924469679032886620636843764760;
            6'd23: xpb[163] = 1024'd50141234866462607617232029253219307468110517559071510710341690399371793872435057512140056434221051530531182694698804289135677609450726367606014179888518857451675775474464229452868712065272453839275525517561091409030036433800263156274032246610941775161341234663519842864021768693914548575090625996722663434461;
            6'd24: xpb[163] = 1024'd63109696876667481113528980734212706292349968507355983708889751291951167113611289483103978123940025450071073195116795209061495230804342325724115676841613680900330433066360171371483024693459708851531869897314811891715199830941222143326379611218654847930688236467509145425945021947904627471148365372808483104162;
            6'd25: xpb[163] = 1024'd76078158886872354609825932215206105116589419455640456707437812184530540354787521454067899813658999369610963695534786128987312852157958283842217173794708504348985090658256113290097337321646963863788214277068532374400363228082181130378726975826367920700035238271498447987868275201894706367206104748894302773863;
            6'd26: xpb[163] = 1024'd89046620897077228106122883696199503940828870403924929705985873077109913595963753425031821503377973289150854195952777048913130473511574241960318670747803327797639748250152055208711649949834218876044558656822252857085526625223140117431074340434080993469382240075487750549791528455884785263263844124980122443564;
            6'd27: xpb[163] = 1024'd102015082907282101602419835177192902765068321352209402704533933969689286837139985395995743193096947208690744696370767968838948094865190200078420167700898151246294405842047997127325962578021473888300903036575973339770690022364099104483421705041794066238729241879477053111714781709874864159321583501065942113265;
            6'd28: xpb[163] = 1024'd114983544917486975098716786658186301589307772300493875703081994862268660078316217366959664882815921128230635196788758888764765716218806158196521664653992974694949063433943939045940275206208728900557247416329693822455853419505058091535769069649507139008076243683466355673638034963864943055379322877151761782966;
            6'd29: xpb[163] = 1024'd3885311243567107196214810734365267668848796123042664573498200689871137982183310427908515357877220738327376289749256374111519496731201781759463036590756757209913046456268663626924348642878778191503394187696174458776655966425120305623137864573990762510603342073338600205454760143926388934318372426611986968336;
            6'd30: xpb[163] = 1024'd16853773253771980692511762215358666493088247071327137572046261582450511223359542398872437047596194657867266790167247294037337118084817739877564533543851580658567704048164605545538661271066033203759738567449894941461819363566079292675485229181703835279950343877327902767378013397916467830376111802697806638037;
            6'd31: xpb[163] = 1024'd29822235263976854188808713696352065317327698019611610570594322475029884464535774369836358737315168577407157290585238213963154739438433697995666030496946404107222361640060547464152973899253288216016082947203615424146982760707038279727832593789416908049297345681317205329301266651906546726433851178783626307738;
            6'd32: xpb[163] = 1024'd42790697274181727685105665177345464141567148967896083569142383367609257705712006340800280427034142496947047791003229133888972360792049656113767527450041227555877019231956489382767286527440543228272427326957335906832146157847997266780179958397129980818644347485306507891224519905896625622491590554869445977439;
            6'd33: xpb[163] = 1024'd55759159284386601181402616658338862965806599916180556567690444260188630946888238311764202116753116416486938291421220053814789982145665614231869024403136051004531676823852431301381599155627798240528771706711056389517309554988956253832527323004843053587991349289295810453147773159886704518549329930955265647140;
            6'd34: xpb[163] = 1024'd68727621294591474677699568139332261790046050864465029566238505152768004188064470282728123806472090336026828791839210973740607603499281572349970521356230874453186334415748373219995911783815053252785116086464776872202472952129915240884874687612556126357338351093285113015071026413876783414607069307041085316841;
            6'd35: xpb[163] = 1024'd81696083304796348173996519620325660614285501812749502564786566045347377429240702253692045496191064255566719292257201893666425224852897530468072018309325697901840992007644315138610224412002308265041460466218497354887636349270874227937222052220269199126685352897274415576994279667866862310664808683126904986542;
            6'd36: xpb[163] = 1024'd94664545315001221670293471101319059438524952761033975563334626937926750670416934224655967185910038175106609792675192813592242846206513488586173515262420521350495649599540257057224537040189563277297804845972217837572799746411833214989569416827982271896032354701263718138917532921856941206722548059212724656243;
            6'd37: xpb[163] = 1024'd107633007325206095166590422582312458262764403709318448561882687830506123911593166195619888875629012094646500293093183733518060467560129446704275012215515344799150307191436198975838849668376818289554149225725938320257963143552792202041916781435695344665379356505253020700840786175847020102780287435298544325944;
            6'd38: xpb[163] = 1024'd120601469335410968662887374063305857087003854657602921560430748723085497152769398166583810565347986014186390793511174653443878088913745404822376509168610168247804964783332140894453162296564073301810493605479658802943126540693751189094264146043408417434726358309242323262764039429837098998838026811384363995645;
            6'd39: xpb[163] = 1024'd9503235661491100760385398139484823166544878480151710430846954550687975056636491227532661040409285624283131886471672138790631869426141028385317881105373950762768947805656865475437235733234122592756640376846139439263929087613813403181632940967892040937253456699114567794580764609898544877777076360844589181015;
            6'd40: xpb[163] = 1024'd22471697671695974256682349620478221990784329428436183429395015443267348297812723198496582730128259543823022386889663058716449490779756986503419378058468774211423605397552807394051548361421377605012984756599859921949092484754772390233980305575605113706600458503103870356504017863888623773834815736930408850716;
            6'd41: xpb[163] = 1024'd35440159681900847752979301101471620815023780376720656427943076335846721538988955169460504419847233463362912887307653978642267112133372944621520875011563597660078262989448749312665860989608632617269329136353580404634255881895731377286327670183318186475947460307093172918427271117878702669892555113016228520417;
            6'd42: xpb[163] = 1024'd48408621692105721249276252582465019639263231325005129426491137228426094780165187140424426109566207382902803387725644898568084733486988902739622371964658421108732920581344691231280173617795887629525673516107300887319419279036690364338675034791031259245294462111082475480350524371868781565950294489102048190118;
            6'd43: xpb[163] = 1024'd61377083702310594745573204063458418463502682273289602425039198121005468021341419111388347799285181302442693888143635818493902354840604860857723868917753244557387578173240633149894486245983142641782017895861021370004582676177649351391022399398744332014641463915071778042273777625858860462008033865187867859819;
            6'd44: xpb[163] = 1024'd74345545712515468241870155544451817287742133221574075423587259013584841262517651082352269489004155221982584388561626738419719976194220818975825365870848068006042235765136575068508798874170397654038362275614741852689746073318608338443369764006457404783988465719061080604197030879848939358065773241273687529520;
            6'd45: xpb[163] = 1024'd87314007722720341738167107025445216111981584169858548422135319906164214503693883053316191178723129141522474888979617658345537597547836777093926862823942891454696893357032516987123111502357652666294706655368462335374909470459567325495717128614170477553335467523050383166120284133839018254123512617359507199221;
            6'd46: xpb[163] = 1024'd100282469732925215234464058506438614936221035118143021420683380798743587744870115024280112868442103061062365389397608578271355218901452735212028359777037714903351550948928458905737424130544907678551051035122182818060072867600526312548064493221883550322682469327039685728043537387829097150181251993445326868922;
            6'd47: xpb[163] = 1024'd113250931743130088730761009987432013760460486066427494419231441691322960986046346995244034558161076980602255889815599498197172840255068693330129856730132538352006208540824400824351736758732162690807395414875903300745236264741485299600411857829596623092029471131028988289966790641819176046238991369531146538623;
            6'd48: xpb[163] = 1024'd2152698069210220828259034063610979840001509888976283289647647518925438889913440056192885033222376590698996982776096983543926620767464316893071228666896320866970191563149125405335810195402211981753542186242383937066038811661547513687780652754080246594556569520901232821783515821880621925178040918991371723993;
            6'd49: xpb[163] = 1024'd15121160079415094324555985544604378664240960837260756288195708411504812131089672027156806722941350510238887483194087903469744242121080275011172725619991144315624849155045067323950122823589466994009886565996104419751202208802506500740128017361793319363903571324890535383706769075870700821235780295077191393694;
            6'd50: xpb[163] = 1024'd28089622089619967820852937025597777488480411785545229286743769304084185372265903998120728412660324429778777983612078823395561863474696233129274222573085967764279506746941009242564435451776722006266230945749824902436365605943465487792475381969506392133250573128879837945630022329860779717293519671163011063395;
            6'd51: xpb[163] = 1024'd41058084099824841317149888506591176312719862733829702285291830196663558613442135969084650102379298349318668484030069743321379484828312191247375719526180791212934164338836951161178748079963977018522575325503545385121529003084424474844822746577219464902597574932869140507553275583850858613351259047248830733096;
            6'd52: xpb[163] = 1024'd54026546110029714813446839987584575136959313682114175283839891089242931854618367940048571792098272268858558984448060663247197106181928149365477216479275614661588821930732893079793060708151232030778919705257265867806692400225383461897170111184932537671944576736858443069476528837840937509408998423334650402797;
            6'd53: xpb[163] = 1024'd66995008120234588309743791468577973961198764630398648282387951981822305095794599911012493481817246188398449484866051583173014727535544107483578713432370438110243479522628834998407373336338487043035264085010986350491855797366342448949517475792645610441291578540847745631399782091831016405466737799420470072498;
            6'd54: xpb[163] = 1024'd79963470130439461806040742949571372785438215578683121280936012874401678336970831881976415171536220107938339985284042503098832348889160065601680210385465261558898137114524776917021685964525742055291608464764706833177019194507301436001864840400358683210638580344837048193323035345821095301524477175506289742199;
            6'd55: xpb[163] = 1024'd92931932140644335302337694430564771609677666526967594279484073766981051578147063852940336861255194027478230485702033423024649970242776023719781707338560085007552794706420718835635998592712997067547952844518427315862182591648260423054212205008071755979985582148826350755246288599811174197582216551592109411900;
            6'd56: xpb[163] = 1024'd105900394150849208798634645911558170433917117475252067278032134659560424819323295823904258550974167947018120986120024342950467591596391981837883204291654908456207452298316660754250311220900252079804297224272147798547345988789219410106559569615784828749332583952815653317169541853801253093639955927677929081601;
            6'd57: xpb[163] = 1024'd118868856161054082294931597392551569258156568423536540276580195552139798060499527794868180240693141866558011486538015262876285212950007939955984701244749731904862109890212602672864623849087507092060641604025868281232509385930178397158906934223497901518679585756804955879092795107791331989697695303763748751302;
            6'd58: xpb[163] = 1024'd7770622487134214392429621468730535337697592246085329146996401379742275964366620855817030715754441476654752579498512748223038993462403563518926073181513514419826092912537327253848697285757556383006788375392348917553311932850240611246275729147981525021206684146677200410909520287852777868636744853223973936672;
            6'd59: xpb[163] = 1024'd20739084497339087888726572949723934161937043194369802145544462272321649205542852826780952405473415396194643079916503668148856614816019521637027570134608337868480750504433269172463009913944811395263132755146069400238475329991199598298623093755694597790553685950666502972832773541842856764694484229309793606373;
            6'd60: xpb[163] = 1024'd33707546507543961385023524430717332986176494142654275144092523164901022446719084797744874095192389315734533580334494588074674236169635479755129067087703161317135408096329211091077322542132066407519477134899789882923638727132158585350970458363407670559900687754655805534756026795832935660752223605395613276074;
            6'd61: xpb[163] = 1024'd46676008517748834881320475911710731810415945090938748142640584057480395687895316768708795784911363235274424080752485508000491857523251437873230564040797984765790065688225153009691635170319321419775821514653510365608802124273117572403317822971120743329247689558645108096679280049823014556809962981481432945775;
            6'd62: xpb[163] = 1024'd59644470527953708377617427392704130634655396039223221141188644950059768929071548739672717474630337154814314581170476427926309478876867395991332060993892808214444723280121094928305947798506576432032165894407230848293965521414076559455665187578833816098594691362634410658602533303813093452867702357567252615476;
            6'd63: xpb[163] = 1024'd72612932538158581873914378873697529458894846987507694139736705842639142170247780710636639164349311074354205081588467347852127100230483354109433557946987631663099380872017036846920260426693831444288510274160951330979128918555035546508012552186546888867941693166623713220525786557803172348925441733653072285177;
        endcase
    end

    always_comb begin
        case(flag[54][16:12])
            5'd0: xpb[164] = 1024'd0;
            5'd1: xpb[164] = 1024'd85581394548363455370211330354690928283134297935792167138284766735218515411424012681600560854068284993894095582006458267777944721584099312227535054900082455111754038463912978765534573054881086456544854653914671813664292315695994533560359916794259961637288694970613015782449039811793251244983181109738891954878;
            5'd2: xpb[164] = 1024'd47096093412602169341623733304567423821570168745848650148437678405460135485538886453186050493478895678345041756555423100976825602326978289899909984783833869289817402358254740193438906918244967191779511699442103780964223781171092294155741263905290474007757486527108973534791551549657869472847672392852189425425;
            5'd3: xpb[164] = 1024'd8610792276840883313036136254443919360006039555905133158590590075701755559653760224771540132889506362795987931104387934175706483069857267572284914667585283467880766252596501621343240781608847927014168744969535748264155246646190054751122611016320986378226278083604931287134063287522487700712163675965486895972;
            5'd4: xpb[164] = 1024'd94192186825204338683247466609134847643140337491697300296875356810920270971077772906372100986957791356690083513110846201953651204653956579799819969567667738579634804716509480386877813836489934383559023398884207561928447562342184588311482527810580948015514973054217947069583103099315738945695344785704378850850;
            5'd5: xpb[164] = 1024'd55706885689443052654659869559011343181576208301753783307028268481161891045192646677957590626368402041141029687659811035152532085396835557472194899451419152757698168610851241814782147699853815118793680444411639529228379027817282348906863874921611460385983764610713904821925614837180357173559836068817676321397;
            5'd6: xpb[164] = 1024'd17221584553681766626072272508887838720012079111810266317181180151403511119307520449543080265779012725591975862208775868351412966139714535144569829335170566935761532505193003242686481563217695854028337489939071496528310493292380109502245222032641972756452556167209862574268126575044975401424327351930973791944;
            5'd7: xpb[164] = 1024'd102802979102045221996283602863578767003146377047602433455465946886622026530731533131143641119847297719486071444215234136129357687723813847372104884235253022047515570969105982008221054618098782310573192143853743310192602808988374643062605138826901934393741251137822878356717166386838226646407508461669865746822;
            5'd8: xpb[164] = 1024'd64317677966283935967696005813455262541582247857658916465618858556863646604846406902729130759257908403937017618764198969328238568466692825044479814119004436225578934863447743436125388481462663045807849189381175277492534274463472403657986485937932446764210042694318836109059678124702844874271999744783163217369;
            5'd9: xpb[164] = 1024'd25832376830522649939108408763331758080018118667715399475771770227105266678961280674314620398668519088387963793313163802527119449209571802716854744002755850403642298757789504864029722344826543781042506234908607244792465739938570164253367833048962959134678834250814793861402189862567463102136491027896460687916;
            5'd10: xpb[164] = 1024'd111413771378886105309319739118022686363152416603507566614056536962323782090385293355915181252736804082282059375319622070305064170793671114944389798902838305515396337221702483629564295399707630237587360888823279058456758055634564697813727749843222920771967529221427809643851229674360714347119672137635352642794;
            5'd11: xpb[164] = 1024'd72928470243124819280732142067899181901588287413564049624209448632565402164500167127500670892147414766733005549868586903503945051536550092616764728786589719693459701116044245057468629263071510972822017934350711025756689521109662458409109096954253433142436320777923767396193741412225332574984163420748650113341;
            5'd12: xpb[164] = 1024'd34443169107363533252144545017775677440024158223620532634362360302807022238615040899086160531558025451183951724417551736702825932279429070289139658670341133871523065010386006485372963126435391708056674979878142993056620986584760219004490444065283945512905112334419725148536253150089950802848654703861947583888;
            5'd13: xpb[164] = 1024'd120024563655726988622355875372466605723158456159412699772647127038025537650039053580686721385626310445078047306424010004480770653863528382516674713570423588983277103474298985250907536181316478164601529633792814806720913302280754752564850360859543907150193807305032740930985292961883202047831835813600839538766;
            5'd14: xpb[164] = 1024'd81539262519965702593768278322343101261594326969469182782800038708267157724153927352272211025036921129528993480972974837679651534606407360189049643454175003161340467368640746678811870044680358899836186679320246774020844767755852513160231707970574419520662598861528698683327804699747820275696327096714137009313;
            5'd15: xpb[164] = 1024'd43053961384204416565180681272219596800030197779525665792952950378508777798268801123857700664447531813979939655521939670878532415349286337861424573337926417339403831262982508106716203908044239635070843724847678741320776233230950273755613055081604931891131390418024656435670316437612438503560818379827434479860;
            5'd16: xpb[164] = 1024'd4568660248443130536593084222096092338466068589582148803105862048750397872383674895443190303858142498430885830070904504077413296092165315533799503221677831517467195157324269534620537771408120370305500770375110708620707698706048034350994402192635444261600181974520614188012828175477056731425309662940731950407;
            5'd17: xpb[164] = 1024'd90150054796806585906804414576787020621600366525374315941390628783968913283807687577043751157926427492324981412077362771855358017676264627761334558121760286629221233621237248300155110826289206826850355424289782522285000014402042567911354318986895405898888876945133629970461867987270307976408490772679623905285;
            5'd18: xpb[164] = 1024'd51664753661045299878216817526663516160036237335430798951543540454210533357922561348629240797337038176775927586626327605054238898419143605433709488005511700807284597515579009728059444689653087562085012469817214489584931479877140328506735666097925918269357668501629587722804379725134926204272982055792921375832;
            5'd19: xpb[164] = 1024'd13179452525284013849629220476540011698472108145487281961696452124452153432037435120214730436747648861226873761175292438253119779162022583106084417889263114985347961409920771155963778553016968297319669515344646456884862945352238089102117013208956430639826460058125545475146891462999544432137473338906218846379;
            5'd20: xpb[164] = 1024'd98760847073647469219840550831230939981606406081279449099981218859670668843461447801815291290815933855120969343181750706031064500746121895333619472789345570097101999873833749921498351607898054753864524169259318270549155261048232622662476930003216392277115155028738561257595931274792795677120654448645110801257;
            5'd21: xpb[164] = 1024'd60275545937886183191252953781107435520042276891335932110134130529912288917576321573400780930226544539571915517730715539229945381489000873005994402673096984275165363768175511349402685471261935489099181214786750237849086726523330383257858277114246904647583946585234519009938443012657413904985145731758408271804;
            5'd22: xpb[164] = 1024'd21790244802124897162665356730983931058478147701392415120287042200153908991691195344986270569637155224022861692279680372428826262231879850678369332556848398453228727662517272777307019334625816224333838260314182205149018191998428143853239624225277417018052738141730476762280954750522032132849637014871705742351;
            5'd23: xpb[164] = 1024'd107371639350488352532876687085674859341612445637184582258571808935372424403115208026586831423705440217916957274286138640206770983815979162905904387456930853564982766126430251542841592389506902680878692914228854018813310507694422677413599541019537378655341433112343492544729994562315283377832818124610597697229;
            5'd24: xpb[164] = 1024'd68886338214727066504289090035551354880048316447241065268724720605614044477230081798172321063116050902367903448835103473405651864558858140578279317340682267743046130020772012970745926252870783416113349959756285986113241973169520438008980888130567891025810224668839450297072506300179901605697309407723895167776;
            5'd25: xpb[164] = 1024'd30401037078965780475701492985427850418484187257297548278877632275855664551344955569757810702526661586818849623384068306604532745301737118250654247224433681921109493915113774398650260116234664151348007005283717953413173438644618198604362235241598403396279016225335408049415018038044519833561800690837192638323;
            5'd26: xpb[164] = 1024'd115982431627329235845912823340118778701618485193089715417162399011074179962768968251358371556594946580712945205390526574382477466885836430478189302124516137032863532379026753164184833171115750607892861659198389767077465754340612732164722152035858365033567711195948423831864057849837771078544981800576084593201;
            5'd27: xpb[164] = 1024'd77497130491567949817325226289995274240054356003146198427315310681315800036883842022943861196005557265163891379939491407581358347628715408150564232008267551210926896273368514592089167034479631343127518704725821734377397219815710492760103499146888877404036502752444381584206569587702389306409473083689382063748;
            5'd28: xpb[164] = 1024'd39011829355806663788737629239871769778490226813202681437468222351557420110998715794529350835416167949614837554488456240780239228371594385822939161892018965388990260167710276019993500897843512078362175750253253701677328685290808253355484846257919389774505294308940339336549081325567007534273964366802679534295;
            5'd29: xpb[164] = 1024'd526528220045377760150032189748265316926097623259164447621134021799040185113589566114840474826778634065783729037421073979120109114473363495314091775770379567053624062052037447897834761207392813596832795780685668977260150765906013950866193368949902144974085865436297088891593063431625762138455649915977004842;
            5'd30: xpb[164] = 1024'd86107922768408833130361362544439193600060395559051331585905900757017555596537602247715401328895063627959879311043879341757064830698572675722849146675852834678807662525965016213432407816088479270141687449695357482641552466461900547511226110163209863782262780836049312871340632875224877007121636759654868959720;
            5'd31: xpb[164] = 1024'd47622621632647547101773765494315689138496266369107814596058812427259175670652476019300890968305674312410825485592844174955945711441451653395224076559604248856871026420306777641336741679452360005376344495222789449941483931936998308106607457274240376152731572392545270623683144613089495234986128042768166430267;
        endcase
    end

    always_comb begin
        case(flag[55][5:0])
            6'd0: xpb[165] = 1024'd0;
            6'd1: xpb[165] = 1024'd4568660248443130536593084222096092338466068589582148803105862048750397872383674895443190303858142498430885830070904504077413296092165315533799503221677831517467195157324269534620537771408120370305500770375110708620707698706048034350994402192635444261600181974520614188012828175477056731425309662940731950407;
            6'd2: xpb[165] = 1024'd9137320496886261073186168444192184676932137179164297606211724097500795744767349790886380607716284996861771660141809008154826592184330631067599006443355663034934390314648539069241075542816240740611001540750221417241415397412096068701988804385270888523200363949041228376025656350954113462850619325881463900814;
            6'd3: xpb[165] = 1024'd13705980745329391609779252666288277015398205768746446409317586146251193617151024686329570911574427495292657490212713512232239888276495946601398509665033494552401585471972808603861613314224361110916502311125332125862123096118144103052983206577906332784800545923561842564038484526431170194275928988822195851221;
            6'd4: xpb[165] = 1024'd18274640993772522146372336888384369353864274358328595212423448195001591489534699581772761215432569993723543320283618016309653184368661262135198012886711326069868780629297078138482151085632481481222003081500442834482830794824192137403977608770541777046400727898082456752051312701908226925701238651762927801628;
            6'd5: xpb[165] = 1024'd22843301242215652682965421110480461692330342947910744015529310243751989361918374477215951519290712492154429150354522520387066480460826577668997516108389157587335975786621347673102688857040601851527503851875553543103538493530240171754972010963177221308000909872603070940064140877385283657126548314703659752035;
            6'd6: xpb[165] = 1024'd27411961490658783219558505332576554030796411537492892818635172292502387234302049372659141823148854990585314980425427024464479776552991893202797019330066989104803170943945617207723226628448722221833004622250664251724246192236288206105966413155812665569601091847123685128076969052862340388551857977644391702442;
            6'd7: xpb[165] = 1024'd31980621739101913756151589554672646369262480127075041621741034341252785106685724268102332127006997489016200810496331528541893072645157208736596522551744820622270366101269886742343764399856842592138505392625774960344953890942336240456960815348448109831201273821644299316089797228339397119977167640585123652849;
            6'd8: xpb[165] = 1024'd36549281987545044292744673776768738707728548716657190424846896390003182979069399163545522430865139987447086640567236032619306368737322524270396025773422652139737561258594156276964302171264962962444006163000885668965661589648384274807955217541083554092801455796164913504102625403816453851402477303525855603256;
            6'd9: xpb[165] = 1024'd41117942235988174829337757998864831046194617306239339227952758438753580851453074058988712734723282485877972470638140536696719664829487839804195528995100483657204756415918425811584839942673083332749506933375996377586369288354432309158949619733718998354401637770685527692115453579293510582827786966466587553663;
            6'd10: xpb[165] = 1024'd45686602484431305365930842220960923384660685895821488031058620487503978723836748954431903038581424984308858300709045040774132960921653155337995032216778315174671951573242695346205377714081203703055007703751107086207076987060480343509944021926354442616001819745206141880128281754770567314253096629407319504070;
            6'd11: xpb[165] = 1024'd50255262732874435902523926443057015723126754485403636834164482536254376596220423849875093342439567482739744130779949544851546257013818470871794535438456146692139146730566964880825915485489324073360508474126217794827784685766528377860938424118989886877602001719726756068141109930247624045678406292348051454477;
            6'd12: xpb[165] = 1024'd54823922981317566439117010665153108061592823074985785637270344585004774468604098745318283646297709981170629960850854048928959553105983786405594038660133978209606341887891234415446453256897444443666009244501328503448492384472576412211932826311625331139202183694247370256153938105724680777103715955288783404884;
            6'd13: xpb[165] = 1024'd59392583229760696975710094887249200400058891664567934440376206633755172340987773640761473950155852479601515790921758553006372849198149101939393541881811809727073537045215503950066991028305564813971510014876439212069200083178624446562927228504260775400802365668767984444166766281201737508529025618229515355291;
            6'd14: xpb[165] = 1024'd63961243478203827512303179109345292738524960254150083243482068682505570213371448536204664254013994978032401620992663057083786145290314417473193045103489641244540732202539773484687528799713685184277010785251549920689907781884672480913921630696896219662402547643288598632179594456678794239954335281170247305698;
            6'd15: xpb[165] = 1024'd68529903726646958048896263331441385076991028843732232046587930731255968085755123431647854557872137476463287451063567561161199441382479733006992548325167472762007927359864043019308066571121805554582511555626660629310615480590720515264916032889531663924002729617809212820192422632155850971379644944110979256105;
            6'd16: xpb[165] = 1024'd73098563975090088585489347553537477415457097433314380849693792780006365958138798327091044861730279974894173281134472065238612737474645048540792051546845304279475122517188312553928604342529925924888012326001771337931323179296768549615910435082167108185602911592329827008205250807632907702804954607051711206512;
            6'd17: xpb[165] = 1024'd77667224223533219122082431775633569753923166022896529652799654828756763830522473222534235165588422473325059111205376569316026033566810364074591554768523135796942317674512582088549142113938046295193513096376882046552030878002816583966904837274802552447203093566850441196218078983109964434230264269992443156919;
            6'd18: xpb[165] = 1024'd82235884471976349658675515997729662092389234612478678455905516877507161702906148117977425469446564971755944941276281073393439329658975679608391057990200967314409512831836851623169679885346166665499013866751992755172738576708864618317899239467437996708803275541371055384230907158587021165655573932933175107326;
            6'd19: xpb[165] = 1024'd86804544720419480195268600219825754430855303202060827259011378926257559575289823013420615773304707470186830771347185577470852625751140995142190561211878798831876707989161121157790217656754287035804514637127103463793446275414912652668893641660073440970403457515891669572243735334064077897080883595873907057733;
            6'd20: xpb[165] = 1024'd91373204968862610731861684441921846769321371791642976062117240975007957447673497908863806077162849968617716601418090081548265921843306310675990064433556630349343903146485390692410755428162407406110015407502214172414153974120960687019888043852708885232003639490412283760256563509541134628506193258814639008140;
            6'd21: xpb[165] = 1024'd95941865217305741268454768664017939107787440381225124865223103023758355320057172804306996381020992467048602431488994585625679217935471626209789567655234461866811098303809660227031293199570527776415516177877324881034861672827008721370882446045344329493603821464932897948269391685018191359931502921755370958547;
            6'd22: xpb[165] = 1024'd100510525465748871805047852886114031446253508970807273668328965072508753192440847699750186684879134965479488261559899089703092514027636941743589070876912293384278293461133929761651830970978648146721016948252435589655569371533056755721876848237979773755204003439453512136282219860495248091356812584696102908954;
            6'd23: xpb[165] = 1024'd105079185714192002341640937108210123784719577560389422471434827121259151064824522595193376988737277463910374091630803593780505810119802257277388574098590124901745488618458199296272368742386768517026517718627546298276277070239104790072871250430615218016804185413974126324295048035972304822782122247636834859361;
            6'd24: xpb[165] = 1024'd109647845962635132878234021330306216123185646149971571274540689170009548937208197490636567292595419962341259921701708097857919106211967572811188077320267956419212683775782468830892906513794888887332018489002657006896984768945152824423865652623250662278404367388494740512307876211449361554207431910577566809768;
            6'd25: xpb[165] = 1024'd114216506211078263414827105552402308461651714739553720077646551218759946809591872386079757596453562460772145751772612601935332402304132888344987580541945787936679878933106738365513444285203009257637519259377767715517692467651200858774860054815886106540004549363015354700320704386926418285632741573518298760175;
            6'd26: xpb[165] = 1024'd118785166459521393951420189774498400800117783329135868880752413267510344681975547281522947900311704959203031581843517106012745698396298203878787083763623619454147074090431007900133982056611129627943020029752878424138400166357248893125854457008521550801604731337535968888333532562403475017058051236459030710582;
            6'd27: xpb[165] = 1024'd123353826707964524488013273996594493138583851918718017683858275316260742554359222176966138204169847457633917411914421610090158994488463519412586586985301450971614269247755277434754519828019249998248520800127989132759107865063296927476848859201156995063204913312056583076346360737880531748483360899399762660989;
            6'd28: xpb[165] = 1024'd3855791272282913625807430813876152732351493382564482358832282300034245089433758162394257293370315646621653834527832679588508449739408500391225965190648241555390789835508329631744818407910164647243823962115859995015454713548448188862864691710562990057985191872460139234252660839428955462789980735714900127065;
            6'd29: xpb[165] = 1024'd8424451520726044162400515035972245070817561972146631161938144348784642961817433057837447597228458145052539664598737183665921745831573815925025468412326073072857984992832599166365356179318285017549324732490970703636162412254496223213859093903198434319585373846980753422265489014906012194215290398655632077472;
            6'd30: xpb[165] = 1024'd12993111769169174698993599258068337409283630561728779965044006397535040834201107953280637901086600643483425494669641687743335041923739131458824971634003904590325180150156868700985893950726405387854825502866081412256870110960544257564853496095833878581185555821501367610278317190383068925640600061596364027879;
            6'd31: xpb[165] = 1024'd17561772017612305235586683480164429747749699151310928768149868446285438706584782848723828204944743141914311324740546191820748338015904446992624474855681736107792375307481138235606431722134525758160326273241192120877577809666592291915847898288469322842785737796021981798291145365860125657065909724537095978286;
            6'd32: xpb[165] = 1024'd22130432266055435772179767702260522086215767740893077571255730495035836578968457744167018508802885640345197154811450695898161634108069762526423978077359567625259570464805407770226969493542646128465827043616302829498285508372640326266842300481104767104385919770542595986303973541337182388491219387477827928693;
            6'd33: xpb[165] = 1024'd26699092514498566308772851924356614424681836330475226374361592543786234451352132639610208812661028138776082984882355199975574930200235078060223481299037399142726765622129677304847507264950766498771327813991413538118993207078688360617836702673740211365986101745063210174316801716814239119916529050418559879100;
            6'd34: xpb[165] = 1024'd31267752762941696845365936146452706763147904920057375177467454592536632323735807535053399116519170637206968814953259704052988226292400393594022984520715230660193960779453946839468045036358886869076828584366524246739700905784736394968831104866375655627586283719583824362329629892291295851341838713359291829507;
            6'd35: xpb[165] = 1024'd35836413011384827381959020368548799101613973509639523980573316641287030196119482430496589420377313135637854645024164208130401522384565709127822487742393062177661155936778216374088582807767007239382329354741634955360408604490784429319825507059011099889186465694104438550342458067768352582767148376300023779914;
            6'd36: xpb[165] = 1024'd40405073259827957918552104590644891440080042099221672783679178690037428068503157325939779724235455634068740475095068712207814818476731024661621990964070893695128351094102485908709120579175127609687830125116745663981116303196832463670819909251646544150786647668625052738355286243245409314192458039240755730321;
            6'd37: xpb[165] = 1024'd44973733508271088455145188812740983778546110688803821586785040738787825940886832221382970028093598132499626305165973216285228114568896340195421494185748725212595546251426755443329658350583247979993330895491856372601824001902880498021814311444281988412386829643145666926368114418722466045617767702181487680728;
            6'd38: xpb[165] = 1024'd49542393756714218991738273034837076117012179278385970389890902787538223813270507116826160331951740630930512135236877720362641410661061655729220997407426556730062741408751024977950196121991368350298831665866967081222531700608928532372808713636917432673987011617666281114380942594199522777043077365122219631135;
            6'd39: xpb[165] = 1024'd54111054005157349528331357256933168455478247867968119192996764836288621685654182012269350635809883129361397965307782224440054706753226971263020500629104388247529936566075294512570733893399488720604332436242077789843239399314976566723803115829552876935587193592186895302393770769676579508468387028062951581542;
            6'd40: xpb[165] = 1024'd58679714253600480064924441479029260793944316457550267996102626885039019558037856907712540939668025627792283795378686728517468002845392286796820003850782219764997131723399564047191271664807609090909833206617188498463947098021024601074797518022188321197187375566707509490406598945153636239893696691003683531949;
            6'd41: xpb[165] = 1024'd63248374502043610601517525701125353132410385047132416799208488933789417430421531803155731243526168126223169625449591232594881298937557602330619507072460051282464326880723833581811809436215729461215333976992299207084654796727072635425791920214823765458787557541228123678419427120630692971319006353944415482356;
            6'd42: xpb[165] = 1024'd67817034750486741138110609923221445470876453636714565602314350982539815302805206698598921547384310624654055455520495736672294595029722917864419010294137882799931522038048103116432347207623849831520834747367409915705362495433120669776786322407459209720387739515748737866432255296107749702744316016885147432763;
            6'd43: xpb[165] = 1024'd72385694998929871674703694145317537809342522226296714405420213031290213175188881594042111851242453123084941285591400240749707891121888233398218513515815714317398717195372372651052884979031970201826335517742520624326070194139168704127780724600094653981987921490269352054445083471584806434169625679825879383170;
            6'd44: xpb[165] = 1024'd76954355247373002211296778367413630147808590815878863208526075080040611047572556489485302155100595621515827115662304744827121187214053548932018016737493545834865912352696642185673422750440090572131836288117631332946777892845216738478775126792730098243588103464789966242457911647061863165594935342766611333577;
            6'd45: xpb[165] = 1024'd81523015495816132747889862589509722486274659405461012011631937128791008919956231384928492458958738119946712945733209248904534483306218864465817519959171377352333107510020911720293960521848210942437337058492742041567485591551264772829769528985365542505188285439310580430470739822538919897020245005707343283984;
            6'd46: xpb[165] = 1024'd86091675744259263284482946811605814824740727995043160814737799177541406792339906280371682762816880618377598775804113752981947779398384179999617023180849208869800302667345181254914498293256331312742837828867852750188193290257312807180763931178000986766788467413831194618483567998015976628445554668648075234391;
            6'd47: xpb[165] = 1024'd90660335992702393821076031033701907163206796584625309617843661226291804664723581175814873066675023116808484605875018257059361075490549495533416526402527040387267497824669450789535036064664451683048338599242963458808900988963360841531758333370636431028388649388351808806496396173493033359870864331588807184798;
            6'd48: xpb[165] = 1024'd95228996241145524357669115255797999501672865174207458420949523275042202537107256071258063370533165615239370435945922761136774371582714811067216029624204871904734692981993720324155573836072572053353839369618074167429608687669408875882752735563271875289988831362872422994509224348970090091296173994529539135205;
            6'd49: xpb[165] = 1024'd99797656489588654894262199477894091840138933763789607224055385323792600409490930966701253674391308113670256266016827265214187667674880126601015532845882703422201888139317989858776111607480692423659340139993184876050316386375456910233747137755907319551589013337393037182522052524447146822721483657470271085612;
            6'd50: xpb[165] = 1024'd104366316738031785430855283699990184178605002353371756027161247372542998281874605862144443978249450612101142096087731769291600963767045442134815036067560534939669083296642259393396649378888812793964840910368295584671024085081504944584741539948542763813189195311913651370534880699924203554146793320411003036019;
            6'd51: xpb[165] = 1024'd108934976986474915967448367922086276517071070942953904830267109421293396154258280757587634282107593110532027926158636273369014259859210757668614539289238366457136278453966528928017187150296933164270341680743406293291731783787552978935735942141178208074789377286434265558547708875401260285572102983351734986426;
            6'd52: xpb[165] = 1024'd113503637234918046504041452144182368855537139532536053633372971470043794026641955653030824585965735608962913756229540777446427555951376073202414042510916197974603473611290798462637724921705053534575842451118517001912439482493601013286730344333813652336389559260954879746560537050878317016997412646292466936833;
            6'd53: xpb[165] = 1024'd118072297483361177040634536366278461194003208122118202436478833518794191899025630548474014889823878107393799586300445281523840852043541388736213545732594029492070668768615067997258262693113173904881343221493627710533147181199649047637724746526449096597989741235475493934573365226355373748422722309233198887240;
            6'd54: xpb[165] = 1024'd122640957731804307577227620588374553532469276711700351239584695567544589771409305443917205193682020605824685416371349785601254148135706704270013048954271861009537863925939337531878800464521294275186843991868738419153854879905697081988719148719084540859589923209996108122586193401832430479848031972173930837647;
            6'd55: xpb[165] = 1024'd3142922296122696715021777405656213126236918175546815914558702551318092306483841429345324282882488794812421838984760855099603603386651685248652427159618651593314384513692389728869099044412208924182147153856609281410201728390848343374734981228490535854370201770399664280492493503380854194154651808489068303723;
            6'd56: xpb[165] = 1024'd7711582544565827251614861627752305464702986765128964717664564600068490178867516324788514586740631293243307669055665359177016899478817000782451930381296483110781579671016659263489636815820329294487647924231719990030909427096896377725729383421125980115970383744920278468505321678857910925579961471429800254130;
            6'd57: xpb[165] = 1024'd12280242793008957788207945849848397803169055354711113520770426648818888051251191220231704890598773791674193499126569863254430195570982316316251433602974314628248774828340928798110174587228449664793148694606830698651617125802944412076723785613761424377570565719440892656518149854334967657005271134370532204537;
            6'd58: xpb[165] = 1024'd16848903041452088324801030071944490141635123944293262323876288697569285923634866115674895194456916290105079329197474367331843491663147631850050936824652146145715969985665198332730712358636570035098649464981941407272324824508992446427718187806396868639170747693961506844530978029812024388430580797311264154944;
            6'd59: xpb[165] = 1024'd21417563289895218861394114294040582480101192533875411126982150746319683796018541011118085498315058788535965159268378871409256787755312947383850440046329977663183165142989467867351250130044690405404150235357052115893032523215040480778712589999032312900770929668482121032543806205289081119855890460251996105351;
            6'd60: xpb[165] = 1024'd25986223538338349397987198516136674818567261123457559930088012795070081668402215906561275802173201286966850989339283375486670083847478262917649943268007809180650360300313737401971787901452810775709651005732162824513740221921088515129706992191667757162371111643002735220556634380766137851281200123192728055758;
            6'd61: xpb[165] = 1024'd30554883786781479934580282738232767157033329713039708733193874843820479540785890802004466106031343785397736819410187879564083379939643578451449446489685640698117555457638006936592325672860931146015151776107273533134447920627136549480701394384303201423971293617523349408569462556243194582706509786133460006165;
            6'd62: xpb[165] = 1024'd35123544035224610471173366960328859495499398302621857536299736892570877413169565697447656409889486283828622649481092383641496676031808893985248949711363472215584750614962276471212863444269051516320652546482384241755155619333184583831695796576938645685571475592043963596582290731720251314131819449074191956572;
            6'd63: xpb[165] = 1024'd39692204283667741007766451182424951833965466892204006339405598941321275285553240592890846713747628782259508479551996887718909972123974209519048452933041303733051945772286546005833401215677171886626153316857494950375863318039232618182690198769574089947171657566564577784595118907197308045557129112014923906979;
        endcase
    end

    always_comb begin
        case(flag[55][11:6])
            6'd0: xpb[166] = 1024'd0;
            6'd1: xpb[166] = 1024'd44260864532110871544359535404521044172431535481786155142511460990071673157936915488334037017605771280690394309622901391796323268216139525052847956154719135250519140929610815540453938987085292256931654087232605658996571016745280652533684600962209534208771839541085191972607947082674364776982438774955655857386;
            6'd2: xpb[166] = 1024'd88521729064221743088719070809042088344863070963572310285022921980143346315873830976668074035211542561380788619245802783592646536432279050105695912309438270501038281859221631080907877974170584513863308174465211317993142033490561305067369201924419068417543679082170383945215894165348729553964877549911311714772;
            6'd3: xpb[166] = 1024'd8715897912207873234279678808748699772596179319622781299402527905238124136501607554987039838159639532628033521411210740809905963807198240603383743447826364817866748219261229283731577769738671049484764653310577130625352200014945184636075233203399153359495615209138517887717313174094461313828626498241373087827;
            6'd4: xpb[166] = 1024'd52976762444318744778639214213269743945027714801408936441913988895309797294438523043321076855765410813318427831034112132606229232023337765656231699602545500068385889148872044824185516756823963306416418740543182789621923216760225837169759834165608687568267454750223709860325260256768826090811065273197028945213;
            6'd5: xpb[166] = 1024'd97237626976429616322998749617790788117459250283195091584425449885381470452375438531655113873371182094008822140657013524402552500239477290709079655757264635318905030078482860364639455743909255563348072827775788448618494233505506489703444435127818221777039294291308901832933207339443190867793504048152684802599;
            6'd6: xpb[166] = 1024'd17431795824415746468559357617497399545192358639245562598805055810476248273003215109974079676319279065256067042822421481619811927614396481206767486895652729635733496438522458567463155539477342098969529306621154261250704400029890369272150466406798306718991230418277035775434626348188922627657252996482746175654;
            6'd7: xpb[166] = 1024'd61692660356526618012918893022018443717623894121031717741316516800547921430940130598308116693925050345946461352445322873416135195830536006259615443050371864886252637368133274107917094526562634355901183393853759920247275416775171021805835067369007840927763069959362227748042573430863287404639691771438402033040;
            6'd8: xpb[166] = 1024'd105953524888637489557278428426539487890055429602817872883827977790619594588877046086642153711530821626636855662068224265212458464046675531312463399205091000136771778297744089648371033513647926612832837481086365579243846433520451674339519668331217375136534909500447419720650520513537652181622130546394057890426;
            6'd9: xpb[166] = 1024'd26147693736623619702839036426246099317788537958868343898207583715714372409504822664961119514478918597884100564233632222429717891421594721810151230343479094453600244657783687851194733309216013148454293959931731391876056600044835553908225699610197460078486845627415553663151939522283383941485879494724119263481;
            6'd10: xpb[166] = 1024'd70408558268734491247198571830767143490220073440654499040719044705786045567441738153295156532084689878574494873856533614226041159637734246862999186498198229704119385587394503391648672296301305405385948047164337050872627616790116206441910300572406994287258685168500745635759886604957748718468318269679775120867;
            6'd11: xpb[166] = 1024'd114669422800845362791558107235288187662651608922440654183230505695857718725378653641629193549690461159264889183479435006022364427853873771915847142652917364954638526517005318932102611283386597662317602134396942709869198633535396858975594901534616528496030524709585937608367833687632113495450757044635430978253;
            6'd12: xpb[166] = 1024'd34863591648831492937118715234994799090384717278491125197610111620952496546006430219948159352638558130512134085644842963239623855228792962413534973791305459271466992877044917134926311078954684197939058613242308522501408800059780738544300932813596613437982460836554071550869252696377845255314505992965492351308;
            6'd13: xpb[166] = 1024'd79124456180942364481478250639515843262816252760277280340121572611024169703943345708282196370244329411202528395267744355035947123444932487466382929946024594521986133806655732675380250066039976454870712700474914181497979816805061391077985533775806147646754300377639263523477199779052210032296944767921148208694;
            6'd14: xpb[166] = 1024'd123385320713053236025837786044036887435247788242063435482633033601095842861880261196616233387850100691892922704890645746832270391661072012519230886100743729772505274736266548215834189053125268711802366787707519840494550833550342043611670134738015681855526139918724455496085146861726574809279383542876804066080;
            6'd15: xpb[166] = 1024'd43579489561039366171398394043743498862980896598113906497012639526190620682508037774935199190798197663140167607056053704049529819035991203016918717239131824089333741096306146418657888848693355247423823266552885653126761000074725923180376166016995766797478076045692589438586565870472306569143132491206865439135;
            6'd16: xpb[166] = 1024'd87840354093150237715757929448264543035412432079900061639524100516262293840444953263269236208403968943830561916678955095845853087252130728069766673393850959339852882025916961959111827835778647504355477353785491312123332016820006575714060766979205301006249915586777781411194512953146671346125571266162521296521;
            6'd17: xpb[166] = 1024'd8034522941136367861318537447971154463145540435950532653903706441357071661072729841588202011352065915077806818844363053063112514627049918567454504532239053656681348385956560161935527631346734039976933832630857124755542183344390455282766798258185385948201851713745915353695931961892403105989320214492582669576;
            6'd18: xpb[166] = 1024'd52295387473247239405678072852492198635577075917736687796415167431428744819009645329922239028957837195768201128467264444859435782843189443620302460686958188907200489315567375702389466618432026296908587919863462783752113200089671107816451399220394920156973691254831107326303879044566767882971758989448238526962;
            6'd19: xpb[166] = 1024'd96556252005358110950037608257013242808008611399522842938926628421500417976946560818256276046563608476458595438090165836655759051059328968673150416841677324157719630245178191242843405605517318553840242007096068442748684216834951760350136000182604454365745530795916299298911826127241132659954197764403894384348;
            6'd20: xpb[166] = 1024'd16750420853344241095598216256719854235741719755573313953306234346595195797574337396575241849511705447705840340255573793873018478434248159170838247980065418474548096605217789445667105401085405089461698485941434255380894383359335639918842031461584539307697466922884433241413245135986864419817946712733955757403;
            6'd21: xpb[166] = 1024'd61011285385455112639957751661240898408173255237359469095817695336666868955511252884909278867117476728396234649878475185669341746650387684223686204134784553725067237534828604986121044388170697346393352573174039914377465400104616292452526632423794073516469306463969625214021192218661229196800385487689611614789;
            6'd22: xpb[166] = 1024'd105272149917565984184317287065761942580604790719145624238329156326738542113448168373243315884723248009086628959501376577465665014866527209276534160289503688975586378464439420526574983375255989603325006660406645573374036416849896944986211233386003607725241146005054817186629139301335593973782824262645267472175;
            6'd23: xpb[166] = 1024'd25466318765552114329877895065468554008337899075196095252708762251833319934075944951562281687671344980333873861666784534682924442241446399774221991427891783292414844824479018729398683170824076138946463139252011386006246583374280824554917264664983692667193082132022951129130558310081325733646573210975328845230;
            6'd24: xpb[166] = 1024'd69727183297662985874237430469989598180769434556982250395220223241904993092012860439896318705277116261024268171289685926479247710457585924827069947582610918542933985754089834269852622157909368395878117226484617045002817600119561477088601865627193226875964921673108143101738505392755690510629011985930984702616;
            6'd25: xpb[166] = 1024'd113988047829773857418596965874510642353200970038768405537731684231976666249949775928230355722882887541714662480912587318275570978673725449879917903737330053793453126683700649810306561144994660652809771313717222703999388616864842129622286466589402761084736761214193335074346452475430055287611450760886640560002;
            6'd26: xpb[166] = 1024'd34182216677759987564157573874217253780934078394818876552111290157071444070577552506549321525830984512961907383077995275492830406048644640377605734875718148110281593043740248013130260940562747188431227792562588516631598783389226009190992497868382846026688697341161469016847871484175787047475199709216701933057;
            6'd27: xpb[166] = 1024'd78443081209870859108517109278738297953365613876605031694622751147143117228514467994883358543436755793652301692700896667289153674264784165430453691030437283360800733973351063553584199927648039445362881879795194175628169800134506661724677098830592380235460536882246660989455818566850151824457638484172357790443;
            6'd28: xpb[166] = 1024'd122703945741981730652876644683259342125797149358391186837134212137214790386451383483217395561042527074342696002323798059085476942480923690483301647185156418611319874902961879094038138914733331702294535967027799834624740816879787314258361699792801914444232376423331852962063765649524516601440077259128013647829;
            6'd29: xpb[166] = 1024'd42898114589967860798437252682965953553530257714441657851513818062309568207079160061536361363990624045589940904489206016302736369855842880980989478323544512928148341263001477296861838710301418237915992445873165647256950983404171193827067731071781999386184312550299986904565184658270248361303826207458075020884;
            6'd30: xpb[166] = 1024'd87158979122078732342796788087486997725961793196227812994025279052381241365016075549870398381596395326280335214112107408099059638071982406033837434478263648178667482192612292837315777697386710494847646533105771306253522000149451846360752332033991533594956152091385178877173131740944613138286264982413730878270;
            6'd31: xpb[166] = 1024'd7353147970064862488357396087193609153694901552278284008404884977476019185643852128189364184544492297527580116277515365316319065446901596531525265616651742495495948552651891040139477492954797030469103011951137118885732166673835725929458363312971618536908088218353312819674550749690344898150013930743792251325;
            6'd32: xpb[166] = 1024'd51614012502175734032716931491714653326126437034064439150916345967547692343580767616523401202150263578217974425900416757112642333663041121584373221771370877746015089482262706580593416480040089287400757099183742777882303183419116378463142964275181152745679927759438504792282497832364709675132452705699448108711;
            6'd33: xpb[166] = 1024'd95874877034286605577076466896235697498557972515850594293427806957619365501517683104857438219756034858908368735523318148908965601879180646637221177926090012996534230411873522121047355467125381544332411186416348436878874200164397030996827565237390686954451767300523696764890444915039074452114891480655103966097;
            6'd34: xpb[166] = 1024'd16069045882272735722637074895942308926291080871901065307807412882714143322145459683176404022704131830155613637688726106126225029254099837134909009064478107313362696771913120323871055262693468079953867665261714249511084366688780910565533596516370771896403703427491830707391863923784806211978640428985165339152;
            6'd35: xpb[166] = 1024'd60329910414383607266996610300463353098722616353687220450318873872785816480082375171510441040309903110846007947311627497922548297470239362187756965219197242563881837701523935864324994249778760336885521752494319908507655383434061563099218197478580306105175542968577022679999811006459170988961079203940821196538;
            6'd36: xpb[166] = 1024'd104590774946494478811356145704984397271154151835473375592830334862857489638019290659844478057915674391536402256934528889718871565686378887240604921373916377814400978631134751404778933236864052593817175839726925567504226400179342215632902798440789840313947382509662214652607758089133535765943517978896477053924;
            6'd37: xpb[166] = 1024'd24784943794480608956916753704691008698887260191523846607209940787952267458647067238163443860863771362783647159099936846936130993061298077738292752512304472131229444991174349607602633032432139129438632318572291380136436566703726095201608829719769925255899318636630348595109177097879267525807266927226538426979;
            6'd38: xpb[166] = 1024'd69045808326591480501276289109212052871318795673310001749721401778023940616583982726497480878469542643474041468722838238732454261277437602791140708667023607381748585920785165148056572019517431386370286405804897039133007583449006747735293430681979459464671158177715540567717124180553632302789705702182194284365;
            6'd39: xpb[166] = 1024'd113306672858702352045635824513733097043750331155096156892232862768095613774520898214831517896075313924164435778345739630528777529493577127843988664821742742632267726850395980688510511006602723643301940493037502698129578600194287400268978031644188993673442997718800732540325071263227997079772144477137850141751;
            6'd40: xpb[166] = 1024'd33500841706688482191196432513439708471483439511146627906612468693190391595148674793150483699023410895411680680511147587746036956868496318341676495960130836949096193210435578891334210802170810178923396971882868510761788766718671279837684062923169078615394933845768866482826490271973728839635893425467911514806;
            6'd41: xpb[166] = 1024'd77761706238799353735555967917960752643914974992932783049123929683262064753085590281484520716629182176102074990134048979542360225084635843394524452114849972199615334140046394431788149789256102435855051059115474169758359783463951932371368663885378612824166773386854058455434437354648093616618332200423567372192;
            6'd42: xpb[166] = 1024'd122022570770910225279915503322481796816346510474718938191635390673333737911022505769818557734234953456792469299756950371338683493300775368447372408269569107450134475069657209972242088776341394692786705146348079828754930800209232584905053264847588147032938612927939250428042384437322458393600770975379223229578;
            6'd43: xpb[166] = 1024'd42216739618896355425476111322188408244079618830769409206014996598428515731650282348137523537183050428039714201922358328555942920675694558945060239407957201766962941429696808175065788571909481228408161625193445641387140966733616464473759296126568231974890549054907384370543803446068190153464519923709284602633;
            6'd44: xpb[166] = 1024'd86477604151007226969835646726709452416511154312555564348526457588500188889587197836471560554788821708730108511545259720352266188891834083997908195562676337017482082359307623715519727558994773485339815712426051300383711983478897117007443897088777766183662388595992576343151750528742554930446958698664940460019;
            6'd45: xpb[166] = 1024'd6671772998993357115396254726416063844244262668606035362906063513594966710214974414790526357736918679977353413710667677569525616266753274495596026701064431334310548719347221918343427354562860020961272191271417113015922150003280996576149928367757851125614324722960710285653169537488286690310707646995001833074;
            6'd46: xpb[166] = 1024'd50932637531104228659755790130937108016675798150392190505417524503666639868151889903124563375342689960667747723333569069365848884482892799548443982855783566584829689648958037458797366341648152277892926278504022772012493166748561649109834529329967385334386164264045902258261116620162651467293146421950657690460;
            6'd47: xpb[166] = 1024'd95193502063215100204115325535458152189107333632178345647928985493738313026088805391458600392948461241358142032956470461162172152699032324601291939010502701835348830578568852999251305328733444534824580365736628431009064183493842301643519130292176919543158003805131094230869063702837016244275585196906313547846;
            6'd48: xpb[166] = 1024'd15387670911201230349675933535164763616840441988228816662308591418833090846716581969777566195896558212605386935121878418379431580073951515098979770148890796152177296938608451202075005124301531070446036844581994243641274350018226181212225161571157004485109939932099228173370482711582748004139334145236374920901;
            6'd49: xpb[166] = 1024'd59648535443312101894035468939685807789271977470014971804820052408904764004653497458111603213502329493295781244744779810175754848290091040151827726303609931402696437868219266742528944111386823327377690931814599902637845366763506833745909762533366538693881779473184420145978429794257112781121772920192030778287;
            6'd50: xpb[166] = 1024'd103909399975422973438395004344206851961703512951801126947331513398976437162590412946445640231108100773986175554367681201972078116506230565204675682458329066653215578797830082282982883098472115584309345019047205561634416383508787486279594363495576072902653619014269612118586376876931477558104211695147686635673;
            6'd51: xpb[166] = 1024'd24103568823409103583955612343913463389436621307851597961711119324071214983218189524764606034056197745233420456533089159189337543881149755702363513596717160970044045157869680485806582894040202119930801497892571374266626550033171365848300394774556157844605555141237746061087795885677209317967960643477748008728;
            6'd52: xpb[166] = 1024'd68364433355519975128315147748434507561868156789637753104222580314142888141155105013098643051661969025923814766155990550985660812097289280755211469751436296220563186087480496026260521881125494376862455585125177033263197566778452018381984995736765692053377394682322938033695742968351574094950399418433403866114;
            6'd53: xpb[166] = 1024'd112625297887630846672674683152955551734299692271423908246734041304214561299092020501432680069267740306614209075778891942781984080313428805808059425906155431471082327017091311566714460868210786633794109672357782692259768583523732670915669596698975226262149234223408130006303690051025938871932838193389059723500;
            6'd54: xpb[166] = 1024'd32819466735616976818235291152662163162032800627474379261113647229309339119719797079751645872215837277861453977944299899999243507688347996305747257044543525787910793377130909769538160663778873169415566151203148504891978750048116550484375627977955311204101170350376263948805109059771670631796587141719121096555;
            6'd55: xpb[166] = 1024'd77080331267727848362594826557183207334464336109260534403625108219381012277656712568085682889821608558551848287567201291795566775904487521358595213199262661038429934306741725309992099650864165426347220238435754163888549766793397203018060228940164845412873009891461455921413056142446035408779025916674776953941;
            6'd56: xpb[166] = 1024'd121341195799838719906954361961704251506895871591046689546136569209452685435593628056419719907427379839242242597190102683591890044120627046411443169353981796288949075236352540850446038637949457683278874325668359822885120783538677855551744829902374379621644849432546647894021003225120400185761464691630432811327;
            6'd57: xpb[166] = 1024'd41535364647824850052514969961410862934628979947097160560516175134547463256221404634738685710375476810489487499355510640809149471495546236909131000492369890605777541596392139053269738433517544218900330804513725635517330950063061735120450861181354464563596785559514781836522422233866131945625213639960494184382;
            6'd58: xpb[166] = 1024'd85796229179935721596874505365931907107060515428883315703027636124619136414158320123072722727981248091179881808978412032605472739711685761961978956647089025856296682526002954593723677420602836475831984891746331294513901966808342387654135462143563998772368625100599973809130369316540496722607652414916150041768;
            6'd59: xpb[166] = 1024'd5990398027921851742435113365638518534793623784933786717407242049713914234786096701391688530929345062427126711143819989822732167086604952459666787785477120173125148886042552796547377216170923011453441370591697107146112133332726267222841493422544083714320561227568107751631788325286228482471401363246211414823;
            6'd60: xpb[166] = 1024'd50251262560032723286794648770159562707225159266719941859918703039785587392723012189725725548535116343117521020766721381619055435302744477512514743940196255423644289815653368337001316203256215268385095457824302766142683150078006919756526094384753617923092400768653299724239735407960593259453840138201867272209;
            6'd61: xpb[166] = 1024'd94512127092143594831154184174680606879656694748506097002430164029857260550659927678059762566140887623807915330389622773415378703518884002565362700094915390674163430745264183877455255190341507525316749545056908425139254166823287572290210695346963152131864240309738491696847682490634958036436278913157523129595;
            6'd62: xpb[166] = 1024'd14706295940129724976714792174387218307389803104556568016809769954952038371287704256378728369088984595055160232555030730632638130893803193063050531233303484990991897105303782080278954985909594060938206023902274237771464333347671451858916726625943237073816176436706625639349101499380689796300027861487584502650;
            6'd63: xpb[166] = 1024'd58967160472240596521074327578908262479821338586342723159321230945023711529224619744712765386694755875745554542177932122428961399109942718115898487388022620241511038034914597620732893972994886317869860111134879896768035350092952104392601327588152771282588015977791817611957048582055054573282466636443240360036;
        endcase
    end

    always_comb begin
        case(flag[55][16:12])
            5'd0: xpb[167] = 1024'd0;
            5'd1: xpb[167] = 1024'd103228025004351468065433862983429306652252874068128878301832691935095384687161535233046802404300527156435948851800833514225284667326082243168746443542741755492030178964525413161186832960080178574801514198367485555764606366838232756926285928550362305491359855518877009584564995664729419350264905411398896217422;
            5'd2: xpb[167] = 1024'd82389354324578194732068798562044180559807321010522072475533528805213874037013931556078533593943380003428748296144173593871505493810944151782332762069152470050369683359479608984743426728643151428292830788347731265164851883455568740887593287417495161715899807623636961139023463255530205683411120996172197950513;
            5'd3: xpb[167] = 1024'd61550683644804921398703734140659054467361767952915266649234365675332363386866327879110264783586232850421547740487513673517726320295806060395919080595563184608709187754433804808300020497206124281784147378327976974565097400072904724848900646284628017940439759728396912693481930846330992016557336580945499683604;
            5'd4: xpb[167] = 1024'd40712012965031648065338669719273928374916214895308460822935202545450852736718724202141995973229085697414347184830853753163947146780667969009505399121973899167048692149388000631856614265769097135275463968308222683965342916690240708810208005151760874164979711833156864247940398437131778349703552165718801416695;
            5'd5: xpb[167] = 1024'd19873342285258374731973605297888802282470661837701654996636039415569342086571120525173727162871938544407146629174193832810167973265529877623091717648384613725388196544342196455413208034332069988766780558288468393365588433307576692771515364018893730389519663937916815802398866027932564682849767750492103149786;
            5'd6: xpb[167] = 1024'd123101367289609842797407468281318108934723535905830533298468731350664726773732655758220529567172465700843095480975027347035452640591612120791838161191126369217418375508867609616600040994412248563568294756655953949130194800145809449697801292569256035880879519456793825386963861692661984033114673161890999367208;
            5'd7: xpb[167] = 1024'd102262696609836569464042403859932982842277982848223727472169568220783216123585052081252260756815318547835894925318367426681673467076474029405424479717537083775757879903821805440156634762975221417059611346636199658530440316763145433659108651436388892105419471561553776941422329283462770366260888746664301100299;
            5'd8: xpb[167] = 1024'd81424025930063296130677339438547856749832429790616921645870405090901705473437448404283991946458171394828694369661707506327894293561335938019010798243947798334097384298776001263713228531538194270550927936616445367930685833380481417620416010303521748329959423666313728495880796874263556699407104331437602833390;
            5'd9: xpb[167] = 1024'd60585355250290022797312275017162730657386876733010115819571241961020194823289844727315723136101024241821493814005047585974115120046197846632597116770358512892436888693730197087269822300101167124042244526596691077330931349997817401581723369170654604554499375771073680050339264465064343032553319916210904566481;
            5'd10: xpb[167] = 1024'd39746684570516749463947210595777604564941323675403309993272078831138684173142241050347454325743877088814293258348387665620335946531059755246183435296769227450776393088684392910826416068664139977533561116576936786731176866615153385543030728037787460779039327875833631604797732055865129365699535500984206299572;
            5'd11: xpb[167] = 1024'd18908013890743476130582146174392478472495770617796504166972915701257173522994637373379185515386729935807092702691727745266556773015921663859769753823179942009115897483638588734383009837227112831024877706557182496131422383232489369504338086904920317003579279980593583159256199646665915698845751085757508032663;
            5'd12: xpb[167] = 1024'd122136038895094944196016009157821785124748644685925382468805607636352558210156172606425987919687257092243041554492561259491841440342003907028516197365921697501146076448164001895569842797307291405826391904924668051896028750070722126430624015455282622494939135499470592743821195311395335049110656497156404250085;
            5'd13: xpb[167] = 1024'd101297368215321670862650944736436659032303091628318576642506444506471047560008568929457719109330109939235840998835901339138062266826865815642102515892332412059485580843118197719126436565870264259317708494904913761296274266688058110391931374322415478719479087604230544298279662902196121382256872081929705983176;
            5'd14: xpb[167] = 1024'd80458697535548397529285880315051532939857538570711770816207281376589536909860965252489450298972962786228640443179241418784283093311727724255688834418743126617825085238072393542683030334433237112809025084885159470696519783305394094353238733189548334944019039708990495852738130492996907715403087666703007716267;
            5'd15: xpb[167] = 1024'd59620026855775124195920815893666406847411985513104964989908118246708026259713361575521181488615815633221439887522581498430503919796589632869275152945153841176164589633026589366239624102996209966300341674865405180096765299922730078314546092056681191168558991813750447407196598083797694048549303251476309449358;
            5'd16: xpb[167] = 1024'd38781356176001850862555751472281280754966432455498159163608955116826515609565757898552912678258668480214239331865921578076724746281451541482861471471564555734504094027980785189796217871559182819791658264845650889497010816540066062275853450923814047393098943918510398961655065674598480381695518836249611182449;
            5'd17: xpb[167] = 1024'd17942685496228577529190687050896154662520879397891353337309791986945004959418154221584643867901521327207038776209261657722945572766313450096447789997975270292843598422934981013352811640122155673282974854825896598897256333157402046237160809790946903617638896023270350516113533265399266714841734421022912915540;
            5'd18: xpb[167] = 1024'd121170710500580045594624550034325461314773753466020231639142483922040389646579689454631446272202048483642987628010095171948230240092395693265194233540717025784873777387460394174539644600202334248084489053193382154661862699995634803163446738341309209108998751542147360100678528930128686065106639832421809132962;
            5'd19: xpb[167] = 1024'd100332039820806772261259485612940335222328200408413425812843320792158878996432085777663177461844901330635787072353435251594451066577257601878780552067127740343213281782414589998096238368765307101575805643173627864062108216612970787124754097208442065333538703646907311655136996520929472398252855417195110866053;
            5'd20: xpb[167] = 1024'd79493369141033498927894421191555209129882647350806619986544157662277368346284482100694908651487754177628586516696775331240671893062119510492366870593538454901552786177368785821652832137328279955067122233153873573462353733230306771086061456075574921558078655751667263209595464111730258731399071001968412599144;
            5'd21: xpb[167] = 1024'd58654698461260225594529356770170083037437094293199814160244994532395857696136878423726639841130607024621385961040115410886892719546981419105953189119949169459892290572322981645209425905891252808558438823134119282862599249847642755047368814942707777782618607856427214764053931702531045064545286586741714332235;
            5'd22: xpb[167] = 1024'd37816027781486952261164292348784956944991541235593008333945831402514347045989274746758371030773459871614185405383455490533113546031843327719539507646359884018231794967277177468766019674454225662049755413114364992262844766464978739008676173809840634007158559961187166318512399293331831397691502171515016065326;
            5'd23: xpb[167] = 1024'd16977357101713678927799227927399830852545988177986202507646668272632836395841671069790102220416312718606984849726795570179334372516705236333125826172770598576571299362231373292322613443017198515541072003094610701663090283082314722969983532676973490231698512065947117872970866884132617730837717756288317798417;
            5'd24: xpb[167] = 1024'd120205382106065146993233090910829137504798862246115080809479360207728221083003206302836904624716839875042933701527629084404619039842787479501872269715512354068601478326756786453509446403097377090342586201462096257427696649920547479896269461227335795723058367584824127457535862548862037081102623167687214015839;
            5'd25: xpb[167] = 1024'd99366711426291873659868026489444011412353309188508274983180197077846710432855602625868635814359692722035733145870969164050839866327649388115458588241923068626940982721710982277066040171660349943833902791442341966827942166537883463857576820094468651947598319689584079011994330139662823414248838752460515748930;
            5'd26: xpb[167] = 1024'd78528040746518600326502962068058885319907756130901469156881033947965199782707998948900367004002545569028532590214309243697060692812511296729044906768333783185280487116665178100622633940223322797325219381422587676228187683155219447818884178961601508172138271794344030566452797730463609747395054337233817482021;
            5'd27: xpb[167] = 1024'd57689370066745326993137897646673759227462203073294663330581870818083689132560395271932098193645398416021332034557649323343281519297373205342631225294744497743619991511619373924179227708786295650816535971402833385628433199772555431780191537828734364396678223899103982120911265321264396080541269922007119215112;
            5'd28: xpb[167] = 1024'd36850699386972053659772833225288633135016650015687857504282707688202178482412791594963829383288251263014131478900989402989502345782235113956217543821155212301959495906573569747735821477349268504307852561383079095028678716389891415741498896695867220621218176003863933675369732912065182413687485506780420948203;
            5'd29: xpb[167] = 1024'd16012028707198780326407768803903507042571096958081051677983544558320667832265187917995560572931104110006930923244329482635723172267097022569803862347565926860299000301527765571292415245912241357799169151363324804428924233007227399702806255563000076845758128108623885229828200502865968746833701091553722681294;
            5'd30: xpb[167] = 1024'd119240053711550248391841631787332813694823971026209929979816236493416052519426723151042362977231631266442879775045162996861007839593179265738550305890307682352329179266053178732479248205992419932600683349730810360193530599845460156629092184113362382337117983627500894814393196167595388097098606502952618898716;
            5'd31: xpb[167] = 1024'd98401383031776975058476567365947687602378417968603124153517073363534541869279119474074094166874484113435679219388503076507228666078041174352136624416718396910668683661007374556035841974555392786091999939711056069593776116462796140590399542980495238561657935732260846368851663758396174430244822087725920631807;
        endcase
    end

    always_comb begin
        case(flag[56][5:0])
            6'd0: xpb[168] = 1024'd0;
            6'd1: xpb[168] = 1024'd38781356176001850862555751472281280754966432455498159163608955116826515609565757898552912678258668480214239331865921578076724746281451541482861471471564555734504094027980785189796217871559182819791658264845650889497010816540066062275853450923814047393098943918510398961655065674598480381695518836249611182449;
            6'd2: xpb[168] = 1024'd77562712352003701725111502944562561509932864910996318327217910233653031219131515797105825356517336960428478663731843156153449492562903082965722942943129111469008188055961570379592435743118365639583316529691301778994021633080132124551706901847628094786197887837020797923310131349196960763391037672499222364898;
            6'd3: xpb[168] = 1024'd116344068528005552587667254416843842264899297366494477490826865350479546828697273695658738034776005440642717995597764734230174238844354624448584414414693667203512282083942355569388653614677548459374974794536952668491032449620198186827560352771442142179296831755531196884965197023795441145086556508748833547347;
            6'd4: xpb[168] = 1024'd31058729019882662051424078484310690275167302696256952526303965402329167100953892684196579498376999611413807920006192877727835144284585831376285760869927182004325701542351923421554632294719525557856435450995363711623682415939367476138435234012026740305575872259924537816513734624465288509663385518372850245465;
            6'd5: xpb[168] = 1024'd69840085195884512913979829956591971030133735151755111689912920519155682710519650582749492176635668091628047251872114455804559890566037372859147232341491737738829795570332708611350850166278708377648093715841014601120693232479433538414288684935840787698674816178434936778168800299063768891358904354622461427914;
            6'd6: xpb[168] = 1024'd108621441371886363776535581428873251785100167607253270853521875635982198320085408481302404854894336571842286583738036033881284636847488914342008703813056293473333889598313493801147068037837891197439751980686665490617704049019499600690142135859654835091773760096945335739823865973662249273054423190872072610363;
            6'd7: xpb[168] = 1024'd23336101863763473240292405496340099795368172937015745888998975687831818592342027469840246318495330742613376508146464177378945542287720121269710050268289808274147309056723061653313046717879868295921212637145076533750354015338668890001017017100239433218052800601338676671372403574332096637631252200496089308481;
            6'd8: xpb[168] = 1024'd62117458039765324102848156968621380550334605392513905052607930804658334201907785368393158996753999222827615840012385755455670288569171662752571521739854364008651403084703846843109264589439051115712870901990727423247364831878734952276870468024053480611151744519849075633027469248930577019326771036745700490930;
            6'd9: xpb[168] = 1024'd100898814215767174965403908440902661305301037848012064216216885921484849811473543266946071675012667703041855171878307333532395034850623204235432993211418919743155497112684632032905482460998233935504529166836378312744375648418801014552723918947867528004250688438359474594682534923529057401022289872995311673379;
            6'd10: xpb[168] = 1024'd15613474707644284429160732508369509315569043177774539251693985973334470083730162255483913138613661873812945096286735477030055940290854411163134339666652434543968916571094199885071461141040211033985989823294789355877025614737970303863598800188452126130529728942752815526231072524198904765599118882619328371497;
            6'd11: xpb[168] = 1024'd54394830883646135291716483980650790070535475633272698415302941090160985693295920154036825816872330354027184428152657055106780686572305952645995811138216990278473010599074985074867679012599393853777648088140440245374036431278036366139452251112266173523628672861263214487886138198797385147294637718868939553946;
            6'd12: xpb[168] = 1024'd93176187059647986154272235452932070825501908088770857578911896206987501302861678052589738495130998834241423760018578633183505432853757494128857282609781546012977104627055770264663896884158576673569306352986091134871047247818102428415305702036080220916727616779773613449541203873395865528990156555118550736395;
            6'd13: xpb[168] = 1024'd7890847551525095618029059520398918835769913418533332614388996258837121575118297041127579958731993005012513684427006776681166338293988701056558629065015060813790524085465338116829875564200553772050767009444502178003697214137271717726180583276664819043006657284166954381089741474065712893566985564742567434513;
            6'd14: xpb[168] = 1024'd46672203727526946480584810992680199590736345874031491777997951375663637184684054939680492636990661485226753016292928354757891084575440242539420100536579616548294618113446123306626093435759736591842425274290153067500708030677337780002034034200478866436105601202677353342744807148664193275262504400992178616962;
            6'd15: xpb[168] = 1024'd85453559903528797343140562464961480345702778329529650941606906492490152794249812838233405315249329965440992348158849932834615830856891784022281572008144172282798712141426908496422311307318919411634083539135803956997718847217403842277887485124292913829204545121187752304399872823262673656958023237241789799411;
            6'd16: xpb[168] = 1024'd168220395405906806897386532428328355970783659292125977084006544339773066506431826771246778850324136212082272567278076332276736297122990949982918463377687083612131599836476348588289987360896510115544195594215000130368813536573131588762366364877511955483585625581093235948410423932521021534852246865806497529;
            6'd17: xpb[168] = 1024'd38949576571407757669453138004709609110937216114790285140692961661166288676072189725324159457108992616426321604433199654409001482578574532432844389934942242818116225627817261538384507858920079329907202460439865889627379630076639193864615817288691559348582529544091492197603476098531001403230371083115417679978;
            6'd18: xpb[168] = 1024'd77730932747409608532008889476990889865903648570288444304301916777992804285637947623877072135367661096640560936299121232485726228860026073915705861406506798552620319655798046728180725730479262149698860725285516779124390446616705256140469268212505606741681473462601891159258541773129481784925889919365028862427;
            6'd19: xpb[168] = 1024'd116512288923411459394564640949272170620870081025786603467910871894819319895203705522429984813626329576854800268165042810562450975141477615398567332878071354287124413683778831917976943602038444969490518990131167668621401263156771318416322719136319654134780417381112290120913607447727962166621408755614640044876;
            6'd20: xpb[168] = 1024'd31226949415288568858321465016739018631138086355549078503387971946668940167460324510967826277227323747625890192573470954060111880581708822326268679333304869087937833142188399770142922282080422067971979646589578711754051229475940607727197600376904252261059457885505631052462145048397809531198237765238656742994;
            6'd21: xpb[168] = 1024'd70008305591290419720877216489020299386104518811047237666996927063495455777026082409520738955485992227840129524439392532136836626863160363809130150804869424822441927170169184959939140153639604887763637911435229601251062046016006670003051051300718299654158401804016030014117210722996289912893756601488267925443;
            6'd22: xpb[168] = 1024'd108789661767292270583432967961301580141070951266545396830605882180321971386591840308073651633744660708054368856305314110213561373144611905291991622276433980556946021198149970149735358025198787707555296176280880490748072862556072732278904502224532347047257345722526428975772276397594770294589275437737879107892;
            6'd23: xpb[168] = 1024'd23504322259169380047189792028768428151338956596307871866082982232171591658848459296611493097345654878825458780713742253711222278584843112219692968731667495357759440656559538001901336705240764806036756832739291533880722828875242021589779383465116945173536386226919769907320813998264617659166104447361895806010;
            6'd24: xpb[168] = 1024'd62285678435171230909745543501049708906305389051806031029691937348998107268414217195164405775604323359039698112579663831787947024866294653702554440203232051092263534684540323191697554576799947625828415097584942423377733645415308083865632834388930992566635330145430168868975879672863098040861623283611506988459;
            6'd25: xpb[168] = 1024'd101067034611173081772301294973330989661271821507304190193300892465824622877979975093717318453862991839253937444445585409864671771147746195185415911674796606826767628712521108381493772448359130445620073362430593312874744461955374146141486285312745039959734274063940567830630945347461578422557142119861118170908;
            6'd26: xpb[168] = 1024'd15781695103050191236058119040797837671539826837066665228777992517674243150236594082255159917463986010025027368854013553362332676587977402113117258130030121627581048170930676233659751128401107544101534018889004356007394428274543435452361166553329638086013314568333908762179482948131425787133971129485134869026;
            6'd27: xpb[168] = 1024'd54563051279052042098613870513079118426506259292564824392386947634500758759802351980808072595722654490239266700719935131439057422869428943595978729601594677362085142198911461423455968999960290363893192283734655245504405244814609497728214617477143685479112258486844307723834548622729906168829489965734746051475;
            6'd28: xpb[168] = 1024'd93344407455053892961169621985360399181472691748062983555995902751327274369368109879360985273981322970453506032585856709515782169150880485078840201073159233096589236226892246613252186871519473183684850548580306135001416061354675560004068068400957732872211202405354706685489614297328386550525008801984357233924;
            6'd29: xpb[168] = 1024'd8059067946931002424926446052827247191740697077825458591473002803176894641624728867898826737582317141224595956994284853013443074591111692006541547528392747897402655685301814465418165551561450282166311205038717178134066027673844849314942949641542330998490242909748047617038151897998233915101837811608373932042;
            6'd30: xpb[168] = 1024'd46840424122932853287482197525108527946707129533323617755081957920003410251190486766451739415840985621438835288860206431090167820872563233489403018999957303631906749713282599655214383423120633101957969469884368067631076844213910911590796400565356378391589186828258446578693217572596714296797356647857985114491;
            6'd31: xpb[168] = 1024'd85621780298934704150037948997389808701673561988821776918690913036829925860756244665004652094099654101653074620726128009166892567154014774972264490471521859366410843741263384845010601294679815921749627734730018957128087660753976973866649851489170425784688130746768845540348283247195194678492875484107596296940;
            6'd32: xpb[168] = 1024'd336440790811813613794773064856656711941567318584251954168013088679546133012863653542493557700648272424164545134556152664553472594245981899965836926755374167224263199672952697176579974721793020231088391188430000260737627073146263177524732729755023910967171251162186471896820847865042043069704493731612995058;
            6'd33: xpb[168] = 1024'd39117796966813664476350524537137937466907999774082411117776968205506061742578621552095406235959316752638403877000477730741278218875697523382827308398319929901728357227653737886972797846280975840022746656034080889757748443613212325453378183653569071304066115169672585433551886522463522424765223329981224177507;
            6'd34: xpb[168] = 1024'd77899153142815515338906276009419218221874432229580570281385923322332577352144379450648318914217985232852643208866399308818002965157149064865688779869884485636232451255634523076769015717840158659814404920879731779254759260153278387729231634577383118697165059088182984395206952197062002806460742166230835359956;
            6'd35: xpb[168] = 1024'd116680509318817366201462027481700498976840864685078729444994878439159092961710137349201231592476653713066882540732320886894727711438600606348550251341449041370736545283615308266565233589399341479606063185725382668751770076693344450005085085501197166090264003006693383356862017871660483188156261002480446542405;
            6'd36: xpb[168] = 1024'd31395169810694475665218851549167346987108870014841204480471978491008713233966756337739073056077647883837972465140749030392388616878831813276251597796682556171549964742024876118731212269441318578087523842183793711884420043012513739315959966741781764216543043511086724288410555472330330552733090012104463240523;
            6'd37: xpb[168] = 1024'd70176525986696326527774603021448627742075302470339363644080933607835228843532514236291985734336316364052211797006670608469113363160283354759113069268247111906054058770005661308527430141000501397879182107029444601381430859552579801591813417665595811609641987429597123250065621146928810934428608848354074422972;
            6'd38: xpb[168] = 1024'd108957882162698177390330354493729908497041734925837522807689888724661744453098272134844898412594984844266451128872592186545838109441734896241974540739811667640558152797986446498323648012559684217670840371875095490878441676092645863867666868589409859002740931348107522211720686821527291316124127684603685605421;
            6'd39: xpb[168] = 1024'd23672542654575286854087178561196756507309740255599997843166988776511364725354891123382739876195979015037541053281020330043499014881966103169675887195045182441371572256396014350489626692601661316152301028333506534011091642411815153178541749829994457129019971852500863143269224422197138680700956694227702303539;
            6'd40: xpb[168] = 1024'd62453898830577137716642930033478037262276172711098157006775943893337880334920649021935652554454647495251780385146941908120223761163417644652537358666609738175875666284376799540285844564160844135943959293179157423508102458951881215454395200753808504522118915771011262104924290096795619062396475530477313485988;
            6'd41: xpb[168] = 1024'd101235255006578988579198681505759318017242605166596316170384899010164395944486406920488565232713315975466019717012863486196948507444869186135398830138174293910379760312357584730082062435720026955735617558024808313005113275491947277730248651677622551915217859689521661066579355771394099444091994366726924668437;
            6'd42: xpb[168] = 1024'd15949915498456098042955505573226166027510610496358791205861999062014016216743025909026406696314310146237109641421291629694609412885100393063100176593407808711193179770767152582248041115762004054217078214483219356137763241811116567041123532918207150041496900193915001998127893372063946808668823376350941366555;
            6'd43: xpb[168] = 1024'd54731271674457948905511257045507446782477042951856950369470954178840531826308783807579319374572978626451348973287213207771334159166551934545961648064972364445697273798747937772044258987321186874008736479328870245634774058351182629316976983842021197434595844112425400959782959046662427190364342212600552549004;
            6'd44: xpb[168] = 1024'd93512627850459799768067008517788727537443475407355109533079909295667047435874541706132232052831647106665588305153134785848058905448003476028823119536536920180201367826728722961840476858880369693800394744174521135131784874891248691592830434765835244827694788030935799921438024721260907572059861048850163731453;
            6'd45: xpb[168] = 1024'd8227288342336909231823832585255575547711480737117584568557009347516667708131160694670073516432641277436678229561562929345719810888234682956524465991770434981014787285138290814006455538922346792281855400632932178264434841210417980903705316006419842953973828535329140852986562321930754936636690058474180429571;
            6'd46: xpb[168] = 1024'd47008644518338760094379584057536856302677913192615743732165964464343183317696918593222986194691309757650917561427484507422444557169686224439385937463334990715518881313119076003802673410481529612073513665478583067761445657750484043179558766930233890347072772453839539814641627996529235318332208894723791612020;
            6'd47: xpb[168] = 1024'd85790000694340610956935335529818137057644345648113902895774919581169698927262676491775898872949978237865156893293406085499169303451137765922247408934899546450022975341099861193598891282040712431865171930324233957258456474290550105455412217854047937740171716372349938776296693671127715700027727730973402794469;
            6'd48: xpb[168] = 1024'd504661186217720420692159597284985067912350977876377931252019633019319199519295480313740336550972408636246817701834228996830208891368972849948755390133061250836394799509429045764869962082689530346632586782645000391106440609719394766287099094632535866450756876743279707845231271797563064604556740597419492587;
            6'd49: xpb[168] = 1024'd39286017362219571283247911069566265822878783433374537094860974749845834809085053378866653014809640888850486149567755807073554955172820514332810226861697616985340488827490214235561087833641872350138290851628295889888117257149785457042140550018446583259549700795253678669500296946396043446300075576847030675036;
            6'd50: xpb[168] = 1024'd78067373538221422145803662541847546577845215888872696258469929866672350418650811277419565693068309369064725481433677385150279701454272055815671698333262172719844582855470999425357305705201055169929949116473946779385128073689851519317994000942260630652648644713764077631155362620994523827995594413096641857485;
            6'd51: xpb[168] = 1024'd116848729714223273008359414014128827332811648344370855422078884983498866028216569175972478371326977849278964813299598963227004447735723597298533169804826728454348676883451784615153523576760237989721607381319597668882138890229917581593847451866074678045747588632274476592810428295593004209691113249346253039934;
            6'd52: xpb[168] = 1024'd31563390206100382472116238081595675343079653674133330457555985035348486300473188164510319834927972020050054737708027106724665353175954804226234516260060243255162096341861352467319502256802215088203068037778008712014788856549086870904722333106659276172026629136667817524358965896262851574267942258970269738052;
            6'd53: xpb[168] = 1024'd70344746382102233334671989553876956098046086129631489621164940152175001910038946063063232513186640500264294069573948684801390099457406345709095987731624798989666190369842137657115720128361397907994726302623659601511799673089152933180575784030473323565125573055178216486014031570861331955963461095219880920501;
            6'd54: xpb[168] = 1024'd109126102558104084197227741026158236853012518585129648784773895269001517519604703961616145191445308980478533401439870262878114845738857887191957459203189354724170284397822922846911937999920580727786384567469310491008810489629218995456429234954287370958224516973688615447669097245459812337658979931469492102950;
            6'd55: xpb[168] = 1024'd23840763049981193660984565093625084863280523914892123820250995320851137791861322950153986655046303151249623325848298406375775751179089094119658805658422869524983703856232490699077916679962557826267845223927721534141460455948388284767304116194871969084503557478081956379217634846129659702235808941093508801068;
            6'd56: xpb[168] = 1024'd62622119225983044523540316565906365618246956370390282983859950437677653401427080848706899333304971631463862657714219984452500497460540635602520277129987425259487797884213275888874134551521740646059503488773372423638471272488454347043157567118686016477602501396592355340872700520728140083931327777343119983517;
            6'd57: xpb[168] = 1024'd101403475401984895386096068038187646373213388825888442147468905554504169010992838747259812011563640111678101989580141562529225243741992177085381748601551980993991891912194061078670352423080923465851161753619023313135482089028520409319011018042500063870701445315102754302527766195326620465626846613592731165966;
            6'd58: xpb[168] = 1024'd16118135893862004849852892105654494383481394155650917182946005606353789283249457735797653475164634282449191913988569706026886149182223384013083095056785495794805311370603628930836331103122900564332622410077434356268132055347689698629885899283084661996980485819496095234076303795996467830203675623216747864084;
            6'd59: xpb[168] = 1024'd54899492069863855712408643577935775138447826611149076346554960723180304892815215634350566153423302762663431245854491284103610895463674925495944566528350051529309405398584414120632548974682083384124280674923085245765142871887755760905739350206898709390079429738006494195731369470594948211899194459466359046533;
            6'd60: xpb[168] = 1024'd93680848245865706574964395050217055893414259066647235510163915840006820502380973532903478831681971242877670577720412862180335641745126466978806037999914607263813499426565199310428766846241266203915938939768736135262153688427821823181592801130712756783178373656516893157386435145193428593594713295715970228982;
            6'd61: xpb[168] = 1024'd8395508737742816038721219117683903903682264396409710545641015891856440774637592521441320295282965413648760502128841005677996547185357673906507384455148122064626918884974767162594745526283243302397399596227147178394803654746991112492467682371297354909457414160910234088934972745863275958171542305339986927100;
            6'd62: xpb[168] = 1024'd47176864913744666901276970589965184658648696851907869709249971008682956384203350419994232973541633893862999833994762583754721293466809215389368855926712677799131012912955552352390963397842426122189057861072798067891814471287057174768321133295111402302556358079420633050590038420461756339867061141589598109549;
            6'd63: xpb[168] = 1024'd85958221089746517763832722062246465413615129307406028872858926125509471993769108318547145651800302374077239165860684161831446039748260756872230327398277233533635106940936337542187181269401608941980716125918448957388825287827123237044174584218925449695655301997931032012245104095060236721562579977839209291998;
        endcase
    end

    always_comb begin
        case(flag[56][11:6])
            6'd0: xpb[169] = 1024'd0;
            6'd1: xpb[169] = 1024'd672881581623627227589546129713313423883134637168503908336026177359092266025727307084987115401296544848329090269112305329106945188491963799931673853510748334448526399345905394353159949443586040462176782376860000521475254146292526355049465459510047821934342502324372943793641695730084086139408987463225990116;
            6'd2: xpb[169] = 1024'd1345763163247254455179092259426626847766269274337007816672052354718184532051454614169974230802593089696658180538224610658213890376983927599863347707021496668897052798691810788706319898887172080924353564753720001042950508292585052710098930919020095643868685004648745887587283391460168172278817974926451980232;
            6'd3: xpb[169] = 1024'd2018644744870881682768638389139940271649403911505511725008078532077276798077181921254961346203889634544987270807336915987320835565475891399795021560532245003345579198037716183059479848330758121386530347130580001564425762438877579065148396378530143465803027506973118831380925087190252258418226962389677970348;
            6'd4: xpb[169] = 1024'd2691526326494508910358184518853253695532538548674015633344104709436369064102909228339948461605186179393316361076449221316427780753967855199726695414042993337794105597383621577412639797774344161848707129507440002085901016585170105420197861838040191287737370009297491775174566782920336344557635949852903960464;
            6'd5: xpb[169] = 1024'd3364407908118136137947730648566567119415673185842519541680130886795461330128636535424935577006482724241645451345561526645534725942459818999658369267553741672242631996729526971765799747217930202310883911884300002607376270731462631775247327297550239109671712511621864718968208478650420430697044937316129950580;
            6'd6: xpb[169] = 1024'd4037289489741763365537276778279880543298807823011023450016157064154553596154363842509922692407779269089974541614673831974641671130951782799590043121064490006691158396075432366118959696661516242773060694261160003128851524877755158130296792757060286931606055013946237662761850174380504516836453924779355940696;
            6'd7: xpb[169] = 1024'd4710171071365390593126822907993193967181942460179527358352183241513645862180091149594909807809075813938303631883786137303748616319443746599521716974575238341139684795421337760472119646105102283235237476638020003650326779024047684485346258216570334753540397516270610606555491870110588602975862912242581930812;
            6'd8: xpb[169] = 1024'd5383052652989017820716369037706507391065077097348031266688209418872738128205818456679896923210372358786632722152898442632855561507935710399453390828085986675588211194767243154825279595548688323697414259014880004171802033170340210840395723676080382575474740018594983550349133565840672689115271899705807920928;
            6'd9: xpb[169] = 1024'd6055934234612645048305915167419820814948211734516535175024235596231830394231545763764884038611668903634961812422010747961962506696427674199385064681596735010036737594113148549178439544992274364159591041391740004693277287316632737195445189135590430397409082520919356494142775261570756775254680887169033911044;
            6'd10: xpb[169] = 1024'd6728815816236272275895461297133134238831346371685039083360261773590922660257273070849871154012965448483290902691123053291069451884919637999316738535107483344485263993459053943531599494435860404621767823768600005214752541462925263550494654595100478219343425023243729437936416957300840861394089874632259901160;
            6'd11: xpb[169] = 1024'd7401697397859899503485007426846447662714481008853542991696287950950014926283000377934858269414261993331619992960235358620176397073411601799248412388618231678933790392804959337884759443879446445083944606145460005736227795609217789905544120054610526041277767525568102381730058653030924947533498862095485891276;
            6'd12: xpb[169] = 1024'd8074578979483526731074553556559761086597615646022046900032314128309107192308727685019845384815558538179949083229347663949283342261903565599180086242128980013382316792150864732237919393323032485546121388522320006257703049755510316260593585514120573863212110027892475325523700348761009033672907849558711881392;
            6'd13: xpb[169] = 1024'd8747460561107153958664099686273074510480750283190550808368340305668199458334454992104832500216855083028278173498459969278390287450395529399111760095639728347830843191496770126591079342766618526008298170899180006779178303901802842615643050973630621685146452530216848269317342044491093119812316837021937871508;
            6'd14: xpb[169] = 1024'd9420342142730781186253645815986387934363884920359054716704366483027291724360182299189819615618151627876607263767572274607497232638887493199043433949150476682279369590842675520944239292210204566470474953276040007300653558048095368970692516433140669507080795032541221213110983740221177205951725824485163861624;
            6'd15: xpb[169] = 1024'd10093223724354408413843191945699701358247019557527558625040392660386383990385909606274806731019448172724936354036684579936604177827379456998975107802661225016727895990188580915297399241653790606932651735652900007822128812194387895325741981892650717329015137534865594156904625435951261292091134811948389851740;
            6'd16: xpb[169] = 1024'd10766105305978035641432738075413014782130154194696062533376418837745476256411636913359793846420744717573265444305796885265711123015871420798906781656171973351176422389534486309650559191097376647394828518029760008343604066340680421680791447352160765150949480037189967100698267131681345378230543799411615841856;
            6'd17: xpb[169] = 1024'd11438986887601662869022284205126328206013288831864566441712445015104568522437364220444780961822041262421594534574909190594818068204363384598838455509682721685624948788880391704003719140540962687857005300406620008865079320486972948035840912811670812972883822539514340044491908827411429464369952786874841831972;
            6'd18: xpb[169] = 1024'd12111868469225290096611830334839641629896423469033070350048471192463660788463091527529768077223337807269923624844021495923925013392855348398770129363193470020073475188226297098356879089984548728319182082783480009386554574633265474390890378271180860794818165041838712988285550523141513550509361774338067822088;
            6'd19: xpb[169] = 1024'd12784750050848917324201376464552955053779558106201574258384497369822753054488818834614755192624634352118252715113133801253031958581347312198701803216704218354522001587572202492710039039428134768781358865160340009908029828779558000745939843730690908616752507544163085932079192218871597636648770761801293812204;
            6'd20: xpb[169] = 1024'd13457631632472544551790922594266268477662692743370078166720523547181845320514546141699742308025930896966581805382246106582138903769839275998633477070214966688970527986918107887063198988871720809243535647537200010429505082925850527100989309190200956438686850046487458875872833914601681722788179749264519802320;
            6'd21: xpb[169] = 1024'd14130513214096171779380468723979581901545827380538582075056549724540937586540273448784729423427227441814910895651358411911245848958331239798565150923725715023419054386264013281416358938315306849705712429914060010950980337072143053456038774649711004260621192548811831819666475610331765808927588736727745792436;
            6'd22: xpb[169] = 1024'd14803394795719799006970014853692895325428962017707085983392575901900029852566000755869716538828523986663239985920470717240352794146823203598496824777236463357867580785609918675769518887758892890167889212290920011472455591218435579811088240109221052082555535051136204763460117306061849895066997724190971782552;
            6'd23: xpb[169] = 1024'd15476276377343426234559560983406208749312096654875589891728602079259122118591728062954703654229820531511569076189583022569459739335315167398428498630747211692316107184955824070122678837202478930630065994667780011993930845364728106166137705568731099904489877553460577707253759001791933981206406711654197772668;
            6'd24: xpb[169] = 1024'd16149157958967053462149107113119522173195231292044093800064628256618214384617455370039690769631117076359898166458695327898566684523807131198360172484257960026764633584301729464475838786646064971092242777044640012515406099511020632521187171028241147726424220055784950651047400697522018067345815699117423762784;
            6'd25: xpb[169] = 1024'd16822039540590680689738653242832835597078365929212597708400654433977306650643182677124677885032413621208227256727807633227673629712299094998291846337768708361213159983647634858828998736089651011554419559421500013036881353657313158876236636487751195548358562558109323594841042393252102153485224686580649752900;
            6'd26: xpb[169] = 1024'd17494921122214307917328199372546149020961500566381101616736680611336398916668909984209665000433710166056556346996919938556780574900791058798223520191279456695661686382993540253182158685533237052016596341798360013558356607803605685231286101947261243370292905060433696538634684088982186239624633674043875743016;
            6'd27: xpb[169] = 1024'd18167802703837935144917745502259462444844635203549605525072706788695491182694637291294652115835006710904885437266032243885887520089283022598155194044790205030110212782339445647535318634976823092478773124175220014079831861949898211586335567406771291192227247562758069482428325784712270325764042661507101733132;
            6'd28: xpb[169] = 1024'd18840684285461562372507291631972775868727769840718109433408732966054583448720364598379639231236303255753214527535144549214994465277774986398086867898300953364558739181685351041888478584420409132940949906552080014601307116096190737941385032866281339014161590065082442426221967480442354411903451648970327723248;
            6'd29: xpb[169] = 1024'd19513565867085189600096837761686089292610904477886613341744759143413675714746091905464626346637599800601543617804256854544101410466266950198018541751811701699007265581031256436241638533863995173403126688928940015122782370242483264296434498325791386836095932567406815370015609176172438498042860636433553713364;
            6'd30: xpb[169] = 1024'd20186447448708816827686383891399402716494039115055117250080785320772767980771819212549613462038896345449872708073369159873208355654758913997950215605322450033455791980377161830594798483307581213865303471305800015644257624388775790651483963785301434658030275069731188313809250871902522584182269623896779703480;
            6'd31: xpb[169] = 1024'd20859329030332444055275930021112716140377173752223621158416811498131860246797546519634600577440192890298201798342481465202315300843250877797881889458833198367904318379723067224947958432751167254327480253682660016165732878535068317006533429244811482479964617572055561257602892567632606670321678611360005693596;
            6'd32: xpb[169] = 1024'd21532210611956071282865476150826029564260308389392125066752837675490952512823273826719587692841489435146530888611593770531422246031742841597813563312343946702352844779068972619301118382194753294789657036059520016687208132681360843361582894704321530301898960074379934201396534263362690756461087598823231683712;
            6'd33: xpb[169] = 1024'd22205092193579698510455022280539342988143443026560628975088863852850044778849001133804574808242785979994859978880706075860529191220234805397745237165854695036801371178414878013654278331638339335251833818436380017208683386827653369716632360163831578123833302576704307145190175959092774842600496586286457673828;
            6'd34: xpb[169] = 1024'd22877973775203325738044568410252656412026577663729132883424890030209137044874728440889561923644082524843189069149818381189636136408726769197676911019365443371249897577760783408007438281081925375714010600813240017730158640973945896071681825623341625945767645079028680088983817654822858928739905573749683663944;
            6'd35: xpb[169] = 1024'd23550855356826952965634114539965969835909712300897636791760916207568229310900455747974549039045379069691518159418930686518743081597218732997608584872876191705698423977106688802360598230525511416176187383190100018251633895120238422426731291082851673767701987581353053032777459350552943014879314561212909654060;
            6'd36: xpb[169] = 1024'd24223736938450580193223660669679283259792846938066140700096942384927321576926183055059536154446675614539847249688042991847850026785710696797540258726386940040146950376452594196713758179969097456638364165566960018773109149266530948781780756542361721589636330083677425976571101046283027101018723548676135644176;
            6'd37: xpb[169] = 1024'd24896618520074207420813206799392596683675981575234644608432968562286413842951910362144523269847972159388176339957155297176956971974202660597471932579897688374595476775798499591066918129412683497100540947943820019294584403412823475136830222001871769411570672586001798920364742742013111187158132536139361634292;
            6'd38: xpb[169] = 1024'd25569500101697834648402752929105910107559116212403148516768994739645506108977637669229510385249268704236505430226267602506063917162694624397403606433408436709044003175144404985420078078856269537562717730320680019816059657559116001491879687461381817233505015088326171864158384437743195273297541523602587624408;
            6'd39: xpb[169] = 1024'd26242381683321461875992299058819223531442250849571652425105020917004598375003364976314497500650565249084834520495379907835170862351186588197335280286919185043492529574490310379773238028299855578024894512697540020337534911705408527846929152920891865055439357590650544807952026133473279359436950511065813614524;
            6'd40: xpb[169] = 1024'd26915263264945089103581845188532536955325385486740156333441047094363690641029092283399484616051861793933163610764492213164277807539678551997266954140429933377941055973836215774126397977743441618487071295074400020859010165851701054201978618380401912877373700092974917751745667829203363445576359498529039604640;
            6'd41: xpb[169] = 1024'd27588144846568716331171391318245850379208520123908660241777073271722782907054819590484471731453158338781492701033604518493384752728170515797198627993940681712389582373182121168479557927187027658949248077451260021380485419997993580557028083839911960699308042595299290695539309524933447531715768485992265594756;
            6'd42: xpb[169] = 1024'd28261026428192343558760937447959163803091654761077164150113099449081875173080546897569458846854454883629821791302716823822491697916662479597130301847451430046838108772528026562832717876630613699411424859828120021901960674144286106912077549299422008521242385097623663639332951220663531617855177473455491584872;
            6'd43: xpb[169] = 1024'd28933908009815970786350483577672477226974789398245668058449125626440967439106274204654445962255751428478150881571829129151598643105154443397061975700962178381286635171873931957185877826074199739873601642204980022423435928290578633267127014758932056343176727599948036583126592916393615703994586460918717574988;
            6'd44: xpb[169] = 1024'd29606789591439598013940029707385790650857924035414171966785151803800059705132001511739433077657047973326479971840941434480705588293646407196993649554472926715735161571219837351539037775517785780335778424581840022944911182436871159622176480218442104165111070102272409526920234612123699790133995448381943565104;
            6'd45: xpb[169] = 1024'd30279671173063225241529575837099104074741058672582675875121177981159151971157728818824420193058344518174809062110053739809812533482138370996925323407983675050183687970565742745892197724961371820797955206958700023466386436583163685977225945677952151987045412604596782470713876307853783876273404435845169555220;
            6'd46: xpb[169] = 1024'd30952552754686852469119121966812417498624193309751179783457204158518244237183456125909407308459641063023138152379166045138919478670630334796856997261494423384632214369911648140245357674404957861260131989335560023987861690729456212332275411137462199808979755106921155414507518003583867962412813423308395545336;
            6'd47: xpb[169] = 1024'd31625434336310479696708668096525730922507327946919683691793230335877336503209183432994394423860937607871467242648278350468026423859122298596788671115005171719080740769257553534598517623848543901722308771712420024509336944875748738687324876596972247630914097609245528358301159699313952048552222410771621535452;
            6'd48: xpb[169] = 1024'd32298315917934106924298214226239044346390462584088187600129256513236428769234910740079381539262234152719796332917390655797133369047614262396720344968515920053529267168603458928951677573292129942184485554089280025030812199022041265042374342056482295452848440111569901302094801395044036134691631398234847525568;
            6'd49: xpb[169] = 1024'd32971197499557734151887760355952357770273597221256691508465282690595521035260638047164368654663530697568125423186502961126240314236106226196652018822026668387977793567949364323304837522735715982646662336466140025552287453168333791397423807515992343274782782613894274245888443090774120220831040385698073515684;
            6'd50: xpb[169] = 1024'd33644079081181361379477306485665671194156731858425195416801308867954613301286365354249355770064827242416454513455615266455347259424598189996583692675537416722426319967295269717657997472179302023108839118843000026073762707314626317752473272975502391096717125116218647189682084786504204306970449373161299505800;
            6'd51: xpb[169] = 1024'd34316960662804988607066852615378984618039866495593699325137335045313705567312092661334342885466123787264783603724727571784454204613090153796515366529048165056874846366641175112011157421622888063571015901219860026595237961460918844107522738435012438918651467618543020133475726482234288393109858360624525495916;
            6'd52: xpb[169] = 1024'd34989842244428615834656398745092298041923001132762203233473361222672797833337819968419330000867420332113112693993839877113561149801582117596447040382558913391323372765987080506364317371066474104033192683596720027116713215607211370462572203894522486740585810120867393077269368177964372479249267348087751486032;
            6'd53: xpb[169] = 1024'd35662723826052243062245944874805611465806135769930707141809387400031890099363547275504317116268716876961441784262952182442668094990074081396378714236069661725771899165332985900717477320510060144495369465973580027638188469753503896817621669354032534562520152623191766021063009873694456565388676335550977476148;
            6'd54: xpb[169] = 1024'd36335605407675870289835491004518924889689270407099211050145413577390982365389274582589304231670013421809770874532064487771775040178566045196310388089580410060220425564678891295070637269953646184957546248350440028159663723899796423172671134813542582384454495125516138964856651569424540651528085323014203466264;
            6'd55: xpb[169] = 1024'd37008486989299497517425037134232238313572405044267714958481439754750074631415001889674291347071309966658099964801176793100881985367058008996242061943091158394668951964024796689423797219397232225419723030727300028681138978046088949527720600273052630206388837627840511908650293265154624737667494310477429456380;
            6'd56: xpb[169] = 1024'd37681368570923124745014583263945551737455539681436218866817465932109166897440729196759278462472606511506429055070289098429988930555549972796173735796601906729117478363370702083776957168840818265881899813104160029202614232192381475882770065732562678028323180130164884852443934960884708823806903297940655446496;
            6'd57: xpb[169] = 1024'd38354250152546751972604129393658865161338674318604722775153492109468259163466456503844265577873903056354758145339401403759095875744041936596105409650112655063566004762716607478130117118284404306344076595481020029724089486338674002237819531192072725850257522632489257796237576656614792909946312285403881436612;
            6'd58: xpb[169] = 1024'd39027131734170379200193675523372178585221808955773226683489518286827351429492183810929252693275199601203087235608513709088202820932533900396037083503623403398014531162062512872483277067727990346806253377857880030245564740484966528592868996651582773672191865134813630740031218352344876996085721272867107426728;
            6'd59: xpb[169] = 1024'd39700013315794006427783221653085492009104943592941730591825544464186443695517911118014239808676496146051416325877626014417309766121025864195968757357134151732463057561408418266836437017171576387268430160234740030767039994631259054947918462111092821494126207637138003683824860048074961082225130260330333416844;
            6'd60: xpb[169] = 1024'd40372894897417633655372767782798805432988078230110234500161570641545535961543638425099226924077792690899745416146738319746416711309517827995900431210644900066911583960754323661189596966615162427730606942611600031288515248777551581302967927570602869316060550139462376627618501743805045168364539247793559406960;
            6'd61: xpb[169] = 1024'd41045776479041260882962313912512118856871212867278738408497596818904628227569365732184214039479089235748074506415850625075523656498009791795832105064155648401360110360100229055542756916058748468192783724988460031809990502923844107658017393030112917137994892641786749571412143439535129254503948235256785397076;
            6'd62: xpb[169] = 1024'd41718658060664888110551860042225432280754347504447242316833622996263720493595093039269201154880385780596403596684962930404630601686501755595763778917666396735808636759446134449895916865502334508654960507365320032331465757070136634013066858489622964959929235144111122515205785135265213340643357222720011387192;
            6'd63: xpb[169] = 1024'd42391539642288515338141406171938745704637482141615746225169649173622812759620820346354188270281682325444732686954075235733737546874993719395695452771177145070257163158792039844249076814945920549117137289742180032852941011216429160368116323949133012781863577646435495458999426830995297426782766210183237377308;
        endcase
    end

    always_comb begin
        case(flag[56][16:12])
            5'd0: xpb[170] = 1024'd0;
            5'd1: xpb[170] = 1024'd43064421223912142565730952301652059128520616778784250133505675350981905025646547653439175385682978870293061777223187541062844492063485683195627126624687893404705689558137945238602236764389506589579314072119040033374416265362721686723165789408643060603797920148759868402793068526725381512922175197646463367424;
            5'd2: xpb[170] = 1024'd86128842447824285131461904603304118257041233557568500267011350701963810051293095306878350771365957740586123554446375082125688984126971366391254253249375786809411379116275890477204473528779013179158628144238080066748832530725443373446331578817286121207595840297519736805586137053450763025844350395292926734848;
            5'd3: xpb[170] = 1024'd5126567987611686298393929500141744640863423210617066272385170987968819739630504050302454942391262301436035924212069188609469635349236715031721254857732639280426394104842618378176471101651314047427744607969880253758887945867268287204518798542699732544573857032162547178272677506247511521647835766313795617941;
            5'd4: xpb[170] = 1024'd48190989211523828864124881801793803769384039989401316405890846338950724765277051703741630328074241171729097701435256729672314127412722398227348381482420532685132083662980563616778707866040820637007058680088920287133304211229989973927684587951342793148371777180922415581065746032972893034570010963960258985365;
            5'd5: xpb[170] = 1024'd91255410435435971429855834103445862897904656768185566539396521689932629790923599357180805713757220042022159478658444270735158619476208081422975508107108426089837773221118508855380944630430327226586372752207960320507720476592711660650850377359985853752169697329682283983858814559698274547492186161606722352789;
            5'd6: xpb[170] = 1024'd10253135975223372596787859000283489281726846421234132544770341975937639479261008100604909884782524602872071848424138377218939270698473430063442509715465278560852788209685236756352942203302628094855489215939760507517775891734536574409037597085399465089147714064325094356545355012495023043295671532627591235882;
            5'd7: xpb[170] = 1024'd53317557199135515162518811301935548410247463200018382678276017326919544504907555754044085270465503473165133625647325918281783762761959113259069636340153171965558477767823181994955178967692134684434803288058800540892192157097258261132203386494042525692945634213084962759338423539220404556217846730274054603306;
            5'd8: xpb[170] = 1024'd96381978423047657728249763603587607538768079978802632811781692677901449530554103407483260656148482343458195402870513459344628254825444796454696762964841065370264167325961127233557415732081641274014117360177840574266608422459979947855369175902685586296743554361844831162131492065945786069140021927920517970730;
            5'd9: xpb[170] = 1024'd15379703962835058895181788500425233922590269631851198817155512963906459218891512150907364827173786904308107772636207565828408906047710145095163764573197917841279182314527855134529413304953942142283233823909640761276663837601804861613556395628099197633721571096487641534818032518742534564943507298941386853823;
            5'd10: xpb[170] = 1024'd58444125186747201460912740802077293051110886410635448950661188314888364244538059804346540212856765774601169549859395106891253398111195828290790891197885811245984871872665800373131650069343448731862547896028680794651080102964526548336722185036742258237519491245247509937611101045467916077865682496587850221247;
            5'd11: xpb[170] = 1024'd101508546410659344026643693103729352179631503189419699084166863665870269270184607457785715598539744644894231327082582647954097890174681511486418017822573704650690561430803745611733886833732955321441861968147720828025496368327248235059887974445385318841317411394007378340404169572193297590787857694234313588671;
            5'd12: xpb[170] = 1024'd20506271950446745193575718000566978563453692842468265089540683951875278958522016201209819769565049205744143696848276754437878541396946860126885019430930557121705576419370473512705884406605256189710978431879521015035551783469073148818075194170798930178295428128650188713090710024990046086591343065255182471764;
            5'd13: xpb[170] = 1024'd63570693174358887759306670302219037691974309621252515223046359302857183984168563854648995155248028076037205474071464295500723033460432543322512146055618450526411265977508418751308121170994762779290292503998561048409968048831794835541240983579441990782093348277410057115883778551715427599513518262901645839188;
            5'd14: xpb[170] = 1024'd106635114398271030325037622603871096820494926400036765356552034653839089009815111508088170540931006946330267251294651836563567525523918226518139272680306343931116955535646363989910357935384269368869606576117601081784384314194516522264406772988085051385891268426169925518676847078440809112435693460548109206612;
            5'd15: xpb[170] = 1024'd25632839938058431491969647500708723204317116053085331361925854939844098698152520251512274711956311507180179621060345943047348176746183575158606274288663196402131970524213091890882355508256570237138723039849401268794439729336341436022593992713498662722869285160812735891363387531237557608239178831568978089705;
            5'd16: xpb[170] = 1024'd68697261161970574057700599802360782332837732831869581495431530290826003723799067904951450097639290377473241398283533484110192668809669258354233400913351089806837660082351037129484592272646076826718037111968441302168855994699063122745759782122141723326667205309572604294156456057962939121161354029215441457129;
            5'd17: xpb[170] = 1024'd111761682385882716623431552104012841461358349610653831628937205641807908749445615558390625483322269247766303175506721025173037160873154941549860527538038983211543349640488982368086829037035583416297351184087481335543272260061784809468925571530784783930465125458332472696949524584688320634083529226861904824553;
            5'd18: xpb[170] = 1024'd30759407925670117790363577000850467845180539263702397634311025927812918437783024301814729654347573808616215545272415131656817812095420290190327529146395835682558364629055710269058826609907884284566467647819281522553327675203609723227112791256198395267443142192975283069636065037485069129887014597882773707646;
            5'd19: xpb[170] = 1024'd73823829149582260356094529302502526973701156042486647767816701278794823463429571955253905040030552678909277322495602672719662304158905973385954655771083729087264054187193655507661063374297390874145781719938321555927743940566331409950278580664841455871241062341735151472429133564210450642809189795529237075070;
            5'd20: xpb[170] = 1024'd116888250373494402921825481604154586102221772821270897901322376629776728489076119608693080425713531549202339099718790213782506796222391656581581782395771622491969743745331600746263300138686897463725095792057361589302160205929053096673444370073484516475038982490495019875222202090935832155731364993175700442494;
            5'd21: xpb[170] = 1024'd35885975913281804088757506500992212486043962474319463906696196915781738177413528352117184596738836110052251469484484320266287447444657005222048784004128474962984758733898328647235297711559198331994212255789161776312215621070878010431631589798898127812016999225137830247908742543732580651534850364196569325587;
            5'd22: xpb[170] = 1024'd78950397137193946654488458802644271614564579253103714040201872266763643203060076005556359982421814980345313246707671861329131939508142688417675910628816368367690448292036273885837534475948704921573526327908201809686631886433599697154797379207541188415814919373897698650701811070457962164457025561843032693011;
            5'd23: xpb[170] = 1024'd122014818361106089220219411104296330743085196031887964173707547617745548228706623658995535368104793850638375023930859402391976431571628371613303037253504261772396137850174219124439771240338211511152840400027241843061048151796321383877963168616184249019612839522657567053494879597183343677379200759489496060435;
            5'd24: xpb[170] = 1024'd41012543900893490387151436001133957126907385684936530179081367903750557917044032402419639539130098411488287393696553508875757082793893720253770038861861114243411152838740947025411768813210512379421956863759042030071103566938146297636150388341597860356590856257300377426181420049980092173182686130510364943528;
            5'd25: xpb[170] = 1024'd84076965124805632952882388302786016255428002463720780312587043254732462942690580055858814924813077281781349170919741049938601574857379403449397165486549007648116842396878892264014005577600018969001270935878082063445519832300867984359316177750240920960388776406060245828974488576705473686104861328156828310952;
            5'd26: xpb[170] = 1024'd3074690664593034119814413199623642639250192116769346317960863540737472631027988799282919095838381842631261540685435156422382226079644752089864167094905860119131857385445620164986003150472319837270387399609882250455575247442692898117503397475654532297366793140703056201661029029502222181908346699177697194045;
            5'd27: xpb[170] = 1024'd46139111888505176685545365501275701767770808895553596451466538891719377656674536452722094481521360712924323317908622697485226718143130435285491293719593753523837546943583565403588239914861826426849701471728922283829991512805414584840669186884297592901164713289462924604454097556227603694830521896824160561469;
            5'd28: xpb[170] = 1024'd89203533112417319251276317802927760896291425674337846584972214242701282682321084106161269867204339583217385095131810238548071210206616118481118420344281646928543236501721510642190476679251333016429015543847962317204407778168136271563834976292940653504962633438222793007247166082952985207752697094470623928893;
            5'd29: xpb[170] = 1024'd8201258652204720418208342699765387280113615327386412590346034528706292370658492849585374038229644144067297464897504345031851861428881467121585421952638499399558251490288238543162474252123633884698132007579762504214463193309961185322022196018354264841940650172865603379933706535749733703556182465491492811986;
            5'd30: xpb[170] = 1024'd51265679876116862983939295001417446408634232106170662723851709879688197396305040503024549423912623014360359242120691886094696353492367150317212548577326392804263941048426183781764711016513140474277446079698802537588879458672682872045187985426997325445738570321625471782726775062475115216478357663137956179410;
            5'd31: xpb[170] = 1024'd94330101100029005549670247303069505537154848884954912857357385230670102421951588156463724809595601884653421019343879427157540845555852833512839675202014286208969630606564129020366947780902647063856760151817842570963295724035404558768353774835640386049536490470385340185519843589200496729400532860784419546834;
        endcase
    end

    always_comb begin
        case(flag[57][5:0])
            6'd0: xpb[171] = 1024'd0;
            6'd1: xpb[171] = 1024'd68697261161970574057700599802360782332837732831869581495431530290826003723799067904951450097639290377473241398283533484110192668809669258354233400913351089806837660082351037129484592272646076826718037111968441302168855994699063122745759782122141723326667205309572604294156456057962939121161354029215441457129;
            6'd2: xpb[171] = 1024'd13327826639816406716602272199907131920977038538003478862731205516675112110288996899887828980620906445503333389109573533641321496778118182153306676810371138679984645595130856921338945353774947932125876615549642757973351139177229472526540994561053997386514507205028150558206384041997245225204018231805288429927;
            6'd3: xpb[171] = 1024'd82025087801786980774302872002267914253814771369873060358162735807501115834088064804839279078260196822976574787393107017751514165587787440507540077723722228486822305677481894050823537626421024758843913727518084060142207133876292595272300776683195720713181712514600754852362840099960184346365372261020729887056;
            6'd4: xpb[171] = 1024'd26655653279632813433204544399814263841954077076006957725462411033350224220577993799775657961241812891006666778219147067282642993556236364306613353620742277359969291190261713842677890707549895864251753231099285515946702278354458945053081989122107994773029014410056301116412768083994490450408036463610576859854;
            6'd5: xpb[171] = 1024'd95352914441603387490905144202175046174791809907876539220893941324176227944377061704727108058881103268479908176502680551392835662365905622660846754534093367166806951272612750972162482980195972690969790343067726818115558273053522067798841771244249718099696219719628905410569224141957429571569390492826018316983;
            6'd6: xpb[171] = 1024'd39983479919449220149806816599721395762931115614010436588193616550025336330866990699663486941862719336510000167328720600923964490334354546459920030431113416039953936785392570764016836061324843796377629846648928273920053417531688417579622983683161992159543521615084451674619152125991735675612054695415865289781;
            6'd7: xpb[171] = 1024'd108680741081419794207507416402082178095768848445880018083625146840851340054666058604614937039502009713983241565612254085034157159144023804814153431344464505846791596867743607893501428333970920623095666958617369576088909412230751540325382765805303715486210726924657055968775608183954674796773408724631306746910;
            6'd8: xpb[171] = 1024'd53311306559265626866409088799628527683908154152013915450924822066700448441155987599551315922483625782013333556438294134565285987112472728613226707241484554719938582380523427685355781415099791728503506462198571031893404556708917890106163978244215989546058028820112602232825536167988980900816072927221153719708;
            6'd9: xpb[171] = 1024'd122008567721236200924109688601989310016745886983883496946356352357526452164955055504502766020122916159486574954721827618675478655922141986967460108154835644526776242462874464814840373687745868555221543574167012334062260551407981012851923760366357712872725234129685206526981992225951920021977426956436595176837;
            6'd10: xpb[171] = 1024'd66639133199082033583011360999535659604885192690017394313656027583375560551444984499439144903104532227516666945547867668206607483890590910766533384051855693399923227975654284606694726768874739660629383077748213789866755695886147362632704972805269986932572536025140752791031920209986226126020091159026442149635;
            6'd11: xpb[171] = 1024'd11269698676927866241913033397082009193024498396151291680955702809224668937934913494375523786086148295546758936373907717737736311859039834565606659948875742273070213488434104398549079850003610766037222581329415245671250840364313712413486185244182260992419837920596299055081848194020532230062755361616289122433;
            6'd12: xpb[171] = 1024'd79966959838898440299613633199442791525862231228020873176387233100050672661733981399326973883725438673020000334657441201847928980668709092919840060862226832079907873570785141528033672122649687592755259693297856547840106835063376835159245967366323984319087043230168903349238304251983471351224109390831730579562;
            6'd13: xpb[171] = 1024'd24597525316744272958515305596989141114001536934154770543686908325899781048223910394263352766707054741050092325483481251379057808637158016718913336759246880953054859083564961319888025203778558698163099196879058003644601979541543184940027179805236258378934345125624449613288232236017777455266773593421577552360;
            6'd14: xpb[171] = 1024'd93294786478714847016215905399349923446839269766024352039118438616725784772022978299214802864346345118523333723767014735489250477446827275073146737672597970759892519165915998449372617476424635524881136308847499305813457974240606307685786961927377981705601550435197053907444688293980716576428127622637019009489;
            6'd15: xpb[171] = 1024'd37925351956560679675117577796896273034978575472158249406418113842574893158512907294151181747327961186553425714593054785020379305415276198872220013569618019633039504678695818241226970557553506630288975812428700761617953118718772657466568174366290255765448852330652600171494616278015022680470791825226865982287;
            6'd16: xpb[171] = 1024'd106622613118531253732818177599257055367816308304027830901849644133400896882311975199102631844967251564026667112876588269130571974224945457226453414482969109439877164761046855370711562830199583457007012924397142063786809113417835780212327956488431979092116057640225204465651072335977961801632145854442307439416;
            6'd17: xpb[171] = 1024'd51253178596377086391719849996803404955955614010161728269149319359250005268801904194039010727948867632056759103702628318661700802193394381025526690379989158313024150273826675162565915911328454562414852427978343519591304257896002129993109168927344253151963359535680750729701000320012267905674810057032154412214;
            6'd18: xpb[171] = 1024'd119950439758347660449420449799164187288793346842031309764580849650076008992600972098990460825588158009530000501986161802771893471003063639379760091293340248119861810356177712292050508183974531389132889539946784821760160252595065252738868951049485976478630564845253355023857456377975207026836164086247595869343;
            6'd19: xpb[171] = 1024'd64581005236193493108322122196710536876932652548165207131880524875925117379090901093926839708569774077560092492812201852303022298971512563178833367190360296993008795868957532083904861265103402494540729043527986277564655397073231602519650163488398250538477866740708901287907384362009513130878828288837442842141;
            6'd20: xpb[171] = 1024'd9211570714039325767223794594256886465071958254299104499180200101774225765580830088863218591551390145590184483638241901834151126939961486977906643087380345866155781381737351875759214346232273599948568547109187733369150541551397952300431375927310524598325168636164447551957312346043819234921492491427289814939;
            6'd21: xpb[171] = 1024'd77908831876009899824924394396617668797909691086168685994611730392600229489379897993814668689190680523063425881921775385944343795749630745332140044000731435672993441464088389005243806618878350426666605659077629035538006536250461075046191158049452247924992373945737051846113768404006758356082846520642731272068;
            6'd22: xpb[171] = 1024'd22539397353855732483826066794164018386048996792302583361911405618449337875869826988751047572172296591093517872747815435475472623718079669131213319897751484546140426976868208797098159700007221532074445162658830491342501680728627424826972370488364521984839675841192598110163696388041064460125510723232578244866;
            6'd23: xpb[171] = 1024'd91236658515826306541526666596524800718886729624172164857342935909275341599668894893702497669811586968566759271031348919585665292527748927485446720811102574352978087059219245926582751972653298358792482274627271793511357675427690547572732152610506245311506881150765202404320152446004003581286864752448019701995;
            6'd24: xpb[171] = 1024'd35867223993672139200428338994071150307026035330306062224642611135124449986158823888638876552793203036596851261857388969116794120496197851284519996708122623226125072571999065718437105053782169464200321778208473249315852819905856897353513365049418519371354183046220748668370080430038309685329528955037866674793;
            6'd25: xpb[171] = 1024'd104564485155642713258128938796431932639863768162175643720074141425950453709957891793590326650432493414070092660140922453226986789305867109638753397621473713032962732654350102847921697326428246290918358890176914551484708814604920020099273147171560242698021388355793352962526536488001248806490882984253308131922;
            6'd26: xpb[171] = 1024'd49195050633488545917030611193978282228003073868309541087373816651799562096447820788526705533414109482100184650966962502758115617274316033437826673518493761906109718167129922639776050407557117396326198393758116007289203959083086369880054359610472516757868690251248899226576464472035554910533547186843155104720;
            6'd27: xpb[171] = 1024'd117892311795459119974731210996339064560840806700179122582805346942625565820246888693478155631053399859573426049250495986868308286083985291792060074431844851712947378249480959769260642680203194223044235505726557309458059953782149492625814141732614240084535895560821503520732920529998494031694901216058596561849;
            6'd28: xpb[171] = 1024'd62522877273304952633632883393885414148980112406313019950105022168474674206736817688414534514035015927603518040076536036399437114052434215591133350328864900586094363762260779561114995761332065328452075009307758765262555098260315842406595354171526514144383197456277049784782848514032800135737565418648443534647;
            6'd29: xpb[171] = 1024'd7153442751150785292534555791431763737119418112446917317404697394323782593226746683350913397016631995633610030902576085930565942020883139390206626225884949459241349275040599352969348842460936433859914512888960221067050242738482192187376566610438788204230499351732596048832776498067106239780229621238290507445;
            6'd30: xpb[171] = 1024'd75850703913121359350235155593792546069957150944316498812836227685149786317025814588302363494655922373106851429186109570040758610830552397744440027139236039266079009357391636482453941115107013260577951624857401523235906237437545314933136348732580511530897704661305200342989232556030045360941583650453731964574;
            6'd31: xpb[171] = 1024'd20481269390967192009136827991338895658096456650450396180135902910998894703515743583238742377637538441136943420012149619571887438799001321543513303036256088139225994870171456274308294196235884365985791128438602979040401381915711664713917561171492785590745006556760746607039160540064351464984247853043578937372;
            6'd32: xpb[171] = 1024'd89178530552937766066837427793699677990934189482319977675567433201824898427314811488190192475276828818610184818295683103682080107608670579897746703949607177946063654952522493403792886468881961192703828240407044281209257376614774787459677343293634508917412211866333350901195616598027290586145601882259020394501;
            6'd33: xpb[171] = 1024'd33809096030783598725739100191246027579073495188453875042867108427674006813804740483126571358258444886640276809121723153213208935577119503696819979846627226819210640465302313195647239550010832298111667743988245737013752521092941137240458555732546782977259513761788897165245544582061596690188266084848867367299;
            6'd34: xpb[171] = 1024'd102506357192754172783439699993606809911911228020323456538298638718500010537603808388078021455897735264113518207405256637323401604386788762051053380759978316626048300547653350325131831822656909124829704855956687039182608515792004259986218337854688506303926719071361501459402000640024535811349620114064308824428;
            6'd35: xpb[171] = 1024'd47136922670600005442341372391153159500050533726457353905598313944349118924093737383014400338879351332143610198231296686854530432355237685850126656656998365499195286060433170116986184903785780230237544359537888494987103660270170609766999550293600780363774020966817047723451928624058841915392284316654155797226;
            6'd36: xpb[171] = 1024'd115834183832570579500041972193513941832888266558326935401029844235175122647892805287965850436518641709616851596514830170964723101164906944204360057570349455306032946142784207246470777176431857056955581471506329797155959654969233732512759332415742503690441226276389652017608384682021781036553638345869597254355;
            6'd37: xpb[171] = 1024'd60464749310416412158943644591060291421027572264460832768329519461024231034382734282902229319500257777646943587340870220495851929133355868003433333467369504179179931655564027038325130257560728162363420975087531252960454799447400082293540544854654777750288528171845198281658312666056087140596302548459444227153;
            6'd38: xpb[171] = 1024'd5095314788262244817845316988606641009166877970594730135629194686873339420872663277838608202481873845677035578166910270026980757101804791802506609364389553052326917168343846830179483338689599267771260478668732708764949943925566432074321757293567051810135830067300744545708240650090393244638966751049291199951;
            6'd39: xpb[171] = 1024'd73792575950232818875545916790967423342004610802464311631060724977699343144671731182790058300121164223150276976450443754137173425911474050156740010277740642859164577250694883959664075611335676094489297590637174010933805938624629554820081539415708775136803035376873348839864696708053332365800320780264732657080;
            6'd40: xpb[171] = 1024'd18423141428078651534447589188513772930143916508598208998360400203548451531161660177726437183102780291180368967276483803668302253879922973955813286174760691732311562763474703751518428692464547199897137094218375466738301083102795904600862751854621049196650337272328895103914624692087638469842984982854579629878;
            6'd41: xpb[171] = 1024'd87120402590049225592148188990874555262981649340467790493791930494374455254960728082677887280742070668653610365560017287778494922689592232310046687088111781539149222845825740881003020965110624026615174206186816768907157077801859027346622533976762772523317542581901499398071080750050577591004339012070021087007;
            6'd42: xpb[171] = 1024'd31750968067895058251049861388420904851120955046601687861091605720223563641450657077614266163723686736683702356386057337309623750658041156109119962985131830412296208358605560672857374046239495132023013709768018224711652222280025377127403746415675046583164844477357045662121008734084883695047003214659868059805;
            6'd43: xpb[171] = 1024'd100448229229865632308750461190781687183958687878471269356523136011049567365249724982565716261362977114156943754669590821419816419467710414463353363898482920219133868440956597802341966318885571958741050821736459526880508216979088499873163528537816769909832049786929649956277464792047822816208357243875309516934;
            6'd44: xpb[171] = 1024'd45078794707711464967652133588328036772097993584605166723822811236898675751739653977502095144344593182187035745495630870950945247436159338262426639795502969092280853953736417594196319400014443064148890325317660982685003361457254849653944740976729043969679351682385196220327392776082128920251021446465156489732;
            6'd45: xpb[171] = 1024'd113776055869682039025352733390688819104935726416474748219254341527724679475538721882453545241983883559660277143779164355061137916245828596616660040708854058899118514036087454723680911672660519890866927437286102284853859356156317972399704523098870767296346556991957800514483848834045068041412375475680597946861;
            6'd46: xpb[171] = 1024'd58406621347527871684254405788235168693075032122608645586554016753573787862028650877389924124965499627690369134605204404592266744214277520415733316605874107772265499548867274515535264753789390996274766940867303740658354500634484322180485735537783041356193858887413346778533776818079374145455039678270444919659;
            6'd47: xpb[171] = 1024'd3037186825373704343156078185781518281214337828742542953853691979422896248518579872326303007947115695720461125431244454123395572182726444214806592502894156645412485061647094307389617834918262101682606444448505196462849645112650671961266947976695315416041160782868893042583704802113680249497703880860291892457;
            6'd48: xpb[171] = 1024'd71734447987344278400856677988142300614052070660612124449285222270248899972317647777277753105586406073193702523714777938233588240992395702569039993416245246452250145143998131436874210107564338928400643556416946498631705639811713794707026730098837038742708366092441497336740160860076619370659057910075733349586;
            6'd49: xpb[171] = 1024'd16365013465190111059758350385688650202191376366746021816584897496098008358807576772214131988568022141223794514540817987764717068960844626368113269313265295325397130656777951228728563188693210033808483059998147954436200784289880144487807942537749312802555667987897043600790088844110925474701722112665580322384;
            6'd50: xpb[171] = 1024'd85062274627160685117458950188049432535029109198615603312016427786924012082606644677165582086207312518697035912824351471874909737770513884722346670226616385132234790739128988358213155461339286860526520171966589256605056778988943267233567724659891036129222873297469647894946544902073864595863076141881021779513;
            6'd51: xpb[171] = 1024'd29692840105006517776360622585595782123168414904749500679316103012773120469096573672101960969188928586727127903650391521406038565738962808521419946123636434005381776251908808150067508542468157965934359675547790712409551923467109617014348937098803310189070175192925194158996472886108170699905740344470868752311;
            6'd52: xpb[171] = 1024'd98390101266977091834061222387956564456006147736619082174747633303599124192895641577053411066828218964200369301933925005516231234548632066875653347036987523812219436334259845279552100815114234792652396787516232014578407918166172739760108719220945033515737380502497798453152928944071109821067094373686310209440;
            6'd53: xpb[171] = 1024'd43020666744822924492962894785502914044145453442752979542047308529448232579385570571989789949809835032230461292759965055047360062517080990674726622934007572685366421847039665071406453896243105898060236291097433470382903062644339089540889931659857307575584682397953344717202856928105415925109758576276157182238;
            6'd54: xpb[171] = 1024'd111717927906793498550663494587863696376983186274622561037478838820274236303184638476941240047449125409703702691043498539157552731326750249028960023847358662492204081929390702200891046168889182724778273403065874772551759057343402212286649713781999030902251887707525949011359312986068355046271112605491598639367;
            6'd55: xpb[171] = 1024'd56348493384639331209565166985410045965122491980756458404778514046123344689674567471877618930430741477733794681869538588688681559295199172828033299744378711365351067442170521992745399250018053830186112906647076228356254201821568562067430926220911304962099189602981495275409240970102661150313776808081445612165;
            6'd56: xpb[171] = 1024'd979058862485163868466839382956395553261797686890355772078189271972453076164496466813997813412357545763886672695578638219810387263648096627106575641398760238498052954950341784599752331146924935593952410228277684160749346299734911848212138659823579021946491498437041539459168954136967254356441010671292584963;
            6'd57: xpb[171] = 1024'd69676320024455737926167439185317177886099530518759937267509719562798456799963564371765447911051647923237128070979112122330003056073317354981339976554749850045335713037301378914084344603793001762311989522196718986329605340998798034593971920781965302348613696808009645833615625012099906375517795039886734042092;
            6'd58: xpb[171] = 1024'd14306885502301570585069111582863527474238836224893834634809394788647565186453493366701826794033263991267220061805152171861131884041766278780413252451769898918482698550081198705938697684921872867719829025777920442134100485476964384374753133220877576408460998703465192097665552996134212479560459242476581014890;
            6'd59: xpb[171] = 1024'd83004146664272144642769711385224309807076569056763416130240925079473568910252561271653276891672554368740461460088685655971324552851435537134646653365120988725320358632432235835423289957567949694437866137746361744302956480176027507120512915343019299735128204013037796391822009054097151600721813271692022472019;
            6'd60: xpb[171] = 1024'd27634712142117977301671383782770659395215874762897313497540600305322677296742490266589655774654170436770553450914725705502453380819884460933719929262141037598467344145212055627277643038696820799845705641327563200107451624654193856901294127781931573794975505908493342655871937038131457704764477474281869444817;
            6'd61: xpb[171] = 1024'd96331973304088551359371983585131441728053607594766894992972130596148681020541558171541105872293460814243794849198259189612646049629553719287953330175492127405305004227563092756762235311342897626563742753296004502276307619353256979647053909904073297121642711218065946950028393096094396825925831503497310901946;
            6'd62: xpb[171] = 1024'd40962538781934384018273655982677791316192913300900792360271805821997789407031487166477484755275076882273886840024299239143774877598002643087026606072512176278451989740342912548616588392471768731971582256877205958080802763831423329427835122342985571181490013113521493214078321080128702929968495706087157874744;
            6'd63: xpb[171] = 1024'd109659799943904958075974255785038573649030646132770373855703336112823793130830555071428934852914367259747128238307832723253967546407671901441260006985863266085289649822693949678101180665117845558689619368845647260249658758530486452173594904465127294508157218423094097508234777138091642051129849735302599331873;
        endcase
    end

    always_comb begin
        case(flag[57][11:6])
            6'd0: xpb[172] = 1024'd0;
            6'd1: xpb[172] = 1024'd54290365421750790734875928182584923237169951838904271223003011338672901517320484066365313735895983327777220229133872772785096374376120825240333282882883314958436635335473769469955533746246716664097458872426848716054153903008652801954376116904039568568004520318549643772284705122125948155172513937892446304671;
            6'd2: xpb[172] = 1024'd108580730843501581469751856365169846474339903677808542446006022677345803034640968132730627471791966655554440458267745545570192748752241650480666565765766629916873270670947538939911067492493433328194917744853697432108307806017305603908752233808079137136009040637099287544569410244251896310345027875784892609342;
            6'd3: xpb[172] = 1024'd38804400581127630805828857142940336966811428390977129540877178951041809214652313289080869993030275673888511279944124883776225282287142141165839723632318903941619231436850091072236362047222944270982179008893306301798100858805061632898149781028889256437193657541531873286747587292449211448398851987051744429682;
            6'd4: xpb[172] = 1024'd93094766002878421540704785325525260203981380229881400763880190289714710731972797355446183728926259001665731509077997656561321656663262966406173006515202218900055866772323860542191895793469660935079637881320155017852254761813714434852525897932928825005198177860081517059032292414575159603571365924944190734353;
            6'd5: xpb[172] = 1024'd23318435740504470876781786103295750696452904943049987858751346563410716911984142511796426250164568019999802330754376994767354190198163457091346164381754492924801827538226412674517190348199171877866899145359763887542047814601470463841923445153738944306382794764514102801210469462772474741625190036211042554693;
            6'd6: xpb[172] = 1024'd77608801162255261611657714285880673933622856781954259081754357902083618429304626578161739986060551347777022559888249767552450564574284282331679447264637807883238462873700182144472724094445888541964358017786612603596201717610123265796299562057778512874387315083063746573495174584898422896797703974103488859364;
            6'd7: xpb[172] = 1024'd7832470899881310947734715063651164426094381495122846176625514175779624609315971734511982507298860366111093381564629105758483098109184773016852605131190081907984423639602734276798018649175399484751619281826221473285994770397879294785697109278588632175571931987496332315673351633095738034851528085370340679704;
            6'd8: xpb[172] = 1024'd62122836321632101682610643246236087663264333334027117399628525514452526126636455800877296243194843693888313610698501878543579472485305598257185888014073396866421058975076503746753552395422116148849078154253070189340148673406532096740073226182628200743576452306045976087958056755221686190024042023262786984375;
            6'd9: xpb[172] = 1024'd116413201743382892417486571428821010900434285172931388622631536853125427643956939867242609979090827021665533839832374651328675846861426423497519170896956711824857694310550273216709086141668832812946537026679918905394302576415184898694449343086667769311580972624595619860242761877347634345196555961155233289046;
            6'd10: xpb[172] = 1024'd46636871481008941753563572206591501392905809886099975717502693126821433823968285023592852500329136039999604661508753989534708380396326914182692328763508985849603655076452825349034380696398343755733798290719527775084095629202940927683846890307477888612765589529028205602420938925544949483250380072422085109386;
            6'd11: xpb[172] = 1024'd100927236902759732488439500389176424630075761725004246940505704465494335341288769089958166236225119367776824890642626762319804754772447739423025611646392300808040290411926594818989914442645060419831257163146376491138249532211593729638223007211517457180770109847577849374705644047670897638422894010314531414057;
            6'd12: xpb[172] = 1024'd31150906640385781824516501166946915122547286438172834035376860739190341521300114246308408757463428386110895712319006100525837288307348230108198769512944574832786251177829146951315208997374571362618518427185985360828042584999349758627620554432327576481954726752010435116883821095868212776476718121581383234397;
            6'd13: xpb[172] = 1024'd85441272062136572559392429349531838359717238277077105258379872077863243038620598312673722493359411713888115941452878873310933662683469055348532052395827889791222886513302916421270742743621288026715977299612834076882196488008002560581996671336367145049959247070560078889168526217994160931649232059473829539068;
            6'd14: xpb[172] = 1024'd15664941799762621895469430127302328852188762990245692353251028351559249218631943469023965014597720732222186763129258211516966196218369546033705210262380163815968847279205468553596037298350798969503238563652442946571989540795758589571394218557177264351143863974992664631346703266191476069703056170740681359408;
            6'd15: xpb[172] = 1024'd69955307221513412630345358309887252089358714829149963576254039690232150735952427535389278750493704059999406992263130984302062570594490371274038493145263478774405482614679238023551571044597515633600697436079291662626143443804411391525770335461216832919148384293542308403631408388317424224875570108633127664079;
            6'd16: xpb[172] = 1024'd178976959139461966422359087657742581830239542318550671125195963928156915963772691739521271732013078333477813939510322508095104129390861959211651011815752799151443380581790155876865599327026576387958700118900532315936496592167420515167882682026952220333001197974894145809585436514739362929394219899979484419;
            6'd17: xpb[172] = 1024'd54469342380890252701298287270242665819000191381222821894128207302601058433284256758104835007627996406110698043073383095293191478505511687199544933894699067757588078716055559625832399345573743240485417572545749248370090399600820222469543999586066520788337521516524537918094290558640687518101908157792425789090;
            6'd18: xpb[172] = 1024'd108759707802641043436174215452827589056170143220127093117131218641273959950604740824470148743523979733887918272207255868078287852881632512439878216777582382716024714051529329095787933091820459904582876444972597964424244302609473024423920116490106089356342041835074181690378995680766635673274422095684872093761;
            6'd19: xpb[172] = 1024'd38983377540267092772251216230598079548641667933295680212002374914969966130616085980820391264762288752221989093883635206284320386416533003125051374644134656740770674817431881228113227646549970847370137709012206834114037355397229053413317663710916208657526658739506767432557172728963950811328246206951723914101;
            6'd20: xpb[172] = 1024'd93273742962017883507127144413183002785811619772199951435005386253642867647936570047185705000658272079999209323017507979069416760792653828365384657527017971699207310152905650698068761392796687511467596581439055550168191258405881855367693780614955777225531179058056411204841877851089898966500760144844170218772;
            6'd21: xpb[172] = 1024'd23497412699643932843204145190953493278283144485368538529876542527338873827947915203535947521896581098333280144693887317275449294327554319050557815393570245723953270918808202830394055947526198454254857845478664419857984311193637884357091327835765896526715795962488996947020054899287214104554584256111022039112;
            6'd22: xpb[172] = 1024'd77787778121394723578080073373538416515453096324272809752879553866011775345268399269901261257792564426110500373827760090060545668703675144290891098276453560682389906254281972300349589693772915118352316717905513135912138214202290686311467444739805465094720316281038640719304760021413162259727098194003468343783;
            6'd23: xpb[172] = 1024'd8011447859020772914157074151308907007924621037441396847750710139707781525279744426251503779030873444444571195504139428266578202238575634976064256143005834707135867020184524432674884248502426061139577981945122005601931266990046715300864991960615584395904933185471226461482937069610477397780922305270320164123;
            6'd24: xpb[172] = 1024'd62301813280771563649033002333893830245094572876345668070753721478380683042600228492616817514926856772221791424638012201051674576614696460216397539025889149665572502355658293902630417994749142725237036854371970721656085169998699517255241108864655152963909453504020870233767642191736425552953436243162766468794;
            6'd25: xpb[172] = 1024'd116592178702522354383908930516478753482264524715249939293756732817053584559920712558982131250822840099999011653771884973836770950990817285456730821908772464624009137691132063372585951740995859389334495726798819437710239073007352319209617225768694721531913973822570514006052347313862373708125950181055212773465;
            6'd26: xpb[172] = 1024'd46815848440148403719985931294249243974736049428418526388627889090749590739932057715332373772061149118333082475448264312042803484525717776141903979775324738648755098457034615504911246295725370332121756990838428307400032125795108348199014772989504840833098590727003099748230524362059688846179774292322064593805;
            6'd27: xpb[172] = 1024'd101106213861899194454861859476834167211906001267322797611630900429422492257252541781697687507957132446110302704582137084827899858901838601382237262658208053607191733792508384974866780041972086996219215863265277023454186028803761150153390889893544409401103111045552743520515229484185637001352288230214510898476;
            6'd28: xpb[172] = 1024'd31329883599525243790938860254604657704377525980491384706502056703118498437263886938047930029195441464444373526258516423033932392436739092067410420524760327631937694558410937107192074596701597939006477127304885893143979081591517179142788437114354528702287727949985329262693406532382952139406112341481362718816;
            6'd29: xpb[172] = 1024'd85620249021276034525814788437189580941547477819395655929505068041791399954584371004413243765091424792221593755392389195819028766812859917307743703407643642590374329893884706577147608342948314603103935999731734609198132984600169981097164554018394097270292248268534973034978111654508900294578626279373809023487;
            6'd30: xpb[172] = 1024'd15843918758902083861891789214960071434019002532564243024376224315487406134595716160763486286329733810555664577068768534025061300347760407992916861274195916615120290659787258709472902897677825545891197263771343478887926037387926010086562101239204216571476865172967558777156288702706215432632450390640660843827;
            6'd31: xpb[172] = 1024'd70134284180652874596767717397544994671188954371468514247379235654160307651916200227128800022225717138332884806202641306810157674723881233233250144157079231573556925995261028179428436643924542209988656136198192194942079940396578812040938218143243785139481385491517202549440993824832163587804964328533107148498;
            6'd32: xpb[172] = 1024'd357953918278923932844718175315485163660479084637101342250391927856313831927545383479042543464026156666955627879020645016190208258781723918423302023631505598302886761163580311753731198654053152775917400237801064631872993184334841030335765364053904440666002395949788291619170873029478725858788439799958968838;
            6'd33: xpb[172] = 1024'd54648319340029714667720646357900408400830430923541372565253403266529215349248029449844356279360009484444175857012893417801286582634902549158756584906514820556739522096637349781709264944900769816873376272664649780686026896192987642984711882268093473008670522714499432063903875995155426881031302377692405273509;
            6'd34: xpb[172] = 1024'd108938684761780505402596574540485331638000382762445643788256414605202116866568513516209670015255992812221396086146766190586382957011023374399089867789398135515176157432111119251664798691147486480970835145091498496740180799201640444939087999172133041576675043033049075836188581117281375036203816315584851578180;
            6'd35: xpb[172] = 1024'd39162354499406554738673575318255822130471907475614230883127570878898123046579858672559912536494301830555466907823145528792415490545923865084263025655950409539922118198013671383990093245876997423758096409131107366429973851989396473928485546392943160877859659937481661578366758165478690174257640426851703398520;
            6'd36: xpb[172] = 1024'd93452719921157345473549503500840745367641859314518502106130582217571024563900342738925226272390285158332687136957018301577511864922044690324596308538833724498358753533487440853945626992123714087855555281557956082484127754998049275882861663296982729445864180256031305350651463287604638329430154364744149703191;
            6'd37: xpb[172] = 1024'd23676389658783394809626504278611235860113384027687089201001738491267030743911687895275468793628594176666757958633397639783544398456945181009769466405385998523104714299389992986270921546853225030642816545597564952173920807785805304872259210517792848747048797160463891092829640335801953467483978476011001523531;
            6'd38: xpb[172] = 1024'd77966755080534185544502432461196159097283335866591360424004749829939932261232171961640782529524577504443978187767270412568640772833066006250102749288269313481541349634863762456226455293099941694740275418024413668228074710794458106826635327421832417315053317479013534865114345457927901622656492413903447828202;
            6'd39: xpb[172] = 1024'd8190424818160234880579433238966649589754860579759947518875906103635938441243517117991025050762886522778049009443649750774673306367966496935275907154821587506287310400766314588551749847829452637527536682064022537917867763582214135816032874642642536616237934383446120607292522506125216760710316525170299648542;
            6'd40: xpb[172] = 1024'd62480790239911025615455361421551572826924812418664218741878917442308839958564001184356338786658869850555269238577522523559769680744087322175609190037704902464723945736240084058507283594076169301624995554490871253972021666590866937770408991546682105184242454701995764379577227628251164915882830463062745953213;
            6'd41: xpb[172] = 1024'd116771155661661816350331289604136496064094764257568489964881928780981741475884485250721652522554853178332489467711395296344866055120208147415942472920588217423160581071713853528462817340322885965722454426917719970026175569599519739724785108450721673752246975020545408151861932750377113071055344400955192257884;
            6'd42: xpb[172] = 1024'd46994825399287865686408290381906986556566288970737077059753085054677747655895830407071895043793162196666560289387774634550898588655108638101115630787140491447906541837616405660788111895052396908509715690957328839715968622387275768714182655671531793053431591924977993894040109798574428209109168512222044078224;
            6'd43: xpb[172] = 1024'd101285190821038656421284218564491909793736240809641348282756096393350649173216314473437208779689145524443780518521647407335994963031229463341448913670023806406343177173090175130743645641299113572607174563384177555770122525395928570668558772575571361621436112243527637666324814920700376364281682450114490382895;
            6'd44: xpb[172] = 1024'd31508860558664705757361219342262400286207765522809935377627252667046655353227659629787451300927454542777851340198026745542027496566129954026622071536576080431089137938992727263068940196028624515394435827423786425459915578183684599657956319796381480922620729147960223408502991968897691502335506561381342203235;
            6'd45: xpb[172] = 1024'd85799225980415496492237147524847323523377717361714206600630264005719556870548143696152765036823437870555071569331899518327123870942250779266955354419459395389525773274466496733024473942275341179491894699850635141514069481192337401612332436700421049490625249466509867180787697091023639657508020499273788507906;
            6'd46: xpb[172] = 1024'd16022895718041545828314148302617814015849242074882793695501420279415563050559488852503007558061746888889142391008278856533156404477151269952128512286011669414271734040369048865349768497004852122279155963890244011203862533980093430601729983921231168791809866370942452922965874139220954795561844610540640328246;
            6'd47: xpb[172] = 1024'd70313261139792336563190076485202737253019193913787064918504431618088464567879972918868321293957730216666362620142151629318252778853272095192461795168894984372708369375842818335305302243251568786376614836317092727258016436988746232556106100825270737359814386689492096695250579261346902950734358548433086632917;
            6'd48: xpb[172] = 1024'd536930877418385899267077262973227745490718626955652013375587891784470747891318075218563815196039235000433441818530967524285312388172585877634953035447258397454330141745370467630596797981079729163876100356701596947809489776502261545503648046080856660999003593924682437428756309544218088788182659699938453257;
            6'd49: xpb[172] = 1024'd54827296299169176634143005445558150982660670465859923236378599230457372265211802141583877551092022562777653670952403740309381686764293411117968235918330573355890965477219139937586130544227796393261334972783550313001963392785155063499879764950120425229003523912474326209713461431670166243960696597592384757928;
            6'd50: xpb[172] = 1024'd109117661720919967369018933628143074219830622304764194459381610569130273782532286207949191286988005890554873900086276513094478061140414236358301518801213888314327600812692909407541664290474513057358793845210399029056117295793807865454255881854159993797008044231023969981998166553796114399133210535484831062599;
            6'd51: xpb[172] = 1024'd39341331458546016705095934405913564712302147017932781554252766842826279962543631364299433808226314908888944721762655851300510594675314727043474676667766162339073561578595461539866958845204024000146055109250007898745910348581563894443653429074970113098192661135456555724176343601993429537187034646751682882939;
            6'd52: xpb[172] = 1024'd93631696880296807439971862588498487949472098856837052777255778181499181479864115430664747544122298236666164950896528624085606969051435552283807959550649477297510196914069231009822492591450740664243513981676856614800064251590216696398029545979009681666197181454006199496461048724119377692359548584644129187610;
            6'd53: xpb[172] = 1024'd23855366617922856776048863366268978441943623570005639872126934455195187659875460587014990065360607255000235772572907962291639502586336042968981117417201751322256157679971783142147787146180251607030775245716465484489857304377972725387427093199819800967381798358438785238639225772316692830413372695910981007950;
            6'd54: xpb[172] = 1024'd78145732039673647510924791548853901679113575408909911095129945793868089177195944653380303801256590582777456001706780735076735876962456868209314400300085066280692793015445552612103320892426968271128234118143314200544011207386625527341803210103859369535386318676988429010923930894442640985585886633803427312621;
            6'd55: xpb[172] = 1024'd8369401777299696847001792326624392171585100122078498190001102067564095357207289809730546322494899601111526823383160073282768410497357358894487558166637340305438753781348104744428615447156479213915495382182923070233804260174381556331200757324669488836570935581421014753102107942639956123639710745070279132961;
            6'd56: xpb[172] = 1024'd62659767199050487581877720509209315408755051960982769413004113406236996874527773876095860058390882928888747052517032846067864784873478184134820841049520655263875389116821874214384149193403195878012954254609771786287958163183034358285576874228709057404575455899970658525386813064765904278812224682962725437632;
            6'd57: xpb[172] = 1024'd116950132620801278316753648691794238645925003799887040636007124744909898391848257942461173794286866256665967281650905618852961159249599009375154123932403970222312024452295643684339682939649912542110413127036620502342112066191687160239952991132748625972579976218520302297671518186891852433984738620855171742303;
            6'd58: xpb[172] = 1024'd47173802358427327652830649469564729138396528513055627730878281018605904571859603098811416315525175275000038103327284957058993692784499500060327281798956244247057985218198195816664977494379423484897674391076229372031905118979443189229350538353558745273764593122952888039849695235089167572038562732122023562643;
            6'd59: xpb[172] = 1024'd101464167780178118387706577652149652375566480351959898953881292357278806089180087165176730051421158602777258332461157729844090067160620325300660564681839559205494620553671965286620511240626140148995133263503078088086059021988095991183726655257598313841769113441502531812134400357215115727211076670014469867314;
            6'd60: xpb[172] = 1024'd31687837517804167723783578429920142868038005065128486048752448630974812269191432321526972572659467621111329154137537068050122600695520815985833722548391833230240581319574517418945805795355651091782394527542686957775852074775852020173124202478408433142953730345935117554312577405412430865264900781281321687654;
            6'd61: xpb[172] = 1024'd85978202939554958458659506612505066105207956904032757271755459969647713786511916387892286308555450948888549383271409840835218975071641641226167005431275148188677216655048286888901339541602367755879853399969535673830005977784504822127500319382448001710958250664484761326597282527538379020437414719173767992325;
            6'd62: xpb[172] = 1024'd16201872677181007794736507390275556597679481617201344366626616243343719966523261544242528829793759967222620204947789179041251508606542131911340163297827422213423177420950839021226634096331878698667114664009144543519799030572260851116897866603258121012142867568917347068775459575735694158491238830440619812665;
            6'd63: xpb[172] = 1024'd70492238098931798529612435572860479834849433456105615589629627582016621483843745610607842565689743294999840434081661951826347882982662957151673446180710737171859812756424608491182167842578595362764573536435993259573952933580913653071273983507297689580147387887466990841060164697861642313663752768333066117336;
        endcase
    end

    always_comb begin
        case(flag[57][16:12])
            5'd0: xpb[173] = 1024'd0;
            5'd1: xpb[173] = 1024'd715907836557847865689436350630970327320958169274202684500783855712627663855090766958085086928052313333911255758041290032380416517563447836846604047263011196605773522327160623507462397308106305551834800475602129263745986368669682060671530728107808881332004791899576583238341746058957451717576879599917937676;
            5'd2: xpb[173] = 1024'd1431815673115695731378872701261940654641916338548405369001567711425255327710181533916170173856104626667822511516082580064760833035126895673693208094526022393211547044654321247014924794616212611103669600951204258527491972737339364121343061456215617762664009583799153166476683492117914903435153759199835875352;
            5'd3: xpb[173] = 1024'd2147723509673543597068309051892910981962874507822608053502351567137882991565272300874255260784156940001733767274123870097141249552690343510539812141789033589817320566981481870522387191924318916655504401426806387791237959106009046182014592184323426643996014375698729749715025238176872355152730638799753813028;
            5'd4: xpb[173] = 1024'd2863631346231391462757745402523881309283832677096810738003135422850510655420363067832340347712209253335645023032165160129521666070253791347386416189052044786423094089308642494029849589232425222207339201902408517054983945474678728242686122912431235525328019167598306332953366984235829806870307518399671750704;
            5'd5: xpb[173] = 1024'd3579539182789239328447181753154851636604790846371013422503919278563138319275453834790425434640261566669556278790206450161902082587817239184233020236315055983028867611635803117537311986540531527759174002378010646318729931843348410303357653640539044406660023959497882916191708730294787258587884397999589688380;
            5'd6: xpb[173] = 1024'd4295447019347087194136618103785821963925749015645216107004703134275765983130544601748510521568313880003467534548247740194282499105380687021079624283578067179634641133962963741044774383848637833311008802853612775582475918212018092364029184368646853287992028751397459499430050476353744710305461277599507626056;
            5'd7: xpb[173] = 1024'd5011354855904935059826054454416792291246707184919418791505486989988393646985635368706595608496366193337378790306289030226662915622944134857926228330841078376240414656290124364552236781156744138862843603329214904846221904580687774424700715096754662169324033543297036082668392222412702162023038157199425563732;
            5'd8: xpb[173] = 1024'd5727262692462782925515490805047762618567665354193621476006270845701021310840726135664680695424418506671290046064330320259043332140507582694772832378104089572846188178617284988059699178464850444414678403804817034109967890949357456485372245824862471050656038335196612665906733968471659613740615036799343501408;
            5'd9: xpb[173] = 1024'd6443170529020630791204927155678732945888623523467824160507054701413648974695816902622765782352470820005201301822371610291423748658071030531619436425367100769451961700944445611567161575772956749966513204280419163373713877318027138546043776552970279931988043127096189249145075714530617065458191916399261439084;
            5'd10: xpb[173] = 1024'd7159078365578478656894363506309703273209581692742026845007838557126276638550907669580850869280523133339112557580412900323804165175634478368466040472630111966057735223271606235074623973081063055518348004756021292637459863686696820606715307281078088813320047918995765832383417460589574517175768795999179376760;
            5'd11: xpb[173] = 1024'd7874986202136326522583799856940673600530539862016229529508622412838904302405998436538935956208575446673023813338454190356184581693197926205312644519893123162663508745598766858582086370389169361070182805231623421901205850055366502667386838009185897694652052710895342415621759206648531968893345675599097314436;
            5'd12: xpb[173] = 1024'd8590894038694174388273236207571643927851498031290432214009406268551531966261089203497021043136627760006935069096495480388564998210761374042159248567156134359269282267925927482089548767697275666622017605707225551164951836424036184728058368737293706575984057502794918998860100952707489420610922555199015252112;
            5'd13: xpb[173] = 1024'd9306801875252022253962672558202614255172456200564634898510190124264159630116179970455106130064680073340846324854536770420945414728324821879005852614419145555875055790253088105597011165005381972173852406182827680428697822792705866788729899465401515457316062294694495582098442698766446872328499434798933189788;
            5'd14: xpb[173] = 1024'd10022709711809870119652108908833584582493414369838837583010973979976787293971270737413191216992732386674757580612578060453325831245888269715852456661682156752480829312580248729104473562313488277725687206658429809692443809161375548849401430193509324338648067086594072165336784444825404324046076314398851127464;
            5'd15: xpb[173] = 1024'd10738617548367717985341545259464554909814372539113040267511757835689414957826361504371276303920784700008668836370619350485706247763451717552699060708945167949086602834907409352611935959621594583277522007134031938956189795530045230910072960921617133219980071878493648748575126190884361775763653193998769065140;
            5'd16: xpb[173] = 1024'd11454525384925565851030981610095525237135330708387242952012541691402042621681452271329361390848837013342580092128660640518086664281015165389545664756208179145692376357234569976119398356929700888829356807609634068219935781898714912970744491649724942101312076670393225331813467936943319227481230073598687002816;
            5'd17: xpb[173] = 1024'd12170433221483413716720417960726495564456288877661445636513325547114670285536543038287446477776889326676491347886701930550467080798578613226392268803471190342298149879561730599626860754237807194381191608085236197483681768267384595031416022377832750982644081462292801915051809683002276679198806953198604940492;
            5'd18: xpb[173] = 1024'd12886341058041261582409854311357465891777247046935648321014109402827297949391633805245531564704941640010402603644743220582847497316142061063238872850734201538903923401888891223134323151545913499933026408560838326747427754636054277092087553105940559863976086254192378498290151429061234130916383832798522878168;
            5'd19: xpb[173] = 1024'd13602248894599109448099290661988436219098205216209851005514893258539925613246724572203616651632993953344313859402784510615227913833705508900085476897997212735509696924216051846641785548854019805484861209036440456011173741004723959152759083834048368745308091046091955081528493175120191582633960712398440815844;
            5'd20: xpb[173] = 1024'd14318156731156957313788727012619406546419163385484053690015677114252553277101815339161701738561046266678225115160825800647608330351268956736932080945260223932115470446543212470149247946162126111036696009512042585274919727373393641213430614562156177626640095837991531664766834921179149034351537591998358753520;
            5'd21: xpb[173] = 1024'd15034064567714805179478163363250376873740121554758256374516460969965180940956906106119786825489098580012136370918867090679988746868832404573778684992523235128721243968870373093656710343470232416588530809987644714538665713742063323274102145290263986507972100629891108248005176667238106486069114471598276691196;
            5'd22: xpb[173] = 1024'd15749972404272653045167599713881347201061079724032459059017244825677808604811996873077871912417150893346047626676908380712369163386395852410625289039786246325327017491197533717164172740778338722140365610463246843802411700110733005334773676018371795389304105421790684831243518413297063937786691351198194628872;
            5'd23: xpb[173] = 1024'd16465880240830500910857036064512317528382037893306661743518028681390436268667087640035956999345203206679958882434949670744749579903959300247471893087049257521932791013524694340671635138086445027692200410938848973066157686479402687395445206746479604270636110213690261414481860159356021389504268230798112566548;
            5'd24: xpb[173] = 1024'd17181788077388348776546472415143287855702996062580864428018812537103063932522178406994042086273255520013870138192990960777129996421522748084318497134312268718538564535851854964179097535394551333244035211414451102329903672848072369456116737474587413151968115005589837997720201905414978841221845110398030504224;
            5'd25: xpb[173] = 1024'd17897695913946196642235908765774258183023954231855067112519596392815691596377269173952127173201307833347781393951032250809510412939086195921165101181575279915144338058179015587686559932702657638795870011890053231593649659216742051516788268202695222033300119797489414580958543651473936292939421989997948441900;
            5'd26: xpb[173] = 1024'd18613603750504044507925345116405228510344912401129269797020380248528319260232359940910212260129360146681692649709073540841890829456649643758011705228838291111750111580506176211194022330010763944347704812365655360857395645585411733577459798930803030914632124589388991164196885397532893744656998869597866379576;
            5'd27: xpb[173] = 1024'd19329511587061892373614781467036198837665870570403472481521164104240946924087450707868297347057412460015603905467114830874271245974213091594858309276101302308355885102833336834701484727318870249899539612841257490121141631954081415638131329658910839795964129381288567747435227143591851196374575749197784317252;
            5'd28: xpb[173] = 1024'd20045419423619740239304217817667169164986828739677675166021947959953574587942541474826382433985464773349515161225156120906651662491776539431704913323364313504961658625160497458208947124626976555451374413316859619384887618322751097698802860387018648677296134173188144330673568889650808648092152628797702254928;
            5'd29: xpb[173] = 1024'd20761327260177588104993654168298139492307786908951877850522731815666202251797632241784467520913517086683426416983197410939032079009339987268551517370627324701567432147487658081716409521935082861003209213792461748648633604691420779759474391115126457558628138965087720913911910635709766099809729508397620192604;
            5'd30: xpb[173] = 1024'd21477235096735435970683090518929109819628745078226080535023515671378829915652723008742552607841569400017337672741238700971412495526903435105398121417890335898173205669814818705223871919243189166555044014268063877912379591060090461820145921843234266439960143756987297497150252381768723551527306387997538130280;
            5'd31: xpb[173] = 1024'd22193142933293283836372526869560080146949703247500283219524299527091457579507813775700637694769621713351248928499279991003792912044466882942244725465153347094778979192141979328731334316551295472106878814743666007176125577428760143880817452571342075321292148548886874080388594127827681003244883267597456067956;
        endcase
    end

    always_comb begin
        case(flag[58][5:0])
            6'd0: xpb[174] = 1024'd0;
            6'd1: xpb[174] = 1024'd11454525384925565851030981610095525237135330708387242952012541691402042621681452271329361390848837013342580092128660640518086664281015165389545664756208179145692376357234569976119398356929700888829356807609634068219935781898714912970744491649724942101312076670393225331813467936943319227481230073598687002816;
            6'd2: xpb[174] = 1024'd22909050769851131702061963220191050474270661416774485904025083382804085243362904542658722781697674026685160184257321281036173328562030330779091329512416358291384752714469139952238796713859401777658713615219268136439871563797429825941488983299449884202624153340786450663626935873886638454962460147197374005632;
            6'd3: xpb[174] = 1024'd34363576154776697553092944830286575711405992125161728856037625074206127865044356813988084172546511040027740276385981921554259992843045496168636994268624537437077129071703709928358195070789102666488070422828902204659807345696144738912233474949174826303936230011179675995440403810829957682443690220796061008448;
            6'd4: xpb[174] = 1024'd45818101539702263404123926440382100948541322833548971808050166765608170486725809085317445563395348053370320368514642562072346657124060661558182659024832716582769505428938279904477593427718803555317427230438536272879743127594859651882977966598899768405248306681572901327253871747773276909924920294394748011264;
            6'd5: xpb[174] = 1024'd57272626924627829255154908050477626185676653541936214760062708457010213108407261356646806954244185066712900460643303202590433321405075826947728323781040895728461881786172849880596991784648504444146784038048170341099678909493574564853722458248624710506560383351966126659067339684716596137406150367993435014080;
            6'd6: xpb[174] = 1024'd68727152309553395106185889660573151422811984250323457712075250148412255730088713627976168345093022080055480552771963843108519985686090992337273988537249074874154258143407419856716390141578205332976140845657804409319614691392289477824466949898349652607872460022359351990880807621659915364887380441592122016896;
            6'd7: xpb[174] = 1024'd80181677694478960957216871270668676659947314958710700664087791839814298351770165899305529735941859093398060644900624483626606649967106157726819653293457254019846634500641989832835788498507906221805497653267438477539550473291004390795211441548074594709184536692752577322694275558603234592368610515190809019712;
            6'd8: xpb[174] = 1024'd91636203079404526808247852880764201897082645667097943616100333531216340973451618170634891126790696106740640737029285124144693314248121323116365318049665433165539010857876559808955186855437607110634854460877072545759486255189719303765955933197799536810496613363145802654507743495546553819849840588789496022528;
            6'd9: xpb[174] = 1024'd103090728464330092659278834490859727134217976375485186568112875222618383595133070441964252517639533120083220829157945764662779978529136488505910982805873612311231387215111129785074585212367307999464211268486706613979422037088434216736700424847524478911808690033539027986321211432489873047331070662388183025344;
            6'd10: xpb[174] = 1024'd114545253849255658510309816100955252371353307083872429520125416914020426216814522713293613908488370133425800921286606405180866642810151653895456647562081791456923763572345699761193983569297008888293568076096340682199357818987149129707444916497249421013120766703932253318134679369433192274812300735986870028160;
            6'd11: xpb[174] = 1024'd1933083550056482962541870306236344863790210666523988344006103540445573501186836074607904084679532837325231605957773611119889466249946484729842187301958929668925465360009052399683142734709504055812727275318734904054932750664967269713210838463744913847612939960208420619841619232447878485174840982959962546645;
            6'd12: xpb[174] = 1024'd13387608934982048813572851916331870100925541374911231296018645231847616122868288345937265475528369850667811698086434251637976130530961650119387852058167108814617841717243622375802541091639204944642084082928368972274868532563682182683955330113469855948925016630601645951655087169391197712656071056558649549461;
            6'd13: xpb[174] = 1024'd24842134319907614664603833526427395338060872083298474248031186923249658744549740617266626866377206864010391790215094892156062794811976815508933516814375287960310218074478192351921939448568905833471440890538003040494804314462397095654699821763194798050237093300994871283468555106334516940137301130157336552277;
            6'd14: xpb[174] = 1024'd36296659704833180515634815136522920575196202791685717200043728614651701366231192888595988257226043877352971882343755532674149459092991980898479181570583467106002594431712762328041337805498606722300797698147637108714740096361112008625444313412919740151549169971388096615282023043277836167618531203756023555093;
            6'd15: xpb[174] = 1024'd47751185089758746366665796746618445812331533500072960152056270306053743987912645159925349648074880890695551974472416173192236123374007146288024846326791646251694970788947332304160736162428307611130154505757271176934675878259826921596188805062644682252861246641781321947095490980221155395099761277354710557909;
            6'd16: xpb[174] = 1024'd59205710474684312217696778356713971049466864208460203104068811997455786609594097431254711038923717904038132066601076813710322787655022311677570511082999825397387347146181902280280134519358008499959511313366905245154611660158541834566933296712369624354173323312174547278908958917164474622580991350953397560725;
            6'd17: xpb[174] = 1024'd70660235859609878068727759966809496286602194916847446056081353688857829231275549702584072429772554917380712158729737454228409451936037477067116175839208004543079723503416472256399532876287709388788868120976539313374547442057256747537677788362094566455485399982567772610722426854107793850062221424552084563541;
            6'd18: xpb[174] = 1024'd82114761244535443919758741576905021523737525625234689008093895380259871852957001973913433820621391930723292250858398094746496116217052642456661840595416183688772099860651042232518931233217410277618224928586173381594483223955971660508422280011819508556797476652960997942535894791051113077543451498150771566357;
            6'd19: xpb[174] = 1024'd93569286629461009770789723187000546760872856333621931960106437071661914474638454245242795211470228944065872342987058735264582780498067807846207505351624362834464476217885612208638329590147111166447581736195807449814419005854686573479166771661544450658109553323354223274349362727994432305024681571749458569173;
            6'd20: xpb[174] = 1024'd105023812014386575621820704797096071998008187042009174912118978763063957096319906516572156602319065957408452435115719375782669444779082973235753170107832541980156852575120182184757727947076812055276938543805441518034354787753401486449911263311269392759421629993747448606162830664937751532505911645348145571989;
            6'd21: xpb[174] = 1024'd116478337399312141472851686407191597235143517750396417864131520454465999718001358787901517993167902970751032527244380016300756109060098138625298834864040721125849228932354752160877126304006512944106295351415075586254290569652116399420655754960994334860733706664140673937976298601881070759987141718946832574805;
            6'd22: xpb[174] = 1024'd3866167100112965925083740612472689727580421333047976688012207080891147002373672149215808169359065674650463211915547222239778932499892969459684374603917859337850930720018104799366285469419008111625454550637469808109865501329934539426421676927489827695225879920416841239683238464895756970349681965919925093290;
            6'd23: xpb[174] = 1024'd15320692485038531776114722222568214964715752041435219640024748772293189624055124420545169560207902687993043304044207862757865596780908134849230039360126038483543307077252674775485683826348709000454811358247103876329801283228649452397166168577214769796537956590810066571496706401839076197830912039518612096106;
            6'd24: xpb[174] = 1024'd26775217869964097627145703832663740201851082749822462592037290463695232245736576691874530951056739701335623396172868503275952261061923300238775704116334217629235683434487244751605082183278409889284168165856737944549737065127364365367910660226939711897850033261203291903310174338782395425312142113117299098922;
            6'd25: xpb[174] = 1024'd38229743254889663478176685442759265438986413458209705544049832155097274867418028963203892341905576714678203488301529143794038925342938465628321368872542396774928059791721814727724480540208110778113524973466372012769672847026079278338655151876664653999162109931596517235123642275725714652793372186715986101738;
            6'd26: xpb[174] = 1024'd49684268639815229329207667052854790676121744166596948496062373846499317489099481234533253732754413728020783580430189784312125589623953631017867033628750575920620436148956384703843878897137811666942881781076006080989608628924794191309399643526389596100474186601989742566937110212669033880274602260314673104554;
            6'd27: xpb[174] = 1024'd61138794024740795180238648662950315913257074874984191448074915537901360110780933505862615123603250741363363672558850424830212253904968796407412698384958755066312812506190954679963277254067512555772238588685640149209544410823509104280144135176114538201786263272382967898750578149612353107755832333913360107370;
            6'd28: xpb[174] = 1024'd72593319409666361031269630273045841150392405583371434400087457229303402732462385777191976514452087754705943764687511065348298918185983961796958363141166934212005188863425524656082675610997213444601595396295274217429480192722224017250888626825839480303098339942776193230564046086555672335237062407512047110186;
            6'd29: xpb[174] = 1024'd84047844794591926882300611883141366387527736291758677352099998920705445354143838048521337905300924768048523856816171705866385582466999127186504027897375113357697565220660094632202073967926914333430952203904908285649415974620938930221633118475564422404410416613169418562377514023498991562718292481110734113002;
            6'd30: xpb[174] = 1024'd95502370179517492733331593493236891624663067000145920304112540612107487975825290319850699296149761781391103948944832346384472246748014292576049692653583292503389941577894664608321472324856615222260309011514542353869351756519653843192377610125289364505722493283562643894190981960442310790199522554709421115818;
            6'd31: xpb[174] = 1024'd106956895564443058584362575103332416861798397708533163256125082303509530597506742591180060686998598794733684041073492986902558911029029457965595357409791471649082317935129234584440870681786316111089665819124176422089287538418368756163122101775014306607034569953955869226004449897385630017680752628308108118634;
            6'd32: xpb[174] = 1024'd118411420949368624435393556713427942098933728416920406208137623994911573219188194862509422077847435808076264133202153627420645575310044623355141022165999650794774694292363804560560269038716016999919022626733810490309223320317083669133866593424739248708346646624349094557817917834328949245161982701906795121450;
            6'd33: xpb[174] = 1024'd5799250650169448887625610918709034591370631999571965032018310621336720503560508223823712254038598511975694817873320833359668398749839454189526561905876789006776396080027157199049428204128512167438181825956204712164798251994901809139632515391234741542838819880625261859524857697343635455524522948879887639935;
            6'd34: xpb[174] = 1024'd17253776035095014738656592528804559828505962707959207984030852312738763125241960495153073644887435525318274910001981473877755063030854619579072226662084968152468772437261727175168826561058213056267538633565838780384734033893616722110377007040959683644150896551018487191338325634286954683005753022478574642751;
            6'd35: xpb[174] = 1024'd28708301420020580589687574138900085065641293416346450936043394004140805746923412766482435035736272538660855002130642114395841727311869784968617891418293147298161148794496297151288224917987913945096895441175472848604669815792331635081121498690684625745462973221411712523151793571230273910486983096077261645567;
            6'd36: xpb[174] = 1024'd40162826804946146440718555748995610302776624124733693888055935695542848368604865037811796426585109552003435094259302754913928391592884950358163556174501326443853525151730867127407623274917614833926252248785106916824605597691046548051865990340409567846775049891804937854965261508173593137968213169675948648383;
            6'd37: xpb[174] = 1024'd51617352189871712291749537359091135539911954833120936840068477386944890990286317309141157817433946565346015186387963395432015055873900115747709220930709505589545901508965437103527021631847315722755609056394740985044541379589761461022610481990134509948087126562198163186778729445116912365449443243274635651199;
            6'd38: xpb[174] = 1024'd63071877574797278142780518969186660777047285541508179792081019078346933611967769580470519208282783578688595278516624035950101720154915281137254885686917684735238277866200007079646419988777016611584965864004375053264477161488476373993354973639859452049399203232591388518592197382060231592930673316873322654015;
            6'd39: xpb[174] = 1024'd74526402959722843993811500579282186014182616249895422744093560769748976233649221851799880599131620592031175370645284676468188384435930446526800550443125863880930654223434577055765818345706717500414322671614009121484412943387191286964099465289584394150711279902984613850405665319003550820411903390472009656831;
            6'd40: xpb[174] = 1024'd85980928344648409844842482189377711251317946958282665696106102461151018855330674123129241989980457605373755462773945316986275048716945611916346215199334043026623030580669147031885216702636418389243679479223643189704348725285906199934843956939309336252023356573377839182219133255946870047893133464070696659647;
            6'd41: xpb[174] = 1024'd97435453729573975695873463799473236488453277666669908648118644152553061477012126394458603380829294618716335554902605957504361712997960777305891879955542222172315406937903717008004615059566119278073036286833277257924284507184621112905588448589034278353335433243771064514032601192890189275374363537669383662463;
            6'd42: xpb[174] = 1024'd108889979114499541546904445409568761725588608375057151600131185843955104098693578665787964771678131632058915647031266598022448377278975942695437544711750401318007783295138286984124013416495820166902393094442911326144220289083336025876332940238759220454647509914164289845846069129833508502855593611268070665279;
            6'd43: xpb[174] = 1024'd120344504499425107397935427019664286962723939083444394552143727535357146720375030937117326162526968645401495739159927238540535041559991108084983209467958580463700159652372856960243411773425521055731749902052545394364156070982050938847077431888484162555959586584557515177659537066776827730336823684866757668095;
            6'd44: xpb[174] = 1024'd7732334200225931850167481224945379455160842666095953376024414161782294004747344298431616338718131349300926423831094444479557864999785938919368749207835718675701861440036209598732570938838016223250909101274939616219731002659869078852843353854979655390451759840833682479366476929791513940699363931839850186580;
            6'd45: xpb[174] = 1024'd19186859585151497701198462835040904692296173374483196328036955853184336626428796569760977729566968362643506515959755084997644529280801104308914413964043897821394237797270779574851969295767717112080265908884573684439666784558583991823587845504704597491763836511226907811179944866734833168180594005438537189396;
            6'd46: xpb[174] = 1024'd30641384970077063552229444445136429929431504082870439280049497544586379248110248841090339120415805375986086608088415725515731193561816269698460078720252076967086614154505349550971367652697418000909622716494207752659602566457298904794332337154429539593075913181620133142993412803678152395661824079037224192212;
            6'd47: xpb[174] = 1024'd42095910355002629403260426055231955166566834791257682232062039235988421869791701112419700511264642389328666700217076366033817857842831435088005743476460256112778990511739919527090766009627118889738979524103841820879538348356013817765076828804154481694387989852013358474806880740621471623143054152635911195028;
            6'd48: xpb[174] = 1024'd53550435739928195254291407665327480403702165499644925184074580927390464491473153383749061902113479402671246792345737006551904522123846600477551408232668435258471366868974489503210164366556819778568336331713475889099474130254728730735821320453879423795700066522406583806620348677564790850624284226234598197844;
            6'd49: xpb[174] = 1024'd65004961124853761105322389275423005640837496208032168136087122618792507113154605655078423292962316416013826884474397647069991186404861765867097072988876614404163743226209059479329562723486520667397693139323109957319409912153443643706565812103604365897012143192799809138433816614508110078105514299833285200660;
            6'd50: xpb[174] = 1024'd76459486509779326956353370885518530877972826916419411088099664310194549734836057926407784683811153429356406976603058287588077850685876931256642737745084793549856119583443629455448961080416221556227049946932744025539345694052158556677310303753329307998324219863193034470247284551451429305586744373431972203476;
            6'd51: xpb[174] = 1024'd87914011894704892807384352495614056115108157624806654040112206001596592356517510197737146074659990442698987068731718928106164514966892096646188402501292972695548495940678199431568359437345922445056406754542378093759281475950873469648054795403054250099636296533586259802060752488394748533067974447030659206292;
            6'd52: xpb[174] = 1024'd99368537279630458658415334105709581352243488333193896992124747692998634978198962469066507465508827456041567160860379568624251179247907262035734067257501151841240872297912769407687757794275623333885763562152012161979217257849588382618799287052779192200948373203979485133874220425338067760549204520629346209108;
            6'd53: xpb[174] = 1024'd110823062664556024509446315715805106589378819041581139944137289384400677599880414740395868856357664469384147252989040209142337843528922427425279732013709330986933248655147339383807156151205324222715120369761646230199153039748303295589543778702504134302260449874372710465687688362281386988030434594228033211924;
            6'd54: xpb[174] = 1024'd122277588049481590360477297325900631826514149749968382896149831075802720221561867011725230247206501482726727345117700849660424507809937592814825396769917510132625625012381909359926554508135025111544477177371280298419088821647018208560288270352229076403572526544765935797501156299224706215511664667826720214740;
            6'd55: xpb[174] = 1024'd9665417750282414812709351531181724318951053332619941720030517702227867505934180373039520423397664186626158029788868055599447331249732423649210936509794648344627326800045261998415713673547520279063636376593674520274663753324836348566054192318724569238064699801042103099208096162239392425874204914799812733225;
            6'd56: xpb[174] = 1024'd21119943135207980663740333141277249556086384041007184672043059393629910127615632644368881814246501199968738121917528696117533995530747589038756601266002827490319703157279831974535112030477221167892993184203308588494599535223551261536798683968449511339376776471435328431021564099182711653355434988398499736041;
            6'd57: xpb[174] = 1024'd32574468520133546514771314751372774793221714749394427624055601085031952749297084915698243205095338213311318214046189336635620659811762754428302266022211006636012079514514401950654510387406922056722349991812942656714535317122266174507543175618174453440688853141828553762835032036126030880836665061997186738857;
            6'd58: xpb[174] = 1024'd44028993905059112365802296361468300030357045457781670576068142776433995370978537187027604595944175226653898306174849977153707324092777919817847930778419185781704455871748971926773908744336622945551706799422576724934471099020981087478287667267899395542000929812221779094648499973069350108317895135595873741673;
            6'd59: xpb[174] = 1024'd55483519289984678216833277971563825267492376166168913528080684467836037992659989458356965986793012239996478398303510617671793988373793085207393595534627364927396832228983541902893307101266323834381063607032210793154406880919696000449032158917624337643313006482615004426461967910012669335799125209194560744489;
            6'd60: xpb[174] = 1024'd66938044674910244067864259581659350504627706874556156480093226159238080614341441729686327377641849253339058490432171258189880652654808250596939260290835544073089208586218111879012705458196024723210420414641844861374342662818410913419776650567349279744625083153008229758275435846955988563280355282793247747305;
            6'd61: xpb[174] = 1024'd78392570059835809918895241191754875741763037582943399432105767850640123236022894001015688768490686266681638582560831898707967316935823415986484925047043723218781584943452681855132103815125725612039777222251478929594278444717125826390521142217074221845937159823401455090088903783899307790761585356391934750121;
            6'd62: xpb[174] = 1024'd89847095444761375769926222801850400978898368291330642384118309542042165857704346272345050159339523280024218674689492539226053981216838581376030589803251902364473961300687251831251502172055426500869134029861112997814214226615840739361265633866799163947249236493794680421902371720842627018242815429990621752937;
            6'd63: xpb[174] = 1024'd101301620829686941620957204411945926216033698999717885336130851233444208479385798543674411550188360293366798766818153179744140645497853746765576254559460081510166337657921821807370900528985127389698490837470747066034150008514555652332010125516524106048561313164187905753715839657785946245724045503589308755753;
        endcase
    end

    always_comb begin
        case(flag[58][11:6])
            6'd0: xpb[175] = 1024'd0;
            6'd1: xpb[175] = 1024'd112756146214612507471988186022041451453169029708105128288143392924846251101067250815003772941037197306709378858946813820262227309778868912155121919315668260655858714015156391783490298885914828278527847645080381134254085790413270565302754617166249048149873389834581131085529307594729265473205275577187995758569;
            6'd2: xpb[175] = 1024'd101445596745100273545177444639268470161639632290474572448154930784715606864825362719992474667416720303975608310436134205945390778716517489755083713615005480378026753460741566229350358580312450835745497681773522422143810730605644357640530664649268647032926876255045204140952087115529897929291861327750397032807;
            6'd3: xpb[175] = 1024'd90135047275588039618366703256495488870110234872844016608166468644584962628583474624981176393796243301241837761925454591628554247654166067355045507914342700100194792906326740675210418274710073392963147718466663710033535670798018149978306712132288245915980362675509277196374866636330530385378447078312798307045;
            6'd4: xpb[175] = 1024'd78824497806075805691555961873722507578580837455213460768178006504454318392341586529969878120175766298508067213414774977311717716591814644955007302213679919822362832351911915121070477969107695950180797755159804997923260610990391942316082759615307844799033849095973350251797646157131162841465032828875199581283;
            6'd5: xpb[175] = 1024'd67513948336563571764745220490949526287051440037582904928189544364323674156099698434958579846555289295774296664904095362994881185529463222554969096513017139544530871797497089566930537663505318507398447791852946285812985551182765734653858807098327443682087335516437423307220425677931795297551618579437600855521;
            6'd6: xpb[175] = 1024'd56203398867051337837934479108176544995522042619952349088201082224193029919857810339947281572934812293040526116393415748678044654467111800154930890812354359266698911243082264012790597357902941064616097828546087573702710491375139526991634854581347042565140821936901496362643205198732427753638204330000002129759;
            6'd7: xpb[175] = 1024'd44892849397539103911123737725403563703992645202321793248212620084062385683615922244935983299314335290306755567882736134361208123404760377754892685111691578988866950688667438458650657052300563621833747865239228861592435431567513319329410902064366641448194308357365569418065984719533060209724790080562403403997;
            6'd8: xpb[175] = 1024'd33582299928026869984312996342630582412463247784691237408224157943931741447374034149924685025693858287572985019372056520044371592342408955354854479411028798711034990134252612904510716746698186179051397901932370149482160371759887111667186949547386240331247794777829642473488764240333692665811375831124804678235;
            6'd9: xpb[175] = 1024'd22271750458514636057502254959857601120933850367060681568235695803801097211132146054913386752073381284839214470861376905727535061280057532954816273710366018433203029579837787350370776441095808736269047938625511437371885311952260904004962997030405839214301281198293715528911543761134325121897961581687205952473;
            6'd10: xpb[175] = 1024'd10961200989002402130691513577084619829404452949430125728247233663670452974890257959902088478452904282105443922350697291410698530217706110554778068009703238155371069025422961796230836135493431293486697975318652725261610252144634696342739044513425438097354767618757788584334323281934957577984547332249607226711;
            6'd11: xpb[175] = 1024'd123717347203614909602679699599126071282573482657535254016390626588516704075957508774905861419490101588814822781297511111672925839996575022709899987325371498811229783040579353579721135021408259572014545620399033859515696042557905261645493661679674486247228157453338919669863630876664223051189822909437602985280;
            6'd12: xpb[175] = 1024'd112406797734102675675868958216353089991044085239904698176402164448386059839715620679894563145869624586081052232786831497356089308934223600309861781624708718533397822486164528025581194715805882129232195657092175147405420982750279053983269709162694085130281643873802992725286410397464855507276408660000004259518;
            6'd13: xpb[175] = 1024'd101096248264590441749058216833580108699514687822274142336413702308255415603473732584883264872249147583347281684276151883039252777871872177909823575924045938255565861931749702471441254410203504686449845693785316435295145922942652846321045756645713684013335130294267065780709189918265487963362994410562405533756;
            6'd14: xpb[175] = 1024'd89785698795078207822247475450807127407985290404643586496425240168124771367231844489871966598628670580613511135765472268722416246809520755509785370223383157977733901377334876917301314104601127243667495730478457723184870863135026638658821804128733282896388616714731138836131969439066120419449580161124806807994;
            6'd15: xpb[175] = 1024'd78475149325565973895436734068034146116455892987013030656436778027994127130989956394860668325008193577879740587254792654405579715747169333109747164522720377699901940822920051363161373798998749800885145767171599011074595803327400430996597851611752881779442103135195211891554748959866752875536165911687208082232;
            6'd16: xpb[175] = 1024'd67164599856053739968625992685261164824926495569382474816448315887863482894748068299849370051387716575145970038744113040088743184684817910709708958822057597422069980268505225809021433493396372358102795803864740298964320743519774223334373899094772480662495589555659284946977528480667385331622751662249609356470;
            6'd17: xpb[175] = 1024'd55854050386541506041815251302488183533397098151751918976459853747732838658506180204838071777767239572412199490233433425771906653622466488309670753121394817144238019714090400254881493187793994915320445840557881586854045683712148015672149946577792079545549075976123358002400308001468017787709337412812010630708;
            6'd18: xpb[175] = 1024'd44543500917029272115004509919715202241867700734121363136471391607602194422264292109826773504146762569678428941722753811455070122560115065909632547420732036866406059159675574700741552882191617472538095877251022874743770623904521808009925994060811678428602562396587431057823087522268650243795923163374411904946;
            6'd19: xpb[175] = 1024'd33232951447517038188193768536942220950338303316490807296482929467471550186022404014815475230526285566944658393212074197138233591497763643509594341720069256588574098605260749146601612576589240029755745913944164162633495564096895600347702041543831277311656048817051504113245867043069282699882508913936813179184;
            6'd20: xpb[175] = 1024'd21922401978004804261383027154169239658808905898860251456494467327340905949780515919804176956905808564210887844701394582821397060435412221109556136019406476310742138050845923592461672270986862586973395950637305450523220504289269392685478089026850876194709535237515577168668646563869915155969094664499214453422;
            6'd21: xpb[175] = 1024'd10611852508492570334572285771396258367279508481229695616506005187210261713538627824792878683285331561477117296190714968504560529373060798709517930318743696032910177496431098038321731965384485144191045987330446738412945444481643185023254136509870475077763021657979650224091426084670547612055680415061615727660;
            6'd22: xpb[175] = 1024'd123367998723105077806560471793437709820448538189334823904649398112056512814605878639796651624322528868186496155137528788766787839151929710864639849634411956688768891511587489821812030851299313422718893632410827872667031234894913750326008753676119523227636411492560781309620733679399813085260955992249611486229;
            6'd23: xpb[175] = 1024'd112057449253592843879749730410664728528919140771704268064660935971925868578363990544785353350702051865452725606626849174449951308089578288464601643933749176410936930957172664267672090545696935979936543669103969160556756175087287542663784801159139122110689897913024854365043513200200445541347541742812012760467;
            6'd24: xpb[175] = 1024'd100746899784080609952938989027891747237389743354073712224672473831795224342122102449774055077081574862718955058116169560133114777027226866064563438233086396133104970402757838713532150240094558537154193705797110448446481115279661335001560848642158720993743384333488927420466292721001077997434127493374414034705;
            6'd25: xpb[175] = 1024'd89436350314568376026128247645118765945860345936443156384684011691664580105880214354762756803461097859985184509605489945816278245964875443664525232532423615855273009848343013159392209934492181094371843742490251736336206055472035127339336896125178319876796870753953000475889072241801710453520713243936815308943;
            6'd26: xpb[175] = 1024'd78125800845056142099317506262345784654330948518812600544695549551533935869638326259751458529840620857251413961094810331499441714902524021264487026831760835577441049293928187605252269628889803651589493779183393024225930995664408919677112943608197918759850357174417073531311851762602342909607298994499216583181;
            6'd27: xpb[175] = 1024'd66815251375543908172506764879572803362801551101182044704707087411403291633396438164740160256220143854517643412584130717182605183840172598864448821131098055299609088739513362051112329323287426208807143815876534312115655935856782712014888991091217517642903843594881146586734631283402975365693884745061617857419;
            6'd28: xpb[175] = 1024'd55504701906031674245696023496799822071272153683551488864718625271272647397154550069728861982599666851783872864073451102865768652777821176464410615430435275021777128185098536496972389017685048766024793852569675600005380876049156504352665038574237116525957330015345219642157410804203607821780470495624019131657;
            6'd29: xpb[175] = 1024'd44194152436519440318885282114026840779742756265920933024730163131142003160912661974717563708979189849050102315562771488548932121715469754064372409729772494743945167630683710942832448712082671323242443889262816887895105816241530296690441086057256715409010816435809292697580190325004240277867056246186420405895;
            6'd30: xpb[175] = 1024'd32883602967007206392074540731253859488213358848290377184741700991011358924670773879706265435358712846316331767052091874232095590653118331664334204029109714466113207076268885388692508406480293880460093925955958175784830756433904089028217133540276314292064302856273365753002969845804872733953641996748821680133;
            6'd31: xpb[175] = 1024'd21573053497494972465263799348480878196683961430659821344753238850880714688428885784694967161738235843582561218541412259915259059590766909264295998328446934188281246521854059834552568100877916437677743962649099463674555696626277881365993181023295913175117789276737438808425749366605505190040227747311222954371;
            6'd32: xpb[175] = 1024'd10262504027982738538453057965707896905154564013029265504764776710750070452186997689683668888117758840848790670030732645598422528528415486864257792627784153910449285967439234280412627795275538994895393999342240751564280636818651673703769228506315512058171275697201511863848528887406137646126813497873624228609;
            6'd33: xpb[175] = 1024'd123018650242595246010441243987749348358323593721134393792908169635596321553254248504687441829154956147558169528977546465860649838307284399019379711943452414566307999982595626063902926681190367273423241644422621885818366427231922239006523845672564560208044665531782642949377836482135403119332089075061619987178;
            6'd34: xpb[175] = 1024'd111708100773083012083630502604976367066794196303503837952919707495465677317012360409676143555534479144824398980466866851543813307244932976619341506242789634288476039428180800509762986375587989830640891681115763173708091367424296031344299893155584159091098151952246716004800616002936035575418674825624021261416;
            6'd35: xpb[175] = 1024'd100397551303570778156819761222203385775264798885873282112931245355335033080770472314664845281914002142090628431956187237226976776182581554219303300542126854010644078873765974955623046069985612387858541717808904461597816307616669823682075940638603757974151638372710789060223395523736668031505260576186422535654;
            6'd36: xpb[175] = 1024'd89087001834058544230009019839430404483735401468242726272942783215204388844528584219653547008293525139356857883445507622910140245120230131819265094841464073732812118319351149401483105764383234945076191754502045749487541247809043616019851988121623356857205124793174862115646175044537300487591846326748823809892;
            6'd37: xpb[175] = 1024'd77776452364546310303198278456657423192206004050612170432954321075073744608286696124642248734673048136623087334934828008593303714057878709419226889140801293454980157764936323847343165458780857502293841791195187037377266188001417408357628035604642955740258611213638935171068954565337932943678432077311225084130;
            6'd38: xpb[175] = 1024'd66465902895034076376387537073884441900676606632981614592965858934943100372044808029630950461052571133889316786424148394276467182995527287019188683440138513177148197210521498293203225153178480059511491827888328325266991128193791200695404083087662554623312097634103008226491734086138565399765017827873626358368;
            6'd39: xpb[175] = 1024'd55155353425521842449576795691111460609147209215351058752977396794812456135802919934619652187432094131155546237913468779959630651933175864619150477739475732899316236656106672739063284847576102616729141864581469613156716068386164993033180130570682153506365584054567081281914513606939197855851603578436027632606;
            6'd40: xpb[175] = 1024'd43844803956009608522766054308338479317617811797720502912988934654681811899561031839608353913811617128421775689402789165642794120870824442219112272038812952621484276101691847184923344541973725173946791901274610901046441008578538785370956178053701752389419070475031154337337293127739830311938189328998428906844;
            6'd41: xpb[175] = 1024'd32534254486497374595955312925565498026088414380089947073000472514551167663319143744597055640191140125688005140892109551325957589808473019819074066338150172343652315547277021630783404236371347731164441937967752188936165948770912577708732225536721351272472556895495227392760072648540462768024775079560830181082;
            6'd42: xpb[175] = 1024'd21223705016985140669144571542792516734559016962459391233012010374420523427077255649585757366570663122954234592381429937009121058746121597419035860637487392065820354992862196076643463930768970288382091974660893476825890888963286370046508273019740950155526043315959300448182852169341095224111360830123231455320;
            6'd43: xpb[175] = 1024'd9913155547472906742333830160019535443029619544828835393023548234289879190835367554574459092950186120220464043870750322692284527683770175018997654936824611787988394438447370522503523625166592845599742011354034764715615829155660162384284320502760549038579529736423373503605631690141727680197946580685632729558;
            6'd44: xpb[175] = 1024'd122669301762085414214322016182060986896198649252933963681166941159136130291902618369578232033987383426929842902817564142954511837462639087174119574252492872443847108453603762305993822511081421124127589656434415898969701619568930727687038937669009597188452919571004504589134939284870993153403222157873628488127;
            6'd45: xpb[175] = 1024'd111358752292573180287511274799288005604669251835303407841178479019005486055660730274566933760366906424196072354306884528637675306400287664774081368551830092166015147899188936751853882205479043681345239693127557186859426559761304520024814985152029196071506405991468577644557718805671625609489807908436029762365;
            6'd46: xpb[175] = 1024'd100048202823060946360700533416515024313139854417672852001190016878874841819418842179555635486746429421462301805796204914320838775337936242374043162851167311888183187344774111197713941899876666238562889729820698474749151499953678312362591032635048794954559892411932650699980498326472258065576393658998431036603;
            6'd47: xpb[175] = 1024'd88737653353548712433889792033742043021610457000042296161201554738744197583176954084544337213125952418728531257285525300004002244275584819974004957150504531610351226790359285643574001594274288795780539766513839762638876440146052104700367080118068393837613378832396723755403277847272890521662979409560832310841;
            6'd48: xpb[175] = 1024'd77427103884036478507079050650969061730081059582411740321213092598613553346935065989533038939505475415994760708774845685687165713213233397573966751449841751332519266235944460089434061288671911352998189803206981050528601380338425897038143127601087992720666865252860796810826057368073522977749565160123233585079;
            6'd49: xpb[175] = 1024'd66116554414524244580268309268196080438551662164781184481224630458482909110693177894521740665884998413260990160264166071370329182150881975173928545749178971054687305681529634535294120983069533910215839839900122338418326320530799689375919175084107591603720351673324869866248836888874155433836150910685634859317;
            6'd50: xpb[175] = 1024'd54806004945012010653457567885423099147022264747150628641236168318352264874451289799510442392264521410527219611753486457053492651088530552773890340048516190776855345127114808981154180677467156467433489876593263626308051260723173481713695222567127190486773838093788942921671616409674787889922736661248036133555;
            6'd51: xpb[175] = 1024'd43495455475499776726646826502650117855492867329520072801247706178221620638209401704499144118644044407793449063242806842736656120026179130373852134347853410499023384572699983427014240371864779024651139913286404914197776200915547274051471270050146789369827324514253015977094395930475420346009322411810437407793;
            6'd52: xpb[175] = 1024'd32184906005987542799836085119877136563963469911889516961259244038090976401967513609487845845023567405059678514732127228419819588963827707973813928647190630221191424018285157872874300066262401581868789949979546202087501141107921066389247317533166388252880810934717089032517175451276052802095908162372838682031;
            6'd53: xpb[175] = 1024'd20874356536475308873025343737104155272434072494258961121270781897960332165725625514476547571403090402325907966221447614102983057901476285573775722946527849943359463463870332318734359760660024139086439986672687489977226081300294858727023365016185987135934297355181162087939954972076685258182493912935239956269;
            6'd54: xpb[175] = 1024'd9563807066963074946214602354331173980904675076628405281282319757829687929483737419465249297782613399592137417710767999786146526839124863173737517245865069665527502909455506764594419455057646696304090023365828777866951021492668651064799412499205586018987783775645235143362734492877317714269079663497641230507;
            6'd55: xpb[175] = 1024'd122319953281575582418202788376372625434073704784733533569425712682675939030550988234469022238819810706301516276657581820048373836617993775328859436561533330321386216924611898548084718340972474974831937668446209912121036811905939216367554029665454634168861173610226366228892042087606583187474355240685636989076;
            6'd56: xpb[175] = 1024'd111009403812063348491392046993599644142544307367102977729437250542545294794309100139457723965199333703567745728146902205731537305555642352928821230860870550043554256370197072993944778035370097532049587705139351200010761752098313008705330077148474233051914660030690439284314821608407215643560940991248038263314;
            6'd57: xpb[175] = 1024'd99698854342551114564581305610826662851014909949472421889448788402414650558067212044446425691578856700833975179636222591414700774493290930528783025160207769765722295815782247439804837729767720089267237741832492487900486692290686801043106124631493831934968146451154512339737601129207848099647526741810439537552;
            6'd58: xpb[175] = 1024'd88388304873038880637770564228053681559485512531841866049460326262284006321825323949435127417958379698100204631125542977097864243430939508128744819459544989487890335261367421885664897424165342646484887778525633775790211632483060593380882172114513430818021632871618585395160380650008480555734112492372840811790;
            6'd59: xpb[175] = 1024'd77077755403526646710959822845280700267956115114211310209471864122153362085583435854423829144337902695366434082614863362781027712368588085728706613758882209210058374706952596331524957118562965203702537815218775063679936572675434385718658219597533029701075119292082658450583160170809113011820698242935242086028;
            6'd60: xpb[175] = 1024'd65767205934014412784149081462507718976426717696580754369483401982022717849341547759412530870717425692632663534104183748464191181306236663328668408058219428932226414152537770777385016812960587760920187851911916351569661512867808178056434267080552628584128605712546731506005939691609745467907283993497643360266;
            6'd61: xpb[175] = 1024'd54456656464502178857338340079734737684897320278950198529494939841892073613099659664401232597096948689898892985593504134147354650243885240928630202357556648654394453598122945223245076507358210318137837888605057639459386453060181970394210314563572227467182092133010804561428719212410377923993869744060044634504;
            6'd62: xpb[175] = 1024'd43146106994989944930527598696961756393367922861319642689506477701761429376857771569389934323476471687165122437082824519830518119181533818528591996656893868376562493043708119669105136201755832875355487925298198927349111393252555762731986362046591826350235578553474877616851498733211010380080455494622445908742;
            6'd63: xpb[175] = 1024'd31835557525477711003716857314188775101838525443689086849518015561630785140615883474378636049855994684431351888572144905513681588119182396128553790956231088098730532489293294114965195896153455432573137961991340215238836333444929555069762409529611425233289064973938950672274278254011642836167041245184847182980;
        endcase
    end

    always_comb begin
        case(flag[58][16:12])
            5'd0: xpb[176] = 1024'd0;
            5'd1: xpb[176] = 1024'd20525008055965477076906115931415793810309128026058531009529553421500140904373995379367337776235517681697581340061465291196845057056830973728515585255568307820898571934878468560825255590551077989790787998684481503128561273637303347407538457012631024116342551394403023727697057774812275292253626995747248457218;
            5'd2: xpb[176] = 1024'd41050016111930954153812231862831587620618256052117062019059106843000281808747990758734675552471035363395162680122930582393690114113661947457031170511136615641797143869756937121650511181102155979581575997368963006257122547274606694815076914025262048232685102788806047455394115549624550584507253991494496914436;
            5'd3: xpb[176] = 1024'd61575024167896431230718347794247381430927384078175593028588660264500422713121986138102013328706553045092744020184395873590535171170492921185546755766704923462695715804635405682475766771653233969372363996053444509385683820911910042222615371037893072349027654183209071183091173324436825876760880987241745371654;
            5'd4: xpb[176] = 1024'd82100032223861908307624463725663175241236512104234124038118213686000563617495981517469351104942070726790325360245861164787380228227323894914062341022273231283594287739513874243301022362204311959163151994737926012514245094549213389630153828050524096465370205577612094910788231099249101169014507982988993828872;
            5'd5: xpb[176] = 1024'd102625040279827385384530579657078969051545640130292655047647767107500704521869976896836688881177588408487906700307326455984225285284154868642577926277841539104492859674392342804126277952755389948953939993422407515642806368186516737037692285063155120581712756972015118638485288874061376461268134978736242286090;
            5'd6: xpb[176] = 1024'd123150048335792862461436695588494762861854768156351186057177320529000845426243972276204026657413106090185488040368791747181070342340985842371093511533409846925391431609270811364951533543306467938744727992106889018771367641823820084445230742075786144698055308366418142366182346648873651753521761974483490743308;
            5'd7: xpb[176] = 1024'd19608360707633598139543884115096123927465469056674032938575018885524090993308828745556293218990949462439919972972763603798851558556596481544448971772647113812599328974578062588146549942340340207225318382404130675535568065240226658887790629405187719547577956346704108063772876349757294028656699143605144716195;
            5'd8: xpb[176] = 1024'd40133368763599075216450000046511917737774597082732563948104572307024231897682824124923630995226467144137501313034228894995696615613427455272964557028215421633497900909456531148971805532891418197016106381088612178664129338877530006295329086417818743663920507741107131791469934124569569320910326139352393173413;
            5'd9: xpb[176] = 1024'd60658376819564552293356115977927711548083725108791094957634125728524372802056819504290968771461984825835082653095694186192541672670258429001480142283783729454396472844334999709797061123442496186806894379773093681792690612514833353702867543430449767780263059135510155519166991899381844613163953135099641630631;
            5'd10: xpb[176] = 1024'd81183384875530029370262231909343505358392853134849625967163679150024513706430814883658306547697502507532663993157159477389386729727089402729995727539352037275295044779213468270622316713993574176597682378457575184921251886152136701110406000443080791896605610529913179246864049674194119905417580130846890087849;
            5'd11: xpb[176] = 1024'd101708392931495506447168347840759299168701981160908156976693232571524654610804810263025644323933020189230245333218624768586231786783920376458511312794920345096193616714091936831447572304544652166388470377142056688049813159789440048517944457455711816012948161924316202974561107449006395197671207126594138545067;
            5'd12: xpb[176] = 1024'd122233400987460983524074463772175092979011109186966687986222785993024795515178805642392982100168537870927826673280090059783076843840751350187026898050488652917092188648970405392272827895095730156179258375826538191178374433426743395925482914468342840129290713318719226702258165223818670489924834122341387002285;
            5'd13: xpb[176] = 1024'd18691713359301719202181652298776454044621810087289534867620484349548041082243662111745248661746381243182258605884061916400858060056361989360382358289725919804300086014277656615467844294129602424659848766123779847942574856843149970368042801797744414978813361299005192399848694924702312765059771291463040975172;
            5'd14: xpb[176] = 1024'd39216721415267196279087768230192247854930938113348065877150037771048181986617657491112586437981898924879839945945527207597703117113192963088897943545294227625198657949156125176293099884680680414450636764808261351071136130480453317775581258810375439095155912693408216127545752699514588057313398287210289432390;
            5'd15: xpb[176] = 1024'd59741729471232673355993884161608041665240066139406596886679591192548322890991652870479924214217416606577421286006992498794548174170023936817413528800862535446097229884034593737118355475231758404241424763492742854199697404117756665183119715823006463211498464087811239855242810474326863349567025282957537889608;
            5'd16: xpb[176] = 1024'd80266737527198150432900000093023835475549194165465127896209144614048463795365648249847261990452934288275002626068457789991393231226854910545929114056430843266995801818913062297943611065782836394032212762177224357328258677755060012590658172835637487327841015482214263582939868249139138641820652278704786346826;
            5'd17: xpb[176] = 1024'd100791745583163627509806116024439629285858322191523658905738698035548604699739643629214599766688451969972583966129923081188238288283685884274444699311999151087894373753791530858768866656333914383823000760861705860456819951392363359998196629848268511444183566876617287310636926023951413934074279274452034804044;
            5'd18: xpb[176] = 1024'd121316753639129104586712231955855423096167450217582189915268251457048745604113639008581937542923969651670165306191388372385083345340516858002960284567567458908792945688669999419594122246884992373613788759546187363585381225029666707405735086860899535560526118271020311038333983798763689226327906270199283261262;
            5'd19: xpb[176] = 1024'd17775066010969840264819420482456784161778151117905036796665949813571991171178495477934204104501813023924597238795360229002864561556127497176315744806804725796000843053977250642789138645918864642094379149843429020349581648446073281848294974190301110410048766251306276735924513499647331501462843439320937234149;
            5'd20: xpb[176] = 1024'd38300074066935317341725536413872577972087279143963567806195503235072132075552490857301541880737330705622178578856825520199709618612958470904831330062373033616899414988855719203614394236469942631885167148527910523478142922083376629255833431202932134526391317645709300463621571274459606793716470435068185691367;
            5'd21: xpb[176] = 1024'd58825082122900794418631652345288371782396407170022098815725056656572272979926486236668879656972848387319759918918290811396554675669789444633346915317941341437797986923734187764439649827021020621675955147212392026606704195720679976663371888215563158642733869040112324191318629049271882085970097430815434148585;
            5'd22: xpb[176] = 1024'd79350090178866271495537768276704165592705535196080629825254610078072413884300481616036217433208366069017341258979756102593399732726620418361862500573509649258696558858612656325264905417572098611466743145896873529735265469357983324070910345228194182759076420434515347919015686824084157378223724426562682605803;
            5'd23: xpb[176] = 1024'd99875098234831748572443884208119959403014663222139160834784163499572554788674476995403555209443883750714922599041221393790244789783451392090378085829077957079595130793491124886090161008123176601257531144581355032863826742995286671478448802240825206875418971828918371646712744598896432670477351422309931063021;
            5'd24: xpb[176] = 1024'd120400106290797225649350000139535753213323791248197691844313716921072695693048472374770892985679401432412503939102686684987089846840282365818893671084646264900493702728369593446915416598674254591048319143265836535992388016632590018885987259253456230991761523223321395374409802373708707962730978418057179520239;
            5'd25: xpb[176] = 1024'd16858418662637961327457188666137114278934492148520538725711415277595941260113328844123159547257244804666935871706658541604871063055893004992249131323883531787701600093676844670110432997708126859528909533563078192756588440048996593328547146582857805841284171203607361072000332074592350237865915587178833493126;
            5'd26: xpb[176] = 1024'd37383426718603438404363304597552908089243620174579069735240968699096082164487324223490497323492762486364517211768123832801716120112723978720764716579451839608600172028555313230935688588259204849319697532247559695885149713686299940736085603595488829957626722598010384799697389849404625530119542582926081950344;
            5'd27: xpb[176] = 1024'd57908434774568915481269420528968701899552748200637600744770522120596223068861319602857835099728280168062098551829589123998561177169554952449280301835020147429498743963433781791760944178810282839110485530932041199013710987323603288143624060608119854073969273992413408527394447624216900822373169578673330407562;
            5'd28: xpb[176] = 1024'd78433442830534392558175536460384495709861876226696131754300075542096363973235314982225172875963797849759679891891054415195406234226385926177795887090588455250397315898312250352586199769361360828901273529616522702142272260960906635551162517620750878190311825386816432255091505399029176114626796574420578864780;
            5'd29: xpb[176] = 1024'd98958450886499869635081652391800289520171004252754662763829628963596504877609310361592510652199315531457261231952519706392251291283216899906311472346156763071295887833190718913411455359912438818692061528301004205270833534598209982958700974633381902306654376781219455982788563173841451406880423570167827321998;
            5'd30: xpb[176] = 1024'd119483458942465346711987768323216083330480132278813193773359182385096645781983305740959848428434833213154842572013984997589096348340047873634827057601725070892194459768069187474236710950463516808482849526985485708399394808235513330366239431646012926422996928175622479710485620948653726699134050565915075779216;
            5'd31: xpb[176] = 1024'd15941771314306082390094956849817444396090833179136040654756880741619891349048162210312114990012676585409274504617956854206877564555658512808182517840962337779402357133376438697431727349497389076963439917282727365163595231651919904808799318975414501272519576155908445408076150649537368974268987735036729752103;
        endcase
    end

    always_comb begin
        case(flag[59][5:0])
            6'd0: xpb[177] = 1024'd0;
            6'd1: xpb[177] = 1024'd80266737527198150432900000093023835475549194165465127896209144614048463795365648249847261990452934288275002626068457789991393231226854910545929114056430843266995801818913062297943611065782836394032212762177224357328258677755060012590658172835637487327841015482214263582939868249139138641820652278704786346826;
            6'd2: xpb[177] = 1024'd36466779370271559467001072781233238206399961205194571664286434163120032253422157589679452766248194267106855844679422145403722621612489486536698103096530645600300929068254907258256982940048467066754227915967208868292156505289223252216337775988045525388862127550311469135773208424349644266522614730783978209321;
            6'd3: xpb[177] = 1024'd116733516897469709899901072874257073681949155370659699560495578777168496048787805839526714756701128555381858470747879935395115852839344397082627217152961488867296730887167969556200594005831303460786440678144433225620415183044283264806995948823683012716703143032525732718713076673488782908343267009488764556147;
            6'd4: xpb[177] = 1024'd72933558740543118934002145562466476412799922410389143328572868326240064506844315179358905532496388534213711689358844290807445243224978973073396206193061291200601858136509814516513965880096934133508455831934417736584313010578446504432675551976091050777724255100622938271546416848699288533045229461567956418642;
            6'd5: xpb[177] = 1024'd29133600583616527968103218250675879143650689450118587096650157875311632964900824519191096308291648513045564907969808646219774633610613549064165195233161093533906985385851659476827337754362564806230470985724402247548210838112609744058355155128499088838745367168720143824379757023909794157747191913647148281137;
            6'd6: xpb[177] = 1024'd109400338110814678401003218343699714619199883615583714992859302489360096760266472769038358298744582801320567534038266436211167864837468459610094309289591936800902787204764721774770948820145401200262683747901626604876469515867669756649013327964136576166586382650934407407319625273048932799567844192351934627963;
            6'd7: xpb[177] = 1024'd65600379953888087435104291031909117350050650655313158760936592038431665218322982108870549074539842780152420752649230791623497255223103035600863298329691739134207914454106566735084320694411031872984698901691611115840367343401832996274692931116544614227607494719031612960152965448259438424269806644431126490458;
            6'd8: xpb[177] = 1024'd21800421796961496469205363720118520080901417695042602529013881587503233676379491448702739850335102758984273971260195147035826645608737611591632287369791541467513041703448411695397692568676662545706714055481595626804265170935996235900372534268952652288628606787128818512986305623469944048971769096510318352953;
            6'd9: xpb[177] = 1024'd102067159324159646902105363813142355556450611860507730425223026201551697471745139698550001840788037047259276597328652937027219876835592522137561401426222384734508843522361473993341303634459498939738926817658819984132523848691056248491030707104590139616469622269343082095926173872609082690792421375215104699779;
            6'd10: xpb[177] = 1024'd58267201167233055936206436501351758287301378900237174193300315750623265929801649038382192616583297026091129815939617292439549267221227098128330390466322187067813970771703318953654675508725129612460941971448804495096421676225219488116710310256998177677490734337440287648759514047819588315494383827294296562274;
            6'd11: xpb[177] = 1024'd14467243010306464970307509189561161018152145939966617961377605299694834387858158378214383392378557004922983034550581647851878657606861674119099379506421989401119098021045163913968047382990760285182957125238789006060319503759382727742389913409406215738511846405537493201592854223030093940196346279373488424769;
            6'd12: xpb[177] = 1024'd94733980537504615403207509282584996493701340105431745857586749913743298183223806628061645382831491293197985660619039437843271888833716584665028493562852832668114899839958226211911658448773596679215169887416013363388578181514442740333048086245043703066352861887751756784532722472169232582016998558078274771595;
            6'd13: xpb[177] = 1024'd50934022380578024437308581970794399224552107145161189625664039462814866641280315967893836158626751272029838879230003793255601279219351160655797482602952635001420027089300071172225030323039227351937185041205997874352476009048605979958727689397451741127373973955848962337366062647379738206718961010157466634090;
            6'd14: xpb[177] = 1024'd7134064223651433471409654659003801955402874184890633393741329011886435099336825307726026934422011250861692097840968148667930669604985736646566471643052437334725154338641916132538402197304858024659200194995982385316373836582769219584407292549859779188395086023946167890199402822590243831420923462236658496585;
            6'd15: xpb[177] = 1024'd87400801750849583904309654752027637430952068350355761289950473625934898894702473557573288924874945539136694723909425938659323900831840647192495585699483280601720956157554978430482013263087694418691412957173206742644632514337829232175065465385497266516236101506160431473139271071729382473241575740941444843411;
            6'd16: xpb[177] = 1024'd43600843593922992938410727440237040161802835390085205058027763175006467352758982897405479700670205517968547942520390294071653291217475223183264574739583082935026083406896823390795385137353325091413428110963191253608530341871992471800745068537905304577257213574257637025972611246939888097943538193020636705906;
            6'd17: xpb[177] = 1024'd123867581121121143371310727533260875637352029555550332954236907789054931148124631147252741691123139806243550568588848084063046522444330133729193688796013926202021885225809885688738996203136161485445640873140415610936789019627052484391403241373542791905098229056471900608912479496079026739764190471725423052732;
            6'd18: xpb[177] = 1024'd80067622964194552405411800221470278368202796595279776722314197338126499606181140487084932466918399785075403787199812439475375912829964709719962677836113728535327012475151730649052368077401792158167656026930400121900686847161215724017082844525950829966119341124569106161745819671289532364466152923804614915227;
            6'd19: xpb[177] = 1024'd36267664807267961439512872909679681099053563635009220490391486887198068064237649826917123242713659763907257005810776794887705303215599285710731666876213530868632139724493575609365739951667422830889671180720384632864584674695378963642762447678358868027140453192666311714579159846500037989168115375883806777722;
            6'd20: xpb[177] = 1024'd116534402334466111872412873002703516574602757800474348386600631501246531859603298076764385233166594052182259631879234584879098534442454196256660780932644374135627941543406637907309351017450259224921883942897608990192843352450438976233420620513996355354981468674880575297519028095639176630988767654588593124548;
            6'd21: xpb[177] = 1024'd72734444177539520906513945690912919305453524840203792154677921050318100317659807416596576008961854031014112850490198940291427924828088772247429769972744176468933068792748482867622722891715889897643899096687593501156741179984602215859100223666404393416002580742977780850352368270849682255690730106667784987043;
            6'd22: xpb[177] = 1024'd28934486020612929940615018379122322036304291879933235922755210599389668775716316756428766784757114009845966069101163295703757315213723348238198759012843978802238196042090327827936094765981520570365914250477578012120639007518765455484779826818812431477023692811074986403185708446060187880392692558746976849538;
            6'd23: xpb[177] = 1024'd109201223547811080373515018472146157511853486045398363818964355213438132571081965006276028775210048298120968695169621085695150546440578258784127873069274822069233997861003390125879705831764356964398127012654802369448897685273825468075437999654449918804864708293289249986125576695199326522213344837451763196364;
            6'd24: xpb[177] = 1024'd65401265390884489407616091160355560242704253085127807587041644762509701029138474346108219551005308276952821913780585441107479936826212834774896862109374624402539125110345235086193077706029987637120142166444786880412795512807988707701117602806857956865885820361386455538958916870409832146915307289530955058859;
            6'd25: xpb[177] = 1024'd21601307233957898441717163848564962973555020124857251355118934311581269487194983685940410326800568255784675132391549796519809327211847410765665851149474426735844252359687080046506449580295618309842157320234771391376693340342151947326797205959265994926906932429483661091792257045620337771617269741610146921354;
            6'd26: xpb[177] = 1024'd101868044761156048874617163941588798449104214290322379251328078925629733282560631935787672317253502544059677758460007586511202558438702321311594965205905270002840054178600142344450060646078454703874370082411995748704952018097211959917455378794903482254747947911697924674732125294759476413437922020314933268180;
            6'd27: xpb[177] = 1024'd58068086604229457908718236629798201179954981330051823019405368474701301740617141275619863093048762522891530977070971941923531948824336897302363954246005072336145181427941987304763432520344085376596385236201980259668849845631375199543134981947311520315769059979795130227565465469969982038139884472394125130675;
            6'd28: xpb[177] = 1024'd14268128447302866942819309318007603910805748369781266787482658023772870198673650615452053868844022501723384195681936297335861339209971473293132943286104874669450308677283832265076804394609716049318400389991964770632747673165538439168814585099719558376790172047892335780398805645180487662841846924473316993170;
            6'd29: xpb[177] = 1024'd94534865974501017375719309411031439386354942535246394683691802637821333994039298865299315859296956789998386821750394087327254570436826383839062057342535717936446110496196894563020415460392552443350613152169189127961006350920598451759472757935357045704631187530106599363338673894319626304662499203178103339996;
            6'd30: xpb[177] = 1024'd50734907817574426409820382099240842117205709574975838451769092186892902452095808205131506635092216768830240040361358442739583960822460959829831046382635520269751237745538739523333787334658183116072628305959173638924904178454761691385152361087765083765652299598203804916172014069530131929364461655257295202491;
            6'd31: xpb[177] = 1024'd6934949660647835443921454787450244848056476614705282219846381735964470910152317544963697410887476747662093258972322798151913351208095535820600035422735322603056364994880584483647159208923813788794643459749158149888802005988924931010831964240173121826673411666301010469005354244740637554066424107336487064986;
            6'd32: xpb[177] = 1024'd87201687187845985876821454880474080323605670780170410116055526350012934705517965794810959401340411035937095885040780588143306582434950446366529149479166165870052166813793646781590770274706650182826856221926382507217060683743984943601490137075810609154514427148515274051945222493879776195887076386041273411812;
            6'd33: xpb[177] = 1024'd43401729030919394910922527568683483054456437819899853884132815899084503163574475134643150177135671014768949103651744943555635972820585022357298138519265968203357294063135491741904142148972280855548871375716367018180958511278148183227169740228218647215535539216612479604778562669090281820589038838120465274307;
            6'd34: xpb[177] = 1024'd123668466558117545343822527661707318530005631985364981780341960513132966958940123384490412167588605303043951729720202733547029204047439932903227252575696811470353095882048554039847753214755117249581084137893591375509217189033208195817827913063856134543376554698826743187718430918229420462409691116825251621133;
            6'd35: xpb[177] = 1024'd79868508401190954377923600349916721260856399025094425548419250062204535416996632724322602943383865281875804948331167088959358594433074508893996241615796613803658223131390399000161125089020747922303099291683575886473115016567371435443507516216264172604397666766923948740551771093439926087111653568904443483628;
            6'd36: xpb[177] = 1024'd36068550244264363412024673038126123991707166064823869316496539611276103875053142064154793719179125260707658166942131444371687984818709084884765230655896416136963350380732243960474496963286378595025114445473560397437012844101534675069187119368672210665418778835021154293385111268650431711813616020983635346123;
            6'd37: xpb[177] = 1024'd116335287771462513844924673131149959467256360230288997212705684225324567670418790314002055709632059548982660793010589234363081216045563995430694344712327259403959152199645306258418108029069214989057327207650784754765271521856594687659845292204309697993259794317235417876324979517789570353634268299688421692949;
            6'd38: xpb[177] = 1024'd72535329614535922879025745819359362198107127270018440980782973774396136128475299653834246485427319527814514011621553589775410606431198571421463333752427061737264279448987151218731479903334845661779342361440769265729169349390757927285524895356717736054280906385332623429158319693000075978336230751767613555444;
            6'd39: xpb[177] = 1024'd28735371457609331913126818507568764928957894309747884748860263323467704586531808993666437261222579506646367230232517945187739996816833147412232322792526864070569406698328996179044851777600476334501357515230753776693067176924921166911204498509125774115302018453429828981991659868210581603038193203846805417939;
            6'd40: xpb[177] = 1024'd109002108984807482346026818600592600404507088475213012645069407937516168381897457243513699251675513794921369856300975735179133228043688057958161436848957707337565208517242058476988462843383312728533570277407978134021325854679981179501862671344763261443143033935644092564931528117349720244858845482551591764765;
            6'd41: xpb[177] = 1024'd65202150827880891380127891288802003135357855514942456413146697486587736839953966583345890027470773773753223074911940090591462618429322633948930425889057509670870335766583903437301834717648943401255585431197962644985223682214144419127542274497171299504164146003741298117764868292560225869560807934630783627260;
            6'd42: xpb[177] = 1024'd21402192670954300414228963977011405866208622554671900181223987035659305298010475923178080803266033752585076293522904446003792008814957209939699414929157312004175463015925748397615206591914574073977600584987947155949121509748307658753221877649579337565185258071838503670598208467770731494262770386709975489755;
            6'd43: xpb[177] = 1024'd101668930198152450847128964070035241341757816720137028077433131649707769093376124173025342793718968040860078919591362235995185240041812120485628528985588155271171264834838810695558817657697410468009813347165171513277380187503367671343880050485216824893026273554052767253538076716909870136083422665414761836581;
            6'd44: xpb[177] = 1024'd57868972041225859881230036758244644072608583759866471845510421198779337551432633512857533569514228019691932138202326591407514630427446696476397518025687957604476392084180655655872189531963041140731828500955156024241278015037530910969559653637624862954047385622149972806371416892120375760785385117493953699076;
            6'd45: xpb[177] = 1024'd14069013884299268915331109446454046803459350799595915613587710747850906009489142852689724345309487998523785356813290946819844020813081272467166507065787759937781519333522500616185561406228671813453843654745140535205175842571694150595239256790032901015068497690247178359204757067330881385487347569573145561571;
            6'd46: xpb[177] = 1024'd94335751411497419348231109539477882279008544965061043509796855361899369804854791102536986335762422286798787982881748736811237252039936183013095621122218603204777321152435562914129172472011508207486056416922364892533434520326754163185897429625670388342909513172461441942144625316470020027307999848277931908397;
            6'd47: xpb[177] = 1024'd50535793254570828382332182227687285009859312004790487277874144910970938262911300442369177111557682265630641201492713092223566642425570759003864610162318405538082448401777407874442544346277138880208071570712349403497332347860917402811577032778078426403930625240558647494977965491680525652009962300357123770892;
            6'd48: xpb[177] = 1024'd6735835097644237416433254915896687740710079044519931045951434460042506720967809782201367887352942244462494420103677447635896032811205334994633599202418207871387575651119252834755916220542769552930086724502333914461230175395080642437256635930486464464951737308655853047811305666891031276711924752436315633387;
            6'd49: xpb[177] = 1024'd87002572624842387849333255008920523216259273209985058942160579074090970516333458032048629877805876532737497046172135237627289264038060245540562713258849051138383377470032315132699527286325605946962299486679558271789488853150140655027914808766123951792792752790870116630751173916030169918532577031141101980213;
            6'd50: xpb[177] = 1024'd43202614467915796883434327697129925947110040249714502710237868623162538974389967371880820653601136511569350264783099593039618654423694821531331702298948853471688504719374160093012899160591236619684314640469542782753386680684303894653594411918531989853813864858967322183584514091240675543234539483220293842708;
            6'd51: xpb[177] = 1024'd123469351995113947316334327790153761422659234415179630606447013237211002769755615621728082644054070799844352890851557383031011885650549732077260816355379696738684306538287222390956510226374073013716527402646767140081645358439363907244252584754169477181654880341181585766524382340379814185055191761925080189534;
            6'd52: xpb[177] = 1024'd79669393838187356350435400478363164153510001454909074374524302786282571227812124961560273419849330778676206109462521738443341276036184308068029805395479499071989433787629067351269882100639703686438542556436751651045543185973527146869932187906577515242675992409278791319357722515590319809757154214004272052029;
            6'd53: xpb[177] = 1024'd35869435681260765384536473166572566884360768494638518142601592335354139685868634301392464195644590757508059328073486093855670666421818884058798794435579301405294561036970912311583253974905334359160557710226736162009441013507690386495611791058985553303697104477375996872191062690800825434459116666083463914524;
            6'd54: xpb[177] = 1024'd116136173208458915817436473259596402359909962660103646038810736949402603481234282551239726186097525045783061954141943883847063897648673794604727908492010144672290362855883974609526865040688170753192770472403960519337699691262750399086269963894623040631538119959590260455130930939939964076279768944788250261350;
            6'd55: xpb[177] = 1024'd72336215051532324851537545947805805090760729699833089806888026498474171939290791891071916961892785024614915172752908239259393288034308370595496897532109947005595490105225819569840236914953801425914785626193945030301597518796913638711949567047031078692559232027687466007964271115150469700981731396867442123845;
            6'd56: xpb[177] = 1024'd28536256894605733885638618636015207821611496739562533574965316047545740397347301230904107737688045003446768391363872594671722678419942946586265886572209749338900617354567664530153608789219432098636800779983929541265495346331076878337629170199439116753580344095784671560797611290360975325683693848946633986340;
            6'd57: xpb[177] = 1024'd108802994421803884318538618729039043297160690905027661471174460661594204192712949480751369728140979291721771017432330384663115909646797857132195000628640592605896419173480726828097219855002268492669013542161153898593754024086136890928287343035076604081421359577998935143737479539500113967504346127651420333166;
            6'd58: xpb[177] = 1024'd65003036264877293352639691417248446028011457944757105239251750210665772650769458820583560503936239270553624236043294740075445300032432433122963989668740394939201546422822571788410591729267899165391028695951138409557651851620300130553966946187484642142442471646096140696570819714710619592206308579730612195661;
            6'd59: xpb[177] = 1024'd21203078107950702386740764105457848758862224984486549007329039759737341108825968160415751279731499249385477454654259095487774690418067009113732978708840197272506673672164416748723963603533529838113043849741122920521549679154463370179646549339892680203463583714193346249404159889921125216908271031809804058156;
            6'd60: xpb[177] = 1024'd101469815635148852819640764198481684234411419149951676903538184373785804904191616410263013270184433537660480080722716885479167921644921919659662092765271040539502475491077479046667574669316366232145256611918347277849808356909523382770304722175530167531304599196407609832344028139060263858728923310514590404982;
            6'd61: xpb[177] = 1024'd57669857478222261853741836886691086965262186189681120671615473922857373362248125750095204045979693516492333299333681240891497312030556495650431081805370842872807602740419324006980946543581996904867271765708331788813706184443686622395984325327938205592325711264504815385177368314270769483430885762593782267477;
            6'd62: xpb[177] = 1024'd13869899321295670887842909574900489696112953229410564439692763471928941820304635089927394821774953495324186517944645596303826702416191071641200070845470645206112729989761168967294318417847627577589286919498316299777604011977849862021663928480346243653346823332602020938010708489481275108132848214672974129972;
            6'd63: xpb[177] = 1024'd94136636848493821320742909667924325171662147394875692335901908085977405615670283339774656812227887783599189144013103386295219933643045982187129184901901488473108531808674231265237929483630463971621499681675540657105862689732909874612322101315983730981187838814816284520950576738620413749953500493377760476798;
        endcase
    end

    always_comb begin
        case(flag[59][11:6])
            6'd0: xpb[178] = 1024'd0;
            6'd1: xpb[178] = 1024'd50336678691567230354843982356133727902512914434605136103979197635048974073726792679606847588023147762431042362624067741707549324028680558177898173942001290806413659058016076225551301357896094644343514835465525168069760517267073114238001704468391769042208950882913490073783916913830919374655462945456952339293;
            6'd2: xpb[178] = 1024'd100673357383134460709687964712267455805025828869210272207958395270097948147453585359213695176046295524862084725248135483415098648057361116355796347884002581612827318116032152451102602715792189288687029670931050336139521034534146228476003408936783538084417901765826980147567833827661838749310925890913904678586;
            6'd3: xpb[178] = 1024'd26943340390576949665733019663586750962840316178079724183805737840170026883871239128805471549411768977849977680414709790543584131244821339978534396809672831485550302604477011339023664882171078211720346898009335657844920701580322569749026543721945857859806949234623412191245222667564125106847699009745262533548;
            6'd4: xpb[178] = 1024'd77280019082144180020577002019720478865353230612684860287784935475219000957598031808412319137434916740281020043038777532251133455273501898156432570751674122291963961662493087564574966240067172856063861733474860825914681218847395683987028248190337626902015900117536902265029139581395044481503161955202214872841;
            6'd5: xpb[178] = 1024'd3550002089586668976622056971039774023167717921554312263632278045291079694015685578004095510800390193268912998205351839379618938460962121779170619677344372164686946150937946452496028406446061779097178960553146147620080885893572025260051382975499946677404947586333334308706528421297330839039935074033572727803;
            6'd6: xpb[178] = 1024'd53886680781153899331466039327173501925680632356159448367611475680340053767742478257610943098823537955699955360829419581087168262489642679957068793619345662971100605208954022678047329764342156423440693796018671315689841403160645139498053087443891715719613898469246824382490445335128250213695398019490525067096;
            6'd7: xpb[178] = 1024'd104223359472721129686310021683307229828193546790764584471590673315389027841469270937217790686846685718130997723453487322794717586518323238134966967561346953777514264266970098903598631122238251067784208631484196483759601920427718253736054791912283484761822849352160314456274362248959169588350860964947477406389;
            6'd8: xpb[178] = 1024'd30493342480163618642355076634626524986008034099634036447438015885461106577886924706809567060212159171118890678620061629923203069705783461757705016487017203650237248755414957791519693288617139990817525858562481805465001587473894595009077926697445804537211896820956746499951751088861455945887634083778835261351;
            6'd9: xpb[178] = 1024'd80830021171730848997199058990760252888520948534239172551417213520510080651613717386416414648235306933549933041244129371630752393734464019935603190429018494456650907813431034017070994646513234635161040694028006973534762104740967709247079631165837573579420847703870236573735668002692375320543097029235787600644;
            6'd10: xpb[178] = 1024'd7100004179173337953244113942079548046335435843108624527264556090582159388031371156008191021600780386537825996410703678759237876921924243558341239354688744329373892301875892904992056812892123558194357921106292295240161771787144050520102765950999893354809895172666668617413056842594661678079870148067145455606;
            6'd11: xpb[178] = 1024'd57436682870740568308088096298213275948848350277713760631243753725631133461758163835615038609623928148968868359034771420466787200950604801736239413296690035135787551359891969130543358170788218202537872756571817463309922289054217164758104470419391662397018846055580158691196973756425581052735333093524097794899;
            6'd12: xpb[178] = 1024'd107773361562307798662932078654347003851361264712318896735222951360680107535484956515221886197647075911399910721658839162174336524979285359914137587238691325942201210417908045356094659528684312846881387592037342631379682806321290278996106174887783431439227796938493648764980890670256500427390796038981050134192;
            6'd13: xpb[178] = 1024'd34043344569750287618977133605666299009175752021188348711070293930752186271902610284813662571012549364387803676825413469302822008166745583536875636164361575814924194906352904244015721695063201769914704819115627953085082473367466620269129309672945751214616844407290080808658279510158786784927569157812407989154;
            6'd14: xpb[178] = 1024'd84380023261317517973821115961800026911688666455793484815049491565801160345629402964420510159035697126818846039449481211010371332195426141714773810106362866621337853964368980469567023052959296414258219654581153121154842990634539734507131014141337520256825795290203570882442196423989706159583032103269360328447;
            6'd15: xpb[178] = 1024'd10650006268760006929866170913119322069503153764662936790896834135873239082047056734012286532401170579806738994616055518138856815382886365337511859032033116494060838452813839357488085219338185337291536881659438442860242657680716075780154148926499840032214842759000002926119585263891992517119805222100718183409;
            6'd16: xpb[178] = 1024'd60986684960327237284710153269253049972016068199268072894876031770922213155773849413619134120424318342237781357240123259846406139411566923515410032974034407300474497510829915583039386577234279981635051717124963610930003174947789190018155853394891609074423793641913492999903502177722911891775268167557670522702;
            6'd17: xpb[178] = 1024'd111323363651894467639554135625386777874528982633873208998855229405971187229500642093225981708447466104668823719864191001553955463440247481693308206916035698106888156568845991808590687935130374625978566552590488778999763692214862304256157557863283378116632744524826983073687419091553831266430731113014622861995;
            6'd18: xpb[178] = 1024'd37593346659336956595599190576706073032343469942742660974702571976043265965918295862817758081812939557656716675030765308682440946627707705316046255841705947979611141057290850696511750101509263549011883779668774100705163359261038645529180692648445697892021791993623415117364807931456117623967504231845980716957;
            6'd19: xpb[178] = 1024'd87930025350904186950443172932839800934856384377347797078681769611092240039645088542424605669836087320087759037654833050389990270656388263493944429783707238786024800115306926922063051459405358193355398615134299268774923876528111759767182397116837466934230742876536905191148724845287036998622967177302933056250;
            6'd20: xpb[178] = 1024'd14200008358346675906488227884159096092670871686217249054529112181164318776062742312016382043201560773075651992821407357518475753843848487116682478709377488658747784603751785809984113625784247116388715842212584590480323543574288101040205531901999786709619790345333337234826113685189323356159740296134290911212;
            6'd21: xpb[178] = 1024'd64536687049913906261332210240292823995183786120822385158508309816213292849789534991623229631224708535506694355445475099226025077872529045294580652651378779465161443661767862035535414983680341760732230677678109758550084060841361215278207236370391555751828741228246827308610030599020242730815203241591243250505;
            6'd22: xpb[178] = 1024'd114873365741481136616176192596426551897696700555427521262487507451262266923516327671230077219247856297937736718069542840933574401901209603472478826593380070271575102719783938261086716341576436405075745513143634926619844578108434329516208940838783324794037692111160317382393947512851162105470666187048195589798;
            6'd23: xpb[178] = 1024'd41143348748923625572221247547745847055511187864296973238334850021334345659933981440821853592613329750925629673236117148062059885088669827095216875519050320144298087208228797149007778507955325328109062740221920248325244245154610670789232075623945644569426739579956749426071336352753448463007439305879553444760;
            6'd24: xpb[178] = 1024'd91480027440490855927065229903879574958024102298902109342314047656383319733660774120428701180636477513356672035860184889769609209117350385273115049461051610950711746266244873374559079865851419972452577575687445416395004762421683785027233780092337413611635690462870239499855253266584367837662902251336505784053;
            6'd25: xpb[178] = 1024'd17750010447933344883110284855198870115838589607771561318161390226455398470078427890020477554001950966344564991026759196898094692304810608895853098386721860823434730754689732262480142032230308895485894802765730738100404429467860126300256914877499733387024737931666671543532642106486654195199675370167863639015;
            6'd26: xpb[178] = 1024'd68086689139500575237954267211332598018351504042376697422140587861504372543805220569627325142025098728775607353650826938605644016333491167073751272328723151629848389812705808488031443390126403539829409638231255906170164946734933240538258619345891502429233688814580161617316559020317573569855138315624815978308;
            6'd27: xpb[178] = 1024'd118423367831067805592798249567466325920864418476981833526119785496553346617532013249234172730048246491206649716274894680313193340362171725251649446270724442436262048870721884713582744748022498184172924473696781074239925464002006354776260323814283271471442639697493651691100475934148492944510601261081768317601;
            6'd28: xpb[178] = 1024'd44693350838510294548843304518785621078678905785851285501967128066625425353949667018825949103413719944194542671441468987441678823549631948874387495196394692308985033359166743601503806914401387107206241700775066395945325131048182696049283458599445591246831687166290083734777864774050779302047374379913126172563;
            6'd29: xpb[178] = 1024'd95030029530077524903687286874919348981191820220456421605946325701674399427676459698432796691436867706625585034065536729149228147578312507052285669138395983115398692417182819827055108272297481751549756536240591564015085648315255810287285163067837360289040638049203573808561781687881698676702837325370078511856;
            6'd30: xpb[178] = 1024'd21300012537520013859732341826238644139006307529325873581793668271746478164094113468024573064802341159613477989232111036277713630765772730675023718064066232988121676905627678714976170438676370674583073763318876885720485315361432151560308297852999680064429685518000005852239170527783985034239610444201436366818;
            6'd31: xpb[178] = 1024'd71636691229087244214576324182372372041519221963931009685772865906795452237820906147631420652825488922044520351856178777985262954794453288852921892006067523794535335963643754940527471796572465318926588598784402053790245832628505265798310002321391449106638636400913495926023087441614904408895073389658388706111;
            6'd32: xpb[178] = 1024'd121973369920654474569420306538506099944032136398536145789752063541844426311547698827238268240848636684475562714480246519692812278823133847030820065948068814600948995021659831166078773154468559963270103434249927221860006349895578380036311706789783218148847587283826985999807004355445823783550536335115341045404;
            6'd33: xpb[178] = 1024'd48243352928096963525465361489825395101846623707405597765599406111916505047965352596830044614214110137463455669646820826821297762010594070653558114873739064473671979510104690053999835320847448886303420661328212543565406016941754721309334841574945537924236634752623418043484393195348110141087309453946698900366;
            6'd34: xpb[178] = 1024'd98580031619664193880309343845959123004359538142010733869578603746965479121692145276436892202237257899894498032270888568528847086039274628831456288815740355280085638568120766279551136678743543530646935496793737711635166534208827835547336546043337306966445585635536908117268310109179029515742772399403651239659;
            6'd35: xpb[178] = 1024'd24850014627106682836354398797278418162174025450880185845425946317037557858109799046028668575602731352882390987437462875657332569226734852454194337741410605152808623056565625167472198845122432453680252723872023033340566201255004176820359680828499626741834633104333340160945698949081315873279545518235009094621;
            6'd36: xpb[178] = 1024'd75186693318673913191198381153412146064686939885485321949405143952086531931836591725635516163625879115313433350061530617364881893255415410632092511683411895959222282114581701393023500203018527098023767559337548201410326718522077291058361385296891395784043583987246830234729615862912235247935008463691961433914;
            6'd37: xpb[178] = 1024'd1456676326116402147243436104731441222501427194354773925252486522158610668254245495227292536991352568301326305228104924493367376442875634254830560609082145831945266603026560280944562369397416021057084786415833523115726385568253632331384520082053715559432631456043262278407004702814521605471781582523319288876;
            6'd38: xpb[178] = 1024'd51793355017683632502087418460865169125014341628959910029231684157207584741981038174834140125014500330732368667852172666200916700471556192432728734551083436638358925661042636506495863727293510665400599621881358691185486902835326746569386224550445484601641582338956752352190921616645440980127244527980271628169;
            6'd39: xpb[178] = 1024'd102130033709250862856931400816998897027527256063565046133210881792256558815707830854440987713037648093163411030476240407908466024500236750610626908493084727444772584719058712732047165085189605309744114457346883859255247420102399860807387929018837253643850533221870242425974838530476360354782707473437223967462;
            6'd40: xpb[178] = 1024'd28400016716693351812976455768318192185341743372434498109058224362328637552125484624032764086403121546151303985642814715036951507687696974233364957418754977317495569207503571619968227251568494232777431684425169180960647087148576202080411063803999573419239580690666674469652227370378646712319480592268581822424;
            6'd41: xpb[178] = 1024'd78736695408260582167820438124451920087854657807039634213037421997377611625852277303639611674426269308582346348266882456744500831716377532411263131360756268123909228265519647845519528609464588877120946519890694349030407604415649316318412768272391342461448531573580164543436144284209566086974943537725534161717;
            6'd42: xpb[178] = 1024'd5006678415703071123865493075771215245669145115909086188884764567449690362269931073231388047791742761570239303433456763872986314903837756034001180286426517996632212753964506733440590775843477800154263746968979670735807271461825657591435903057553662236837579042376596587113533124111852444511716656556892016679;
            6'd43: xpb[178] = 1024'd55343357107270301478709475431904943148182059550514222292863962202498664435996723752838235635814890524001281666057524505580535638932518314211899354228427808803045871811980582958991892133739572444497778582434504838805567788728898771829437607525945431279046529925290086660897450037942771819167179602013844355972;
            6'd44: xpb[178] = 1024'd105680035798837531833553457788038671050694973985119358396843159837547638509723516432445083223838038286432324028681592247288084962961198872389797528170429099609459530869996659184543193491635667088841293417900030006875328305995971886067439311994337200321255480808203576734681366951773691193822642547470796695265;
            6'd45: xpb[178] = 1024'd31950018806280020789598512739357966208509461293988810372690502407619717246141170202036859597203511739420216983848166554416570446148659096012535577096099349482182515358441518072464255658014556011874610644978315328580727973042148227340462446779499520096644528277000008778358755791675977551359415666302154550227;
            6'd46: xpb[178] = 1024'd82286697497847251144442495095491694111022375728593946476669700042668691319867962881643707185226659501851259346472234296124119770177339654190433751038100640288596174416457594298015557015910650656218125480443840496650488490309221341578464151247891289138853479159913498852142672705506896926014878611759106889520;
            6'd47: xpb[178] = 1024'd8556680505289740100487550046810989268836863037463398452517042612740770056285616651235483558592132954839152301638808603252605253364799877813171799963770890161319158904902453185936619182289539579251442707522125818355888157355397682851487286033053608914242526628709930895820061545409183283551651730590464744482;
            6'd48: xpb[178] = 1024'd58893359196856970455331532402944717171349777472068534556496240247789744130012409330842331146615280717270194664262876344960154577393480435991069973905772180967732817962918529411487920540185634223594957542987650986425648674622470797089488990501445377956451477511623420969603978459240102658207114676047417083775;
            6'd49: xpb[178] = 1024'd109230037888424200810175514759078445073862691906673670660475437882838718203739202010449178734638428479701237026886944086667703901422160994168968147847773471774146477020934605637039221898081728867938472378453176154495409191889543911327490694969837146998660428394536911043387895373071022032862577621504369423068;
            6'd50: xpb[178] = 1024'd35500020895866689766220569710397740231677179215543122636322780452910796940156855780040955108003901932689129982053518393796189384609621217791706196773443721646869461509379464524960284064460617790971789605531461476200808858935720252600513829754999466774049475863333343087065284212973308390399350740335727278030;
            6'd51: xpb[178] = 1024'd85836699587433920121064552066531468134190093650148258740301978087959771013883648459647802696027049695120172344677586135503738708638301775969604370715445012453283120567395540750511585422356712435315304440996986644270569376202793366838515534223391235816258426746246833160849201126804227765054813685792679617323;
            6'd52: xpb[178] = 1024'd12106682594876409077109607017850763292004580959017710716149320658031849750301302229239579069392523148108065299844160442632224191825761999592342419641115262326006105055840399638432647588735601358348621668075271965975969043248969708111538669008553555591647474215043265204526589966706514122591586804624037472285;
            6'd53: xpb[178] = 1024'd62443361286443639431953589373984491194517495393622846820128518293080823824028094908846426657415670910539107662468228184339773515854442557770240593583116553132419764113856475863983948946631696002692136503540797134045729560516042822349540373476945324633856425097956755278310506880537433497247049750080989811578;
            6'd54: xpb[178] = 1024'd112780039978010869786797571730118219097030409828227982924107715928129797897754887588453274245438818672970150025092295926047322839883123115948138767525117843938833423171872552089535250304527790647035651339006322302115490077783115936587542077945337093676065375980870245352094423794368352871902512695537942150871;
            6'd55: xpb[178] = 1024'd39050022985453358742842626681437514254844897137097434899955058498201876634172541358045050618804292125958042980258870233175808323070583339570876816450788093811556407660317410977456312470906679570068968566084607623820889744829292277860565212730499413451454423449666677395771812634270639229439285814369300005833;
            6'd56: xpb[178] = 1024'd89386701677020589097686609037571242157357811571702571003934256133250850707899334037651898206827439888389085342882937974883357647099263897748774990392789384617970066718333487203007613828802774214412483401550132791890650262096365392098566917198891182493663374332580167469555729548101558604094748759826252345126;
            6'd57: xpb[178] = 1024'd15656684684463078053731663988890537315172298880572022979781598703322929444316987807243674580192913341376978298049512282011843130286724121371513039318459634490693051206778346090928675995181663137445800628628418113596049929142541733371590051984053502269052421801376599513233118388003844961631521878657610200088;
            6'd58: xpb[178] = 1024'd65993363376030308408575646345024265217685213315177159083760796338371903518043780486850522168216061103808020660673580023719392454315404679549411213260460925297106710264794422316479977353077757781789315464093943281665810446409614847609591756452445271311261372684290089587017035301834764336286984824114562539381;
            6'd59: xpb[178] = 1024'd116330042067597538763419628701157993120198127749782295187739993973420877591770573166457369756239208866239063023297647765426941778344085237727309387202462216103520369322810498542031278710973852426132830299559468449735570963676687961847593460920837040353470323567203579660800952215665683710942447769571514878674;
            6'd60: xpb[178] = 1024'd42600025075040027719464683652477288278012615058651747163587336543492956328188226936049146129604682319226955978464222072555427261531545461350047436128132465976243353811255357429952340877352741349166147526637753771440970630722864303120616595705999360128859371036000011704478341055567970068479220888402872733636;
            6'd61: xpb[178] = 1024'd92936703766607258074308666008611016180525529493256883267566534178541930401915019615655993717627830081657998341088289814262976585560226019527945610070133756782657012869271433655503642235248835993509662362103278939510731147989937417358618300174391129171068321918913501778262257969398889443134683833859825072929;
            6'd62: xpb[178] = 1024'd19206686774049747030353720959930311338340016802126335243413876748614009138332673385247770090993303534645891296254864121391462068747686243150683658995804006655379997357716292543424704401627724916542979589181564261216130815036113758631641434959553448946457369387709933821939646809301175800671456952691182927891;
            6'd63: xpb[178] = 1024'd69543365465616977385197703316064039240852931236731471347393074383662983212059466064854617679016451297076933658878931863099011392776366801328581832937805297461793656415732368768976005759523819560886494424647089429285891332303186872869643139427945217988666320270623423895723563723132095175326919898148135267184;
        endcase
    end

    always_comb begin
        case(flag[59][16:12])
            5'd0: xpb[179] = 1024'd0;
            5'd1: xpb[179] = 1024'd119880044157184207740041685672197767143365845671336607451372272018711957285786258744461465267039599059507976021502999604806560716805047359506480006879806588268207315473748444994527307117419914205230009260112614597355651849570259987107644843896336987030875271153536913969507480636963014549982382843605087606477;
            5'd2: xpb[179] = 1024'd115693392630243674081284443939581101542033264216937530774612688972447019234263378578907859319421523809572802635548505775034057592768874384457799888743282135602723956377925672651424375043322622689149820911837989348346942848919623201250311118109444524794930638892956769908908433199997396082846075860584580728623;
            5'd3: xpb[179] = 1024'd111506741103303140422527202206964435940700682762538454097853105926182081182740498413354253371803448559637629249594011945261554468732701409409119770606757682937240597282102900308321442969225331173069632563563364099338233848268986415392977392322552062558986006632376625848309385763031777615709768877564073850769;
            5'd4: xpb[179] = 1024'd107320089576362606763769960474347770339368101308139377421093522879917143131217618247800647424185373309702455863639518115489051344696528434360439652470233230271757238186280127965218510895128039656989444215288738850329524847618349629535643666535659600323041374371796481787710338326066159148573461894543566972915;
            5'd5: xpb[179] = 1024'd103133438049422073105012718741731104738035519853740300744333939833652205079694738082247041476567298059767282477685024285716548220660355459311759534333708777606273879090457355622115578821030748140909255867014113601320815846967712843678309940748767138087096742111216337727111290889100540681437154911523060095061;
            5'd6: xpb[179] = 1024'd98946786522481539446255477009114439136702938399341224067574356787387267028171857916693435528949222809832109091730530455944045096624182484263079416197184324940790519994634583279012646746933456624829067518739488352312106846317076057820976214961874675851152109850636193666512243452134922214300847928502553217207;
            5'd7: xpb[179] = 1024'd94760134995541005787498235276497773535370356944942147390814773741122328976648977751139829581331147559896935705776036626171541972588009509214399298060659872275307160898811810935909714672836165108748879170464863103303397845666439271963642489174982213615207477590056049605913196015169303747164540945482046339353;
            5'd8: xpb[179] = 1024'd90573483468600472128740993543881107934037775490543070714055190694857390925126097585586223633713072309961762319821542796399038848551836534165719179924135419609823801802989038592806782598738873592668690822190237854294688845015802486106308763388089751379262845329475905545314148578203685280028233962461539461499;
            5'd9: xpb[179] = 1024'd86386831941659938469983751811264442332705194036143994037295607648592452873603217420032617686094997060026588933867048966626535724515663559117039061787610966944340442707166266249703850524641582076588502473915612605285979844365165700248975037601197289143318213068895761484715101141238066812891926979441032583645;
            5'd10: xpb[179] = 1024'd82200180414719404811226510078647776731372612581744917360536024602327514822080337254479011738476921810091415547912555136854032600479490584068358943651086514278857083611343493906600918450544290560508314125640987356277270843714528914391641311814304826907373580808315617424116053704272448345755619996420525705791;
            5'd11: xpb[179] = 1024'd78013528887778871152469268346031111130040031127345840683776441556062576770557457088925405790858846560156242161958061307081529476443317609019678825514562061613373724515520721563497986376446999044428125777366362107268561843063892128534307586027412364671428948547735473363517006267306829878619313013400018827937;
            5'd12: xpb[179] = 1024'd73826877360838337493712026613414445528707449672946764007016858509797638719034576923371799843240771310221068776003567477309026352407144633970998707378037608947890365419697949220395054302349707528347937429091736858259852842413255342676973860240519902435484316287155329302917958830341211411483006030379511950083;
            5'd13: xpb[179] = 1024'd69640225833897803834954784880797779927374868218547687330257275463532700667511696757818193895622696060285895390049073647536523228370971658922318589241513156282407006323875176877292122228252416012267749080817111609251143841762618556819640134453627440199539684026575185242318911393375592944346699047359005072229;
            5'd14: xpb[179] = 1024'd65453574306957270176197543148181114326042286764148610653497692417267762615988816592264587948004620810350722004094579817764020104334798683873638471104988703616923647228052404534189190154155124496187560732542486360242434841111981770962306408666734977963595051765995041181719863956409974477210392064338498194375;
            5'd15: xpb[179] = 1024'd61266922780016736517440301415564448724709705309749533976738109371002824564465936426710982000386545560415548618140085987991516980298625708824958352968464250951440288132229632191086258080057832980107372384267861111233725840461344985104972682879842515727650419505414897121120816519444356010074085081317991316521;
            5'd16: xpb[179] = 1024'd57080271253076202858683059682947783123377123855350457299978526324737886512943056261157376052768470310480375232185592158219013856262452733776278234831939798285956929036406859847983326005960541464027184035993235862225016839810708199247638957092950053491705787244834753060521769082478737542937778098297484438667;
            5'd17: xpb[179] = 1024'd52893619726135669199925817950331117522044542400951380623218943278472948461420176095603770105150395060545201846231098328446510732226279758727598116695415345620473569940584087504880393931863249947946995687718610613216307839160071413390305231306057591255761154984254608999922721645513119075801471115276977560813;
            5'd18: xpb[179] = 1024'd48706968199195135541168576217714451920711960946552303946459360232208010409897295930050164157532319810610028460276604498674007608190106783678917998558890892954990210844761315161777461857765958431866807339443985364207598838509434627532971505519165129019816522723674464939323674208547500608665164132256470682959;
            5'd19: xpb[179] = 1024'd44520316672254601882411334485097786319379379492153227269699777185943072358374415764496558209914244560674855074322110668901504484153933808630237880422366440289506851748938542818674529783668666915786618991169360115198889837858797841675637779732272666783871890463094320878724626771581882141528857149235963805105;
            5'd20: xpb[179] = 1024'd40333665145314068223654092752481120718046798037754150592940194139678134306851535598942952262296169310739681688367616839129001360117760833581557762285841987624023492653115770475571597709571375399706430642894734866190180837208161055818304053945380204547927258202514176818125579334616263674392550166215456927251;
            5'd21: xpb[179] = 1024'd36147013618373534564896851019864455116714216583355073916180611093413196255328655433389346314678094060804508302413123009356498236081587858532877644149317534958540133557292998132468665635474083883626242294620109617181471836557524269960970328158487742311982625941934032757526531897650645207256243183194950049397;
            5'd22: xpb[179] = 1024'd31960362091433000906139609287247789515381635128955997239421028047148258203805775267835740367060018810869334916458629179583995112045414883484197526012793082293056774461470225789365733561376792367546053946345484368172762835906887484103636602371595280076037993681353888696927484460685026740119936200174443171543;
            5'd23: xpb[179] = 1024'd27773710564492467247382367554631123914049053674556920562661445000883320152282895102282134419441943560934161530504135349811491988009241908435517407876268629627573415365647453446262801487279500851465865598070859119164053835256250698246302876584702817840093361420773744636328437023719408272983629217153936293689;
            5'd24: xpb[179] = 1024'd23587059037551933588625125822014458312716472220157843885901861954618382100760014936728528471823868310998988144549641520038988863973068933386837289739744176962090056269824681103159869413182209335385677249796233870155344834605613912388969150797810355604148729160193600575729389586753789805847322234133429415835;
            5'd25: xpb[179] = 1024'd19400407510611399929867884089397792711383890765758767209142278908353444049237134771174922524205793061063814758595147690266485739936895958338157171603219724296606697174001908760056937339084917819305488901521608621146635833954977126531635425010917893368204096899613456515130342149788171338711015251112922537981;
            5'd26: xpb[179] = 1024'd15213755983670866271110642356781127110051309311359690532382695862088505997714254605621316576587717811128641372640653860493982615900722983289477053466695271631123338078179136416954005264987626303225300553246983372137926833304340340674301699224025431132259464639033312454531294712822552871574708268092415660127;
            5'd27: xpb[179] = 1024'd11027104456730332612353400624164461508718727856960613855623112815823567946191374440067710628969642561193467986686160030721479491864550008240796935330170818965639978982356364073851073190890334787145112204972358123129217832653703554816967973437132968896314832378453168393932247275856934404438401285071908782273;
            5'd28: xpb[179] = 1024'd6840452929789798953596158891547795907386146402561537178863529769558629894668494274514104681351567311258294600731666200948976367828377033192116817193646366300156619886533591730748141116793043271064923856697732874120508832003066768959634247650240506660370200117873024333333199838891315937302094302051401904419;
            5'd29: xpb[179] = 1024'd2653801402849265294838917158931130306053564948162460502103946723293691843145614108960498733733492061323121214777172371176473243792204058143436699057121913634673260790710819387645209042695751754984735508423107625111799831352429983102300521863348044424425567857292880272734152401925697470165787319030895026565;
            5'd30: xpb[179] = 1024'd122533845560033473034880602831128897449419410619499067953476218742005649128931872853421964000773091120831097236280171975983033960597251417649916705936928501902880576264459264382172516160115665960214744768535722222467451680922689970209945365759685031455300839010829794242241633038888712020148170162635982633042;
            5'd31: xpb[179] = 1024'd118347194033092939376123361098512231848086829165099991276716635695740711077408992687868358053155015870895923850325678146210530836561078442601236587800404049237397217168636492039069584086018374444134556420261096973458742680272053184352611639972792569219356206750249650181642585601923093553011863179615475755188;
        endcase
    end

    always_comb begin
        case(flag[60][5:0])
            6'd0: xpb[180] = 1024'd0;
            6'd1: xpb[180] = 1024'd57080271253076202858683059682947783123377123855350457299978526324737886512943056261157376052768470310480375232185592158219013856262452733776278234831939798285956929036406859847983326005960541464027184035993235862225016839810708199247638957092950053491705787244834753060521769082478737542937778098297484438667;
            6'd2: xpb[180] = 1024'd114160542506152405717366119365895566246754247710700914599957052649475773025886112522314752105536940620960750464371184316438027712524905467552556469663879596571913858072813719695966652011921082928054368071986471724450033679621416398495277914185900106983411574489669506121043538164957475085875556196594968877334;
            6'd3: xpb[180] = 1024'd47174118075103867177250251644028916625432944440315687771803723909236764201520029873457056943647736621997976289099283040077977727946137866773674579479488353924180112539649362206319738826364418670771354499592467740310689669211227824777938301595620711208297458320387201151458779173507579611694644468266858831670;
            6'd4: xpb[180] = 1024'd104254389328180070035933311326976699748810068295666145071782250233974650714463086134614432996416206932478351521284875198296991584208590600549952814311428152210137041576056222054303064832324960134798538535585703602535706509021936024025577258688570764700003245565221954211980548255986317154632422566564343270337;
            6'd5: xpb[180] = 1024'd37267964897131531495817443605110050127488765025280918243628921493735641890097003485756737834527002933515577346012973921936941599629822999771070924127036909562403296042891864564656151646768295877515524963191699618396362498611747450308237646098291368924889129395939649242395789264536421680451510838236233224673;
            6'd6: xpb[180] = 1024'd94348236150207734354500503288057833250865888880631375543607447818473528403040059746914113887295473243995952578198566080155955455892275733547349158958976707848360225079298724412639477652728837341542708999184935480621379338422455649555876603191241422416594916640774402302917558347015159223389288936533717663340;
            6'd7: xpb[180] = 1024'd27361811719159195814384635566191183629544585610246148715454119078234519578673977098056418725406269245033178402926664803795905471313508132768467268774585465200626479546134366922992564467172173084259695426790931496482035328012267075838536990600962026641480800471492097333332799355565263749208377208205607617676;
            6'd8: xpb[180] = 1024'd84442082972235398673067695249138966752921709465596606015432645402972406091617033359213794778174739555513553635112256962014919327575960866544745503606525263486583408582541226770975890473132714548286879462784167358707052167822975275086175947693912080133186587716326850393854568438044001292146155306503092056343;
            6'd9: xpb[180] = 1024'd17455658541186860132951827527272317131600406195211379187279316662733397267250950710356099616285535556550779459840355685654869342997193265765863613422134020838849663049376869281328977287576050291003865890390163374567708157412786701368836335103632684358072471547044545424269809446594105817965243578174982010679;
            6'd10: xpb[180] = 1024'd74535929794263062991634887210220100254977530050561836487257842987471283780194006971513475669054005867031154692025947843873883199259645999542141848254073819124806592085783729129312303293536591755031049926383399236792724997223494900616475292196582737849778258791879298484791578529072843360903021676472466449346;
            6'd11: xpb[180] = 1024'd7549505363214524451519019488353450633656226780176609659104514247232274955827924322655780507164801868068380516754046567513833214680878398763259958069682576477072846552619371639665390107979927497748036353989395252653380986813306326899135679606303342074664142622596993515206819537622947886722109948144356403682;
            6'd12: xpb[180] = 1024'd64629776616290727310202079171301233757033350635527066959083040571970161468770980583813156559933272178548755748939638725732847070943331132539538192901622374763029775589026231487648716113940468961775220389982631114878397826624014526146774636699253395566369929867431746575728588620101685429659888046441840842349;
            6'd13: xpb[180] = 1024'd121710047869366930168885138854249016880410474490877524259061566896708047981714036844970532612701742489029130981125230883951860927205783866315816427733562173048986704625433091335632042119901010425802404425975866977103414666434722725394413593792203449058075717112266499636250357702580422972597666144739325281016;
            6'd14: xpb[180] = 1024'd54723623438318391628769271132382367259089171220492297430908238156469039157347954196112837450812538490066356805853329607591810942627016265536934537549170930401252959092268733845985128934344346168519390853581862992964070656024534151677073981201924053282961600942984194666665598711130527498416754416411215235352;
            6'd15: xpb[180] = 1024'd111803894691394594487452330815330150382466295075842754730886764481206925670291010457270213503581008800546732038038921765810824798889468999313212772381110728687209888128675593693968454940304887632546574889575098855189087495835242350924712938294874106774667388187818947727187367793609265041354532514708699674019;
            6'd16: xpb[180] = 1024'd44817470260346055947336463093463500761144991805457527902733435740967916845924927808412518341691804801583957862767020489450774814310701398534330882196719486039476142595511236204321541754748223375263561317181094871049743485425053777207373325704594710999553272018536642757602608802159369567173620786380589628355;
            6'd17: xpb[180] = 1024'd101897741513422258806019522776411283884522115660807985202711962065705803358867984069569894394460275112064333094952612647669788670573154132310609117028659284325433071631918096052304867760708764839290745353174330733274760325235761976455012282797544764491259059263371395818124377884638107110111398884678074067022;
            6'd18: xpb[180] = 1024'd34911317082373720265903655054544634263200812390422758374558633325466794534501901420712199232571071113101558919680711371309738685994386531531727226844268041677699326098753738562657954575152100582007731780780326749135416314825573402737672670207265368716144943094089090848539618893188211635930487156349964021358;
            6'd19: xpb[180] = 1024'd91991588335449923124586714737492417386577936245773215674537159650204681047444957681869575285339541423581934151866303529528752542256839265308005461676207839963656255135160598410641280581112642046034915816773562611360433154636281601985311627300215422207850730338923843909061387975666949178868265254647448460025;
            6'd20: xpb[180] = 1024'd25005163904401384584470847015625767765256632975387988846383830909965672223078875033011880123450337424619159976594402253168702557678071664529123571491816597315922509601996240920994367395555977788751902244379558627221089144226093028267972014709936026432736614169641538939476628984217053704687353526319338414361;
            6'd21: xpb[180] = 1024'd82085435157477587443153906698573550888633756830738446146362357234703558736021931294169256176218807735099535208779994411387716413940524398305401806323756395601879438638403100768977693401516519252779086280372794489446105984036801227515610971802886079924442401414476291999998398066695791247625131624616822853028;
            6'd22: xpb[180] = 1024'd15099010726429048903038038976706901267312453560353219318209028494464549911655848645311561014329603736136761033508093135027666429361756797526519916139365152954145693105238743279330780215959854995496072707978790505306761973626612653798271359212606684149328285245193987030413639075245895773444219896288712807364;
            6'd23: xpb[180] = 1024'd72179281979505251761721098659654684390689577415703676618187554819202436424598904906468937067098074046617136265693685293246680285624209531302798150971304951240102622141645603127314106221920396459523256743972026367531778813437320853045910316305556737641034072490028740090935408157724633316381997994586197246031;
            6'd24: xpb[180] = 1024'd5192857548456713221605230937788034769368274145318449790034226078963427600232822257611241905208870047654362090421784016886630301045441930523916260786913708592368876608481245637667193036363732202240243171578022383392434803027132279328570703715277341865919956320746435121350649166274737842201086266258087200367;
            6'd25: xpb[180] = 1024'd62273128801532916080288290620735817892745398000668907090012752403701314113175878518768617957977340358134737322607376175105644157307894664300194495618853506878325805644888105485650519042324273666267427207571258245617451642837840478576209660808227395357625743565581188181872418248753475385138864364555571639034;
            6'd26: xpb[180] = 1024'd119353400054609118938971350303683601016122521856019364389991278728439200626118934779925994010745810668615112554792968333324658013570347398076472730450793305164282734681294965333633845048284815130294611243564494107842468482648548677823848617901177448849331530810415941242394187331232212928076642462853056077701;
            6'd27: xpb[180] = 1024'd52366975623560580398855482581816951394801218585634137561837949988200191801752852131068298848856606669652338379521067056964608028991579797297590840266402062516548989148130607843986931862728150873011597671170490123703124472238360104106509005310898053074217414641133636272809428339782317453895730734524946032037;
            6'd28: xpb[180] = 1024'd109447246876636783257538542264764734518178342440984594861816476312938078314695908392225674901625076980132713611706659215183621885254032531073869075098341860802505918184537467691970257868688692337038781707163725985928141312049068303354147962403848106565923201885968389333331197422261054996833508832822430470704;
            6'd29: xpb[180] = 1024'd42460822445588244717422674542898084896857039170599368033663147572699069490329825743367979739735872981169939436434757938823571900675264930294987184913950618154772172651373110202323344683132028079755768134769722001788797301638879729636808349813568710790809085716686084363746438430811159522652597104494320425040;
            6'd30: xpb[180] = 1024'd99541093698664447576105734225845868020234163025949825333641673897436956003272882004525355792504343291650314668620350097042585756937717664071265419745890416440729101687779970050306670689092569543782952170762957864013814141449587928884447306906518764282514872961520837424268207513289897065590375202791804863707;
            6'd31: xpb[180] = 1024'd32554669267615909035989866503979218398912859755564598505488345157197947178906799355667660630615139292687540493348448820682535772358950063292383529561499173792995356154615612560659757503535905286499938598368953879874470131039399355167107694316239368507400756792238532454683448521840001591409463474463694818043;
            6'd32: xpb[180] = 1024'd89634940520692111894672926186927001522289983610915055805466871481935833691849855616825036683383609603167915725534040978901549628621402797068661764393438972078952285191022472408643083509496446750527122634362189742099486970850107554414746651409189421999106544037073285515205217604318739134347241572761179256710;
            6'd33: xpb[180] = 1024'd22648516089643573354557058465060351900968680340529828977313542741696824867483772967967341521494405604205141550262139702541499644042635196289779874209047729431218539657858114918996170323939782493244109061968185757960142960439918980697407038818910026223992427867790980545620458612868843660166329844433069211046;
            6'd34: xpb[180] = 1024'd79728787342719776213240118148008135024345804195880286277292069066434711380426829229124717574262875914685516782447731860760513500305087930066058109040987527717175468694264974766979496329900323957271293097961421620185159800250627179945045995911860079715698215112625733606142227695347581203104107942730553649713;
            6'd35: xpb[180] = 1024'd12742362911671237673124250426141485403024500925495059449138740326195702556060746580267022412373671915722742607175830584400463515726320329287176218856596285069441723161100617277332583144343659699988279525567417636045815789840438606227706383321580683940584098943343428636557468703897685728923196214402443604049;
            6'd36: xpb[180] = 1024'd69822634164747440531807310109089268526401624780845516749117266650933589069003802841424398465142142226203117839361422742619477371988773063063454453688536083355398652197507477125315909150304201164015463561560653498270832629651146805475345340414530737432289886188178181697079237786376423271860974312699928042716;
            6'd37: xpb[180] = 1024'd2836209733698901991691442387222618905080321510460289920963937910694580244637720192566703303252938227240343664089521466259427387410005462284572563504144840707664906664343119635668995964747536906732449989166649514131488619240958231758005727824251341657175770018895876727494478794926527797680062584371817997052;
            6'd38: xpb[180] = 1024'd59916480986775104850374502070170402028457445365810747220942464235432466757580776453724079356021408537720718896275113624478441243672458196060850798336084638993621835700749979483652321970708078370759634025159885376356505459051666431005644684917201395148881557263730629788016247877405265340617840682669302435719;
            6'd39: xpb[180] = 1024'd116996752239851307709057561753118185151834569221161204520920990560170353270523832714881455408789878848201094128460705782697455099934910929837129033168024437279578764737156839331635647976668619834786818061153121238581522298862374630253283642010151448640587344508565382848538016959884002883555618780966786874386;
            6'd40: xpb[180] = 1024'd50010327808802769168941694031251535530513265950775977692767661819931344446157750066023760246900674849238319953188804506337405115356143329058247142983633194631845019203992481841988734791111955577503804488759117254442178288452186056535944029419872052865473228339283077878953257968434107409374707052638676828722;
            6'd41: xpb[180] = 1024'd107090599061878972027624753714199318653890389806126434992746188144669230959100806327181136299669145159718695185374396664556418971618596062834525377815572992917801948240399341689972060797072497041530988524752353116667195128262894255783582986512822106357179015584117830939475027050912844952312485150936161267389;
            6'd42: xpb[180] = 1024'd40104174630830433487508885992332669032569086535741208164592859404430222134734723678323441137779941160755921010102495388196368987039828462055643487631181750270068202707234984200325147611515832784247974952358349132527851117852705682066243373922542710582064899414835525969890268059462949478131573422608051221725;
            6'd43: xpb[180] = 1024'd97184445883906636346191945675280452155946210391091665464571385729168108647677779939480817190548411471236296242288087546415382843302281195831921722463121548556025131743641844048308473617476374248275158988351584994752867957663413881313882331015492764073770686659670279030412037141941687021069351520905535660392;
            6'd44: xpb[180] = 1024'd30198021452858097806076077953413802534624907120706438636418056988929099823311697290623122028659207472273522067016186270055332858723513595053039832278730305908291386210477486558661560431919709990992145415957581010613523947253225307596542718425213368298656570490387974060827278150491791546888439792577425614728;
            6'd45: xpb[180] = 1024'd87278292705934300664759137636361585658002030976056895936396583313666986336254753551780498081427677782753897299201778428274346714985966328829318067110670104194248315246884346406644886437880251455019329451950816872838540787063933506844181675518163421790362357735222727121349047232970529089826217890874910053395;
            6'd46: xpb[180] = 1024'd20291868274885762124643269914494936036680727705671669108243254573427977511888670902922802919538473783791123123929877151914296730407198728050436176926278861546514569713719988916997973252323587197736315879556812888699196776653744933126842062927884026015248241565940422151764288241520633615645306162546800007731;
            6'd47: xpb[180] = 1024'd77372139527961964983326329597442719160057851561022126408221780898165864024831727164080178972306944094271498356115469310133310586669651461826714411758218659832471498750126848764981299258284128661763499915550048750924213616464453132374481020020834079506954028810775175212286057323999371158583084260844284446398;
            6'd48: xpb[180] = 1024'd10385715096913426443210461875576069538736548290636899580068452157926855200465644515222483810417740095308724180843568033773260602090883861047832521573827417184737753216962491275334386072727464404480486343156044766784869606054264558657141407430554683731839912641492870242701298332549475684402172532516174400734;
            6'd49: xpb[180] = 1024'd67465986349989629301893521558523852662113672145987356880046978482664741713408700776379859863186210405789099413029160191992274458353336594824110756405767215470694682253369351123317712078688005868507670379149280629009886445864972757904780364523504737223545699886327623303223067415028213227339950630813658839401;
            6'd50: xpb[180] = 1024'd479561918941090761777653836657203040792368875602130051893649742425732889042618127522164701297006406826325237757258915632224473774568994045228866221375972822960936720204993633670798893131341611224656806755276644870542435454784184187440751933225341448431583717045318333638308423578317753159038902485548793737;
            6'd51: xpb[180] = 1024'd57559833172017293620460713519604986164169492730952587351872176067163619401985674388679540754065476717306700469942851073851238330037021727821507101053315771108917865756611853481654124899091883075251840842748512507095559275265492383435079709026175394940137370961880071394160077506057055296096817000783033232404;
            6'd52: xpb[180] = 1024'd114640104425093496479143773202552769287546616586303044651850702391901505914928730649836916806833947027787075702128443232070252186299474461597785335885255569394874794793018713329637450905052424539279024878741748369320576115076200582682718666119125448431843158206714824454681846588535792839034595099080517671071;
            6'd53: xpb[180] = 1024'd47653679994044957939027905480686119666225313315917817823697373651662497090562648000979221644944743028824301526856541955710202201720706860818903445700864326747141049259854355839990537719495760281996011306347744385181232104666012008965379053528846052656729042037432519485097087597085897364853683370752407625407;
            6'd54: xpb[180] = 1024'd104733951247121160797710965163633902789602437171268275123675899976400383603505704262136597697713213339304676759042134113929216057983159594595181680532804125033097978296261215687973863725456301746023195342340980247406248944476720208213018010621796106148434829282267272545618856679564634907791461469049892064074;
            6'd55: xpb[180] = 1024'd37747526816072622257595097441767253168281133900883048295522571236161374779139621613278902535824009340341902583770232837569166073404391993816299790348412882385364232763096858198326950539899637488740181769946976263266904934066531634495678398031516710373320713112984967576034097688114739433610549740721782018410;
            6'd56: xpb[180] = 1024'd94827798069148825116278157124715036291658257756233505595501097560899261292082677874436278588592479650822277815955824995788179929666844727592578025180352680671321161799503718046310276545860178952767365805940212125491921773877239833743317355124466763865026500357819720636555866770593476976548327839019266457077;
            6'd57: xpb[180] = 1024'd27841373638100286576162289402848386670336954485848278767347768820660252467716595225578583426703275651859503640683923719428129945088077126813696134995961438023587416266339360556663363360303514695484352233546208141352577763467051260025977742534187368089912384188537415666971107779143581502367416110691156411413;
            6'd58: xpb[180] = 1024'd84921644891176489434845349085796169793714078341198736067326295145398138980659651486735959479471745962339878872869515877647143801350529860589974369827901236309544345302746220404646689366264056159511536269539444003577594603277759459273616699627137421581618171433372168727492876861622319045305194208988640850080;
            6'd59: xpb[180] = 1024'd17935220460127950894729481363929520172392775070813509239172966405159130156293568837878264317582541963377104697597614601287093816771762259811092479643509993661810599769581862914999776180707391902228522697145440019438250592867570885556277087036858025806504055264089863757908117870172423571124282480660530804416;
            6'd60: xpb[180] = 1024'd75015491713204153753412541046877303295769898926163966539151492729897016669236625099035640370351012273857479929783206759506107673034214993587370714475449791947767528805988722762983102186667933366255706733138675881663267432678279084803916044129808079298209842508924616818429886952651161114062060578958015243083;
            6'd61: xpb[180] = 1024'd8029067282155615213296673325010653674448595655778739710998163989658007844870542450177945208461808274894705754511305483146057688455447392808488824291058549300033783272824365273336189001111269108972693160744671897523923422268090511086576431539528683523095726339642311848845127961201265639881148850629905197419;
            6'd62: xpb[180] = 1024'd65109338535231818071979733007958436797825719511129197010976690314395894357813598711335321261230278585375080986696897641365071544717900126584767059122998347585990712309231225121319515007071810572999877196737907759748940262078798710334215388632478737014801513584477064909366897043680003182818926948927389636086;
            6'd63: xpb[180] = 1024'd122189609788308020930662792690906219921202843366479654310955216639133780870756654972492697313998748895855456218882489799584085400980352860361045293954938145871947641345638084969302841013032352037027061232731143621973957101889506909581854345725428790506507300829311817969888666126158740725756705047224874074753;
        endcase
    end

    always_comb begin
        case(flag[60][11:6])
            6'd0: xpb[181] = 1024'd0;
            6'd1: xpb[181] = 1024'd55203185357259482390546924969039570299881540096094427482801887898894772046390572323635002152109544896892682043610588523224035416401585259582163403770546903224213895812473727479655927827475687779744047660337139637834613091479318335864514733135149394731393184660029513000303907134708845251575793318896764029089;
            6'd2: xpb[181] = 1024'd110406370714518964781093849938079140599763080192188854965603775797789544092781144647270004304219089793785364087221177046448070832803170519164326807541093806448427791624947454959311855654951375559488095320674279275669226182958636671729029466270298789462786369320059026000607814269417690503151586637793528058178;
            6'd3: xpb[181] = 1024'd41542860387653705772841847502304278154946193162547598320273808631707420801862578060889935241670960381234896723374272135093042408363535444191330086295309668738951012867849965101337544290909857617921945372624179067139478424217058234628565629722218734927359650565971480970805193330197902737608690130064697602936;
            6'd4: xpb[181] = 1024'd96746045744913188163388772471343848454827733258642025803075696530602192848253150384524937393780505278127578766984860658317077824765120703773493490065856571963164908680323692580993472118385545397665993032961318704974091515696376570493080362857368129658752835226000993971109100464906747989184483448961461632025;
            6'd5: xpb[181] = 1024'd27882535418047929155136770035568986010010846229000769157745729364520069557334583798144868331232375865577111403137955746962049400325485628800496768820072434253688129923226202723019160754344027456099843084911218496444343756954798133392616526309288075123326116471913448941306479525686960223641586941232631176783;
            6'd6: xpb[181] = 1024'd83085720775307411545683695004608556309892386325095196640547617263414841603725156121779870483341920762469793446748544270186084816727070888382660172590619337477902025735699930202675088581819715235843890745248358134278956848434116469257131259444437469854719301131942961941610386660395805475217380260129395205872;
            6'd7: xpb[181] = 1024'd14222210448442152537431692568833693865075499295453939995217650097332718312806589535399801420793791349919326082901639358831056392287435813409663451344835199768425246978602440344700777217778197294277740797198257925749209089692538032156667422896357415319292582377855416911807765721176017709674483752400564750630;
            6'd8: xpb[181] = 1024'd69425395805701634927978617537873264164957039391548367478019537996227490359197161859034803572903336246812008126512227882055091808689021072991826855115382102992639142791076167824356705045253885074021788457535397563583822181171856368021182156031506810050685767037884929912111672855884862961250277071297328779719;
            6'd9: xpb[181] = 1024'd561885478836375919726615102098401720140152361907110832689570830145367068278595272654734510355206834261540762665322970700063384249385998018830133869597965283162364033978677966382393681212367132455638509485297355054074422430277930920718319483426755515259048283797384882309051916665075195707380563568498324477;
            6'd10: xpb[181] = 1024'd55765070836095858310273540071137972020021692458001538315491458729040139114669167596289736662464751731154222806275911493924098800650971257600993537640144868507376259846452405446038321508688054912199686169822436992888687513909596266785233052618576150246652232943826897882612959051373920447283173882465262353566;
            6'd11: xpb[181] = 1024'd110968256193355340700820465040177542319903232554095965798293346627934911161059739919924738814574296628046904849886500017148134217052556517183156941410691771731590155658926132925694249336163742691943733830159576630723300605388914602649747785753725544978045417603856410882916866186082765698858967201362026382655;
            6'd12: xpb[181] = 1024'd42104745866490081692568462604402679875086345524454709152963379461852787870141173333544669752026167215496437486039595105793105792612921442210160220164907634022113376901828643067719937972122224750377583882109476422193552846647336165549283949205645490442618698849768865853114245246862977933316070693633195927413;
            6'd13: xpb[181] = 1024'd97307931223749564083115387573442250174967885620549136635765267360747559916531745657179671904135712112389119529650183629017141209014506701792323623935454537246327272714302370547375865799597912530121631542446616060028165938126654501413798682340794885174011883509798378853418152381571823184891864012529959956502;
            6'd14: xpb[181] = 1024'd28444420896884305074863385137667387730150998590907879990435300194665436625613179070799602841587582699838652165803278717662112784574871626819326902689670399536850493957204880689401554435556394588555481594396515851498418179385076064313334845792714830638585164755710833823615531442352035419348967504801129501260;
            6'd15: xpb[181] = 1024'd83647606254143787465410310106706958030032538687002307473237188093560208672003751394434604993697127596731334209413867240886148200976456886401490306460217302761064389769678608169057482263032082368299529254733655489333031270864394400177849578927864225369978349415740346823919438577060880670924760823697893530349;
            6'd16: xpb[181] = 1024'd14784095927278528457158307670932095585215651657361050827907220927478085381085184808054535931148998184180866845566962329531119776536821811428493585214433165051587611012581118311083170898990564426733379306683555280803283512122815963077385742379784170834551630661652801794116817637841092905381864315969063075107;
            6'd17: xpb[181] = 1024'd69987281284538010847705232639971665885097191753455478310709108826372857427475757131689538083258543081073548889177550852755155192938407071010656988984980068275801506825054845790739098726466252206477426967020694918637896603602134298941900475514933565565944815321682314794420724772549938156957657634865827104196;
            6'd18: xpb[181] = 1024'd1123770957672751839453230204196803440280304723814221665379141660290734136557190545309469020710413668523081525330645941400126768498771996037660267739195930566324728067957355932764787362424734264911277018970594710108148844860555861841436638966853511030518096567594769764618103833330150391414761127136996648954;
            6'd19: xpb[181] = 1024'd56326956314932234230000155173236373740161844819908649148181029559185506182947762868944471172819958565415763568941234464624162184900357255619823671509742833790538623880431083412420715189900422044655324679307734347942761936339874197705951372102002905761911281227624282764922010968038995642990554446033760678043;
            6'd20: xpb[181] = 1024'd111530141672191716620547080142275944040043384916003076630982917458080278229338335192579473324929503462308445612551822987848197601301942515201987075280289737014752519692904810892076643017376109824399372339644873985777375027819192533570466105237152300493304465887653795765225918102747840894566347764930524707132;
            6'd21: xpb[181] = 1024'd42666631345326457612295077706501081595226497886361819985652950291998154938419768606199404262381374049757978248704918076493169176862307440228990354034505599305275740935807321034102331653334591882833222391594773777247627269077614096470002268689072245957877747133566250735423297163528053129023451257201694251890;
            6'd22: xpb[181] = 1024'd97869816702585940002842002675540651895108037982456247468454838190892926984810340929834406414490918946650660292315506599717204593263892699811153757805052502529489636748281048513758259480810279662577270051931913415082240360556932432334517001824221640689270931793595763735727204298236898380599244576098458280979;
            6'd23: xpb[181] = 1024'd29006306375720680994590000239765789450291150952814990823124871024810803693891774343454337351942789534100192928468601688362176168824257624838157036559268364820012857991183558655783948116768761721011120103881813206552492601815353995234053165276141586153844213039508218705924583359017110615056348068369627825737;
            6'd24: xpb[181] = 1024'd84209491732980163385136925208805359750172691048909418305926758923705575740282346667089339504052334430992874972079190211586211585225842884420320440329815268044226753803657286135439875944244449500755167764218952844387105693294672331098567898411290980885237397699537731706228490493725955866632141387266391854826;
            6'd25: xpb[181] = 1024'd15345981406114904376884922773030497305355804019268161660596791757623452449363780080709270441504205018442407608232285300231183160786207809447323719084031130334749975046559796277465564580202931559189017816168852635857357934553093893998104061863210926349810678945450186676425869554506168101089244879537561399584;
            6'd26: xpb[181] = 1024'd70549166763374386767431847742070067605237344115362589143398679656518224495754352404344272593613749915335089651842873823455218577187793069029487122854578033558963870859033523757121492407678619338933065476505992273691971026032412229862618794998360321081203863605479699676729776689215013352665038198434325428673;
            6'd27: xpb[181] = 1024'd1685656436509127759179845306295205160420457085721332498068712490436101204835785817964203531065620502784622287995968912100190152748157994056490401608793895849487092101936033899147181043637101397366915528455892065162223267290833792762154958450280266545777144851392154646927155749995225587122141690705494973431;
            6'd28: xpb[181] = 1024'd56888841793768610149726770275334775460301997181815759980870600389330873251226358141599205683175165399677304331606557435324225569149743253638653805379340799073700987914409761378803108871112789177110963188793031702996836358770152128626669691585429661277170329511421667647231062884704070838697935009602259002520;
            6'd29: xpb[181] = 1024'd112092027151028092540273695244374345760183537277910187463672488288225645297616930465234207835284710296569986375217145958548260985551328513220817209149887702297914883726883488858459036698588476956855010849130171340831449450249470464491184424720579056008563514171451180647534970019412916090273728328499023031609;
            6'd30: xpb[181] = 1024'd43228516824162833532021692808599483315366650248268930818342521122143522006698363878854138772736580884019519011370241047193232561111693438247820487904103564588438104969785999000484725334546959015288860901080071132301701691507892027390720588172499001473136795417363635617732349080193128324730831820770192576367;
            6'd31: xpb[181] = 1024'd98431702181422315922568617777639053615248190344363358301144409021038294053088936202489140924846125780912201054980829570417267977513278697829983891674650467812652000782259726480140653162022646795032908561417210770136314782987210363255235321307648396204529980077393148618036256214901973576306625139666956605456;
            6'd32: xpb[181] = 1024'd29568191854557056914316615341864191170431303314722101655814441854956170762170369616109071862297996368361733691133924659062239553073643622856987170428866330103175222025162236622166341797981128853466758613367110561606567024245631926154771484759568341669103261323305603588233635275682185810763728631938126150214;
            6'd33: xpb[181] = 1024'd84771377211816539304863540310903761470312843410816529138616329753850942808560941939744074014407541265254415734744513182286274969475228882439150574199413233327389117837635964101822269625456816633210806273704250199441180115724950262019286217894717736400496445983335116588537542410391031062339521950834890179303;
            6'd34: xpb[181] = 1024'd15907866884951280296611537875128899025495956381175272493286362587768819517642375353364004951859411852703948370897608270931246545035593807466153852953629095617912339080538474243847958261415298691644656325654149990911432356983371824918822381346637681865069727229247571558734921471171243296796625443106059724061;
            6'd35: xpb[181] = 1024'd71111052242210762687158462844168469325377496477269699976088250486663591564032947676999007103968956749596630414508196794155281961437179067048317256724175998842126234893012201723503886088890986471388703985991289628746045448462690160783337114481787076596462911889277084559038828605880088548372418762002823753150;
            6'd36: xpb[181] = 1024'd2247541915345503678906460408393606880560609447628443330758283320581468273114381090618938041420827337046163050661291882800253536997543992075320535478391861132649456135914711865529574724849468529822554037941189420216297689721111723682873277933707022061036193135189539529236207666660300782829522254273993297908;
            6'd37: xpb[181] = 1024'd57450727272604986069453385377433177180442149543722870813560171219476240319504953414253940193530372233938845094271880406024288953399129251657483939248938764356863351948388439345185502552325156309566601698278329058050910781200430059547388011068856416792429377795219052529540114801369146034405315573170757326997;
            6'd38: xpb[181] = 1024'd112653912629864468460000310346472747480323689639817298296362059118371012365895525737888942345639917130831527137882468929248324369800714511239647343019485667581077247760862166824841430379800844089310649358615468695885523872679748395411902744204005811523822562455248565529844021936077991285981108892067521356086;
            6'd39: xpb[181] = 1024'd43790402302999209451748307910697885035506802610176041651032091952288889074976959151508873283091787718281059774035564017893295945361079436266650621773701529871600469003764676966867119015759326147744499410565368487355776113938169958311438907655925756988395843701161020500041400996858203520438212384338690900844;
            6'd40: xpb[181] = 1024'd98993587660258691842295232879737455335388342706270469133833979851183661121367531475143875435201332615173741817646152541117331361762664695848814025544248433095814364816238404446523046843235013927488547070902508125190389205417488294175953640791075151719789028361190533500345308131567048772014005703235454929933;
            6'd41: xpb[181] = 1024'd30130077333393432834043230443962592890571455676629212488504012685101537830448964888763806372653203202623274453799247629762302937323029620875817304298464295386337586059140914588548735479193495985922397122852407916660641446675909857075489804242995097184362309607102988470542687192347261006471109195506624474691;
            6'd42: xpb[181] = 1024'd85333262690652915224590155413002163190452995772723639971305900583996309876839537212398808524762748099515956497409836152986338353724614880457980708069011198610551481871614642068204663306669183765666444783189547554495254538155228192940004537378144491915755494267132501470846594327056106258046902514403388503780;
            6'd43: xpb[181] = 1024'd16469752363787656216338152977227300745636108743082383325975933417914186585920970626018739462214618686965489133562931241631309929284979805484983986823227060901074703114517152210230351942627665824100294835139447345965506779413649755839540700830064437380328775513044956441043973387836318492504006006674558048538;
            6'd44: xpb[181] = 1024'd71672937721047138606885077946266871045517648839176810808777821316808958632311542949653741614324163583858171177173519764855345345686565065067147390593773964125288598926990879689886279770103353603844342495476586983800119870892968091704055433965213832111721960173074469441347880522545163744079799325571322077627;
            6'd45: xpb[181] = 1024'd2809427394181879598633075510492008600700761809535554163447854150726835341392976363273672551776034171307703813326614853500316921246929990094150669347989826415811820169893389831911968406061835662278192547426486775270372112151389654603591597417133777576295241418986924411545259583325375978536902817842491622385;
            6'd46: xpb[181] = 1024'd58012612751441361989180000479531578900582301905629981646249742049621607387783548686908674703885579068200385856937203376724352337648515249676314073118536729640025715982367117311567896233537523442022240207763626413104985203630707990468106330552283172307688426079016437411849166718034221230112696136739255651474;
            6'd47: xpb[181] = 1024'd113215798108700844379726925448571149200463842001724409129051629948516379434174121010543676855995123965093067900547791899948387754050100509258477476889083632864239611794840844791223824061013211221766287868100766050939598295110026326332621063687432567039081610739045950412153073852743066481688489455636019680563;
            6'd48: xpb[181] = 1024'd44352287781835585371474923012796286755646954972083152483721662782434256143255554424163607793446994552542600536700886988593359329610465434285480755643299495154762833037743354933249512696971693280200137920050665842409850536368447889232157227139352512503654891984958405382350452913523278716145592947907189225321;
            6'd49: xpb[181] = 1024'd99555473139095067762021847981835857055528495068177579966523550681329028189646126747798609945556539449435282580311475511817394746012050693867644159413846398378976728850217082412905440524447381059944185580387805480244463627847766225096671960274501907235048076644987918382654360048232123967721386266803953254410;
            6'd50: xpb[181] = 1024'd30691962812229808753769845546060994610711608038536323321193583515246904898727560161418540883008410036884815216464570600462366321572415618894647438168062260669499950093119592554931129160405863118378035632337705271714715869106187787996208123726421852699621357890900373352851739109012336202178489759075122799168;
            6'd51: xpb[181] = 1024'd85895148169489291144316770515100564910593148134630750803995471414141676945118132485053543035117954933777497260075159123686401737974000878476810841938609163893713845905593320034587056987881550898122083292674844909549328960585506123860722856861571247431014542550929886353155646243721181453754283077971886828257;
            6'd52: xpb[181] = 1024'd17031637842624032136064768079325702465776261104989494158665504248059553654199565898673473972569825521227029896228254212331373313534365803503814120692825026184237067148495830176612745623840032956555933344624744701019581201843927686760259020313491192895587823796842341323353025304501393688211386570243056373015;
            6'd53: xpb[181] = 1024'd72234823199883514526611693048365272765657801201083921641467392146954325700590138222308476124679370418119711939838842735555408729935951063085977524463371929408450962960969557656268673451315720736299981004961884338854194293323246022624773753448640587626981008456871854323656932439210238939787179889139820402104;
            6'd54: xpb[181] = 1024'd3371312873018255518359690612590410320840914171442664996137424980872202409671571635928407062131241005569244575991937824200380305496315988112980803217587791698974184203872067798294362087274202794733831056911784130324446534581667585524309916900560533091554289702784309293854311499990451174244283381410989946862;
            6'd55: xpb[181] = 1024'd58574498230277737908906615581629980620722454267537092478939312879766974456062143959563409214240785902461926619602526347424415721897901247695144206988134694923188080016345795277950289914749890574477878717248923768159059626060985921388824650035709927822947474362813822294158218634699296425820076700307753975951;
            6'd56: xpb[181] = 1024'd113777683587537220299453540550669550920603994363631519961741200778661746502452716283198411366350330799354608663213114870648451138299486507277307610758681598147401975828819522757606217742225578354221926377586063405993672717540304257253339383170859322554340659022843335294462125769408141677395870019204518005040;
            6'd57: xpb[181] = 1024'd44914173260671961291201538114894688475787107333990263316411233612579623211534149696818342303802201386804141299366209959293422713859851432304310889512897460437925197071722032899631906378184060412655776429535963197463924958798725820152875546622779268018913940268755790264659504830188353911852973511475687549798;
            6'd58: xpb[181] = 1024'd100117358617931443681748463083934258775668647430084690799213121511474395257924722020453344455911746283696823342976798482517458130261436691886474293283444363662139092884195760379287834205659748192399824089873102835298538050278044156017390279757928662750307124928785303264963411964897199163428766830372451578887;
            6'd59: xpb[181] = 1024'd31253848291066184673496460648159396330851760400443434153883154345392271967006155434073275393363616871146355979129893571162429705821801616913477572037660225952662314127098270521313522841618230250833674141823002626768790291536465718916926443209848608214880406174697758235160791025677411397885870322643621123645;
            6'd60: xpb[181] = 1024'd86457033648325667064043385617198966630733300496537861636685042244287044013396727757708277545473161768039038022740482094386465122223386876495640975808207129176876209939571998000969450669093918030577721802160142264603403383015784054781441176344998002946273590834727271235464698160386256649461663641540385152734;
            6'd61: xpb[181] = 1024'd17593523321460408055791383181424104185916413466896604991355075078204920722478161171328208482925032355488570658893577183031436697783751801522644254562422991467399431182474508142995139305052400089011571854110042056073655624274205617680977339796917948410846872080639726205662077221166468883918767133811554697492;
            6'd62: xpb[181] = 1024'd72796708678719890446338308150463674485797953562991032474156962977099692768868733494963210635034577252381252702504165706255472114185337061104807658332969894691613326994948235622651067132528087868755619514447181693908268715753523953545492072932067343142240056740669239205965984355875314135494560452708318726581;
            6'd63: xpb[181] = 1024'd3933198351854631438086305714688812040981066533349775828826995811017569477950166908583141572486447839830785338657260794900443689745701986131810937087185756982136548237850745764676755768486569927189469566397081485378520957011945516445028236383987288606813337986581694176163363416655526369951663944979488271339;
        endcase
    end

    always_comb begin
        case(flag[60][16:12])
            5'd0: xpb[182] = 1024'd0;
            5'd1: xpb[182] = 1024'd59136383709114113828633230683728382340862606629444203311628883709912341524340739232218143724595992736723467382267849318124479106147287245713974340857732660206350444050324473244332683595962257706933517226734221123213134048491263852309542969519136683338206522646611207176467270551364371621527457263876252300428;
            5'd2: xpb[182] = 1024'd118272767418228227657266461367456764681725213258888406623257767419824683048681478464436287449191985473446934764535698636248958212294574491427948681715465320412700888100648946488665367191924515413867034453468442246426268096982527704619085939038273366676413045293222414352934541102728743243054914527752504600856;
            5'd3: xpb[182] = 1024'd53342455443217600087100764646370714277889392762596925806754796064760129235713078786639359959130303900727252739346054519794373477600641402586762897556866939685360657581402202395367811596369567399490354071815423523275041295252894783963650338874180600747799664525716563499295283580164481847463681965003162416953;
            5'd4: xpb[182] = 1024'd112478839152331713915733995330099096618751999392041129118383679774672470760053818018857503683726296637450720121613903837918852583747928648300737238414599599891711101631726675639700495192331825106423871298549644646488175343744158636273193308393317284086006187172327770675762554131528853468991139228879414717381;
            5'd5: xpb[182] = 1024'd47548527177321086345568298609013046214916178895749648301880708419607916947085418341060576193664615064731038096424259721464267849053995559459551454256001219164370871112479931546402939596776877092047190916896625923336948542014525715617757708229224518157392806404821919822123296608964592073399906666130072533478;
            5'd6: xpb[182] = 1024'd106684910886435200174201529292741428555778785525193851613509592129520258471426157573278719918260607801454505478692109039588746955201282805173525795113733879370721315162804404790735623192739134798980708143630847046550082590505789567927300677748361201495599329051433126998590567160328963694927363930006324833906;
            5'd7: xpb[182] = 1024'd41754598911424572604035832571655378151942965028902370797006620774455704658457757895481792428198926228734823453502464923134162220507349716332340010955135498643381084643557660697438067597184186784604027761977828323398855788776156647271865077584268435566985948283927276144951309637764702299336131367256982650003;
            5'd8: xpb[182] = 1024'd100890982620538686432669063255383760492805571658346574108635504484368046182798497127699936152794918965458290835770314241258641326654636962046314351812868158849731528693882133941770751193146444491537544988712049446611989837267420499581408047103405118905192470930538483321418580189129073920863588631133234950431;
            5'd9: xpb[182] = 1024'd35960670645528058862503366534297710088969751162055093292132533129303492369830097449903008662733237392738608810580670124804056591960703873205128567654269778122391298174635389848473195597591496477160864607059030723460763035537787578925972446939312352976579090163032632467779322666564812525272356068383892766528;
            5'd10: xpb[182] = 1024'd95097054354642172691136597218026092429832357791499296603761416839215833894170836682121152387329230129462076192848519442928535698107991118919102908512002438328741742224959863092805879193553754184094381833793251846673897084029051431235515416458449036314785612809643839644246593217929184146799813332260145066956;
            5'd11: xpb[182] = 1024'd30166742379631545120970900496940042025996537295207815787258445484151280081202437004324224897267548556742394167658875326473950963414058030077917124353404057601401511705713118999508323597998806169717701452140233123522670282299418510580079816294356270386172232042137988790607335695364922751208580769510802883053;
            5'd12: xpb[182] = 1024'd89303126088745658949604131180668424366859143924652019098887329194063621605543176236542368621863541293465861549926724644598430069561345275791891465211136717807751955756037592243841007193961063876651218678874454246735804330790682362889622785813492953724378754688749195967074606246729294372736038033387055183481;
            5'd13: xpb[182] = 1024'd24372814113735031379438434459582373963023323428360538282384357838999067792574776558745441131801859720746179524737080528143845334867412186950705681052538337080411725236790848150543451598406115862274538297221435523584577529061049442234187185649400187795765373921243345113435348724165032977144805470637712999578;
            5'd14: xpb[182] = 1024'd83509197822849145208071665143310756303885930057804741594013241548911409316915515790963584856397852457469646907004929846268324441014699432664680021910270997286762169287115321394876135194368373569208055523955656646797711577552313294543730155168536871133971896567854552289902619275529404598672262734513965300006;
            5'd15: xpb[182] = 1024'd18578885847838517637905968422224705900050109561513260777510270193846855503947116113166657366336170884749964881815285729813739706320766343823494237751672616559421938767868577301578579598813425554831375142302637923646484775822680373888294555004444105205358515800348701436263361752965143203081030171764623116103;
            5'd16: xpb[182] = 1024'd77715269556952631466539199105953088240912716190957464089139153903759197028287855345384801090932163621473432264083135047938218812468053589537468578609405276765772382818193050545911263194775683261764892369036859046859618824313944226197837524523580788543565038446959908612730632304329514824608487435640875416531;
            5'd17: xpb[182] = 1024'd12784957581942003896373502384867037837076895694665983272636182548694643215319455667587873600870482048753750238893490931483634077774120500696282794450806896038432152298946306452613707599220735247388211987383840323708392022584311305542401924359488022614951657679454057759091374781765253429017254872891533232628;
            5'd18: xpb[182] = 1024'd71921341291056117725006733068595420177939502324110186584265066258606984739660194899806017325466474785477217621161340249608113183921407746410257135308539556244782596349270779696946391195182992954321729214118061446921526071075575157851944893878624705953158180326065264935558645333129625050544712136767785533056;
            5'd19: xpb[182] = 1024'd6991029316045490154841036347509369774103681827818705767762094903542430926691795222009089835404793212757535595971696133153528449227474657569071351149941175517442365830024035603648835599628044939945048832465042723770299269345942237196509293714531940024544799558559414081919387810565363654953479574018443349153;
            5'd20: xpb[182] = 1024'd66127413025159603983474267031237752114966288457262909079390978613454772451032534454227233560000785949481002978239545451278007555374761903283045692007673835723792809880348508847981519195590302646878566059199263846983433317837206089506052263233668623362751322205170621258386658361929735276480936837894695649581;
            5'd21: xpb[182] = 1024'd1197101050148976413308570310151701711130467960971428262888007258390218638064134776430306069939104376761320953049901334823422820680828814441859907849075454996452579361101764754683963600035354632501885677546245123832206516107573168850616663069575857434137941437664770404747400839365473880889704275145353465678;
            5'd22: xpb[182] = 1024'd60333484759263090241941800993880084051993074590415631574516890968302560162404874008648449794535097113484788335317750652947901926828116060155834248706808115202803023411426237999016647195997612339435402904280466247045340564598837021160159632588712540772344464084275977581214671390729845502417161539021605766106;
            5'd23: xpb[182] = 1024'd119469868468377204070575031677608466392855681219859834886145774678214901686745613240866593519131089850208255717585599971072381032975403305869808589564540775409153467461750711243349330791959870046368920131014687370258474613090100873469702602107849224110550986730887184757681941942094217123944618802897858066534;
            5'd24: xpb[182] = 1024'd54539556493366576500409334956522415989019860723568354069642803323150347873777213563069666029069408277488573692395955854617796298281470217028622805405942394681813236942503967150051775196404922031992239749361668647107247811360467952814267001943756458181937605963381333904042684419529955728353386240148515882631;
            5'd25: xpb[182] = 1024'd113675940202480690329042565640250798329882467353012557381271687033062689398117952795287809753665401014212041074663805172742275404428757462742597146263675054888163680992828440394384458792367179738925756976095889770320381859851731805123809971462893141520144128609992541080509954970894327349880843504024768183059;
            5'd26: xpb[182] = 1024'd48745628227470062758876868919164747926046646856721076564768715677998135585149553117490882263603719441492359049474161056287690669734824373901411362105076674160823450473581696301086903196812231724549076594442871047169155058122098884468374371298800375591530747842486690226870697448330065954289610941275425999156;
            5'd27: xpb[182] = 1024'd107882011936584176587510099602893130266909253486165279876397599387910477109490292349709025988199712178215826431742010374412169775882111619615385702962809334367173894523906169545419586792774489431482593821177092170382289106613362736777917340817937058929737270489097897403337967999694437575817068205151678299584;
            5'd28: xpb[182] = 1024'd42951699961573549017344402881807079863073432989873799059894628032845923296521892671912098498138030605496144406552366257957585041188178530774199918804210953639833664004659425452122031197219541417105913439524073447231062304883729816122481740653844293001123889721592046549698710477130176180225835642402336115681;
            5'd29: xpb[182] = 1024'd102088083670687662845977633565535462203936039619318002371523511742758264820862631904130242222734023342219611788820215576082064147335465776488174259661943613846184108054983898696454714793181799124039430666258294570444196353374993668432024710172980976339330412368203253726165981028494547801753292906278588416109;
            5'd30: xpb[182] = 1024'd37157771695677035275811936844449411800100219123026521555020540387693711007894232226333314732672341769499929763630571459627479412641532687646988475503345233118843877535737154603157159197626851109662750284605275847292969551645360747776589110008888210410717031600697402872526723505930286406162060343529246232206;
            5'd31: xpb[182] = 1024'd96294155404791149104445167528177794140962825752470724866649424097606052532234971458551458457268334506223397145898420777751958518788819933360962816361077893325194321586061627847489842793589108816596267511339496970506103600136624600086132079528024893748923554247308610048993994057294658027689517607405498532634;
        endcase
    end

    always_comb begin
        case(flag[61][5:0])
            6'd0: xpb[183] = 1024'd0;
            6'd1: xpb[183] = 1024'd77715269556952631466539199105953088240912716190957464089139153903759197028287855345384801090932163621473432264083135047938218812468053589537468578609405276765772382818193050545911263194775683261764892369036859046859618824313944226197837524523580788543565038446959908612730632304329514824608487435640875416531;
            6'd2: xpb[183] = 1024'd31363843429780521534279470807091743737127005256179244050146452742541498719266571780754530967206652933503715120708776661297373784094886844519777032202479512597854091066814883754192287198034160802219587129686478247354876798406991679430696479363932127820310173479802759195354736534730396632098285044656156348731;
            6'd3: xpb[183] = 1024'd109079112986733153000818669913044831978039721447136708139285606646300695747554427126139332058138816554977147384791911709235592596562940434057245610811884789363626473885007934300103550392809844063984479498723337294214495622720935905628534003887512916363875211926762667808085368839059911456706772480297031765262;
            6'd4: xpb[183] = 1024'd62727686859561043068558941614183487474254010512358488100292905485082997438533143561509061934413305867007430241417553322594747568189773689039554064404959025195708182133629767508384574396068321604439174259372956494709753596813983358861392958727864255640620346959605518390709473069460793264196570089312312697462;
            6'd5: xpb[183] = 1024'd16376260732388933136299213315322142970468299577580268061300204323865299129511859996878791810687795179037713098043194935953902539816606944021862517998033261027789890382251600716665598399326799144893869020022575695205011570907030812094251913568215594917365481992448368973333577299861675071686367698327593629662;
            6'd6: xpb[183] = 1024'd94091530289341564602838412421275231211381015768537732150439358227624496157799715342263592901619958800511145362126329983892121352284660533559331096607438537793562273200444651262576861594102482406658761389059434742064630395220975038292089438091796383460930520439408277586064209604191189896294855133968469046193;
            6'd7: xpb[183] = 1024'd47740104162169454670578684122413886707595304833759512111446657066406797848778431777633322777894448112541428218751971597251276323911493788541639550200512773625643981449066484470857885597360959947113456149709053942559888369314022491524948392932147722737675655472251128168688313834592071703784652742983749978393;
            6'd8: xpb[183] = 1024'd1388678034997344738318955823552542203809593898981292072453955905189099539757148213003052654168937424571711075377613210610431295538327043523948003793587009457725689697688317679138909600619437487568150910358673143055146343407069944757807347772499062014420790505093978751312418064992953511274450351999030910593;
            6'd9: xpb[183] = 1024'd79103947591949976204858154929505630444722310089938756161593109808948296568045003558387853745101101046045143339460748258548650108006380633061416582402992286223498072515881368225050172795395120749333043279395532189914765167721014170955644872296079850557985828952053887364043050369322468335882937787639906327124;
            6'd10: xpb[183] = 1024'd32752521464777866272598426630644285940936599155160536122600408647730598259023719993757583621375590358075426196086389871907805079633213888043725035996066522055579780764503201433331196798653598289787738040045151390410023141814061624188503827136431189834730963984896737946667154599723350143372735396655187259324;
            6'd11: xpb[183] = 1024'd110467791021730497739137625736597374181849315346118000211739562551489795287311575339142384712307753979548858460169524919846023892101267477581193614605471798821352163582696251979242459993429281551552630409082010437269641966128005850386341351660011978378296002431856646559397786904052864967981222832296062675855;
            6'd12: xpb[183] = 1024'd64116364894558387806877897437736029678063604411339780172746861390272096978290291774512114588582243291579141316795166533205178863728100732563502068198546034653433871831318085187523483996687759092007325169731629637764899940221053303619200306500363317655041137464699497142021891134453746775471020441311343608055;
            6'd13: xpb[183] = 1024'd17764938767386277874618169138874685174277893476561560133754160229054398669269008209881844464856732603609424173420808146564333835354933987545810521791620270485515580079939918395804507999946236632462019930381248838260157914314100756852059261340714656931786272497542347724645995364854628582960818050326624540255;
            6'd14: xpb[183] = 1024'd95480208324338909341157368244827773415190609667519024222893314132813595697556863555266645555788896225082856437503943194502552647822987577083279100401025547251287962898132968941715771194721919894226912299418107885119776738628044983049896785864295445475351310944502256337376627669184143407569305485967499956786;
            6'd15: xpb[183] = 1024'd49128782197166799408897639945966428911404898732740804183900612971595897388535579990636375432063385537113139294129584807861707619449820832065587553994099783083369671146754802149996795197980397434681607060067727085615034712721092436282755740704646784752096445977345106920000731899585025215059103094982780888986;
            6'd16: xpb[183] = 1024'd2777356069994689476637911647105084407619187797962584144907911810378199079514296426006105308337874849143422150755226421220862591076654087047896007587174018915451379395376635358277819201238874975136301820717346286110292686814139889515614695544998124028841581010187957502624836129985907022548900703998061821186;
            6'd17: xpb[183] = 1024'd80492625626947320943177110753058172648531903988920048234047065714137396107802151771390906399270038470616854414838361469159081403544707676585364586196579295681223762213569685904189082396014558236901194189754205332969911511128084115713452220068578912572406619457147866115355468434315421847157388139638937237717;
            6'd18: xpb[183] = 1024'd34141199499775211010917382454196828144746193054141828195054364552919697798780868206760636275544527782647137271464003082518236375171540931567673039789653531513305470462191519112470106399273035777355888950403824533465169485221131568946311174908930251849151754489990716697979572664716303654647185748654218169917;
            6'd19: xpb[183] = 1024'd111856469056727842477456581560149916385658909245099292284193518456678894827068723552145437366476691404120569535547138130456455187639594521105141618399058808279077853280384569658381369594048719039120781319440683580324788309535075795144148699432511040392716792936950625310710204969045818479255673184295093586448;
            6'd20: xpb[183] = 1024'd65505042929555732545196853261288571881873198310321072245200817295461196518047439987515167242751180716150852392172779743815610159266427776087450071992133044111159561529006402866662393597307196579575476080090302780820046283628123248377007654272862379669461927969793475893334309199446700286745470793310374518648;
            6'd21: xpb[183] = 1024'd19153616802383622612937124962427227378087487375542852206208116134243498209026156422884897119025670028181135248798421357174765130893261031069758525585207279943241269777628236074943417600565674120030170840739921981315304257721170701609866609113213718946207063002636326475958413429847582094235268402325655450848;
            6'd22: xpb[183] = 1024'd96868886359336254079476324068380315619000203566500316295347270038002695237314011768269698209957833649654567512881556405112983943361314620607227104194612556709013652595821286620854680795341357381795063209776781028174923082035114927807704133636794507489772101449596235088689045734177096918843755837966530867379;
            6'd23: xpb[183] = 1024'd50517460232164144147216595769518971115214492631722096256354568876784996928292728203639428086232322961684850369507198018472138914988147875589535557787686792541095360844443119829135704798599834922249757970426400228670181056128162381040563088477145846766517236482439085671313149964577978726333553446981811799579;
            6'd24: xpb[183] = 1024'd4166034104992034214956867470657626611428781696943876217361867715567298619271444639009157962506812273715133226132839631831293886614981130571844011380761028373177069093064953037416728801858312462704452731076019429165439030221209834273422043317497186043262371515281936253937254194978860533823351055997092731779;
            6'd25: xpb[183] = 1024'd81881303661944665681496066576610714852341497887901340306501021619326495647559299984393959053438975895188565490215974679769512699083034720109312589990166305138949451911258003583327991996633995724469345100112878476025057854535154060471259567841077974586827409962241844866667886499308375358431838491637968148310;
            6'd26: xpb[183] = 1024'd35529877534772555749236338277749370348555786953123120267508320458108797338538016419763688929713465207218848346841616293128667670709867975091621043583240540971031160159879836791609015999892473264924039860762497676520315828628201513704118522681429313863572544995084695449291990729709257165921636100653249080510;
            6'd27: xpb[183] = 1024'd113245147091725187215775537383702458589468503144080584356647474361867994366825871765148490020645628828692280610924751341066886483177921564629089622192645817736803542978072887337520279194668156526688932229799356723379934652942145739901956047205010102407137583442044604062022623034038771990530123536294124497041;
            6'd28: xpb[183] = 1024'd66893720964553077283515809084841114085682792209302364317654773200650296057804588200518219896920118140722563467550392954426041454804754819611398075785720053568885251226694720545801303197926634067143626990448975923875192627035193193134815002045361441683882718474887454644646727264439653798019921145309405429241;
            6'd29: xpb[183] = 1024'd20542294837380967351256080785979769581897081274524144278662072039432597748783304635887949773194607452752846324176034567785196426431588074593706529378794289400966959475316553754082327201185111607598321751098595124370450601128240646367673956885712780960627853507730305227270831494840535605509718754324686361441;
            6'd30: xpb[183] = 1024'd98257564394333598817795279891932857822809797465481608367801225943191794777071159981272750864126771074226278588259169615723415238899641664131175107988199566166739342293509604299993590395960794869363214120135454171230069425442184872565511481409293569504192891954690213840001463799170050430118206189965561777972;
            6'd31: xpb[183] = 1024'd51906138267161488885535551593071513319024086530703388328808524781974096468049876416642480740401260386256561444884811229082570210526474919113483561581273801998821050542131437508274614399219272409817908880785073371725327399535232325798370436249644908780938026987533064422625568029570932237608003798980842710172;
            6'd32: xpb[183] = 1024'd5554712139989378953275823294210168815238375595925168289815823620756398159028592852012210616675749698286844301510452842441725182153308174095792015174348037830902758790753270716555638402477749950272603641434692572220585373628279779031229391089996248057683162020375915005249672259971814045097801407996123642372;
            6'd33: xpb[183] = 1024'd83269981696942010419815022400163257056151091786882632378954977524515595187316448197397011707607913319760276565593587890379943994621361763633260593783753314596675141608946321262466901597253433212037496010471551619080204197942224005229066915613577036601248200467335823617980304564301328869706288843636999058903;
            6'd34: xpb[183] = 1024'd36918555569769900487555294101301912552365380852104412339962276363297896878295164632766741583882402631790559422219229503739098966248195018615569047376827550428756849857568154470747925600511910752492190771121170819575462172035271458461925870453928375877993335500178674200604408794702210677196086452652279991103;
            6'd35: xpb[183] = 1024'd114633825126722531954094493207255000793278097043061876429101430267057093906583019978151542674814566253263991686302364551677317778716248608153037625986232827194529232675761205016659188795287594014257083140158029866435080996349215684659763394977509164421558373947138582813335041099031725501804573888293155407634;
            6'd36: xpb[183] = 1024'd68282398999550422021834764908393656289492386108283656390108729105839395597561736413521272551089055565294274542928006165036472750343081863135346079579307063026610940924383038224940212798546071554711777900807649066930338970442263137892622349817860503698303508979981433395959145329432607309294371497308436339834;
            6'd37: xpb[183] = 1024'd21930972872378312089575036609532311785706675173505436351116027944621697288540452848891002427363544877324557399553647778395627721969915118117654533172381298858692649173004871433221236801804549095166472661457268267425596944535310591125481304658211842975048644012824283978583249559833489116784169106323717272034;
            6'd38: xpb[183] = 1024'd99646242429330943556114235715485400026619391364462900440255181848380894316828308194275803518295708498797989663636782826333846534437968707655123111781786575624465031991197921979132499996580232356931365030494127314285215768849254817323318829181792631518613682459784192591313881864163003941392656541964592688565;
            6'd39: xpb[183] = 1024'd53294816302158833623854507416624055522833680429684680401262480687163196007807024629645533394570197810828272520262424439693001506064801962637431565374860811456546740239819755187413523999838709897386059791143746514780473742942302270556177784022143970795358817492627043173937986094563885748882454150979873620765;
            6'd40: xpb[183] = 1024'd6943390174986723691594779117762711019047969494906460362269779525945497698785741065015263270844687122858555376888066053052156477691635217619740018967935047288628448488441588395694548003097187437840754551793365715275731717035349723789036738862495310072103952525469893756562090324964767556372251759995154552965;
            6'd41: xpb[183] = 1024'd84658659731939355158133978223715799259960685685863924451408933429704694727073596410400064361776850744331987640971201100990375290159688807157208597577340324054400831306634638941605811197872870699605646920830224762135350541349293949986874263386076098615668990972429802369292722629294282380980739195636029969496;
            6'd42: xpb[183] = 1024'd38307233604767245225874249924854454756174974751085704412416232268486996418052312845769794238051340056362270497596842714349530261786522062139517051170414559886482539555256472149886835201131348240060341681479843962630608515442341403219733218226427437892414126005272652951916826859695164188470536804651310901696;
            6'd43: xpb[183] = 1024'd116022503161719876692413449030807542997087690942043168501555386172246193446340168191154595328983503677835702761679977762287749074254575651676985629779819836652254922373449522695798098395907031501825234050516703009490227339756285629417570742750008226435979164452232561564647459164024679013079024240292186318227;
            6'd44: xpb[183] = 1024'd69671077034547766760153720731946198493301980007264948462562685011028495137318884626524325205257992989865985618305619375646904045881408906659294083372894072484336630622071355904079122399165509042279928811166322209985485313849333082650429697590359565712724299485075412147271563394425560820568821849307467250427;
            6'd45: xpb[183] = 1024'd23319650907375656827893992433084853989516269072486728423569983849810796828297601061894055081532482301896268474931260989006059017508242161641602536965968308316418338870693189112360146402423986582734623571815941410480743287942380535883288652430710904989469434517918262729895667624826442628058619458322748182627;
            6'd46: xpb[183] = 1024'd101034920464328288294433191539037942230428985263444192512709137753569993856585456407278856172464645923369700739014396036944277829976295751179071115575373585082190721688886239658271409597199669844499515940852800457340362112256324762081126176954291693533034472964878171342626299929155957452667106893963623599158;
            6'd47: xpb[183] = 1024'd54683494337156178362173463240176597726643274328665972473716436592352295547564172842648586048739135235399983595640037650303432801603129006161379569168447820914272429937508072866552433600458147384954210701502419657835620086349372215313985131794643032809779607997721021925250404159556839260156904502978904531358;
            6'd48: xpb[183] = 1024'd8332068209984068429913734941315253222857563393887752434723735431134597238542889278018315925013624547430266452265679263662587773229962261143688022761522056746354138186129906074833457603716624925408905462152038858330878060442419668546844086634994372086524743030563872507874508389957721067646702111994185463558;
            6'd49: xpb[183] = 1024'd86047337766936699896452934047268341463770279584845216523862889334893794266830744623403117015945788168903698716348814311600806585698015850681156601370927333512126521004322956620744720798492308187173797831188897905190496884756363894744681611158575160630089781477523781120605140694287235892255189547635060880089;
            6'd50: xpb[183] = 1024'd39695911639764589964193205748406996959984568650066996484870188173676095957809461058772846892220277480933981572974455924959961557324849105663465054964001569344208229252944789829025744801750785727628492591838517105685754858849411347977540565998926499906834916510366631703229244924688117699744987156650341812289;
            6'd51: xpb[183] = 1024'd117411181196717221430732404854360085200897284841024460574009342077435292986097316404157647983152441102407413837057590972898180369792902695200933633573406846109980612071137840374937007996526468989393384960875376152545373683163355574175378090522507288450399954957326540315959877229017632524353474592291217228820;
            6'd52: xpb[183] = 1024'd71059755069545111498472676555498740697111573906246240535016640916217594677076032839527377859426930414437696693683232586257335341419735950183242087166481081942062320319759673583218031999784946529848079721524995353040631657256403027408237045362858627727145089990169390898583981459418514331843272201306498161020;
            6'd53: xpb[183] = 1024'd24708328942373001566212948256637396193325862971468020496023939754999896368054749274897107735701419726467979550308874199616490313046569205165550540759555317774144028568381506791499056003043424070302774482174614553535889631349450480641096000203209967003890225023012241481208085689819396139333069810321779093220;
            6'd54: xpb[183] = 1024'd102423598499325633032752147362590484434238579162425484585163093658759093396342604620281908826633583347941411814392009247554709125514622794703019119368960594539916411386574557337410319197819107332067666851211473600395508455663394706838933524726790755547455263469972150093938717994148910963941557245962654509751;
            6'd55: xpb[183] = 1024'd56072172372153523100492419063729139930452868227647264546170392497541395087321321055651638702908072659971694671017650860913864097141456049685327572962034830371998119635196390545691343201077584872522361611861092800890766429756442160071792479567142094824200398502815000676562822224549792771431354854977935441951;
            6'd56: xpb[183] = 1024'd9720746244981413168232690764867795426667157292869044507177691336323696778300037491021368579182561972001977527643292474273019068768289304667636026555109066204079827883818223753972367204336062412977056372510712001386024403849489613304651434407493434100945533535657851259186926454950674578921152463993216374151;
            6'd57: xpb[183] = 1024'd87436015801934044634771889870820883667579873483826508596316845240082893806587892836406169670114725593475409791726427522211237881236342894205104605164514342969852210702011274299883630399111745674741948741547571048245643228163433839502488958931074222644510571982617759871917558759280189403529639899634091790682;
            6'd58: xpb[183] = 1024'd41084589674761934702512161571959539163794162549048288557324144078865195497566609271775899546389214905505692648352069135570392852863176149187413058757588578801933918950633107508164654402370223215196643502197190248740901202256481292735347913771425561921255707015460610454541662989681071211019437508649372722882;
            6'd59: xpb[183] = 1024'd118799859231714566169051360677912627404706878740005752646463297982624392525854464617160700637321378526979124912435204183508611665331229738724881637366993855567706301768826158054075917597145906476961535871234049295600520026570425518933185438295006350464820745462420519067272295294010586035627924944290248139413;
            6'd60: xpb[183] = 1024'd72448433104542456236791632379051282900921167805227532607470596821406694216833181052530430513595867839009407769060845796867766636958062993707190090960068091399788010017447991262356941600404384017416230631883668496095778000663472972166044393135357689741565880495263369649896399524411467843117722553305529071613;
            6'd61: xpb[183] = 1024'd26097006977370346304531904080189938397135456870449312568477895660188995907811897487900160389870357151039690625686487410226921608584896248689498544553142327231869718266069824470637965603662861557870925392533287696591035974756520425398903347975709029018311015528106220232520503754812349650607520162320810003813;
            6'd62: xpb[183] = 1024'd103812276534322977771071103186143026638048173061406776657617049563948192936099752833284961480802520772513122889769622458165140421052949838226967123162547603997642101084262875016549228798438544819635817761570146743450654799070464651596740872499289817561876053975066128845251136059141864475216007597961685420344;
            6'd63: xpb[183] = 1024'd57460850407150867838811374887281682134262462126628556618624348402730494627078469268654691357077010084543405746395264071524295392679783093209275576755621839829723809332884708224830252801697022360090512522219765943945912773163512104829599827339641156838621189007908979427875240289542746282705805206976966352544;
        endcase
    end

    always_comb begin
        case(flag[61][11:6])
            6'd0: xpb[184] = 1024'd0;
            6'd1: xpb[184] = 1024'd11109424279978757906551646588420337630476751191850336579631647241512796318057185704024421233351499396573688603020905684883450364306616348191584030348696075661805517581506541433111276804955499900545207282869385144441170747256559558062458782179992496115366324040751830010499344519943628090195602815992247284744;
            6'd2: xpb[184] = 1024'd22218848559957515813103293176840675260953502383700673159263294483025592636114371408048842466702998793147377206041811369766900728613232696383168060697392151323611035163013082866222553609910999801090414565738770288882341494513119116124917564359984992230732648081503660020998689039887256180391205631984494569488;
            6'd3: xpb[184] = 1024'd33328272839936273719654939765261012891430253575551009738894941724538388954171557112073263700054498189721065809062717054650351092919849044574752091046088226985416552744519624299333830414866499701635621848608155433323512241769678674187376346539977488346098972122255490031498033559830884270586808447976741854232;
            6'd4: xpb[184] = 1024'd44437697119915031626206586353681350521907004767401346318526588966051185272228742816097684933405997586294754412083622739533801457226465392766336121394784302647222070326026165732445107219821999602180829131477540577764682989026238232249835128719969984461465296163007320041997378079774512360782411263968989138976;
            6'd5: xpb[184] = 1024'd55547121399893789532758232942101688152383755959251682898158236207563981590285928520122106166757496982868443015104528424417251821533081740957920151743480378309027587907532707165556384024777499502726036414346925722205853736282797790312293910899962480576831620203759150052496722599718140450978014079961236423720;
            6'd6: xpb[184] = 1024'd66656545679872547439309879530522025782860507151102019477789883449076777908343114224146527400108996379442131618125434109300702185839698089149504182092176453970833105489039248598667660829732999403271243697216310866647024483539357348374752693079954976692197944244510980062996067119661768541173616895953483708464;
            6'd7: xpb[184] = 1024'd77765969959851305345861526118942363413337258342952356057421530690589574226400299928170948633460495776015820221146339794184152550146314437341088212440872529632638623070545790031778937634688499303816450980085696011088195230795916906437211475259947472807564268285262810073495411639605396631369219711945730993208;
            6'd8: xpb[184] = 1024'd88875394239830063252413172707362701043814009534802692637053177932102370544457485632195369866811995172589508824167245479067602914452930785532672242789568605294444140652052331464890214439643999204361658262955081155529365978052476464499670257439939968922930592326014640083994756159549024721564822527937978277952;
            6'd9: xpb[184] = 1024'd99984818519808821158964819295783038674290760726653029216684825173615166862514671336219791100163494569163197427188151163951053278759547133724256273138264680956249658233558872898001491244599499104906865545824466299970536725309036022562129039619932465038296916366766470094494100679492652811760425343930225562696;
            6'd10: xpb[184] = 1024'd111094242799787579065516465884203376304767511918503365796316472415127963180571857040244212333514993965736886030209056848834503643066163481915840303486960756618055175815065414331112768049554999005452072828693851444411707472565595580624587821799924961153663240407518300104993445199436280901956028159922472847440;
            6'd11: xpb[184] = 1024'd122203667079766336972068112472623713935244263110353702375948119656640759498629042744268633566866493362310574633229962533717954007372779830107424333835656832279860693396571955764224044854510498905997280111563236588852878219822155138687046603979917457269029564448270130115492789719379908992151630975914720132184;
            6'd12: xpb[184] = 1024'd9246395675620353479820831656229618821022587176468354827447911833176660479377089538277983585560318449441113828793374784022340530838175843743848239168021867007975536408507279859705082467948793085232289786045381886929688116857817923784526816476680504117575985074904902095885606165394904065228543965281372932597;
            6'd13: xpb[184] = 1024'd20355819955599111386372478244649956451499338368318691407079559074689456797434275242302404818911817846014802431814280468905790895144792191935432269516717942669781053990013821292816359272904292985777497068914767031370858864114377481846985598656673000232942309115656732106384950685338532155424146781273620217341;
            6'd14: xpb[184] = 1024'd31465244235577869292924124833070294081976089560169027986711206316202253115491460946326826052263317242588491034835186153789241259451408540127016299865414018331586571571520362725927636077859792886322704351784152175812029611370937039909444380836665496348308633156408562116884295205282160245619749597265867502085;
            6'd15: xpb[184] = 1024'd42574668515556627199475771421490631712452840752019364566342853557715049433548646650351247285614816639162179637856091838672691623758024888318600330214110093993392089153026904159038912882815292786867911634653537320253200358627496597971903163016657992463674957197160392127383639725225788335815352413258114786829;
            6'd16: xpb[184] = 1024'd53684092795535385106027418009910969342929591943869701145974500799227845751605832354375668518966316035735868240876997523556141988064641236510184360562806169655197606734533445592150189687770792687413118917522922464694371105884056156034361945196650488579041281237912222137882984245169416426010955229250362071573;
            6'd17: xpb[184] = 1024'd64793517075514143012579064598331306973406343135720037725606148040740642069663018058400089752317815432309556843897903208439592352371257584701768390911502245317003124316039987025261466492726292587958326200392307609135541853140615714096820727376642984694407605278664052148382328765113044516206558045242609356317;
            6'd18: xpb[184] = 1024'd75902941355492900919130711186751644603883094327570374305237795282253438387720203762424510985669314828883245446918808893323042716677873932893352421260198320978808641897546528458372743297681792488503533483261692753576712600397175272159279509556635480809773929319415882158881673285056672606402160861234856641061;
            6'd19: xpb[184] = 1024'd87012365635471658825682357775171982234359845519420710884869442523766234705777389466448932219020814225456934049939714578206493080984490281084936451608894396640614159479053069891484020102637292389048740766131077898017883347653734830221738291736627976925140253360167712169381017805000300696597763677227103925805;
            6'd20: xpb[184] = 1024'd98121789915450416732234004363592319864836596711271047464501089765279031023834575170473353452372313622030622652960620263089943445291106629276520481957590472302419677060559611324595296907592792289593948049000463042459054094910294388284197073916620473040506577400919542179880362324943928786793366493219351210549;
            6'd21: xpb[184] = 1024'd109231214195429174638785650952012657495313347903121384044132737006791827341891760874497774685723813018604311255981525947973393809597722977468104512306286547964225194642066152757706573712548292190139155331869848186900224842166853946346655856096612969155872901441671372190379706844887556876988969309211598495293;
            6'd22: xpb[184] = 1024'd120340638475407932545337297540432995125790099094971720623764384248304623659948946578522195919075312415177999859002431632856844173904339325659688542654982623626030712223572694190817850517503792090684362614739233331341395589423413504409114638276605465271239225482423202200879051364831184967184572125203845780037;
            6'd23: xpb[184] = 1024'd7383367071261949053090016724038900011568423161086373075264176424840524640696993372531545937769137502308539054565843883161230697369735339296112447987347658354145555235508018286298888130942086269919372289221378629418205486459076289506594850773368512119785646109057974181271867810846180040261485114570498580450;
            6'd24: xpb[184] = 1024'd18492791351240706959641663312459237642045174352936709654895823666353320958754179076555967171120636898882227657586749568044681061676351687487696478336043734015951072817014559719410164935897586170464579572090763773859376233715635847569053632953361008235151970149809804191771212330789808130457087930562745865194;
            6'd25: xpb[184] = 1024'd29602215631219464866193309900879575272521925544787046234527470907866117276811364780580388404472136295455916260607655252928131425982968035679280508684739809677756590398521101152521441740853086071009786854960148918300546980972195405631512415133353504350518294190561634202270556850733436220652690746554993149938;
            6'd26: xpb[184] = 1024'd40711639911198222772744956489299912902998676736637382814159118149378913594868550484604809637823635692029604863628560937811581790289584383870864539033435885339562107980027642585632718545808585971554994137829534062741717728228754963693971197313346000465884618231313464212769901370677064310848293562547240434682;
            6'd27: xpb[184] = 1024'd51821064191176980679296603077720250533475427928487719393790765390891709912925736188629230871175135088603293466649466622695032154596200732062448569382131961001367625561534184018743995350764085872100201420698919207182888475485314521756429979493338496581250942272065294223269245890620692401043896378539487719426;
            6'd28: xpb[184] = 1024'd62930488471155738585848249666140588163952179120338055973422412632404506230982921892653652104526634485176982069670372307578482518902817080254032599730828036663173143143040725451855272155719585772645408703568304351624059222741874079818888761673330992696617266312817124233768590410564320491239499194531735004170;
            6'd29: xpb[184] = 1024'd74039912751134496492399896254560925794428930312188392553054059873917302549040107596678073337878133881750670672691277992461932883209433428445616630079524112324978660724547266884966548960675085673190615986437689496065229969998433637881347543853323488811983590353568954244267934930507948581435102010523982288914;
            6'd30: xpb[184] = 1024'd85149337031113254398951542842981263424905681504038729132685707115430098867097293300702494571229633278324359275712183677345383247516049776637200660428220187986784178306053808318077825765630585573735823269307074640506400717254993195943806326033315984927349914394320784254767279450451576671630704826516229573658;
            6'd31: xpb[184] = 1024'd96258761311092012305503189431401601055382432695889065712317354356942895185154479004726915804581132674898047878733089362228833611822666124828784690776916263648589695887560349751189102570586085474281030552176459784947571464511552754006265108213308481042716238435072614265266623970395204761826307642508476858402;
            6'd32: xpb[184] = 1024'd107368185591070770212054836019821938685859183887739402291949001598455691503211664708751337037932632071471736481753995047112283976129282473020368721125612339310395213469066891184300379375541585374826237835045844929388742211768112312068723890393300977158082562475824444275765968490338832852021910458500724143146;
            6'd33: xpb[184] = 1024'd118477609871049528118606482608242276316335935079589738871580648839968487821268850412775758271284131468045425084774900731995734340435898821211952751474308414972200731050573432617411656180497085275371445117915230073829912959024671870131182672573293473273448886516576274286265313010282460942217513274492971427890;
            6'd34: xpb[184] = 1024'd5520338466903544626359201791848181202114259145704391323080441016504388802016897206785108289977956555175964280338312982300120863901294834848376656806673449700315574062508756712892693793935379454606454792397375371906722856060334655228662885070056520121995307143211046266658129456297456015294426263859624228303;
            6'd35: xpb[184] = 1024'd16629762746882302532910848380268518832591010337554727902712088258017185120074082910809529523329455951749652883359218667183571228207911183039960687155369525362121091644015298146003970598890879355151662075266760516347893603316894213291121667250049016237361631183962876277157473976241084105490029079851871513047;
            6'd36: xpb[184] = 1024'd27739187026861060439462494968688856463067761529405064482343735499529981438131268614833950756680955348323341486380124352067021592514527531231544717504065601023926609225521839579115247403846379255696869358136145660789064350573453771353580449430041512352727955224714706287656818496184712195685631895844118797791;
            6'd37: xpb[184] = 1024'd38848611306839818346014141557109194093544512721255401061975382741042777756188454318858371990032454744897030089401030036950471956821143879423128747852761676685732126807028381012226524208801879156242076641005530805230235097830013329416039231610034008468094279265466536298156163016128340285881234711836366082535;
            6'd38: xpb[184] = 1024'd49958035586818576252565788145529531724021263913105737641607029982555574074245640022882793223383954141470718692421935721833922321127760227614712778201457752347537644388534922445337801013757379056787283923874915949671405845086572887478498013790026504583460603306218366308655507536071968376076837527828613367279;
            6'd39: xpb[184] = 1024'd61067459866797334159117434733949869354498015104956074221238677224068370392302825726907214456735453538044407295442841406717372685434376575806296808550153828009343161970041463878449077818712878957332491206744301094112576592343132445540956795970019000698826927346970196319154852056015596466272440343820860652023;
            6'd40: xpb[184] = 1024'd72176884146776092065669081322370206984974766296806410800870324465581166710360011430931635690086952934618095898463747091600823049740992923997880838898849903671148679551548005311560354623668378857877698489613686238553747339599692003603415578150011496814193251387722026329654196575959224556468043159813107936767;
            6'd41: xpb[184] = 1024'd83286308426754849972220727910790544615451517488656747380501971707093963028417197134956056923438452331191784501484652776484273414047609272189464869247545979332954197133054546744671631428623878758422905772483071382994918086856251561665874360330003992929559575428473856340153541095902852646663645975805355221511;
            6'd42: xpb[184] = 1024'd94395732706733607878772374499210882245928268680507083960133618948606759346474382838980478156789951727765473104505558461367723778354225620381048899596242054994759714714561088177782908233579378658968113055352456527436088834112811119728333142509996489044925899469225686350652885615846480736859248791797602506255;
            6'd43: xpb[184] = 1024'd105505156986712365785324021087631219876405019872357420539765266190119555664531568543004899390141451124339161707526464146251174142660841968572632929944938130656565232296067629610894185038534878559513320338221841671877259581369370677790791924689988985160292223509977516361152230135790108827054851607789849790999;
            6'd44: xpb[184] = 1024'd116614581266691123691875667676051557506881771064207757119396913431632351982588754247029320623492950520912850310547369831134624506967458316764216960293634206318370749877574171044005461843490378460058527621091226816318430328625930235853250706869981481275658547550729346371651574655733736917250454423782097075743;
            6'd45: xpb[184] = 1024'd3657309862545140199628386859657462392660095130322409570896705608168252963336801041038670642186775608043389506110782081439011030432854330400640865625999241046485592889509495139486499456928672639293537295573372114395240225661593020950730919366744528124204968177364118352044391101748731990327367413148749876156;
            6'd46: xpb[184] = 1024'd14766734142523898106180033448077800023136846322172746150528352849681049281393986745063091875538275004617078109131687766322461394739470678592224895974695316708291110471016036572597776261884172539838744578442757258836410972918152579013189701546737024239571292218115948362543735621692360080522970229140997160900;
            6'd47: xpb[184] = 1024'd25876158422502656012731680036498137653613597514023082730160000091193845599451172449087513108889774401190766712152593451205911759046087026783808926323391392370096628052522578005709053066839672440383951861312142403277581720174712137075648483726729520354937616258867778373043080141635988170718573045133244445644;
            6'd48: xpb[184] = 1024'd36985582702481413919283326624918475284090348705873419309791647332706641917508358153111934342241273797764455315173499136089362123352703374975392956672087468031902145634029119438820329871795172340929159144181527547718752467431271695138107265906722016470303940299619608383542424661579616260914175861125491730388;
            6'd49: xpb[184] = 1024'd48095006982460171825834973213338812914567099897723755889423294574219438235565543857136355575592773194338143918194404820972812487659319723166976987020783543693707663215535660871931606676750672241474366427050912692159923214687831253200566048086714512585670264340371438394041769181523244351109778677117739015132;
            6'd50: xpb[184] = 1024'd59204431262438929732386619801759150545043851089574092469054941815732234553622729561160776808944272590911832521215310505856262851965936071358561017369479619355513180797042202305042883481706172142019573709920297836601093961944390811263024830266707008701036588381123268404541113701466872441305381493109986299876;
            6'd51: xpb[184] = 1024'd70313855542417687638938266390179488175520602281424429048686589057245030871679915265185198042295771987485521124236216190739713216272552419550145047718175695017318698378548743738154160286661672042564780992789682981042264709200950369325483612446699504816402912421875098415040458221410500531500984309102233584620;
            6'd52: xpb[184] = 1024'd81423279822396445545489912978599825805997353473274765628318236298757827189737100969209619275647271384059209727257121875623163580579168767741729078066871770679124215960055285171265437091617171943109988275659068125483435456457509927387942394626692000931769236462626928425539802741354128621696587125094480869364;
            6'd53: xpb[184] = 1024'd92532704102375203452041559567020163436474104665125102207949883540270623507794286673234040508998770780632898330278027560506613944885785115933313108415567846340929733541561826604376713896572671843655195558528453269924606203714069485450401176806684497047135560503378758436039147261297756711892189941086728154108;
            6'd54: xpb[184] = 1024'd103642128382353961358593206155440501066950855856975438787581530781783419825851472377258461742350270177206586933298933245390064309192401464124897138764263922002735251123068368037487990701528171744200402841397838414365776950970629043512859958986676993162501884544130588446538491781241384802087792757078975438852;
            6'd55: xpb[184] = 1024'd114751552662332719265144852743860838697427607048825775367213178023296216143908658081282882975701769573780275536319838930273514673499017812316481169112959997664540768704574909470599267506483671644745610124267223558806947698227188601575318741166669489277868208584882418457037836301185012892283395573071222723596;
            6'd56: xpb[184] = 1024'd1794281258186735772897571927466743583205931114940427818712970199832117124656704875292232994395594660910814731883251180577901196964413825952905074445325032392655611716510233566080305119921965823980619798749368856883757595262851386672798953663432536126414629211517190437430652747200007965360308562437875524009;
            6'd57: xpb[184] = 1024'd12903705538165493679449218515887081213682682306790764398344617441344913442713890579316654227747094057484503334904156865461351561271030174144489104794021108054461129298016774999191581924877465724525827081618754001324928342519410944735257735843425032241780953252269020447929997267143636055555911378430122808753;
            6'd58: xpb[184] = 1024'd24013129818144251586000865104307418844159433498641100977976264682857709760771076283341075461098593454058191937925062550344801925577646522336073135142717183716266646879523316432302858729832965625071034364488139145766099089775970502797716518023417528357147277293020850458429341787087264145751514194422370093497;
            6'd59: xpb[184] = 1024'd35122554098123009492552511692727756474636184690491437557607911924370506078828261987365496694450092850631880540945968235228252289884262870527657165491413259378072164461029857865414135534788465525616241647357524290207269837032530060860175300203410024472513601333772680468928686307030892235947117010414617378241;
            6'd60: xpb[184] = 1024'd46231978378101767399104158281148094105112935882341774137239559165883302396885447691389917927801592247205569143966873920111702654190879218719241195840109335039877682042536399298525412339743965426161448930226909434648440584289089618922634082383402520587879925374524510479428030826974520326142719826406864662985;
            6'd61: xpb[184] = 1024'd57341402658080525305655804869568431735589687074192110716871206407396098714942633395414339161153091643779257746987779604995153018497495566910825226188805410701683199624042940731636689144699465326706656213096294579089611331545649176985092864563395016703246249415276340489927375346918148416338322642399111947729;
            6'd62: xpb[184] = 1024'd68450826938059283212207451457988769366066438266042447296502853648908895032999819099438760394504591040352946350008685289878603382804111915102409256537501486363488717205549482164747965949654965227251863495965679723530782078802208735047551646743387512818612573456028170500426719866861776506533925458391359232473;
            6'd63: xpb[184] = 1024'd79560251218038041118759098046409106996543189457892783876134500890421691351057004803463181627856090436926634953029590974762053747110728263293993286886197562025294234787056023597859242754610465127797070778835064867971952826058768293110010428923380008933978897496780000510926064386805404596729528274383606517217;
        endcase
    end

    always_comb begin
        case(flag[61][16:12])
            5'd0: xpb[185] = 1024'd0;
            5'd1: xpb[185] = 1024'd90669675498016799025310744634829444627019940649743120455766148131934487669114190507487602861207589833500323556050496659645504111417344611485577317234893637687099752368562565030970519559565965028342278061704450012413123573315327851172469211103372505049345221537531830521425408906749032686925131090375853801961;
            5'd2: xpb[185] = 1024'd57272655311908856651822561864844456509341454173750556783400441198892080000919242104960134507757505357557497704643499884711944381993468888415994509453456234440508830167553912724310799927614724335374358515021660178461886296409758929379959852523515560831870539660946603012744289739569432356731572354126113119591;
            5'd3: xpb[185] = 1024'd23875635125800914278334379094859468391662967697757993111034734265849672332724293702432666154307420881614671853236503109778384652569593165346411701672018831193917907966545260417651080295663483642406438968338870344510649019504190007587450493943658616614395857784361375504063170572389832026538013617876372437221;
            5'd4: xpb[185] = 1024'd114545310623817713303645123729688913018682908347501113566800882397784160001838484209920269015515010715114995409286999769423888763986937776831989018906912468881017660335107825448621599855229448670748717030043320356923772592819517858759919705047031121663741079321893206025488579479138864713463144708252226239182;
            5'd5: xpb[185] = 1024'd81148290437709770930156940959703924901004421871508549894435175464741752333643535807392800662064926239172169557880002994490329034563062053762406211125475065634426738134099173141961880223278207977780797483360530522972535315913948936967410346467174177446266397445307978516807460311959264383269585972002485556812;
            5'd6: xpb[185] = 1024'd47751270251601828556668758189718936783325935395515986222069468531699344665448587404865332308614841763229343706473006219556769305139186330692823403344037662387835815933090520835302160591326967284812877936677740689021298039008380015174900987887317233228791715568722751008126341144779664053076027235752744874442;
            5'd7: xpb[185] = 1024'd14354250065493886183180575419733948665647448919523422549703761598656936997253639002337863955164757287286517855066009444623209575715310607623240595562600259141244893732081868528642440959375726591844958389994950855070060762102811093382391629307460289011317033692137523499445221977600063722882468499503004192072;
            5'd8: xpb[185] = 1024'd105023925563510685208491320054563393292667389569266543005469909730591424666367829509825466816372347120786841411116506104268713687132655219108817912797493896828344646100644433559612960518941691620187236451699400867483184335418138944554860840410832794060662255229669354020870630884349096409807599589878857994033;
            5'd9: xpb[185] = 1024'd71626905377402742835003137284578405174988903093273979333104202797549016998172881107297998462922262644844015559709509329335153957708779496039235105016056493581753723899635781252953240886990450927219316905016611033531947058512570022762351481830975849843187573353084126512189511717169496079614040853629117311663;
            5'd10: xpb[185] = 1024'd38229885191294800461514954514593417057310416617281415660738495864506609329977932704770530109472178168901189708302512554401594228284903772969652297234619090335162801698627128946293521255039210234251397358333821199580709781607001100969842123251118905625712891476498899003508392549989895749420482117379376629293;
            5'd11: xpb[185] = 1024'd4832865005186858088026771744608428939631930141288851988372788931464201661782984302243061756022093692958363856895515779468034498861028049900069489453181687088571879497618476639633801623087969541283477811651031365629472504701432179177332764671261961408238209599913671494827273382810295419226923381129635946923;
            5'd12: xpb[185] = 1024'd95502540503203657113337516379437873566651870791031972444138937063398689330897174809730664617229683526458687412946012439113538610278372661385646806688075324775671631866181041670604321182653934569625755873355481378042596078016760030349801975774634466457583431137445502016252682289559328106152054471505489748884;
            5'd13: xpb[185] = 1024'd62105520317095714739849333609452885448973384315039408771773230130356281662702226407203196263779599050515861561539015664179978880854496938316063998906637921529080709665172389363944601550702693876657836326672691544091358801111191108557292617194777522240108749260860274507571563122379727775958495735255749066514;
            5'd14: xpb[185] = 1024'd28708500130987772366361150839467897331294897839046845099407523197313873994507278004675727910329514574573035710132018889246419151430621215246481191125200518282489787464163737057284881918751453183689916779989901710140121524205622186764783258614920578022634067384275046998890443955200127445764936999006008384144;
            5'd15: xpb[185] = 1024'd119378175629004571391671895474297341958314838488789965555173671329248361663621468512163330771537104408073359266182515548891923262847965826732058508360094155969589539832726302088255401478317418212032194841694351722553245097520950037937252469718293083071979288921806877520315852861949160132690068089381862186105;
            5'd16: xpb[185] = 1024'd85981155442896629018183712704312353840636352012797401882807964396205953995426520109635862418087019932130533414775518773958363533424090103662475700578656752722998617631717649781595681846366177519064275295011561888602007820615381116144743111138436138854504607045221650011634733694769559802496509353132121503735;
            5'd17: xpb[185] = 1024'd52584135256788686644695529934327365722957865536804838210442257463163546327231571707108394064636935456187707563368521999024803804000214380592892892797219349476407695430708997474935962214414936826096355748328772054650770543709812194352233752558579194637029925168636422502953614527589959472302950616882380821365;
            5'd18: xpb[185] = 1024'd19187115070680744271207347164342377605279379060812274538076550530121138659036623304580925711186850980244881711961525224091244074576338657523310085015781946229816773229700345168276242582463696133128436201645982220699533266804243272559724393978722250419555243292051194994272495360410359142109391880632640138995;
            5'd19: xpb[185] = 1024'd109856790568697543296518091799171822232299319710555394993842698662055626328150813812068528572394440813745205268012021883736748185993683269008887402250675583916916525598262910199246762142029661161470714263350432233112656840119571123732193605082094755468900464829583025515697904267159391829034522971008493940956;
            5'd20: xpb[185] = 1024'd76459770382589600923029909029186834114620833234562831321476991729013218659955865409541060218944356337802379416605025108803188456569807545939304594469238180670325603397254257892587042510078420468502794716667642399161419563214002201939684246502237811251425782952997798007016785099979791498840964234758753258586;
            5'd21: xpb[185] = 1024'd43062750196481658549541726259201845996942346758570267649111284795970810991760917007013591865494271861859553565198028333869628727145931822869721786687800777423734681196245605585927322878127179775534875169984852565210182286308433280147174887922380867033951101076412570498335665932800191168647405498509012576216;
            5'd22: xpb[185] = 1024'd9665730010373716176053543489216857879263860282577703976745577862928403323565968604486123512044187385916727713791031558936068997722056099800138978906363374177143758995236953279267603246175939082566955623302062731258945009402864358354665529342523922816476419199827342989654546765620590838453846762259271893846;
            5'd23: xpb[185] = 1024'd100335405508390515201364288124046302506283800932320824432511725994862890992680159111973726373251777219417051269841528218581573109139400711285716296141257011864243511363799518310238122805741904110909233685006512743672068582718192209527134740445896427865821640737359173511079955672369623525378977852635125695807;
            5'd24: xpb[185] = 1024'd66938385322282572827876105354061314388605314456328260760146019061820483324485210709446258019801692743474225418434531443648013379715524988216133488359819608617652589162790866003578403173790663417941314138323722909720831305812623287734625381866039483648346958860773946002398836505190023195185419116385385013437;
            5'd25: xpb[185] = 1024'd33541365136174630454387922584076326270926827980335697087780312128778075656290262306918789666351608267531399567027534668714453650291649265146550680578382205371061666961782213696918683541839422724973394591640933075769594028907054365942116023286182539430872276984188718493717717338010422864991860380135644331067;
            5'd26: xpb[185] = 1024'd144344950066688080899739814091338153248341504343133415414605195735667988095313904391321312901523791588573715620537893780893920867773542076967872796944802124470744760773561390258963909888182032005475044958143241818356752001485444149606664706325595213397595107603490985036598170830822534798301643885903648697;
            5'd27: xpb[185] = 1024'd90814020448083487106210484448920782780268282154086253871180753327670155657209504411878924174109113625088897271671034553426398032285118153562545190031838439811570497129336126421229483469454147060347753106662593254231480325316813295322075875809698100262742816645135321506462007077579855221723432734261757450658;
            5'd28: xpb[185] = 1024'd57417000261975544732722301678935794662589795678093690198815046394627747989014556009351455820659029149146071420264037778492838302861242430492962382250401036564979574928327474114569763837502906367379833559979803420280243048411244373529566517229841156045268134768550093997780887910400254891529873998012016768288;
            5'd29: xpb[185] = 1024'd24019980075867602359234118908950806544911309202101126526449339461585340320819607606823987467208944673203245568857041003559278573437366707423379574468963633318388652727318821807910044205551665674411914013297013586329005771505675451737057158649984211827793452891964866489099768743220654561336315261762276085918;
            5'd30: xpb[185] = 1024'd114689655573884401384544863543780251171931249851844246982215487593519827989933798114311590328416534506703569124907537663204782684854711318908956891703857271005488405095881386838880563765117630702754192075001463598742129344821003302909526369753356716877138674429496697010525177649969687248261446352138129887879;
            5'd31: xpb[185] = 1024'd81292635387776459011056680773795263054252763375851683309849780660477420321738849711784121974966450030760743273500540888271222955430835595839374083922419867758897482894872734532220844133166390009786272528318673764790892067915434381117017011173499772659663992552911469501844058482790086918067887615888389205509;
        endcase
    end

    always_comb begin
        case(flag[62][5:0])
            6'd0: xpb[186] = 1024'd0;
            6'd1: xpb[186] = 1024'd85981155442896629018183712704312353840636352012797401882807964396205953995426520109635862418087019932130533414775518773958363533424090103662475700578656752722998617631717649781595681846366177519064275295011561888602007820615381116144743111138436138854504607045221650011634733694769559802496509353132121503735;
            6'd2: xpb[186] = 1024'd47895615201668516637568498003810274936574276899859119637484073727435012653543901309256653621516365554817917422093544113337663226006959872769791276140982464512306560693864082225561124501215149316818352981635883930839654791009865459324507652593642828442189310676326241993162939315610486587874328879638648523139;
            6'd3: xpb[186] = 1024'd9810074960440404256953283303308196032512201786920837392160183058664071311661282508877444824945711177505301429411569452716962918589829641877106851703308176301614503756010514669526567156064121114572430668260205973077301761404349802504272194048849518029874014307430833974691144936451413373252148406145175542543;
            6'd4: xpb[186] = 1024'd95791230403337033275136996007620549873148553799718239274968147454870025307087802618513307243032731109635834844187088226675326452013919745539582552281964929024613121387728164451122249002430298633636705963271767861679309582019730918649015305187285656884378621352652483986325878631220973175748657759277297046278;
            6'd5: xpb[186] = 1024'd57705690162108920894521781307118470969086478686779957029644256786099083965205183818134098446462076732323218851505113566054626144596789514646898127844290640813921064449874596895087691657279270431390783649896089903916956552414215261828779846642492346472063324983757075967854084252061899961126477285783824065682;
            6'd6: xpb[186] = 1024'd19620149920880808513906566606616392065024403573841674784320366117328142623322565017754889649891422355010602858823138905433925837179659283754213703406616352603229007512021029339053134312128242229144861336520411946154603522808699605008544388097699036059748028614861667949382289872902826746504296812290351085086;
            6'd7: xpb[186] = 1024'd105601305363777437532090279310928745905660755586639076667128330513534096618749085127390752067978442287141136273598657679392289370603749387416689403985273105326227625143738679120648816158494419748209136631531973834756611343424080721153287499236135174914252635660083317961017023567672386549000806165422472588821;
            6'd8: xpb[186] = 1024'd67515765122549325151475064610426667001598680473700794421804439844763155276866466327011543271407787909828520280916683018771589063186619156524004979547598817115535568205885111564614258813343391545963214318156295876994258313818565064333052040691341864501937339291187909942545229188513313334378625691928999608225;
            6'd9: xpb[186] = 1024'd29430224881321212770859849909924588097536605360762512176480549175992213934983847526632334474837133532515904288234708358150888755769488925631320555109924528904843511268031544008579701468192363343717292004780617919231905284213049407512816582146548554089622042922292501924073434809354240119756445218435526627629;
            6'd10: xpb[186] = 1024'd115411380324217841789043562614236941938172957373559914059288513572198167930410367636268196892924153464646437703010227132109252289193579029293796255688581281627842128899749193790175383314558540862781567299792179807833913104828430523657559693284984692944126649967514151935708168504123799922252954571567648131364;
            6'd11: xpb[186] = 1024'd77325840082989729408428347913734863034110882260621631813964622903427226588527748835888988096353499087333821710328252471488551981776448798401111831250906993417150071961895626234140825969407512660535644986416501850071560075222914866837324234740191382531811353598618743917236374124964726707630774098074175150768;
            6'd12: xpb[186] = 1024'd39240299841761617027813133213232784130048807147683349568640732234656285246645130035509779299782844710021205717646277810867851674359318567508427406813232705206458015024042058678106268624256484458289722673040823892309207045617399210017088776195398072119496057229723335898764579745805653493008593624580702170172;
            6'd13: xpb[186] = 1024'd1154759600533504647197918512730705225986732034745067323316841565885343904762511235130570503212190332708589724964303150247151366942188336615742982375558416995765958086188491122071711279105456256043800359665145934546854016011883553196853317650604761707180760860827927880292785366646580278386413151087229189576;
            6'd14: xpb[186] = 1024'd87135915043430133665381631217043059066623084047542469206124805962091297900189031344766432921299210264839123139739821924205514900366278440278218682954215169718764575717906140903667393125471633775108075654676707823148861836627264669341596428789040900561685367906049577891927519061416140080882922504219350693311;
            6'd15: xpb[186] = 1024'd49050374802202021284766416516540980162561008934604186960800915293320356558306412544387224124728555887526507147057847263584814592949148209385534258516540881508072518780052573347632835780320605572862153341301029865386508807021749012521360970244247590149370071537154169873455724682257066866260742030725877712715;
            6'd16: xpb[186] = 1024'd10964834560973908904151201816038901258498933821665904715477024624549415216423793744008015328157901510213891154375872602964114285532017978492849834078866593297380461842199005791598278435169577370616231027925351907624155777416233355701125511699454279737054775168258761854983930303097993651638561557232404732119;
            6'd17: xpb[186] = 1024'd96945990003870537922334914520351255099135285834463306598284989020755369211850313853643877746244921442344424569151391376922477818956108082155325534657523346020379079473916655573193960281535754889680506322936913796226163598031614471845868622837890418591559382213480411866618663997867553454135070910364526235854;
            6'd18: xpb[186] = 1024'd58860449762642425541719699819849176195073210721525024352961098351984427869967695053264668949674267065031808576469416716301777511538977851262641110219849057809687022536063088017159402936384726687434584009561235838463810568426098815025633164293097108179244085844585003848146869618708480239512890436871053255258;
            6'd19: xpb[186] = 1024'd20774909521414313161104485119347097291011135608586742107637207683213486528085076252885460153103612687719192583787442055681077204121847620369956685782174769598994965598209520461124845591233698485188661696185557880701457538820583158205397705748303797766928789475689595829675075239549407024890709963377580274662;
            6'd20: xpb[186] = 1024'd106756064964310942179288197823659451131647487621384143990445172079419440523511596362521322571190632619849725998562960829639440737545937724032432386360831522321993583229927170242720527437599876004252936991197119769303465359435964274350140816886739936621433396520911245841309808934318966827387219316509701778397;
            6'd21: xpb[186] = 1024'd68670524723082829798672983123157372227585412508445861745121281410648499181628977562142113774619978242537110005880986169018740430128807493139747961923157234111301526292073602686685970092448847802007014677821441811541112329830448617529905358341946626209118100152015837822838014555159893612765038843016228797801;
            6'd22: xpb[186] = 1024'd30584984481854717418057768422655293323523337395507579499797390741877557839746358761762904978049323865224494013199011508398040122711677262247063537485482945900609469354220035130651412747297819599761092364445763853778759300224932960709669899797153315796802803783120429804366220176000820398142858369522755817205;
            6'd23: xpb[186] = 1024'd116566139924751346436241481126967647164159689408304981382605355138083511835172878871398767396136343797355027427974530282356403656135767365909539238064139698623608086985937684912247094593663997118825367659457325742380767120840314076854413010935589454651307410828342079816000953870770380200639367722654877320940;
            6'd24: xpb[186] = 1024'd78480599683523234055626266426465568260097614295366699137281464469312570493290260071019558599565689420042411435292555621735703348718637135016854813626465410412916030048084117356212537248512968916579445346081647784618414091234798420034177552390796144238992114459446671797529159491611306986017187249161404340344;
            6'd25: xpb[186] = 1024'd40395059442295121675011051725963489356035539182428416891957573800541629151407641270640349802995035042729795442610580961115003041301506904124170389188791122202223973110230549800177979903361940714333523032705969826856061061629282763213942093846002833826676818090551263779057365112452233771395006775667931359748;
            6'd26: xpb[186] = 1024'd2309519201067009294395837025461410451973464069490134646633683131770687809525022470261141006424380665417179449928606300494302733884376673231485964751116833991531916172376982244143422558210912512087600719330291869093708032023767106393706635301209523414361521721655855760585570733293160556772826302174458379152;
            6'd27: xpb[186] = 1024'd88290674643963638312579549729773764292609816082287536529441647527976641804951542579897003424511400597547712864704125074452666267308466776893961665329773586714530533804094632025739104404577090031151876014341853757695715852639148222538449746439645662268866128766877505772220304428062720359269335655306579882887;
            6'd28: xpb[186] = 1024'd50205134402735525931964335029271685388547740969349254284117756859205700463068923779517794627940746220235096872022150413831965959891336546001277240892099298503838476866241064469704547059426061828905953700966175799933362823033632565718214287894852351856550832397982097753748510048903647144647155181813106902291;
            6'd29: xpb[186] = 1024'd12119594161507413551349120328769606484485665856410972038793866190434759121186304979138585831370091842922480879340175753211265652474206315108592816454425010293146419928387496913669989714275033626660031387590497842171009793428116908897978829350059041444235536029086689735276715669744573930024974708319633921695;
            6'd30: xpb[186] = 1024'd98100749604404042569532833033081960325122017869208373921601830586640713116612825088774448249457111775053014294115694527169629185898296418771068517033081763016145037560105146695265671560641211145724306682602059730773017614043498025042721940488495180298740143074308339746911449364514133732521484061451755425430;
            6'd31: xpb[186] = 1024'd60015209363175930188917618332579881421059942756270091676277939917869771774730206288395239452886457397740398301433719866548928878481166187878384092595407474805452980622251579139231114215490182943478384369226381773010664584437982368222486481943701869886424846705412931728439654985355060517899303587958282444834;
            6'd32: xpb[186] = 1024'd21929669121947817808302403632077802516997867643331809430954049249098830432847587488016030656315803020427782308751745205928228571064035956985699668157733186594760923684398011583196556870339154741232462055850703815248311554832466711402251023398908559474109550336517523709967860606195987303277123114464809464238;
            6'd33: xpb[186] = 1024'd107910824564844446826486116336390156357634219656129211313762013645304784428274107597651893074402822952558315723527263979886592104488126060648175368736389939317759541316115661364792238716705332260296737350862265703850319375447847827546994134537344698328614157381739173721602594300965547105773632467596930967973;
            6'd34: xpb[186] = 1024'd69825284323616334445870901635888077453572144543190929068438122976533843086391488797272684277832168575245699730845289319265891797070995829755490944298715651107067484378262093808757681371554304058050815037486587746087966345842332170726758675992551387916298861012843765703130799921806473891151451994103457987377;
            6'd35: xpb[186] = 1024'd31739744082388222065255686935385998549510069430252646823114232307762901744508869996893475481261514197933083738163314658645191489653865598862806519861041362896375427440408526252723124026403275855804892724110909788325613316236816513906523217447758077503983564643948357684659005542647400676529271520609985006781;
            6'd36: xpb[186] = 1024'd117720899525284851083439399639698352390146421443050048705922196703968855739935390106529337899348534130063617152938833432603555023077955702525282220439698115619374045072126176034318805872769453374869168019122471676927621136852197630051266328586194216358488171689170007696293739237416960479025780873742106510516;
            6'd37: xpb[186] = 1024'd79635359284056738702824184939196273486084346330111766460598306035197914398052771306150129102777879752751001160256858771982854715660825471632597796002023827408681988134272608478284248527618425172623245705746793719165268107246681973231030870041400905946172875320274599677821944858257887264403600400248633529920;
            6'd38: xpb[186] = 1024'd41549819042828626322208970238694194582022271217173484215274415366426973056170152505770920306207225375438385167574884111362154408243695240739913371564349539197989931196419040922249691182467396970377323392371115761402915077641166316410795411496607595533857578951379191659350150479098814049781419926755160549324;
            6'd39: xpb[186] = 1024'd3464278801600513941593755538192115677960196104235201969950524697656031714287533705391711509636570998125769174892909450741454100826565009847228947126675250987297874258565473366215133837316368768131401078995437803640562048035650659590559952951814285121542282582483783640878356099939740835159239453261687568728;
            6'd40: xpb[186] = 1024'd89445434244497142959777468242504469518596548117032603852758489093861985709714053815027573927723590930256302589668428224699817634250655113509704647705332003710296491890283123147810815683682546287195676374006999692242569868651031775735303064090250423976046889627705433652513089794709300637655748806393809072463;
            6'd41: xpb[186] = 1024'd51359894003269030579162253542002390614534473004094321607434598425091044367831435014648365131152936552943686596986453564079117326833524882617020223267657715499604434952429555591776258338531518084949754060631321734480216839045516118915067605545457113563731593258810025634041295415550227423033568332900336091867;
            6'd42: xpb[186] = 1024'd13274353762040918198547038841500311710472397891156039362110707756320103025948816214269156334582282175631070604304478903458417019416394651724335798829983427288912378014575988035741700993380489882703831747255643776717863809440000462094832147000663803151416296889914617615569501036391154208411387859406863111271;
            6'd43: xpb[186] = 1024'd99255509204937547216730751545812665551108749903953441244918672152526057021375336323905018752669302107761604019079997677416780552840484755386811499408640180011910995646293637817337382839746667401768107042267205665319871630055381578239575258139099942005920903935136267627204234731160714010907897212538984615006;
            6'd44: xpb[186] = 1024'd61169968963709434836115536845310586647046674791015158999594781483755115679492717523525809956098647730448988026398023016796080245423354524494127074970965891801218938708440070261302825494595639199522184728891527707557518600449865921419339799594306631593605607566240859608732440352001640796285716739045511634410;
            6'd45: xpb[186] = 1024'd23084428722481322455500322144808507742984599678076876754270890814984174337610098723146601159527993353136372033716048356175379938006224293601442650533291603590526881770586502705268268149444610997276262415515849749795165570844350264599104341049513321181290311197345451590260645972842567581663536265552038653814;
            6'd46: xpb[186] = 1024'd109065584165377951473684034849120861583620951690874278637078855211190128333036618832782463577615013285266905448491567130133743471430314397263918351111948356313525499402304152486863949995810788516340537710527411638397173391459731380743847452187949460035794918242567101601895379667612127384160045618684160157549;
            6'd47: xpb[186] = 1024'd70980043924149839093068820148618782679558876577935996391754964542419186991154000032403254781044358907954289455809592469513043164013184166371233926674274068102833442464450584930829392650659760314094615397151733680634820361854215723923611993643156149623479621873671693583423585288453054169537865145190687176953;
            6'd48: xpb[186] = 1024'd32894503682921726712453605448116703775496801464997714146431073873648245649271381232024045984473704530641673463127617808892342856596053935478549502236599779892141385526597017374794835305508732111848693083776055722872467332248700067103376535098362839211164325504776285564951790909293980954915684671697214196357;
            6'd49: xpb[186] = 1024'd118875659125818355730637318152429057616133153477795116029239038269854199644697901341659908402560724462772206877903136582850706390020144039141025202815256532615140003158314667156390517151874909630912968378787617611474475152864081183248119646236798978065668932549997935576586524604063540757412194024829335700092;
            6'd50: xpb[186] = 1024'd80790118884590243350022103451926978712071078364856833783915147601083258302815282541280699605990070085459590885221161922230006082603013808248340778377582244404447946220461099600355959806723881428667046065411939653712122123258565526427884187692005667653353636181102527558114730224904467542790013551335862719496;
            6'd51: xpb[186] = 1024'd42704578643362130969406888751424899808009003251918551538591256932312316960932663740901490809419415708146974892539187261609305775185883577355656353939907956193755889282607532044321402461572853226421123752036261695949769093653049869607648729147212357241038339812207119539642935845745394328167833077842389738900;
            6'd52: xpb[186] = 1024'd4619038402134018588791674050922820903946928138980269293267366263541375619050044940522282012848761330834358899857212600988605467768753346462971929502233667983063832344753964488286845116421825024175201438660583738187416064047534212787413270602419046828723043443311711521171141466586321113545652604348916758304;
            6'd53: xpb[186] = 1024'd90600193845030647606975386755235174744583280151777671176075330659747329614476565050158144430935781262964892314632731374946969001192843450125447630080890420706062449976471614269882526962788002543239476733672145626789423884662915328932156381740855185683227650488533361532805875161355880916042161957481038262039;
            6'd54: xpb[186] = 1024'd52514653603802535226360172054733095840521205038839388930751439990976388272593946249778935634365126885652276321950756714326268693775713219232763205643216132495370393038618046713847969617636974340993554420296467669027070855057399672111920923196061875270912354119637953514334080782196807701419981483987565281443;
            6'd55: xpb[186] = 1024'd14429113362574422845744957354231016936459129925901106685427549322205446930711327449399726837794472508339660329268782053705568386358582988340078781205541844284678336100764479157813412272485946138747632106920789711264717825451884015291685464651268564858597057750742545495862286403037734486797801010494092300847;
            6'd56: xpb[186] = 1024'd100410268805471051863928670058543370777095481938698508568235513718411400926137847559035589255881492440470193744044300827663931919782673092002554481784198597007676953732482128939409094118852123657811907401932351599866725646067265131436428575789704703713101664795964195507497020097807294289294310363626213804582;
            6'd57: xpb[186] = 1024'd62324728564242939483313455358041291873033406825760226322911623049640459584255228758656380459310838063157577751362326167043231612365542861109870057346524308796984896794628561383374536773701095455565985088556673642104372616461749474616193117244911393300786368427068787489025225718648221074672129890132740823986;
            6'd58: xpb[186] = 1024'd24239188323014827102698240657539212968971331712821944077587732380869518242372609958277171662740183685844961758680351506422531304948412630217185632908850020586292839856774993827339979428550067253320062775180995684342019586856233817795957658700118082888471072058173379470553431339489147860049949416639267843390;
            6'd59: xpb[186] = 1024'd110220343765911456120881953361851566809607683725619345960395696777075472237799130067913034080827203617975495173455870280380894838372502733879661333487506773309291457488492643608935661274916244772384338070192557572944027407471614933940700769838554221742975679103395029482188165034258707662546458769771389347125;
            6'd60: xpb[186] = 1024'd72134803524683343740266738661349487905545608612681063715071806108304530895916511267533825284256549240662879180773895619760194530955372502986976909049832485098599400550639076052901103929765216570138415756816879615181674377866099277120465311293760911330660382734499621463716370655099634447924278296277916366529;
            6'd61: xpb[186] = 1024'd34049263283455231359651523960847409001483533499742781469747915439533589554033892467154616487685894863350263188091920959139494223538242272094292484612158196887907343612785508496866546584614188367892493443441201657419321348260583620300229852748967600918345086365604213445244576275940561233302097822784443385933;
            6'd62: xpb[186] = 1024'd120030418726351860377835236665159762842119885512540183352555879835739543549460412576790478905772914795480796602867439733097857756962332375756768185190814949610905961244503158278462228430980365886956768738452763546021329168875964736444972963887403739772849693410825863456879309970710121035798607175916564889668;
            6'd63: xpb[186] = 1024'd81944878485123747997220021964657683938057810399601901107231989166968602207577793776411270109202260418168180610185465072477157449545202144864083760753140661400213904306649590722427671085829337684710846425077085588258976139270449079624737505342610429360534397041930455438407515591551047821176426702423091909072;
        endcase
    end

    always_comb begin
        case(flag[62][11:6])
            6'd0: xpb[187] = 1024'd0;
            6'd1: xpb[187] = 1024'd43859338243895635616604807264155605033995735286663618861908098498197660865695174976032061312631606040855564617503490411856457142128071913971399336315466373189521847368796023166393113740678309482464924111701407630496623109664933422804502046797817118948219100673035047419935721212391974606554246228929618928476;
            6'd2: xpb[187] = 1024'd87718676487791271233209614528311210067991470573327237723816196996395321731390349952064122625263212081711129235006980823712914284256143827942798672630932746379043694737592046332786227481356618964929848223402815260993246219329866845609004093595634237896438201346070094839871442424783949213108492457859237856952;
            6'd3: xpb[187] = 1024'd7511319047562165451015494387652382357288778734255172457592440429616087259776386018081112723237143813123544445052977800990307585542995407359037883930068078634874867536816852161549102030517722726084574726716983045125508478773903495448527570710221907577837398604988084229700635563247290802544048860163262301097;
            6'd4: xpb[187] = 1024'd51370657291457801067620301651807987391284514020918791319500538927813748125471560994113174035868749853979109062556468212846764727671067321330437220245534451824396714905612875327942215771196032208549498838418390675622131588438836918253029617508039026526056499278023131649636356775639265409098295089092881229573;
            6'd5: xpb[187] = 1024'd95229995535353436684225108915963592425280249307582410181408637426011408991166735970145235348500355894834673680059958624703221869799139235301836556561000825013918562274408898494335329511874341691014422950119798306118754698103770341057531664305856145474275599951058179069572077988031240015652541318022500158049;
            6'd6: xpb[187] = 1024'd15022638095124330902030988775304764714577557468510344915184880859232174519552772036162225446474287626247088890105955601980615171085990814718075767860136157269749735073633704323098204061035445452169149453433966090251016957547806990897055141420443815155674797209976168459401271126494581605088097720326524602194;
            6'd7: xpb[187] = 1024'd58881976339019966518635796039460369748573292755173963777092979357429835385247947012194286759105893667102653507609446013837072313214062728689475104175602530459271582442429727489491317801713754934634073565135373720747640067212740413701557188218260934103893897883011215879336992338886556211642343949256143530670;
            6'd8: xpb[187] = 1024'd102741314582915602135240603303615974782569028041837582639001077855627496250943121988226348071737499707958218125112936425693529455342134642660874440491068903648793429811225750655884431542392064417098997676836781351244263176877673836506059235016078053052112998556046263299272713551278530818196590178185762459146;
            6'd9: xpb[187] = 1024'd22533957142686496353046483162957147071866336202765517372777321288848261779329158054243338169711431439370633335158933402970922756628986222077113651790204235904624602610450556484647306091553168178253724180150949135376525436321710486345582712130665722733512195814964252689101906689741872407632146580489786903291;
            6'd10: xpb[187] = 1024'd66393295386582131969651290427112752105862071489429136234685419787045922645024333030275399482343037480226197952662423814827379898757058136048512988105670609094146449979246579651040419832231477660718648291852356765873148545986643909150084758928482841681731296487999300109037627902133847014186392809419405831767;
            6'd11: xpb[187] = 1024'd110252633630477767586256097691268357139857806776092755096593518285243583510719508006307460794974643521081762570165914226683837040885130050019912324421136982283668297348042602817433533572909787143183572403553764396369771655651577331954586805726299960629950397161034347528973349114525821620740639038349024760243;
            6'd12: xpb[187] = 1024'd30045276190248661804061977550609529429155114937020689830369761718464349039105544072324450892948575252494177780211911203961230342171981629436151535720272314539499470147267408646196408122070890904338298906867932180502033915095613981794110282840887630311349594419952336918802542252989163210176195440653049204388;
            6'd13: xpb[187] = 1024'd73904614434144297420666784814765134463150850223684308692277860216662009904800719048356512205580181293349742397715401615817687484300053543407550872035738687729021317516063431812589521862749200386803223018569339810998657024760547404598612329638704749259568695092987384338738263465381137816730441669582668132864;
            6'd14: xpb[187] = 1024'd117763952678039933037271592078920739497146585510347927554185958714859670770495894024388573518211787334205307015218892027674144626428125457378950208351205060918543164884859454978982635603427509869268147130270747441495280134425480827403114376436521868207787795766022431758673984677773112423284687898512287061340;
            6'd15: xpb[187] = 1024'd37556595237810827255077471938261911786443893671275862287962202148080436298881930090405563616185719065617722225264889004951537927714977036795189419650340393174374337684084260807745510152588613630422873633584915225627542393869517477242637853551109537889186993024940421148503177816236454012720244300816311505485;
            6'd16: xpb[187] = 1024'd81415933481706462871682279202417516820439628957939481149870300646278097164577105066437624928817325106473286842768379416807995069843048950766588755965806766363896185052880283974138623893266923112887797745286322856124165503534450900047139900348926656837406093697975468568438899028628428619274490529745930433961;
            6'd17: xpb[187] = 1024'd1208576041477357089488159061758689109736937118867415883646544079498862692963141132454615026791256837885702052814376394085388371129900530182827967264942098619727357852105089802901498442428026874042524248600490640256427762978487549886663377463514326518805290956893457958268092167091770208710046932049954878106;
            6'd18: xpb[187] = 1024'd45067914285372992706092966325914294143732672405531034745554642577696523558658316108486676339422862878741266670317866805941845513257972444154227303580408471809249205220901112969294612183106336356507448360301898270753050872643420972691165424261331445467024391629928505378203813379483744815264293160979573806582;
            6'd19: xpb[187] = 1024'd88927252529268628322697773590069899177728407692194653607462741075894184424353491084518737652054468919596831287821357217798302655386044358125626639895874844998771052589697136135687725923784645838972372472003305901249673982308354395495667471059148564415243492302963552798139534591875719421818539389909192735058;
            6'd20: xpb[187] = 1024'd8719895089039522540503653449411071467025715853122588341238984509114949952739527150535727750028400651009246497867354195075695956672895937541865851195010177254602225388921941964450600472945749600127098975317473685381936241752391045335190948173736234096642689561881542187968727730339061011254095792213217179203;
            6'd21: xpb[187] = 1024'd52579233332935158157108460713566676501021451139786207203147083007312610818434702126567789062660006691864811115370844606932153098800967851513265187510476550444124072757717965130843714213624059082592023087018881315878559351417324468139692994971553353044861790234916589607904448942731035617808342021142836107679;
            6'd22: xpb[187] = 1024'd96438571576830793773713267977722281535017186426449826065055181505510271684129877102599850375291612732720375732874335018788610240929039765484664523825942923633645920126513988297236827954302368565056947198720288946375182461082257890944195041769370471993080890907951637027840170155123010224362588250072455036155;
            6'd23: xpb[187] = 1024'd16231214136601687991519147837063453824314494587377760798831424938731037212515913168616840473265544464132790942920331996066003542215891344900903735125078255889477092925738794125999702503463472326211673702034456730507444720526294540783718518883958141674480088166869626417669363293586351813798144652376479480300;
            6'd24: xpb[187] = 1024'd60090552380497323608123955101219058858310229874041379660739523436928698078211088144648901785897150504988355560423822407922460684343963258872303071440544629078998940294534817292392816244141781808676597813735864361004067830191227963588220565681775260622699188839904673837605084505978326420352390881306098408776;
            6'd25: xpb[187] = 1024'd103949890624392959224728762365374663892305965160704998522647621935126358943906263120680963098528756545843920177927312819778917826472035172843702407756011002268520787663330840458785929984820091291141521925437271991500690939856161386392722612479592379570918289512939721257540805718370301026906637110235717337252;
            6'd26: xpb[187] = 1024'd23742533184163853442534642224715836181603273321632933256423865368347124472292299186697953196502688277256335387973309797056311127758886752259941619055146334524351960462555646287548804533981195052296248428751439775632953199300198036232246089594180049252317486771857710647369998856833642616342193512539741781397;
            6'd27: xpb[187] = 1024'd67601871428059489059139449488871441215599008608296552118331963866544785337987474162730014509134294318111900005476800208912768269886958666231340955370612707713873807831351669453941918274659504534761172540452847406129576308965131459036748136391997168200536587444892758067305720069225617222896439741469360709873;
            6'd28: xpb[187] = 1024'd111461209671955124675744256753027046249594743894960170980240062364742446203682649138762075821765900358967464622980290620769225412015030580202740291686079080903395655200147692620335032015337814017226096652154255036626199418630064881841250183189814287148755688117927805487241441281617591829450685970398979638349;
            6'd29: xpb[187] = 1024'd31253852231726018893550136612368218538892052055888105714016305797963211732068685204779065919739832090379879833026287598046618713301882159618979502985214413159226827999372498449097906564498917778380823155468422820758461678074101531680773660304401956830154885376845794877070634420080933418886242372703004082494;
            6'd30: xpb[187] = 1024'd75113190475621654510154943876523823572887787342551724575924404296160872597763860180811127232371438131235444450529778009903075855429954073590378839300680786348748675368168521615491020305177227260845747267169830451255084787739034954485275707102219075778373986049880842297006355632472908025440488601632623010970;
            6'd31: xpb[187] = 1024'd118972528719517290126759751140679428606883522629215343437832502794358533463459035156843188545003044172091009068033268421759532997558025987561778175616147159538270522736964544781884134045855536743310671378871238081751707897403968377289777753900036194726593086722915889716942076844864882631994734830562241939446;
            6'd32: xpb[187] = 1024'd38765171279288184344565631000020600896180830790143278171608746227579298991845071222860178642976975903503424278079265399036926298844877566978017386915282491794101695536189350610647008595016640504465397882185405865883970156848005027129301231014623864407992283981833879106771269983328224221430291232866266383591;
            6'd33: xpb[187] = 1024'd82624509523183819961170438264176205930176566076806897033516844725776959857540246198892239955608581944358988895582755810893383440972949480949416723230748864983623542904985373777040122335694949986930321993886813496380593266512938449933803277812440983356211384654868926526706991195720198827984537461795885312067;
            6'd34: xpb[187] = 1024'd2417152082954714178976318123517378219473874237734831767293088158997725385926282264909230053582513675771404105628752788170776742259801060365655934529884197239454715704210179605802996884856053748085048497200981280512855525956975099773326754927028653037610581913786915916536184334183540417420093864099909756212;
            6'd35: xpb[187] = 1024'd46276490326850349795581125387672983253469609524398450629201186657195386251621457240941291366214119716626968723132243200027233884387872974337055270845350570428976563073006202772196110625534363230549972608902388911009478635621908522577828801724845771985829682586821963336471905546575515023974340093029528684688;
            6'd36: xpb[187] = 1024'd90135828570745985412185932651828588287465344811062069491109285155393047117316632216973352678845725757482533340635733611883691026515944888308454607160816943618498410441802225938589224366212672713014896720603796541506101745286841945382330848522662890934048783259857010756407626758967489630528586321959147613164;
            6'd37: xpb[187] = 1024'd9928471130516879629991812511169760576762652971990004224885528588613812645702668282990342776819657488894948550681730589161084327802796467724693818459952275874329583241027031767352098915373776474169623223917964325638364004730878595221854325637250560615447980518775000146236819897430831219964142724263172057309;
            6'd38: xpb[187] = 1024'd53787809374412515246596619775325365610758388258653623086793627086811473511397843259022404089451263529750513168185221001017541469930868381696093154775418649063851430609823054933745212656052085956634547335619371956134987114395812018026356372435067679563667081191810047566172541109822805826518388953192790985785;
            6'd39: xpb[187] = 1024'd97647147618308150863201427039480970644754123545317241948701725585009134377093018235054465402082869570606077785688711412873998612058940295667492491090885022253373277978619078100138326396730395439099471447320779586631610224060745440830858419232884798511886181864845094986108262322214780433072635182122409914261;
            6'd40: xpb[187] = 1024'd17439790178079045081007306898822142934051431706245176682477969018229899905479054301071455500056801302018492995734708390151391913345791875083731702390020354509204450777843883928901200945891499200254197950634947370763872483504782090670381896347472468193285379123763084375937455460678122022508191584426434358406;
            6'd41: xpb[187] = 1024'd61299128421974680697612114162977747968047166992908795544386067516427560771174229277103516812688407342874057613238198802007849055473863789055131038705486727698726298146639907095294314686569808682719122062336355001260495593169715513474883943145289587141504479796798131795873176673070096629062437813356053286882;
            6'd42: xpb[187] = 1024'd105158466665870316314216921427133353002042902279572414406294166014625221636869404253135578125320013383729622230741689213864306197601935703026530375020953100888248145515435930261687428427248118165184046174037762631757118702834648936279385989943106706089723580469833179215808897885462071235616684042285672215358;
            6'd43: xpb[187] = 1024'd24951109225641210532022801286474525291340210440500349140070409447845987165255440319152568223293945115142037440787686191141699498888787282442769586320088433144079318314660736090450302976409221926338772677351930415889380962278685586118909467057694375771122777728751168605638091023925412825052240444589696659503;
            6'd44: xpb[187] = 1024'd68810447469536846148627608550630130325335945727163968001978507946043648030950615295184629535925551155997602058291176602998156641016859196414168922635554806333601165683456759256843416717087531408803696789053338046386004071943619008923411513855511494719341878401786216025573812236317387431606486673519315587979;
            6'd45: xpb[187] = 1024'd112669785713432481765232415814785735359331681013827586863886606444241308896645790271216690848557157196853166675794667014854613783144931110385568258951021179523123013052252782423236530457765840891268620900754745676882627181608552431727913560653328613667560979074821263445509533448709362038160732902448934516455;
            6'd46: xpb[187] = 1024'd32462428273203375983038295674126907648628989174755521597662849877462074425031826337233680946531088928265581885840663992132007084431782689801807470250156511778954185851477588251999405006926944652423347404068913461014889441052589081567437037767916283348960176333739252835338726587172703627596289304752958960600;
            6'd47: xpb[187] = 1024'd76321766517099011599643102938282512682624724461419140459570948375659735290727001313265742259162694969121146503344154403988464226559854603773206806565622884968476033220273611418392518747605254134888271515770321091511512550717522504371939084565733402297179277006774300255274447799564678234150535533682577889076;
            6'd48: xpb[187] = 1024'd120181104760994647216247910202438117716620459748082759321479046873857396156422176289297803571794301009976711120847644815844921368687926517744606142881089258157997880589069634584785632488283563617353195627471728722008135660382455927176441131363550521245398377679809347675210169011956652840704781762612196817552;
            6'd49: xpb[187] = 1024'd39973747320765541434053790061779290005917767909010694055255290307078161684808212355314793669768232741389126330893641793122314669974778097160845354180224590413829053388294440413548507037444667378507922130785896506140397919826492577015964608478138190926797574938727337065039362150419994430140338164916221261697;
            6'd50: xpb[187] = 1024'd83833085564661177050658597325934895039913503195674312917163388805275822550503387331346854982399838782244690948397132204978771812102850011132244690495690963603350900757090463579941620778122976860972846242487304136637021029491425999820466655275955309875016675611762384484975083362811969036694584393845840190173;
            6'd51: xpb[187] = 1024'd3625728124432071268464477185276067329210811356602247650939632238496588078889423397363845080373770513657106158443129182256165113389701590548483901794826295859182073556315269408704495327284080622127572745801471920769283288935462649659990132390542979556415872870680373874804276501275310626130140796149864634318;
            6'd52: xpb[187] = 1024'd47485066368327706885069284449431672363206546643265866512847730736694248944584598373395906393005376554512670775946619594112622255517773504519883238110292669048703920925111292575097609067962390104592496857502879551265906398600396072464492179188360098504634973543715421294739997713667285232684387025079483562794;
            6'd53: xpb[187] = 1024'd91344404612223342501674091713587277397202281929929485374755829234891909810279773349427967705636982595368235393450110005969079397645845418491282574425759042238225768293907315741490722808640699587057420969204287181762529508265329495268994225986177217452854074216750468714675718926059259839238633254009102491270;
            6'd54: xpb[187] = 1024'd11137047171994236719479971572928449686499590090857420108532072668112675338665809415444957803610914326780650603496106983246472698932696997907521785724894374494056941093132121570253597357801803348212147472518454965894791767709366145108517703100764887134253271475668458104504912064522601428674189656313126935415;
            6'd55: xpb[187] = 1024'd54996385415889872336084778837084054720495325377521038970440171166310336204360984391477019116242520367636215220999597395102929841060768911878921122040360747683578788461928144736646711098480112830677071584219862596391414877374299567913019749898582006082472372148703505524440633276914576035228435885242745863891;
            6'd56: xpb[187] = 1024'd98855723659785507952689586101239659754491060664184657832348269664507997070056159367509080428874126408491779838503087806959386983188840825850320458355827120873100635830724167903039824839158422313141995695921270226888037987039232990717521796696399125030691472821738552944376354489306550641782682114172364792367;
            6'd57: xpb[187] = 1024'd18648366219556402170495465960580832043788368825112592566124513097728762598442195433526070526848058139904195048549084784236780284475692405266559669654962453128931808629948973731802699388319526074296722199235438011020300246483269640557045273810986794712090670080656542334205547627769892231218238516476389236512;
            6'd58: xpb[187] = 1024'd62507704463452037787100273224736437077784104111776211428032611595926423464137370409558131839479664180759759666052575196093237426603764319237959005970428826318453655998744996898195813128997835556761646310936845641516923356148203063361547320608803913660309770753691589754141268840161866837772484745406008164988;
            6'd59: xpb[187] = 1024'd106367042707347673403705080488892042111779839398439830289940710094124084329832545385590193152111270221615324283556065607949694568731836233209358342285895199507975503367541020064588926869676145039226570422638253272013546465813136486166049367406621032608528871426726637174076990052553841444326730974335627093464;
            6'd60: xpb[187] = 1024'd26159685267118567621510960348233214401077147559367765023716953527344849858218581451607183250085201953027739493602062585227087870018687812625597553585030531763806676166765825893351801418837248800381296925952421056145808725257173136005572844521208702289928068685644626563906183191017183033762287376639651537609;
            6'd61: xpb[187] = 1024'd70019023511014203238115767612388819435072882846031383885625052025542510723913756427639244562716807993883304111105552997083545012146759726596996889900496904953328523535561849059744915159515558282846221037653828686642431834922106558810074891319025821238147169358679673983841904403409157640316533605569270466085;
            6'd62: xpb[187] = 1024'd113878361754909838854720574876544424469068618132695002747533150523740171589608931403671305875348414034738868728609043408940002154274831640568396226215963278142850370904357872226138028900193867765311145149355236317139054944587039981614576938116842940186366270031714721403777625615801132246870779834498889394561;
            6'd63: xpb[187] = 1024'd33671004314680733072526454735885596758365926293622937481309393956960937117994967469688295973322345766151283938655040386217395455561683219984635437515098610398681543703582678054900903449354971526465871652669404101271317204031076631454100415231430609867765467290632710793606818754264473836306336236802913838706;
        endcase
    end

    always_comb begin
        case(flag[62][16:12])
            5'd0: xpb[188] = 1024'd0;
            5'd1: xpb[188] = 1024'd77530342558576368689131262000041201792361661580286556343217492455158597983690142445720357285953951807006848556158530798073852597689755133956034773830564983588203391072378701221294017190033281008930795764370811731767940313696010054258602462029247728815984567963667758213542539966656448442860582465732532767182;
            5'd2: xpb[188] = 1024'd30993989433027995979463596595267970840024896034837428558303129845340300630071145981425643357250229304570547704859568161568641354538289933356909422644798926242716107575186185104957795188549356296551393920354383617171519777171123335552226354375266008365149232513218458396978551859384263868602475104839471050033;
            5'd3: xpb[188] = 1024'd108524331991604364668594858595309172632386557615123984901520622300498898613761288427146000643204181111577396261018098959642493952228045067312944196475363909830919498647564886326251812378582637305482189684725195348939460090867133389810828816404513737181133800476886216610521091826040712311463057570572003817215;
            5'd4: xpb[188] = 1024'd61987978866055991958927193190535941680049792069674857116606259690680601260142291962851286714500458609141095409719136323137282709076579866713818845289597852485432215150372370209915590377098712593102787840708767234343039554342246671104452708750532016730298465026436916793957103718768527737204950209678942100066;
            5'd5: xpb[188] = 1024'd15451625740507619249259527785762710727713026524225729331691897080862303906523295498556572785796736106704794558420173686632071465925114666114693494103831795139944931653179854093579368375614787880723385996692339119746619017817359952398076601096550296279463129575987616977393115611496343162946842848785880382917;
            5'd6: xpb[188] = 1024'd92981968299083987938390789785803912520074688104512285674909389536020901890213437944276930071750687913711643114578704484705924063614869800070728267934396778728148322725558555314873385565648068889654181761063150851514559331513370006656679063125798025095447697539655375190935655578152791605807425314518413150099;
            5'd7: xpb[188] = 1024'd46445615173535615228723124381030681567737922559063157889995026926202604536594441479982216143046965411275342263279741848200712820463404599471602916748630721382661039228366039198537163564164144177274779917046722736918138794988483287950302955471816304644612362089206075374371667470880607031549317953625351432950;
            5'd8: xpb[188] = 1024'd123975957732111983917854386381071883360099584139349714233212519381361202520284583925702573429000917218282190819438272646274565418153159733427637690579195704970864430300744740419831180754197425186205575681417534468686079108684493342208905417501064033460596930052873833587914207437537055474409900419357884200132;
            5'd9: xpb[188] = 1024'd77439604606563611208186720976298652407762818593900586448298156771542905166665587461407859500297194715845889968139310009769354175001694532828512339393429647625377146803552224303494958752713500473826173837401106354089658572159606623502529309847082313009761594602424533771350219330264870900151793058464822482983;
            5'd10: xpb[188] = 1024'd30903251481015238498519055571525421455426053048451458663383794161724607813046590997113145571593472213409589116840347373264142931850229332229386988207663590279889863306359708187158736751229575761446771993384678239493238035634719904796153202193100592558926259151975233954786231222992686325893685697571760765834;
            5'd11: xpb[188] = 1024'd108433594039591607187650317571566623247787714628738015006601286616883205796736733442833502857547424020416437672998878171337995529539984466185421762038228573868093254378738409408452753941262856770377567757755489971261178349330729959054755664222348321374910827115642992168328771189649134768754268163304293533016;
            5'd12: xpb[188] = 1024'd61897240914043234477982652166793392295450949083288887221686924007064908443117736978538788928843701517980136821699915534832784286388519265586296410852462516522605970881545893292116531939778932057998165913739061856664757812805843240348379556568366600924075491665193692351764783082376950194496160802411231815867;
            5'd13: xpb[188] = 1024'd15360887788494861768314986762020161343114183537839759436772561397246611089498740514244075000139979015543835970400952898327573043237054064987171059666696459177118687384353377175780309938295007345618764069722633742068337276280956521642003448914384880473240156214744392535200794975104765620238053441518170098718;
            5'd14: xpb[188] = 1024'd92891230347071230457446248762061363135475845118126315779990053852405209073188882959964432286093930822550684526559483696401425640926809198943205833497261442765322078456732078397074327128328288354549559834093445473836277589976966575900605910943632609289224724178412150748743334941761214063098635907250702865900;
            5'd15: xpb[188] = 1024'd46354877221522857747778583357288132183139079572677187995075691242586911719569886495669718357390208320114383675260521059896214397775343998344080482311495385419834794959539562280738105126844363642170157990077017359239857053452079857194229803289650888838389388727962850932179346834489029488840528546357641148751;
            5'd16: xpb[188] = 1024'd123885219780099226436909845357329333975500741152963744338293183697745509703260028941390075643344160127121232231419051857970066995465099132300115256142060369008038186031918263502032122316877644651100953754447829091007797367148089911452832265318898617654373956691630609145721886801145477931701111012090173915933;
            5'd17: xpb[188] = 1024'd77348866654550853727242179952556103023163975607514616553378821087927212349641032477095361714640437624684931380120089221464855752313633931700989904956294311662550902534725747385695900315393719938721551910431400976411376830623203192746456157664916897203538621241181309329157898693873293357443003651197112198784;
            5'd18: xpb[188] = 1024'd30812513529002481017574514547782872070827210062065488768464458478108914996022036012800647785936715122248630528821126584959644509162168731101864553770528254317063619037533231269359678313909795226342150066414972861814956294098316474040080050010935176752703285790732009512593910586601108783184896290304050481635;
            5'd19: xpb[188] = 1024'd108342856087578849706705776547824073863188871642352045111681950933267512979712178458521005071890666929255479084979657383033497106851923865057899327601093237905267010109911932490653695503943076235272945830785784593582896607794326528298682512040182905568687853754399767726136450553257557226045478756036583248817;
            5'd20: xpb[188] = 1024'd61806502962030476997038111143050842910852106096902917326767588323449215626093181994226291143186944426819178233680694746528285863700458664458773976415327180559779726612719416374317473502459151522893543986769356478986476071269439809592306404386201185117852518303950467909572462445985372651787371395143521531668;
            5'd21: xpb[188] = 1024'd15270149836482104287370445738277611958515340551453789541853225713630918272474185529931577214483221924382877382381732110023074620548993463859648625229561123214292443115526900257981251500975226810514142142752928364390055534744553090885930296732219464667017182853501168093008474338713188077529264034250459814519;
            5'd22: xpb[188] = 1024'd92800492395058472976501707738318813750877002131740345885070718168789516256164327975651934500437173731389725938540262908096927218238748597815683399060126106802495834187905601479275268691008507819444937907123740096157995848440563145144532758761467193483001750817168926306551014305369636520389846499982992581701;
            5'd23: xpb[188] = 1024'd46264139269510100266834042333545582798540236586291218100156355558971218902545331511357220571733451228953425087241300271591715975087283397216558047874360049457008550690713085362939046689524583107065536063107311981561575311915676426438156651107485473032166415366719626489987026198097451946131739139089930864552;
            5'd24: xpb[188] = 1024'd123794481828086468955965304333586784590901898166577774443373848014129816886235473957077577857687403035960273643399831069665568572777038531172592821704925033045211941763091786584233063879557864115996331827478123713329515625611686480696759113136733201848150983330387384703529566164753900388992321604822463631734;
            5'd25: xpb[188] = 1024'd77258128702538096246297638928813553638565132621128646658459485404311519532616477492782863928983680533523972792100868433160357329625573330573467470519158975699724658265899270467896841878073939403616929983461695598733095089086799761990383005482751481397315647879938084886965578057481715814734214243929401914585;
            5'd26: xpb[188] = 1024'd30721775576989723536629973524040322686228367075679518873545122794493222178997481028488150000279958031087671940801905796655146086474108129974342119333392918354237374768706754351560619876590014691237528139445267484136674552561913043284006897828769760946480312429488785070401589950209531240476106883036340197436;
            5'd27: xpb[188] = 1024'd108252118135566092225761235524081524478590028655966075216762615249651820162687623474208507286233909838094520496960436594728998684163863263930376893163957901942440765841085455572854637066623295700168323903816079215904614866257923097542609359858017489762464880393156543283944129916865979683336689348768872964618;
            5'd28: xpb[188] = 1024'd61715765010017719516093570119308293526253263110516947431848252639833522809068627009913793357530187335658219645661473958223787441012398063331251541978191844596953482343892939456518415065139370987788922059799651101308194329733036378836233252204035769311629544942707243467380141809593795109078581987875811247469;
            5'd29: xpb[188] = 1024'd15179411884469346806425904714535062573916497565067819646933890030015225455449630545619079428826464833221918794362511321718576197860932862732126190792425787251466198846700423340182193063655446275409520215783222986711773793208149660129857144550054048860794209492257943650816153702321610534820474626982749530320;
            5'd30: xpb[188] = 1024'd92709754443045715495557166714576264366278159145354375990151382485173823439139772991339436714780416640228767350521042119792428795550687996688160964622990770839669589919079124561476210253688727284340315980154034718479714106904159714388459606579301777676778777455925701864358693668978058977681057092715282297502;
            5'd31: xpb[188] = 1024'd46173401317497342785889501309803033413941393599905248205237019875355526085520776527044722786076694137792466499222079483287217552399222796089035613437224713494182306421886608445139988252204802571960914136137606603883293570379272995682083498925320057225943442005476402047794705561705874403422949731822220580353;
        endcase
    end

    always_comb begin
        case(flag[63][5:0])
            6'd0: xpb[189] = 1024'd0;
            6'd1: xpb[189] = 1024'd123885219780099226436909845357329333975500741152963744338293183697745509703260028941390075643344160127121232231419051857970066995465099132300115256142060369008038186031918263502032122316877644651100953754447829091007797367148089911452832265318898617654373956691630609145721886801145477931701111012090173915933;
            6'd2: xpb[189] = 1024'd123703743876073711475020763309844235206303055180191804548454512330514124069210918972765080072030645944799315055380610281361070150088977930045070387267789697082385697494265309666434005442238083580891709900508418335651233884075283049940685960954567786041928009969144160261337245528362322846283532197554753347535;
            6'd3: xpb[189] = 1024'd123522267972048196513131681262359136437105369207419864758615840963282738435161809004140084500717131762477397879342168704752073304712856727790025518393519025156733208956612355830835888567598522510682466046569007580294670401002476188428539656590236954429482063246657711376952604255579167760865953383019332779137;
            6'd4: xpb[189] = 1024'd123340792068022681551242599214874037667907683234647924968777169596051352801112699035515088929403617580155480703303727128143076459336735525534980649519248353231080720418959401995237771692958961440473222192629596824938106917929669326916393352225906122817036116524171262492567962982796012675448374568483912210739;
            6'd5: xpb[189] = 1024'd123159316163997166589353517167388938898709997261875985178938498228819967167063589066890093358090103397833563527265285551534079613960614323279935780644977681305428231881306448159639654818319400370263978338690186069581543434856862465404247047861575291204590169801684813608183321710012857590030795753948491642341;
            6'd6: xpb[189] = 1024'd122977840259971651627464435119903840129512311289104045389099826861588581533014479098265097786776589215511646351226843974925082768584493121024890911770707009379775743343653494324041537943679839300054734484750775314224979951784055603892100743497244459592144223079198364723798680437229702504613216939413071073943;
            6'd7: xpb[189] = 1024'd122796364355946136665575353072418741360314625316332105599261155494357195898965369129640102215463075033189729175188402398316085923208371918769846042896436337454123254806000540488443421069040278229845490630811364558868416468711248742379954439132913627979698276356711915839414039164446547419195638124877650505545;
            6'd8: xpb[189] = 1024'd122614888451920621703686271024933642591116939343560165809422484127125810264916259161015106644149560850867811999149960821707089077832250716514801174022165665528470766268347586652845304194400717159636246776871953803511852985638441880867808134768582796367252329634225466955029397891663392333778059310342229937147;
            6'd9: xpb[189] = 1024'd122433412547895106741797188977448543821919253370788226019583812759894424630867149192390111072836046668545894823111519245098092232456129514259756305147894993602818277730694632817247187319761156089427002922932543048155289502565635019355661830404251964754806382911739018070644756618880237248360480495806809368749;
            6'd10: xpb[189] = 1024'd122251936643869591779908106929963445052721567398016286229745141392663038996818039223765115501522532486223977647073077668489095387080008312004711436273624321677165789193041678981649070445121595019217759068993132292798726019492828157843515526039921133142360436189252569186260115346097082162942901681271388800351;
            6'd11: xpb[189] = 1024'd122070460739844076818019024882478346283523881425244346439906470025431653362768929255140119930209018303902060471034636091880098541703887109749666567399353649751513300655388725146050953570482033949008515215053721537442162536420021296331369221675590301529914489466766120301875474073313927077525322866735968231953;
            6'd12: xpb[189] = 1024'd121888984835818561856129942834993247514326195452472406650067798658200267728719819286515124358895504121580143294996194515271101696327765907494621698525082977825860812117735771310452836695842472878799271361114310782085599053347214434819222917311259469917468542744279671417490832800530771992107744052200547663555;
            6'd13: xpb[189] = 1024'd121707508931793046894240860787508148745128509479700466860229127290968882094670709317890128787581989939258226118957752938662104850951644705239576829650812305900208323580082817474854719821202911808590027507174900026729035570274407573307076612946928638305022596021793222533106191527747616906690165237665127095157;
            6'd14: xpb[189] = 1024'd121526033027767531932351778740023049975930823506928527070390455923737496460621599349265133216268475756936308942919311362053108005575523502984531960776541633974555835042429863639256602946563350738380783653235489271372472087201600711794930308582597806692576649299306773648721550254964461821272586423129706526759;
            6'd15: xpb[189] = 1024'd121344557123742016970462696692537951206733137534156587280551784556506110826572489380640137644954961574614391766880869785444111160199402300729487091902270962048903346504776909803658486071923789668171539799296078516015908604128793850282784004218266975080130702576820324764336908982181306735855007608594285958361;
            6'd16: xpb[189] = 1024'd121163081219716502008573614645052852437535451561384647490713113189274725192523379412015142073641447392292474590842428208835114314823281098474442223028000290123250857967123955968060369197284228597962295945356667760659345121055986988770637699853936143467684755854333875879952267709398151650437428794058865389963;
            6'd17: xpb[189] = 1024'd120981605315690987046684532597567753668337765588612707700874441822043339558474269443390146502327933209970557414803986632226117469447159896219397354153729618197598369429471002132462252322644667527753052091417257005302781637983180127258491395489605311855238809131847426995567626436614996565019849979523444821565;
            6'd18: xpb[189] = 1024'd120800129411665472084795450550082654899140079615840767911035770454811953924425159474765150931014419027648640238765545055617120624071038693964352485279458946271945880891818048296864135448005106457543808237477846249946218154910373265746345091125274480242792862409360978111182985163831841479602271164988024253167;
            6'd19: xpb[189] = 1024'd120618653507639957122906368502597556129942393643068828121197099087580568290376049506140155359700904845326723062727103479008123778694917491709307616405188274346293392354165094461266018573365545387334564383538435494589654671837566404234198786760943648630346915686874529226798343891048686394184692350452603684769;
            6'd20: xpb[189] = 1024'd120437177603614442161017286455112457360744707670296888331358427720349182656326939537515159788387390663004805886688661902399126933318796289454262747530917602420640903816512140625667901698725984317125320529599024739233091188764759542722052482396612817017900968964388080342413702618265531308767113535917183116371;
            6'd21: xpb[189] = 1024'd120255701699588927199128204407627358591547021697524948541519756353117797022277829568890164217073876480682888710650220325790130087942675087199217878656646930494988415278859186790069784824086423246916076675659613983876527705691952681209906178032281985405455022241901631458029061345482376223349534721381762547973;
            6'd22: xpb[189] = 1024'd120074225795563412237239122360142259822349335724753008751681084985886411388228719600265168645760362298360971534611778749181133242566553884944173009782376258569335926741206232954471667949446862176706832821720203228519964222619145819697759873667951153793009075519415182573644420072699221137931955906846341979575;
            6'd23: xpb[189] = 1024'd119892749891537897275350040312657161053151649751981068961842413618655025754179609631640173074446848116039054358573337172572136397190432682689128140908105586643683438203553279118873551074807301106497588967780792473163400739546338958185613569303620322180563128796928733689259778799916066052514377092310921411177;
            6'd24: xpb[189] = 1024'd119711273987512382313460958265172062283953963779209129172003742251423640120130499663015177503133333933717137182534895595963139551814311480434083272033834914718030949665900325283275434200167740036288345113841381717806837256473532096673467264939289490568117182074442284804875137527132910967096798277775500842779;
            6'd25: xpb[189] = 1024'd119529798083486867351571876217686963514756277806437189382165070884192254486081389694390181931819819751395220006496454019354142706438190278179038403159564242792378461128247371447677317325528178966079101259901970962450273773400725235161320960574958658955671235351955835920490496254349755881679219463240080274381;
            6'd26: xpb[189] = 1024'd119348322179461352389682794170201864745558591833665249592326399516960868852032279725765186360506305569073302830458012442745145861062069075923993534285293570866725972590594417612079200450888617895869857405962560207093710290327918373649174656210627827343225288629469387036105854981566600796261640648704659705983;
            6'd27: xpb[189] = 1024'd119166846275435837427793712122716765976360905860893309802487728149729483217983169757140190789192791386751385654419570866136149015685947873668948665411022898941073484052941463776481083576249056825660613552023149451737146807255111512137028351846296995730779341906982938151721213708783445710844061834169239137585;
            6'd28: xpb[189] = 1024'd118985370371410322465904630075231667207163219888121370012649056782498097583934059788515195217879277204429468478381129289527152170309826671413903796536752227015420995515288509940882966701609495755451369698083738696380583324182304650624882047481966164118333395184496489267336572436000290625426483019633818569187;
            6'd29: xpb[189] = 1024'd118803894467384807504015548027746568437965533915349430222810385415266711949884949819890199646565763022107551302342687712918155324933705469158858927662481555089768506977635556105284849826969934685242125844144327941024019841109497789112735743117635332505887448462010040382951931163217135540008904205098398000789;
            6'd30: xpb[189] = 1024'd118622418563359292542126465980261469668767847942577490432971714048035326315835839851265204075252248839785634126304246136309158479557584266903814058788210883164116018439982602269686732952330373615032881990204917185667456358036690927600589438753304500893441501739523591498567289890433980454591325390562977432391;
            6'd31: xpb[189] = 1024'd118440942659333777580237383932776370899570161969805550643133042680803940681786729882640208503938734657463716950265804559700161634181463064648769189913940211238463529902329648434088616077690812544823638136265506430310892874963884066088443134388973669280995555017037142614182648617650825369173746576027556863993;
            6'd32: xpb[189] = 1024'd118259466755308262618348301885291272130372475997033610853294371313572555047737619914015212932625220475141799774227362983091164788805341862393724321039669539312811041364676694598490499203051251474614394282326095674954329391891077204576296830024642837668549608294550693729798007344867670283756167761492136295595;
            6'd33: xpb[189] = 1024'd118077990851282747656459219837806173361174790024261671063455699946341169413688509945390217361311706292819882598188921406482167943429220660138679452165398867387158552827023740762892382328411690404405150428386684919597765908818270343064150525660312006056103661572064244845413366072084515198338588946956715727197;
            6'd34: xpb[189] = 1024'd117896514947257232694570137790321074591977104051489731273617028579109783779639399976765221789998192110497965422150479829873171098053099457883634583291128195461506064289370786927294265453772129334195906574447274164241202425745463481552004221295981174443657714849577795961028724799301360112921010132421295158799;
            6'd35: xpb[189] = 1024'd117715039043231717732681055742835975822779418078717791483778357211878398145590290008140226218684677928176048246112038253264174252676978255628589714416857523535853575751717833091696148579132568263986662720507863408884638942672656620039857916931650342831211768127091347076644083526518205027503431317885874590401;
            6'd36: xpb[189] = 1024'd117533563139206202770791973695350877053581732105945851693939685844647012511541180039515230647371163745854131070073596676655177407300857053373544845542586851610201087214064879256098031704493007193777418866568452653528075459599849758527711612567319511218765821404604898192259442253735049942085852503350454022003;
            6'd37: xpb[189] = 1024'd117352087235180687808902891647865778284384046133173911904101014477415626877492070070890235076057649563532213894035155100046180561924735851118499976668316179684548598676411925420499914829853446123568175012629041898171511976527042897015565308202988679606319874682118449307874800980951894856668273688815033453605;
            6'd38: xpb[189] = 1024'd117170611331155172847013809600380679515186360160401972114262343110184241243442960102265239504744135381210296717996713523437183716548614648863455107794045507758896110138758971584901797955213885053358931158689631142814948493454236035503419003838657847993873927959632000423490159708168739771250694874279612885207;
            6'd39: xpb[189] = 1024'd116989135427129657885124727552895580745988674187630032324423671742952855609393850133640243933430621198888379541958271946828186871172493446608410238919774835833243621601106017749303681080574323983149687304750220387458385010381429173991272699474327016381427981237145551539105518435385584685833116059744192316809;
            6'd40: xpb[189] = 1024'd116807659523104142923235645505410481976790988214858092534585000375721469975344740165015248362117107016566462365919830370219190025796372244353365370045504163907591133063453063913705564205934762912940443450810809632101821527308622312479126395109996184768982034514659102654720877162602429600415537245208771748411;
            6'd41: xpb[189] = 1024'd116626183619078627961346563457925383207593302242086152744746329008490084341295630196390252790803592834244545189881388793610193180420251042098320501171233491981938644525800110078107447331295201842731199596871398876745258044235815450966980090745665353156536087792172653770336235889819274514997958430673351180013;
            6'd42: xpb[189] = 1024'd116444707715053112999457481410440284438395616269314212954907657641258698707246520227765257219490078651922628013842947217001196335044129839843275632296962820056286155988147156242509330456655640772521955742931988121388694561163008589454833786381334521544090141069686204885951594617036119429580379616137930611615;
            6'd43: xpb[189] = 1024'd116263231811027598037568399362955185669197930296542273165068986274027313073197410259140261648176564469600710837804505640392199489668008637588230763422692148130633667450494202406911213582016079702312711888992577366032131078090201727942687482017003689931644194347199756001566953344252964344162800801602510043217;
            6'd44: xpb[189] = 1024'd116081755907002083075679317315470086900000244323770333375230314906795927439148300290515266076863050287278793661766064063783202644291887435333185894548421476204981178912841248571313096707376518632103468035053166610675567595017394866430541177652672858319198247624713307117182312071469809258745221987067089474819;
            6'd45: xpb[189] = 1024'd115900280002976568113790235267984988130802558350998393585391643539564541805099190321890270505549536104956876485727622487174205798915766233078141025674150804279328690375188294735714979832736957561894224181113755855319004111944588004918394873288342026706752300902226858232797670798686654173327643172531668906421;
            6'd46: xpb[189] = 1024'd115718804098951053151901153220499889361604872378226453795552972172333156171050080353265274934236021922634959309689180910565208953539645030823096156799880132353676201837535340900116862958097396491684980327174345099962440628871781143406248568924011195094306354179740409348413029525903499087910064357996248338023;
            6'd47: xpb[189] = 1024'd115537328194925538190012071173014790592407186405454514005714300805101770537000970384640279362922507740313042133650739333956212108163523828568051287925609460428023713299882387064518746083457835421475736473234934344605877145798974281894102264559680363481860407457253960464028388253120344002492485543460827769625;
            6'd48: xpb[189] = 1024'd115355852290900023228122989125529691823209500432682574215875629437870384902951860416015283791608993557991124957612297757347215262787402626313006419051338788502371224762229433228920629208818274351266492619295523589249313662726167420381955960195349531869414460734767511579643746980337188917074906728925407201227;
            6'd49: xpb[189] = 1024'd115174376386874508266233907078044593054011814459910634426036958070638999268902750447390288220295479375669207781573856180738218417411281424057961550177068116576718736224576479393322512334178713281057248765356112833892750179653360558869809655831018700256968514012281062695259105707554033831657327914389986632829;
            6'd50: xpb[189] = 1024'd114992900482848993304344825030559494284814128487138694636198286703407613634853640478765292648981965193347290605535414604129221572035160221802916681302797444651066247686923525557724395459539152210848004911416702078536186696580553697357663351466687868644522567289794613810874464434770878746239749099854566064431;
            6'd51: xpb[189] = 1024'd114811424578823478342455742983074395515616442514366754846359615336176228000804530510140297077668451011025373429496973027520224726659039019547871812428526772725413759149270571722126278584899591140638761057477291323179623213507746835845517047102357037032076620567308164926489823161987723660822170285319145496033;
            6'd52: xpb[189] = 1024'd114629948674797963380566660935589296746418756541594815056520943968944842366755420541515301506354936828703456253458531450911227881282917817292826943554256100799761270611617617886528161710260030070429517203537880567823059730434939974333370742738026205419630673844821716042105181889204568575404591470783724927635;
            6'd53: xpb[189] = 1024'd114448472770772448418677578888104197977221070568822875266682272601713456732706310572890305935041422646381539077420089874302231035906796615037782074679985428874108782073964664050930044835620469000220273349598469812466496247362133112821224438373695373807184727122335267157720540616421413489987012656248304359237;
            6'd54: xpb[189] = 1024'd114266996866746933456788496840619099208023384596050935476843601234482071098657200604265310363727908464059621901381648297693234190530675412782737205805714756948456293536311710215331927960980907930011029495659059057109932764289326251309078134009364542194738780399848818273335899343638258404569433841712883790839;
            6'd55: xpb[189] = 1024'd114085520962721418494899414793134000438825698623278995687004929867250685464608090635640314792414394281737704725343206721084237345154554210527692336931444085022803804998658756379733811086341346859801785641719648301753369281216519389796931829645033710582292833677362369388951258070855103319151855027177463222441;
            6'd56: xpb[189] = 1024'd113904045058695903533010332745648901669628012650507055897166258500019299830558980667015319221100880099415787549304765144475240499778433008272647468057173413097151316461005802544135694211701785789592541787780237546396805798143712528284785525280702878969846886954875920504566616798071948233734276212642042654043;
            6'd57: xpb[189] = 1024'd113722569154670388571121250698163802900430326677735116107327587132787914196509870698390323649787365917093870373266323567866243654402311806017602599182902741171498827923352848708537577337062224719383297933840826791040242315070905666772639220916372047357400940232389471620181975525288793148316697398106622085645;
            6'd58: xpb[189] = 1024'd113541093250644873609232168650678704131232640704963176317488915765556528562460760729765328078473851734771953197227881991257246809026190603762557730308632069245846339385699894872939460462422663649174054079901416035683678831998098805260492916552041215744954993509903022735797334252505638062899118583571201517247;
            6'd59: xpb[189] = 1024'd113359617346619358647343086603193605362034954732191236527650244398325142928411650761140332507160337552450036021189440414648249963650069401507512861434361397320193850848046941037341343587783102578964810225962005280327115348925291943748346612187710384132509046787416573851412692979722482977481539769035780948849;
            6'd60: xpb[189] = 1024'd113178141442593843685454004555708506592837268759419296737811573031093757294362540792515336935846823370128118845150998838039253118273948199252467992560090725394541362310393987201743226713143541508755566372022594524970551865852485082236200307823379552520063100064930124967028051706939327892063960954500360380451;
            6'd61: xpb[189] = 1024'd112996665538568328723564922508223407823639582786647356947972901663862371660313430823890341364533309187806201669112557261430256272897826996997423123685820053468888873772741033366145109838503980438546322518083183769613988382779678220724054003459048720907617153342443676082643410434156172806646382139964939812053;
            6'd62: xpb[189] = 1024'd112815189634542813761675840460738309054441896813875417158134230296630986026264320855265345793219795005484284493074115684821259427521705794742378254811549381543236385235088079530546992963864419368337078664143773014257424899706871359211907699094717889295171206619957227198258769161373017721228803325429519243655;
            6'd63: xpb[189] = 1024'd112633713730517298799786758413253210285244210841103477368295558929399600392215210886640350221906280823162367317035674108212262582145584592487333385937278709617583896697435125694948876089224858298127834810204362258900861416634064497699761394730387057682725259897470778313874127888589862635811224510894098675257;
        endcase
    end

    always_comb begin
        case(flag[63][11:6])
            6'd0: xpb[190] = 1024'd0;
            6'd1: xpb[190] = 1024'd112452237826491783837897676365768111516046524868331537578456887562168214758166100918015354650592766640840450140997232531603265736769463390232288517063008037691931408159782171859350759214585297227918590956264951503544297933561257636187615090366056226070279313174984329429489486615806707550393645696358678106859;
            6'd2: xpb[190] = 1024'd100837779968858826276996425326721790287394622610927391028781920059359534179023062926015638086527858972237750874536971628627467632697706445909416909109685034450172141749993126381071279237653388734526984304142663160724235016901618499410251611048883002873738722935851600828872445157684782083668601566091761729387;
            6'd3: xpb[190] = 1024'd89223322111225868716095174287675469058742720353523244479106952556550853599880024934015921522462951303635051608076710725651669528625949501586545301156362031208412875340204080902791799260721480241135377652020374817904172100241979362632888131731709779677198132696718872228255403699562856616943557435824845351915;
            6'd4: xpb[190] = 1024'd77608864253592911155193923248629147830090818096119097929431985053742173020736986942016204958398043635032352341616449822675871424554192557263673693203039027966653608930415035424512319283789571747743770999898086475084109183582340225855524652414536556480657542457586143627638362241440931150218513305557928974443;
            6'd5: xpb[190] = 1024'd65994406395959953594292672209582826601438915838714951379757017550933492441593948950016488394333135966429653075156188919700073320482435612940802085249716024724894342520625989946232839306857663254352164347775798132264046266922701089078161173097363333284116952218453415027021320783319005683493469175291012596971;
            6'd6: xpb[190] = 1024'd54379948538326996033391421170536505372787013581310804830082050048124811862450910958016771830268228297826953808695928016724275216410678668617930477296393021483135076110836944467953359329925754760960557695653509789443983350263061952300797693780190110087576361979320686426404279325197080216768425045024096219499;
            6'd7: xpb[190] = 1024'd42765490680694038472490170131490184144135111323906658280407082545316131283307872966017055266203320629224254542235667113748477112338921724295058869343070018241375809701047898989673879352993846267568951043531221446623920433603422815523434214463016886891035771740187957825787237867075154750043380914757179842027;
            6'd8: xpb[190] = 1024'd31151032823061080911588919092443862915483209066502511730732115042507450704164834974017338702138412960621555275775406210772679008267164779972187261389747014999616543291258853511394399376061937774177344391408933103803857516943783678746070735145843663694495181501055229225170196408953229283318336784490263464555;
            6'd9: xpb[190] = 1024'd19536574965428123350687668053397541686831306809098365181057147539698770125021796982017622138073505292018856009315145307796880904195407835649315653436424011757857276881469808033114919399130029280785737739286644760983794600284144541968707255828670440497954591261922500624553154950831303816593292654223347087083;
            6'd10: xpb[190] = 1024'd7922117107795165789786417014351220458179404551694218631382180036890089545878758990017905574008597623416156742854884404821082800123650891326444045483101008516098010471680762554835439422198120787394131087164356418163731683624505405191343776511497217301414001022789772023936113492709378349868248523956430709611;
            6'd11: xpb[190] = 1024'd120374354934286949627684093380119331974225929420025756209839067599058304304044859908033260224601364264256606883852116936424348536893114281558732562546109046208029418631462934414186198636783418015312722043429307921708029617185763041378958866877553443371693314197774101453425600108516085900261894220315108816470;
            6'd12: xpb[190] = 1024'd108759897076653992066782842341073010745574027162621609660164100096249623724901821916033543660536456595653907617391856033448550432821357337235860954592786042966270152221673888935906718659851509521921115391307019578887966700526123904601595387560380220175152723958641372852808558650394160433536850090048192438998;
            6'd13: xpb[190] = 1024'd97145439219021034505881591302026689516922124905217463110489132593440943145758783924033827096471548927051208350931595130472752328749600392912989346639463039724510885811884843457627238682919601028529508739184731236067903783866484767824231908243206996978612133719508644252191517192272234966811805959781276061526;
            6'd14: xpb[190] = 1024'd85530981361388076944980340262980368288270222647813316560814165090632262566615745932034110532406641258448509084471334227496954224677843448590117738686140036482751619402095797979347758705987692535137902087062442893247840867206845631046868428926033773782071543480375915651574475734150309500086761829514359684054;
            6'd15: xpb[190] = 1024'd73916523503755119384079089223934047059618320390409170011139197587823581987472707940034393968341733589845809818011073324521156120606086504267246130732817033240992352992306752501068278729055784041746295434940154550427777950547206494269504949608860550585530953241243187050957434276028384033361717699247443306582;
            6'd16: xpb[190] = 1024'd62302065646122161823177838184887725830966418133005023461464230085014901408329669948034677404276825921243110551550812421545358016534329559944374522779494029999233086582517707022788798752123875548354688782817866207607715033887567357492141470291687327388990363002110458450340392817906458566636673568980526929110;
            6'd17: xpb[190] = 1024'd50687607788489204262276587145841404602314515875600876911789262582206220829186631956034960840211918252640411285090551518569559912462572615621502914826171026757473820172728661544509318775191967054963082130695577864787652117227928220714777990974514104192449772762977729849723351359784533099911629438713610551638;
            6'd18: xpb[190] = 1024'd39073149930856246701375336106795083373662613618196730362114295079397540250043593964035244276147010584037712018630290615593761808390815671298631306872848023515714553762939616066229838798260058561571475478573289521967589200568289083937414511657340880995909182523845001249106309901662607633186585308446694174166;
            6'd19: xpb[190] = 1024'd27458692073223289140474085067748762145010711360792583812439327576588859670900555972035527712082102915435012752170029712617963704319058726975759698919525020273955287353150570587950358821328150068179868826451001179147526283908649947160051032340167657799368592284712272648489268443540682166461541178179777796694;
            6'd20: xpb[190] = 1024'd15844234215590331579572834028702440916358809103388437262764360073780179091757517980035811148017195246832313485709768809642165600247301782652888090966202017032196020943361525109670878844396241574788262174328712836327463367249010810382687553022994434602828002045579544047872226985418756699736497047912861419222;
            6'd21: xpb[190] = 1024'd4229776357957374018671582989656119687706906845984290713089392570971498512614479988036094583952287578229614219249507906666367496175544838330016483012879013790436754533572479631391398867464333081396655522206424493507400450589371673605324073705821211406287411806446815447255185527296831233011452917645945041750;
            6'd22: xpb[190] = 1024'd116682014184449157856569259355424231203753431714315828291546280133139713270780580906051449234545054219070064360246740438269633232945008228562305000075887051482368162693354651490742158082049630309315246478471375997051698384150629309792939164071877437476566724981431144876744672143103538783405098614004623148609;
            6'd23: xpb[190] = 1024'd105067556326816200295668008316377909975101529456911681741871312630331032691637542914051732670480146550467365093786479535293835128873251284239433392122564048240608896283565606012462678105117721815923639826349087654231635467490990173015575684754704214280026134742298416276127630684981613316680054483737706771137;
            6'd24: xpb[190] = 1024'd93453098469183242734766757277331588746449627199507535192196345127522352112494504922052016106415238881864665827326218632318037024801494339916561784169241044998849629873776560534183198128185813322532033174226799311411572550831351036238212205437530991083485544503165687675510589226859687849955010353470790393665;
            6'd25: xpb[190] = 1024'd81838640611550285173865506238285267517797724942103388642521377624713671533351466930052299542350331213261966560865957729342238920729737395593690176215918041757090363463987515055903718151253904829140426522104510968591509634171711899460848726120357767886944954264032959074893547768737762383229966223203874016193;
            6'd26: xpb[190] = 1024'd70224182753917327612964255199238946289145822684699242092846410121904990954208428938052582978285423544659267294405696826366440816657980451270818568262595038515331097054198469577624238174321996335748819869982222625771446717512072762683485246803184544690404364024900230474276506310615836916504922092936957638721;
            6'd27: xpb[190] = 1024'd58609724896284370052063004160192625060493920427295095543171442619096310375065390946052866414220515876056568027945435923390642712586223506947946960309272035273571830644409424099344758197390087842357213217859934282951383800852433625906121767486011321493863773785767501873659464852493911449779877962670041261249;
            6'd28: xpb[190] = 1024'd46995267038651412491161753121146303831842018169890948993496475116287629795922352954053149850155608207453868761485175020414844608514466562625075352355949032031812564234620378621065278220458179348965606565737645940131320884192794489128758288168838098297323183546634773273042423394371985983054833832403124883777;
            6'd29: xpb[190] = 1024'd35380809181018454930260502082099982603190115912486802443821507613478949216779314962053433286090700538851169495024914117439046504442709618302203744402626028790053297824831333142785798243526270855573999913615357597311257967533155352351394808851664875100782593307502044672425381936250060516329789702136208506305;
            6'd30: xpb[190] = 1024'd23766351323385497369359251043053661374538213655082655894146540110670268637636276970053716722025792870248470228564653214463248400370952673979332136449303025548294031415042287664506318266594362362182393261493069254491195050873516215574031329534491651904242003068369316071808340478128135049604745571869292128833;
            6'd31: xpb[190] = 1024'd12151893465752539808458000004007340145886311397678509344471572607861588058493238978054000157960885201645770962104392311487450296299195729656460528495980022306534765005253242186226838289662453868790786609370780911671132134213877078796667850217318428707701412829236587471191299020006209582879701441602375751361;
            6'd32: xpb[190] = 1024'd537435608119582247556748964961018917234409140274362794796605105052907479350200986054283593895977533043071695644131408511652192227438785333588920542657019064775498595464196707947358312730545375399179957248492568851069217554237942019304370900145205511160822590103858870574257561884284116154657311335459373889;
            6'd33: xpb[190] = 1024'd112989673434611366085454425330729130433280934008605900373253492667221122237516301904069638244488744173883521836641363940114917928996902175565877437605665056756706906755246368567298117527315842603317770913513444072395367151115495578206919461266201431581440135765088188300063744177690991666548303007694137480748;
            6'd34: xpb[190] = 1024'd101375215576978408524553174291682809204629031751201753823578525164412441658373263912069921680423836505280822570181103037139119824925145231243005829652342053514947640345457323089018637550383934109926164261391155729575304234455856441429555981949028208384899545525955459699446702719569066199823258877427221103276;
            6'd35: xpb[190] = 1024'd89760757719345450963651923252636487975977129493797607273903557661603761079230225920070205116358928836678123303720842134163321720853388286920134221699019050273188373935668277610739157573452025616534557609268867386755241317796217304652192502631854985188358955286822731098829661261447140733098214747160304725804;
            6'd36: xpb[190] = 1024'd78146299861712493402750672213590166747325227236393460724228590158795080500087187928070488552294021168075424037260581231187523616781631342597262613745696047031429107525879232132459677596520117123142950957146579043935178401136578167874829023314681761991818365047690002498212619803325215266373170616893388348332;
            6'd37: xpb[190] = 1024'd66531842004079535841849421174543845518673324978989314174553622655986399920944149936070771988229113499472724770800320328211725512709874398274391005792373043789669841116090186654180197619588208629751344305024290701115115484476939031097465543997508538795277774808557273897595578345203289799648126486626471970860;
            6'd38: xpb[190] = 1024'd54917384146446578280948170135497524290021422721585167624878655153177719341801111944071055424164205830870025504340059425235927408638117453951519397839050040547910574706301141175900717642656300136359737652902002358295052567817299894320102064680335315598737184569424545296978536887081364332923082356359555593388;
            6'd39: xpb[190] = 1024'd43302926288813620720046919096451203061369520464181021075203687650369038762658073952071338860099298162267326237879798522260129304566360509628647789885727037306151308296512095697621237665724391642968131000779714015474989651157660757542738585363162092402196594330291816696361495428959438866198038226092639215916;
            6'd40: xpb[190] = 1024'd31688468431180663159145668057404881832717618206776874525528720147560358183515035960071622296034390493664626971419537619284331200494603565305776181932404034064392041886723050219341757688792483149576524348657425672654926734498021620765375106045988869205656004091159088095744453970837513399472994095825722838444;
            6'd41: xpb[190] = 1024'd20074010573547705598244417018358560604065715949372727975853752644751677604371997968071905731969482825061927704959276716308533096422846620982904573979081030822632775476934004741062277711860574656184917696535137329834863817838382483988011626728815646009115413852026359495127412512715587932747949965558806460972;
            6'd42: xpb[190] = 1024'd8459552715914748037343165979312239375413813691968581426178785141942997025228959976072189167904575156459228438499015813332734992351089676660032966025758027580873509067144959262782797734928666162793311044412848987014800901178743347210648147411642422812574823612893630894510371054593662466022905835291890083500;
            6'd43: xpb[190] = 1024'd120911790542406531875240842345080350891460338560300119004635672704111211783395060894087543818497341797299678579496248344936000729120553066892321483088766065272804917226927131122133556949513963390711902000677800490559098834740000983398263237777698648882854136787877960323999857670400370016416551531650568190359;
            6'd44: xpb[190] = 1024'd109297332684773574314339591306034029662808436302895972454960705201302531204252022902087827254432434128696979313035987441960202625048796122569449875135443062031045650817138085643854076972582054897320295348555512147739035918080361846620899758460525425686313546548745231723382816212278444549691507401383651812887;
            6'd45: xpb[190] = 1024'd97682874827140616753438340266987708434156534045491825905285737698493850625108984910088110690367526460094280046575726538984404520977039178246578267182120058789286384407349040165574596995650146403928688696433223804918973001420722709843536279143352202489772956309612503122765774754156519082966463271116735435415;
            6'd46: xpb[190] = 1024'd86068416969507659192537089227941387205504631788087679355610770195685170045965946918088394126302618791491580780115465636008606416905282233923706659228797055547527117997559994687295117018718237910537082044310935462098910084761083573066172799826178979293232366070479774522148733296034593616241419140849819057943;
            6'd47: xpb[190] = 1024'd74453959111874701631635838188895065976852729530683532805935802692876489466822908926088677562237711122888881513655204733032808312833525289600835051275474052305767851587770949209015637041786329417145475392188647119278847168101444436288809320509005756096691775831347045921531691837912668149516375010582902680471;
            6'd48: xpb[190] = 1024'd62839501254241744070734587149848744748200827273279386256260835190067808887679870934088960998172803454286182247194943830057010208761768345277963443322151049064008585177981903730736157064854420923753868740066358776458784251441805299511445841191832532900151185592214317320914650379790742682791330880315986302999;
            6'd49: xpb[190] = 1024'd51225043396608786509833336110802423519548925015875239706585867687259128308536832942089244434107895785683482980734682927081212104690011400955091835368828045822249318768192858252456677087922512430362262087944070433638721334782166162734082361874659309703610595353081588720297608921668817216066286750049069925527;
            6'd50: xpb[190] = 1024'd39610585538975828948932085071756102290897022758471093156910900184450447729393794950089527870042988117080783714274422024105414000618254456632220227415505042580490052358403812774177197110990603936970655435821782090818658418122527025956718882557486086507070005113948860119680567463546891749341242619782153548055;
            6'd51: xpb[190] = 1024'd27996127681342871388030834032709781062245120501066946607235932681641767150250756958089811305978080448478084447814161121129615896546497512309348619462182039338730785948614767295897717134058695443579048783699493747998595501462887889179355403240312863310529414874816131519063526005424966282616198489515237170583;
            6'd52: xpb[190] = 1024'd16381669823709913827129582993663459833593218243662800057560965178833086571107718966090094741913172779875385181353900218153817792474740567986477011508859036096971519538825721817618237157126786950187442131577205405178532584803248752401991923923139640113988824635683402918446484547303040815891154359248320793111;
            6'd53: xpb[190] = 1024'd4767211966076956266228331954617138604941315986258653507885997676024405991964680974090378177848265111272685914893639315178019688402983623663605403555536032855212253129036676339338757180194878456795835479454917062358469668143609615624628444605966416917448234396550674317829443089181115349166110228981404415639;
            6'd54: xpb[190] = 1024'd117219449792568740104126008320385250120987840854590191086342885238192620750130781892105732828441031752113136055890871846781285425172447013895893920618544070547143661288818848198689516394780175684714426435719868565902767601704867251812243534972022642987727547571535003747318929704987822899559755925340082522498;
            6'd55: xpb[190] = 1024'd105604991934935782543224757281338928892335938597186044536667917735383940170987743900106016264376124083510436789430610943805487321100690069573022312665221067305384394879029802720410036417848267191322819783597580223082704685045228115034880055654849419791186957332402275146701888246865897432834711795073166145026;
            6'd56: xpb[190] = 1024'd93990534077302824982323506242292607663684036339781897986992950232575259591844705908106299700311216414907737522970350040829689217028933125250150704711898064063625128469240757242130556440916358697931213131475291880262641768385588978257516576337676196594646367093269546546084846788743971966109667664806249767554;
            6'd57: xpb[190] = 1024'd82376076219669867421422255203246286435032134082377751437317982729766579012701667916106583136246308746305038256510089137853891112957176180927279096758575060821865862059451711763851076463984450204539606479353003537442578851725949841480153097020502973398105776854136817945467805330622046499384623534539333390082;
            6'd58: xpb[190] = 1024'd70761618362036909860521004164199965206380231824973604887643015226957898433558629924106866572181401077702338990049828234878093008885419236604407488805252057580106595649662666285571596487052541711147999827230715194622515935066310704702789617703329750201565186615004089344850763872500121032659579404272417012610;
            6'd59: xpb[190] = 1024'd59147160504403952299619753125153643977728329567569458337968047724149217854415591932107150008116493409099639723589567331902294904813662292281535880851929054338347329239873620807292116510120633217756393175108426851802453018406671567925426138386156527005024596375871360744233722414378195565934535274005500635138;
            6'd60: xpb[190] = 1024'd47532702646770994738718502086107322749076427310165311788293080221340537275272553940107433444051585740496940457129306428926496800741905347958664272898606051096588062830084575329012636533188724724364786522986138508982390101747032431148062659068983303808484006136738632143616680956256270099209491143738584257666;
            6'd61: xpb[190] = 1024'd35918244789138037177817251047061001520424525052761165238618112718531856696129515948107716879986678071894241190669045525950698696670148403635792664945283047854828796420295529850733156556256816230973179870863850166162327185087393294370699179751810080611943415897605903542999639498134344632484447013471667880194;
            6'd62: xpb[190] = 1024'd24303786931505079616916000008014680291772622795357018688943145215723176116986477956108000315921770403291541924208784622974900592598391459312921056991960044613069530010506484372453676579324907737581573218741561823342264268427754157593335700434636857415402825658473174942382598040012419165759402883204751502722;
            6'd63: xpb[190] = 1024'd12689329073872122056014748968968359063120720537952872139268177712914495537843439964108283751856862734688842657748523719999102488526634514990049449038637041371310263600717438894174196602392999244189966566619273480522201351768115020815972221117463634218862235419340446341765556581890493699034358752937835125250;
        endcase
    end

    always_comb begin
        case(flag[63][16:12])
            5'd0: xpb[191] = 1024'd0;
            5'd1: xpb[191] = 1024'd1074871216239164495113497929922037834468818280548725589593210210105814958700401972108567187791955066086143391288262817023304384454877570667177841085314038129550997190928393415894716625461090750798359914496985137702138435108475884038608741800290411022321645180207717741148515123768568232309314622670918747778;
            5'd2: xpb[191] = 1024'd2149742432478328990226995859844075668937636561097451179186420420211629917400803944217134375583910132172286782576525634046608768909755141334355682170628076259101994381856786831789433250922181501596719828993970275404276870216951768077217483600580822044643290360415435482297030247537136464618629245341837495556;
            5'd3: xpb[191] = 1024'd3224613648717493485340493789766113503406454841646176768779630630317444876101205916325701563375865198258430173864788451069913153364632712001533523255942114388652991572785180247684149876383272252395079743490955413106415305325427652115826225400871233066964935540623153223445545371305704696927943868012756243334;
            5'd4: xpb[191] = 1024'd4299484864956657980453991719688151337875273122194902358372840840423259834801607888434268751167820264344573565153051268093217537819510282668711364341256152518203988763713573663578866501844363003193439657987940550808553740433903536154434967201161644089286580720830870964594060495074272929237258490683674991112;
            5'd5: xpb[191] = 1024'd5374356081195822475567489649610189172344091402743627947966051050529074793502009860542835938959775330430716956441314085116521922274387853335889205426570190647754985954641967079473583127305453753991799572484925688510692175542379420193043709001452055111608225901038588705742575618842841161546573113354593738890;
            5'd6: xpb[191] = 1024'd6449227297434986970680987579532227006812909683292353537559261260634889752202411832651403126751730396516860347729576902139826306729265424003067046511884228777305983145570360495368299752766544504790159486981910826212830610650855304231652450801742466133929871081246306446891090742611409393855887736025512486668;
            5'd7: xpb[191] = 1024'd7524098513674151465794485509454264841281727963841079127152471470740704710902813804759970314543685462603003739017839719163130691184142994670244887597198266906856980336498753911263016378227635255588519401478895963914969045759331188270261192602032877156251516261454024188039605866379977626165202358696431234446;
            5'd8: xpb[191] = 1024'd8598969729913315960907983439376302675750546244389804716745681680846519669603215776868537502335640528689147130306102536186435075639020565337422728682512305036407977527427147327157733003688726006386879315975881101617107480867807072308869934402323288178573161441661741929188120990148545858474516981367349982224;
            5'd9: xpb[191] = 1024'd9673840946152480456021481369298340510219364524938530306338891890952334628303617748977104690127595594775290521594365353209739460093898136004600569767826343165958974718355540743052449629149816757185239230472866239319245915976282956347478676202613699200894806621869459670336636113917114090783831604038268730002;
            5'd10: xpb[191] = 1024'd10748712162391644951134979299220378344688182805487255895932102101058149587004019721085671877919550660861433912882628170233043844548775706671778410853140381295509971909283934158947166254610907507983599144969851377021384351084758840386087418002904110223216451802077177411485151237685682323093146226709187477780;
            5'd11: xpb[191] = 1024'd11823583378630809446248477229142416179157001086035981485525312311163964545704421693194239065711505726947577304170890987256348229003653277338956251938454419425060969100212327574841882880071998258781959059466836514723522786193234724424696159803194521245538096982284895152633666361454250555402460849380106225558;
            5'd12: xpb[191] = 1024'd12898454594869973941361975159064454013625819366584707075118522521269779504404823665302806253503460793033720695459153804279652613458530848006134093023768457554611966291140720990736599505533089009580318973963821652425661221301710608463304901603484932267859742162492612893782181485222818787711775472051024973336;
            5'd13: xpb[191] = 1024'd13973325811109138436475473088986491848094637647133432664711732731375594463105225637411373441295415859119864086747416621302956997913408418673311934109082495684162963482069114406631316130994179760378678888460806790127799656410186492501913643403775343290181387342700330634930696608991387020021090094721943721114;
            5'd14: xpb[191] = 1024'd15048197027348302931588971018908529682563455927682158254304942941481409421805627609519940629087370925206007478035679438326261382368285989340489775194396533813713960672997507822526032756455270511177038802957791927829938091518662376540522385204065754312503032522908048376079211732759955252330404717392862468892;
            5'd15: xpb[191] = 1024'd16123068243587467426702468948830567517032274208230883843898153151587224380506029581628507816879325991292150869323942255349565766823163560007667616279710571943264957863925901238420749381916361261975398717454777065532076526627138260579131127004356165334824677703115766117227726856528523484639719340063781216670;
            5'd16: xpb[191] = 1024'd17197939459826631921815966878752605351501092488779609433491363361693039339206431553737075004671281057378294260612205072372870151278041130674845457365024610072815955054854294654315466007377452012773758631951762203234214961735614144617739868804646576357146322883323483858376241980297091716949033962734699964448;
            5'd17: xpb[191] = 1024'd18272810676065796416929464808674643185969910769328335023084573571798854297906833525845642192463236123464437651900467889396174535732918701342023298450338648202366952245782688070210182632838542763572118546448747340936353396844090028656348610604936987379467968063531201599524757104065659949258348585405618712226;
            5'd18: xpb[191] = 1024'd19347681892304960912042962738596681020438729049877060612677783781904669256607235497954209380255191189550581043188730706419478920187796272009201139535652686331917949436711081486104899258299633514370478460945732478638491831952565912694957352405227398401789613243738919340673272227834228181567663208076537460004;
            5'd19: xpb[191] = 1024'd20422553108544125407156460668518718854907547330425786202270993992010484215307637470062776568047146255636724434476993523442783304642673842676378980620966724461468946627639474901999615883760724265168838375442717616340630267061041796733566094205517809424111258423946637081821787351602796413876977830747456207782;
            5'd20: xpb[191] = 1024'd21497424324783289902269958598440756689376365610974511791864204202116299174008039442171343755839101321722867825765256340466087689097551413343556821706280762591019943818567868317894332509221815015967198289939702754042768702169517680772174836005808220446432903604154354822970302475371364646186292453418374955560;
            5'd21: xpb[191] = 1024'd22572295541022454397383456528362794523845183891523237381457414412222114132708441414279910943631056387809011217053519157489392073552428984010734662791594800720570941009496261733789049134682905766765558204436687891744907137277993564810783577806098631468754548784362072564118817599139932878495607076089293703338;
            5'd22: xpb[191] = 1024'd23647166757261618892496954458284832358314002172071962971050624622327929091408843386388478131423011453895154608341781974512696458007306554677912503876908838850121938200424655149683765760143996517563918118933673029447045572386469448849392319606389042491076193964569790305267332722908501110804921698760212451116;
            5'd23: xpb[191] = 1024'd24722037973500783387610452388206870192782820452620688560643834832433744050109245358497045319214966519981297999630044791536000842462184125345090344962222876979672935391353048565578482385605087268362278033430658167149184007494945332888001061406679453513397839144777508046415847846677069343114236321431131198894;
            5'd24: xpb[191] = 1024'd25796909189739947882723950318128908027251638733169414150237045042539559008809647330605612507006921586067441390918307608559305226917061696012268186047536915109223932582281441981473199011066178019160637947927643304851322442603421216926609803206969864535719484324985225787564362970445637575423550944102049946672;
            5'd25: xpb[191] = 1024'd26871780405979112377837448248050945861720457013718139739830255252645373967510049302714179694798876652153584782206570425582609611371939266679446027132850953238774929773209835397367915636527268769958997862424628442553460877711897100965218545007260275558041129505192943528712878094214205807732865566772968694450;
            5'd26: xpb[191] = 1024'd27946651622218276872950946177972983696189275294266865329423465462751188926210451274822746882590831718239728173494833242605913995826816837346623868218164991368325926964138228813262632261988359520757357776921613580255599312820372985003827286807550686580362774685400661269861393217982774040042180189443887442228;
            5'd27: xpb[191] = 1024'd29021522838457441368064444107895021530658093574815590919016675672857003884910853246931314070382786784325871564783096059629218380281694408013801709303479029497876924155066622229157348887449450271555717691418598717957737747928848869042436028607841097602684419865608379011009908341751342272351494812114806190006;
            5'd28: xpb[191] = 1024'd30096394054696605863177942037817059365126911855364316508609885882962818843611255219039881258174741850412014956071358876652522764736571978680979550388793067627427921345995015645052065512910541022354077605915583855659876183037324753081044770408131508625006065045816096752158423465519910504660809434785724937784;
            5'd29: xpb[191] = 1024'd31171265270935770358291439967739097199595730135913042098203096093068633802311657191148448445966696916498158347359621693675827149191449549348157391474107105756978918536923409060946782138371631773152437520412568993362014618145800637119653512208421919647327710226023814493306938589288478736970124057456643685562;
            5'd30: xpb[191] = 1024'd32246136487174934853404937897661135034064548416461767687796306303174448761012059163257015633758651982584301738647884510699131533646327120015335232559421143886529915727851802476841498763832722523950797434909554131064153053254276521158262254008712330669649355406231532234455453713057046969279438680127562433340;
            5'd31: xpb[191] = 1024'd33321007703414099348518435827583172868533366697010493277389516513280263719712461135365582821550607048670445129936147327722435918101204690682513073644735182016080912918780195892736215389293813274749157349406539268766291488362752405196870995809002741691971000586439249975603968836825615201588753302798481181118;
        endcase
    end

    always_comb begin
        case(flag[64][5:0])
            6'd0: xpb[192] = 1024'd0;
            6'd1: xpb[192] = 1024'd17197939459826631921815966878752605351501092488779609433491363361693039339206431553737075004671281057378294260612205072372870151278041130674845457365024610072815955054854294654315466007377452012773758631951762203234214961735614144617739868804646576357146322883323483858376241980297091716949033962734699964448;
            6'd2: xpb[192] = 1024'd34395878919653263843631933757505210703002184977559218866982726723386078678412863107474150009342562114756588521224410144745740302556082261349690914730049220145631910109708589308630932014754904025547517263903524406468429923471228289235479737609293152714292645766646967716752483960594183433898067925469399928896;
            6'd3: xpb[192] = 1024'd51593818379479895765447900636257816054503277466338828300474090085079118017619294661211225014013843172134882781836615217118610453834123392024536372095073830218447865164562883962946398022132356038321275895855286609702644885206842433853219606413939729071438968649970451575128725940891275150847101888204099893344;
            6'd4: xpb[192] = 1024'd68791757839306527687263867515010421406004369955118437733965453446772157356825726214948300018685124229513177042448820289491480605112164522699381829460098440291263820219417178617261864029509808051095034527807048812936859846942456578470959475218586305428585291533293935433504967921188366867796135850938799857792;
            6'd5: xpb[192] = 1024'd85989697299133159609079834393763026757505462443898047167456816808465196696032157768685375023356405286891471303061025361864350756390205653374227286825123050364079775274271473271577330036887260063868793159758811016171074808678070723088699344023232881785731614416617419291881209901485458584745169813673499822240;
            6'd6: xpb[192] = 1024'd103187636758959791530895801272515632109006554932677656600948180170158236035238589322422450028027686344269765563673230434237220907668246784049072744190147660436895730329125767925892796044264712076642551791710573219405289770413684867706439212827879458142877937299940903150257451881782550301694203776408199786688;
            6'd7: xpb[192] = 1024'd120385576218786423452711768151268237460507647421457266034439543531851275374445020876159525032698967401648059824285435506610091058946287914723918201555172270509711685383980062580208262051642164089416310423662335422639504732149299012324179081632526034500024260183264387008633693862079642018643237739142899751136;
            6'd8: xpb[192] = 1024'd13516819994488313975728807625206410067310312784501191339799051828567419376342313519881528822712574149583204677440147144403897369383108710843603533903865839648836965869263139896893488867502410380879871447226857779509358843664016383976940380753943161590350679652470812836903407768448100718473581875252005231253;
            6'd9: xpb[192] = 1024'd30714759454314945897544774503959015418811405273280800773290415190260458715548745073618603827383855206961498938052352216776767520661149841518448991268890449721652920924117434551208954874879862393653630079178619982743573805399630528594680249558589737947497002535794296695279649748745192435422615837986705195701;
            6'd10: xpb[192] = 1024'd47912698914141577819360741382711620770312497762060410206781778551953498054755176627355678832055136264339793198664557289149637671939190972193294448633915059794468875978971729205524420882257314406427388711130382185977788767135244673212420118363236314304643325419117780553655891729042284152371649800721405160149;
            6'd11: xpb[192] = 1024'd65110638373968209741176708261464226121813590250840019640273141913646537393961608181092753836726417321718087459276762361522507823217232102868139905998939669867284831033826023859839886889634766419201147343082144389212003728870858817830159987167882890661789648302441264412032133709339375869320683763456105124597;
            6'd12: xpb[192] = 1024'd82308577833794841662992675140216831473314682739619629073764505275339576733168039734829828841397698379096381719888967433895377974495273233542985363363964279940100786088680318514155352897012218431974905975033906592446218690606472962447899855972529467018935971185764748270408375689636467586269717726190805089045;
            6'd13: xpb[192] = 1024'd99506517293621473584808642018969436824815775228399238507255868637032616072374471288566903846068979436474675980501172506268248125773314364217830820728988890012916741143534613168470818904389670444748664606985668795680433652342087107065639724777176043376082294069088232128784617669933559303218751688925505053493;
            6'd14: xpb[192] = 1024'd116704456753448105506624608897722042176316867717178847940747231998725655411580902842303978850740260493852970241113377578641118277051355494892676278094013500085732696198388907822786284911767122457522423238937430998914648614077701251683379593581822619733228616952411715987160859650230651020167785651660205017941;
            6'd15: xpb[192] = 1024'd9835700529149996029641648371660214783119533080222773246106740295441799413478195486025982640753867241788115094268089216434924587488176291012361610442707069224857976683671985139471511727627368748985984262501953355784502725592418623336140892703239746823555036421618141815430573556599109719998129787769310498058;
            6'd16: xpb[192] = 1024'd27033639988976627951457615250412820134620625569002382679598103657134838752684627039763057645425148299166409354880294288807794738766217421687207067807731679297673931738526279793786977735004820761759742894453715559018717687328032767953880761507886323180701359304941625673806815536896201436947163750504010462506;
            6'd17: xpb[192] = 1024'd44231579448803259873273582129165425486121718057781992113089467018827878091891058593500132650096429356544703615492499361180664890044258552362052525172756289370489886793380574448102443742382272774533501526405477762252932649063646912571620630312532899537847682188265109532183057517193293153896197713238710426954;
            6'd18: xpb[192] = 1024'd61429518908629891795089549007918030837622810546561601546580830380520917431097490147237207654767710413922997876104704433553535041322299683036897982537780899443305841848234869102417909749759724787307260158357239965487147610799261057189360499117179475894994005071588593390559299497490384870845231675973410391402;
            6'd19: xpb[192] = 1024'd78627458368456523716905515886670636189123903035341210980072193742213956770303921700974282659438991471301292136716909505926405192600340813711743439902805509516121796903089163756733375757137176800081018790309002168721362572534875201807100367921826052252140327954912077248935541477787476587794265638708110355850;
            6'd20: xpb[192] = 1024'd95825397828283155638721482765423241540624995524120820413563557103906996109510353254711357664110272528679586397329114578299275343878381944386588897267830119588937751957943458411048841764514628812854777422260764371955577534270489346424840236726472628609286650838235561107311783458084568304743299601442810320298;
            6'd21: xpb[192] = 1024'd113023337288109787560537449644175846892126088012900429847054920465600035448716784808448432668781553586057880657941319650672145495156423075061434354632854729661753707012797753065364307771892080825628536054212526575189792496006103491042580105531119204966432973721559044965688025438381660021692333564177510284746;
            6'd22: xpb[192] = 1024'd6154581063811678083554489118114019498928753375944355152414428762316179450614077452170436458795160333993025511096031288465951805593243871181119686981548298800878987498080830382049534587752327117092097077777048932059646607520820862695341404652536332056759393190765470793957739344750118721522677700286615764863;
            6'd23: xpb[192] = 1024'd23352520523638310005370455996866624850429845864723964585905792124009218789820509005907511463466441391371319771708236360838821956871285001855965144346572908873694942552935125036365000595129779129865855709728811135293861569256435007313081273457182908413905716074088954652333981325047210438471711663021315729311;
            6'd24: xpb[192] = 1024'd40550459983464941927186422875619230201930938353503574019397155485702258129026940559644586468137722448749614032320441433211692108149326132530810601711597518946510897607789419690680466602507231142639614341680573338528076530992049151930821142261829484771052038957412438510710223305344302155420745625756015693759;
            6'd25: xpb[192] = 1024'd57748399443291573849002389754371835553432030842283183452888518847395297468233372113381661472809003506127908292932646505584562259427367263205656059076622129019326852662643714344995932609884683155413372973632335541762291492727663296548561011066476061128198361840735922369086465285641393872369779588490715658207;
            6'd26: xpb[192] = 1024'd74946338903118205770818356633124440904933123331062792886379882209088336807439803667118736477480284563506202553544851577957432410705408393880501516441646739092142807717498008999311398617262135168187131605584097744996506454463277441166300879871122637485344684724059406227462707265938485589318813551225415622655;
            6'd27: xpb[192] = 1024'd92144278362944837692634323511877046256434215819842402319871245570781376146646235220855811482151565620884496814157056650330302561983449524555346973806671349164958762772352303653626864624639587180960890237535859948230721416198891585784040748675769213842491007607382890085838949246235577306267847513960115587103;
            6'd28: xpb[192] = 1024'd109342217822771469614450290390629651607935308308622011753362608932474415485852666774592886486822846678262791074769261722703172713261490655230192431171695959237774717827206598307942330632017039193734648869487622151464936377934505730401780617480415790199637330490706373944215191226532669023216881476694815551551;
            6'd29: xpb[192] = 1024'd2473461598473360137467329864567824214737973671665937058722117229190559487749959418314890276836453426197935927923973360496979023698311451349877763520389528376899998312489675624627557447877285485198209893052144508334790489449223102054541916601832917289963749959912799772484905132901127723047225612803921031668;
            6'd30: xpb[192] = 1024'd19671401058299992059283296743320429566239066160445546492213480590883598826956390972051965281507734483576230188536178432869849174976352582024723220885414138449715953367343970278943023455254737497971968525003906711569005451184837246672281785406479493647110072843236283630861147113198219439996259575538620996116;
            6'd31: xpb[192] = 1024'd36869340518126623981099263622073034917740158649225155925704843952576638166162822525789040286179015540954524449148383505242719326254393712699568678250438748522531908422198264933258489462632189510745727156955668914803220412920451391290021654211126070004256395726559767489237389093495311156945293538273320960564;
            6'd32: xpb[192] = 1024'd54067279977953255902915230500825640269241251138004765359196207314269677505369254079526115290850296598332818709760588577615589477532434843374414135615463358595347863477052559587573955470009641523519485788907431118037435374656065535907761523015772646361402718609883251347613631073792402873894327501008020925012;
            6'd33: xpb[192] = 1024'd71265219437779887824731197379578245620742343626784374792687570675962716844575685633263190295521577655711112970372793649988459628810475974049259592980487968668163818531906854241889421477387093536293244420859193321271650336391679680525501391820419222718549041493206735205989873054089494590843361463742720889460;
            6'd34: xpb[192] = 1024'd88463158897606519746547164258330850972243436115563984226178934037655756183782117187000265300192858713089407230984998722361329780088517104724105050345512578740979773586761148896204887484764545549067003052810955524505865298127293825143241260625065799075695364376530219064366115034386586307792395426477420853908;
            6'd35: xpb[192] = 1024'd105661098357433151668363131137083456323744528604343593659670297399348795522988548740737340304864139770467701491597203794734199931366558235398950507710537188813795728641615443550520353492141997561840761684762717727740080259862907969760981129429712375432841687259853702922742357014683678024741429389212120818356;
            6'd36: xpb[192] = 1024'd122859037817259783590179098015836061675245621093123203093161660761041834862194980294474415309535420827845995752209408867107070082644599366073795965075561798886611683696469738204835819499519449574614520316714479930974295221598522114378720998234358951789988010143177186781118598994980769741690463351946820782804;
            6'd37: xpb[192] = 1024'd15990281592961674113196137489774234282048286456167128398521169057757978864092272938196419099549027575781140605364120504900876393081420162193481297424255368025736964181752815521521046315379695866078081340279002287844149333113239486031482297355776078880314429612383612609388312901349228441520807488055926262921;
            6'd38: xpb[192] = 1024'd33188221052788306035012104368526839633549378944946737832012532419451018203298704491933494104220308633159434865976325577273746544359461292868326754789279978098552919236607110175836512322757147878851839972230764491078364294848853630649222166160422655237460752495707096467764554881646320158469841450790626227369;
            6'd39: xpb[192] = 1024'd50386160512614937956828071247279444985050471433726347265503895781144057542505136045670569108891589690537729126588530649646616695637502423543172212154304588171368874291461404830151978330134599891625598604182526694312579256584467775266962034965069231594607075379030580326140796861943411875418875413525326191817;
            6'd40: xpb[192] = 1024'd67584099972441569878644038126032050336551563922505956698995259142837096881711567599407644113562870747916023387200735722019486846915543554218017669519329198244184829346315699484467444337512051904399357236134288897546794218320081919884701903769715807951753398262354064184517038842240503592367909376260026156265;
            6'd41: xpb[192] = 1024'd84782039432268201800460005004784655688052656411285566132486622504530136220917999153144719118234151805294317647812940794392356998193584684892863126884353808317000784401169994138782910344889503917173115868086051100781009180055696064502441772574362384308899721145677548042893280822537595309316943338994726120713;
            6'd42: xpb[192] = 1024'd101979978892094833722275971883537261039553748900065175565977985866223175560124430706881794122905432862672611908425145866765227149471625815567708584249378418389816739456024288793098376352266955929946874500037813304015224141791310209120181641379008960666046044029001031901269522802834687026265977301729426085161;
            6'd43: xpb[192] = 1024'd119177918351921465644091938762289866391054841388844784999469349227916214899330862260618869127576713920050906169037350939138097300749666946242554041614403028462632694510878583447413842359644407942720633131989575507249439103526924353737921510183655537023192366912324515759645764783131778743215011264464126049609;
            6'd44: xpb[192] = 1024'd12309162127623356167108978236228038997857506751888710304828857524632358901228154904340872917590320667986051022192062576931903611186487742362239373963096597601757974996161660764099069175504654234184194155554097864119293215041641725390682809305072664113518786381530941587915478689500237443045355400573231529726;
            6'd45: xpb[192] = 1024'd29507101587449988088924945114980644349358599240668319738320220886325398240434586458077947922261601725364345282804267649304773762464528873037084831328121207674573930051015955418414535182882106246957952787505860067353508176777255870008422678109719240470665109264854425446291720669797329159994389363307931494174;
            6'd46: xpb[192] = 1024'd46705041047276620010740911993733249700859691729447929171811584248018437579641018011815022926932882782742639543416472721677643913742570003711930288693145817747389885105870250072730001190259558259731711419457622270587723138512870014626162546914365816827811432148177909304667962650094420876943423326042631458622;
            6'd47: xpb[192] = 1024'd63902980507103251932556878872485855052360784218227538605302947609711476918847449565552097931604163840120933804028677794050514065020611134386775746058170427820205840160724544727045467197637010272505470051409384473821938100248484159243902415719012393184957755031501393163044204630391512593892457288777331423070;
            6'd48: xpb[192] = 1024'd81100919966929883854372845751238460403861876707007148038794310971404516258053881119289172936275444897499228064640882866423384216298652265061621203423195037893021795215578839381360933205014462285279228683361146677056153061984098303861642284523658969542104077914824877021420446610688604310841491251512031387518;
            6'd49: xpb[192] = 1024'd98298859426756515776188812629991065755362969195786757472285674333097555597260312673026247940946725954877522325253087938796254367576693395736466660788219647965837750270433134035676399212391914298052987315312908880290368023719712448479382153328305545899250400798148360879796688590985696027790525214246731351966;
            6'd50: xpb[192] = 1024'd115496798886583147698004779508743671106864061684566366905777037694790594936466744226763322945618007012255816585865293011169124518854734526411312118153244258038653705325287428689991865219769366310826745947264671083524582985455326593097122022132952122256396723681471844738172930571282787744739559176981431316414;
            6'd51: xpb[192] = 1024'd8628042662285038221021818982681843713666727047610292211136545991506738938364036870485326735631613760190961439020004648962930829291555322530997450501937827177778985810570506006677092035629612602290306970829193440394437096970043964749883321254369249346723143150678270566442644477651246444569903313090536796531;
            6'd52: xpb[192] = 1024'd25825982122111670142837785861434449065167819536389901644627909353199778277570468424222401740302894817569255699632209721335800980569596453205842907866962437250594940865424800660992558043007064615064065602780955643628652058705658109367623190059015825703869466034001754424818886457948338161518937275825236760979;
            6'd53: xpb[192] = 1024'd43023921581938302064653752740187054416668912025169511078119272714892817616776899977959476744974175874947549960244414793708671131847637583880688365231987047323410895920279095315308024050384516627837824234732717846862867020441272253985363058863662402061015788917325238283195128438245429878467971238559936725427;
            6'd54: xpb[192] = 1024'd60221861041764933986469719618939659768170004513949120511610636076585856955983331531696551749645456932325844220856619866081541283125678714555533822597011657396226850975133389969623490057761968640611582866684480050097081982176886398603102927668308978418162111800648722141571370418542521595417005201294636689875;
            6'd55: xpb[192] = 1024'd77419800501591565908285686497692265119671097002728729945101999438278896295189763085433626754316737989704138481468824938454411434403719845230379279962036267469042806029987684623938956065139420653385341498636242253331296943912500543220842796472955554775308434683972205999947612398839613312366039164029336654323;
            6'd56: xpb[192] = 1024'd94617739961418197830101653376444870471172189491508339378593362799971935634396194639170701758988019047082432742081030010827281585681760975905224737327060877541858761084841979278254422072516872666159100130588004456565511905648114687838582665277602131132454757567295689858323854379136705029315073126764036618771;
            6'd57: xpb[192] = 1024'd111815679421244829751917620255197475822673281980287948812084726161664974973602626192907776763659300104460727002693235083200151736959802106580070194692085487614674716139696273932569888079894324678932858762539766659799726867383728832456322534082248707489601080450619173716700096359433796746264107089498736583219;
            6'd58: xpb[192] = 1024'd4946923196946720274934659729135648429475947343331874117444234458381118975499918836629780553672906852395871855847946720993958047396622902699755527040779056753799996624979351249255114895754570970396419786104289016669580978898446204109083833203665834579927499919825599544969810265802255446094451225607842063336;
            6'd59: xpb[192] = 1024'd22144862656773352196750626607888253780977039832111483550935597820074158314706350390366855558344187909774166116460151793366828198674664033374600984405803666826615951679833645903570580903132022983170178418056051219903795940634060348726823702008312410937073822803149083403346052246099347163043485188342542027784;
            6'd60: xpb[192] = 1024'd39342802116599984118566593486640859132478132320891092984426961181767197653912781944103930563015468967152460377072356865739698349952705164049446441770828276899431906734687940557886046910509474995943937050007813423138010902369674493344563570812958987294220145686472567261722294226396438879992519151077241992232;
            6'd61: xpb[192] = 1024'd56540741576426616040382560365393464483979224809670702417918324543460236993119213497841005567686750024530754637684561938112568501230746294724291899135852886972247861789542235212201512917886927008717695681959575626372225864105288637962303439617605563651366468569796051120098536206693530596941553113811941956680;
            6'd62: xpb[192] = 1024'd73738681036253247962198527244146069835480317298450311851409687905153276332325645051578080572358031081909048898296767010485438652508787425399137356500877497045063816844396529866516978925264379021491454313911337829606440825840902782580043308422252140008512791453119534978474778186990622313890587076546641921128;
            6'd63: xpb[192] = 1024'd90936620496079879884014494122898675186981409787229921284901051266846315671532076605315155577029312139287343158908972082858308803786828556073982813865902107117879771899250824520832444932641831034265212945863100032840655787576516927197783177226898716365659114336443018836851020167287714030839621039281341885576;
        endcase
    end

    always_comb begin
        case(flag[64][11:6])
            6'd0: xpb[193] = 1024'd0;
            6'd1: xpb[193] = 1024'd108134559955906511805830461001651280538482502276009530718392414628539355010738508159052230581700593196665637419521177155231178955064869686748828271230926717190695726954105119175147910940019283047038971577814862236074870749312131071815523046031545292722805437219766502695227262147584805747788655002016041850024;
            6'd2: xpb[193] = 1024'd92202424227688282212861994598488128332266577426283377308652974192101814684167877408089389948743512083888125431584860875883294069288519038942496417445522393447700779338639021012665582688521360372767745547242484625785380648403365370666067522379861136178790971025415947360347996221240978478458620177406489215717;
            6'd3: xpb[193] = 1024'd76270288499470052619893528195324976126050652576557223898913533755664274357597246657126549315786430971110613443648544596535409183512168391136164563660118069704705831723172922850183254437023437698496519516670107015495890547494599669516611998728176979634776504831065392025468730294897151209128585352796936581410;
            6'd4: xpb[193] = 1024'd60338152771251823026925061792161823919834727726831070489174093319226734031026615906163708682829349858333101455712228317187524297735817743329832709874713745961710884107706824687700926185525515024225293486097729405206400446585833968367156475076492823090762038636714836690589464368553323939798550528187383947103;
            6'd5: xpb[193] = 1024'd44406017043033593433956595388998671713618802877104917079434652882789193704455985155200868049872268745555589467775912037839639411959467095523500856089309422218715936492240726525218597934027592349954067455525351794916910345677068267217700951424808666546747572442364281355710198442209496670468515703577831312796;
            6'd6: xpb[193] = 1024'd28473881314815363840988128985835519507402878027378763669695212446351653377885354404238027416915187632778077479839595758491754526183116447717169002303905098475720988876774628362736269682529669675682841424952974184627420244768302566068245427773124510002733106248013726020830932515865669401138480878968278678489;
            6'd7: xpb[193] = 1024'd12541745586597134248019662582672367301186953177652610259955772009914113051314723653275186783958106520000565491903279479143869640406765799910837148518500774732726041261308530200253941431031747001411615394380596574337930143859536864918789904121440353458718640053663170685951666589521842131808446054358726044182;
            6'd8: xpb[193] = 1024'd120676305542503646053850123584323647839669455453662140978348186638453468062053231812327417365658699716666202911424456634375048595471635486659665419749427491923421768215413649375401852371051030048450586972195458810412800893171667936734312950152985646181524077273429673381178928737106647879597101056374767894206;
            6'd9: xpb[193] = 1024'd104744169814285416460881657181160495633453530603935987568608746202015927735482601061364576732701618603888690923488140355027163709695284838853333565964023168180426820599947551212919524119553107374179360941623081200123310792262902235584857426501301489637509611079079118046299662810762820610267066231765215259899;
            6'd10: xpb[193] = 1024'd88812034086067186867913190777997343427237605754209834158869305765578387408911970310401736099744537491111178935551824075679278823918934191047001712178618844437431872984481453050437195868055184699908134911050703589833820691354136534435401902849617333093495144884728562711420396884418993340937031407155662625592;
            6'd11: xpb[193] = 1024'd72879898357848957274944724374834191221021680904483680749129865329140847082341339559438895466787456378333666947615507796331393938142583543240669858393214520694436925369015354887954867616557262025636908880478325979544330590445370833285946379197933176549480678690378007376541130958075166071606996582546109991285;
            6'd12: xpb[193] = 1024'd56947762629630727681976257971671039014805756054757527339390424892703306755770708808476054833830375265556154959679191516983509052366232895434338004607810196951441977753549256725472539365059339351365682849905948369254840489536605132136490855546249020005466212496027452041661865031731338802276961757936557356978;
            6'd13: xpb[193] = 1024'd41015626901412498089007791568507886808589831205031373929650984456265766429200078057513214200873294152778642971742875237635624166589882247628006150822405873208447030138083158562990211113561416677094456819333570758965350388627839430987035331894564863461451746301676896706782599105387511532946926933327004722671;
            6'd14: xpb[193] = 1024'd25083491173194268496039325165344734602373906355305220519911544019828226102629447306550373567916213040001130983806558958287739280813531599821674297037001549465452082522617060400507882862063494002823230788761193148675860287719073729837579808242880706917437280107326341371903333179043684263616892108717452088364;
            6'd15: xpb[193] = 1024'd9151355444976038903070858762181582396157981505579067110172103583390685776058816555587532934959131927223618995870242678939854395037180952015342443251597225722457134907150962238025554610565571328552004758188815538386370186810308028688124284591196550373422813912975786037024067252699856994286857284107899454057;
            6'd16: xpb[193] = 1024'd117285915400882550708901319763832862934640483781588597828564518211930040786797324714639763516659725123889256415391419834171033350102050638764170714482523942913152861861256081413173465550584854375590976336003677774461240936122439100503647330622741843096228251132742288732251329400284662742075512286123941304081;
            6'd17: xpb[193] = 1024'd101353779672664321115932853360669710728424558931862444418825077775492500460226693963676922883702644011111744427455103554823148464325699990957838860697119619170157914245789983250691137299086931701319750305431300164171750835213673399354191806971057686552213784938391733397372063473940835472745477461514388669774;
            6'd18: xpb[193] = 1024'd85421643944446091522964386957506558522208634082136291009085637339054960133656063212714082250745562898334232439518787275475263578549349343151507006911715295427162966630323885088208809047589009027048524274858922553882260734304907698204736283319373530008199318744041178062492797547597008203415442636904836035467;
            6'd19: xpb[193] = 1024'd69489508216227861929995920554343406315992709232410137599346196902617419807085432461751241617788481785556720451582470996127378692772998695345175153126310971684168019014857786925726480796091086352777298244286544943592770633396141997055280759667689373464184852549690622727613531621253180934085407812295283401160;
            6'd20: xpb[193] = 1024'd53557372488009632337027454151180254109776784382683984189606756466179879480514801710788400984831400672779208463646154716779493806996648047538843299340906647941173071399391688763244152544593163678506072213714167333303280532487376295905825236016005216920170386355340067392734265694909353664755372987685730766853;
            6'd21: xpb[193] = 1024'd37625236759791402744058987748017101903560859532957830779867316029742339153944170959825560351874319560001696475709838437431608921220297399732511445555502324198178123783925590600761824293095241004234846183141789723013790431578610594756369712364321060376155920160989512057854999768565526395425338163076178132546;
            6'd22: xpb[193] = 1024'd21693101031573173151090521344853949697344934683231677370127875593304798827373540208862719718917238447224184487773522158083724035443946751926179591770098000455183176168459492438279496041597318329963620152569412112724300330669844893606914188712636903832141453966638956722975733842221699126095303338466625498239;
            6'd23: xpb[193] = 1024'd5760965303354943558122054941690797491129009833505523960388435156867258500802909457899879085960157334446672499837205878735839149667596104119847737984693676712188228552993394275797167790099395655692394121997034502434810229761079192457458665060952747288126987772288401388096467915877871856765268513857072863932;
            6'd24: xpb[193] = 1024'd113895525259261455363952515943342078029611512109515054678780849785406613511541417616952109667660750531112309919358383033967018104732465790868676009215620393902883955507098513450945078730118678702731365699811896738509680979073210264272981711092498040010932424992054904083323730063462677604553923515873114713956;
            6'd25: xpb[193] = 1024'd97963389531043225770984049540178925823395587259788901269041409348969073184970786865989269034703669418334797931422066754619133218956115143062344155430216070159889007891632415288462750478620756028460139669239519128220190878164444563123526187440813883466917958797704348748444464137118850335223888691263562079649;
            6'd26: xpb[193] = 1024'd82031253802824996178015583137015773617179662410062747859301968912531532858400156115026428401746588305557285943485750475271248333179764495256012301644811746416894060276166317125980422227122833354188913638667141517930700777255678861974070663789129726922903492603353793413565198210775023065893853866654009445342;
            6'd27: xpb[193] = 1024'd66099118074606766585047116733852621410963737560336594449562528476093992531829525364063587768789507192779773955549434195923363447403413847449680447859407422673899112660700218963498093975624910679917687608094763907641210676346913160824615140137445570378889026409003238078685932284431195796563819042044456811035;
            6'd28: xpb[193] = 1024'd50166982346388536992078650330689469204747812710610441039823088039656452205258894613100747135832426080002261967613117916575478561627063199643348594074003098930904165045234120801015765724126988005646461577522386297351720575438147459675159616485761413834874560214652682743806666358087368527233784217434904176728;
            6'd29: xpb[193] = 1024'd34234846618170307399110183927526316998531887860884287630083647603218911878688263862137906502875344967224749979676801637227593675850712551837016740288598775187909217429768022638533437472629065331375235546950008687062230474529381758525704092834077257290860094020302127408927400431743541257903749392825351542421;
            6'd30: xpb[193] = 1024'd18302710889952077806141717524363164792315963011158134220344207166781371552117633111175065869918263854447237991740485357879708790074361904030684886503194451444914269814301924476051109221131142657104009516377631076772740373620616057376248569182393100746845627825951572074048134505399713988573714568215798908114;
            6'd31: xpb[193] = 1024'd2370575161733848213173251121200012586100038161431980810604766730343831225547002360212225236961182741669726003804169078531823904298011256224353032717790127701919322198835826313568780969633219982832783485805253466483250272711850356226793045530708944202831161631601016739168868579055886719243679743606246273807;
            6'd32: xpb[193] = 1024'd110505135117640360019003712122851293124582540437441511528997181358883186236285510519264455818661775938335363423325346233763002859362880942973181303948716844892615049152940945488716691909652503029871755063620115702558121022023981428042316091562254236925636598851367519434396130726640692467032334745622288123831;
            6'd33: xpb[193] = 1024'd94572999389422130426035245719688140918366615587715358119257740922445645909714879768301615185704694825557851435389029954415117973586530295166849450163312521149620101537474847326234363658154580355600529033047738092268630921115215726892860567910570080381622132657016964099516864800296865197702299921012735489524;
            6'd34: xpb[193] = 1024'd78640863661203900833066779316524988712150690737989204709518300486008105583144249017338774552747613712780339447452713675067233087810179647360517596377908197406625153922008749163752035406656657681329303002475360481979140820206450025743405044258885923837607666462666408764637598873953037928372265096403182855217;
            6'd35: xpb[193] = 1024'd62708727932985671240098312913361836505934765888263051299778860049570565256573618266375933919790532600002827459516397395719348202033828999554185742592503873663630206306542651001269707155158735007058076971902982871689650719297684324593949520607201767293593200268315853429758332947609210659042230271793630220910;
            6'd36: xpb[193] = 1024'd46776592204767441647129846510198684299718841038536897890039419613133024930002987515413093286833451487225315471580081116371463316257478351747853888807099549920635258691076552838787378903660812332786850941330605261400160618388918623444493996955517610749578734073965298094879067021265383389712195447184077586603;
            6'd37: xpb[193] = 1024'd30844456476549212054161380107035532093502916188810744480299979176695484603432356764450252653876370374447803483643764837023578430481127703941522035021695226177640311075610454676305050652162889658515624910758227651110670517480152922295038473303833454205564267879614742759999801094921556120382160622574524952296;
            6'd38: xpb[193] = 1024'd14912320748330982461192913703872379887286991339084591070560538740257944276861726013487412020919289261670291495707448557675693544704777056135190181236290902434645363460144356513822722400664966984244398880185850040821180416571387221145582949652149297661549801685264187425120535168577728851052125797964972317989;
            6'd39: xpb[193] = 1024'd123046880704237494267023374705523660425769493615094121788952953368797299287600234172539642602619882458335928915228625712906872499769646742884018452467217619625341090414249475688970633340684250031283370458000712276896051165883518292961105995683694590384355238905030690120347797316162534598840780799981014168013;
            6'd40: xpb[193] = 1024'd107114744976019264674054908302360508219553568765367968379213512932359758961029603421576801969662801345558416927292309433558987613993296095077686598681813295882346142798783377526488305089186327357012144427428334666606561064974752591811650472032010433840340772710680134785468531389818707329510745975371461533706;
            6'd41: xpb[193] = 1024'd91182609247801035081086441899197356013337643915641814969474072495922218634458972670613961336705720232780904939355993154211102728216945447271354744896408972139351195183317279364005976837688404682740918396855957056317070964065986890662194948380326277296326306516329579450589265463474880060180711150761908899399;
            6'd42: xpb[193] = 1024'd75250473519582805488117975496034203807121719065915661559734632059484678307888341919651120703748639120003392951419676874863217842440594799465022891111004648396356247567851181201523648586190482008469692366283579446027580863157221189512739424728642120752311840321979024115709999537131052790850676326152356265092;
            6'd43: xpb[193] = 1024'd59318337791364575895149509092871051600905794216189508149995191623047137981317711168688280070791558007225880963483360595515332956664244151658691037325600324653361299952385083039041320334692559334198466335711201835738090762248455488363283901076957964208297374127628468780830733610787225521520641501542803630785;
            6'd44: xpb[193] = 1024'd43386202063146346302181042689707899394689869366463354740255751186609597654747080417725439437834476894448368975547044316167448070887893503852359183540196000910366352336918984876558992083194636659927240305138824225448600661339689787213828377425273807664282907933277913445951467684443398252190606676933250996478;
            6'd45: xpb[193] = 1024'd27454066334928116709212576286544747188473944516737201330516310750172057328176449666762598804877395781670856987610728036819563185111542856046027329754791677167371404721452886714076663831696713985656014274566446615159110560430924086064372853773589651120268441738927358111072201758099570982860571852323698362171;
            6'd46: xpb[193] = 1024'd11521930606709887116244109883381594982258019667011047920776870313734517001605818915799758171920314668893344999674411757471678299335192208239695475969387353424376457105986788551594335580198791311384788243994069004869620459522158384914917330121905494576253975544576802776192935831755743713530537027714145727864;
            6'd47: xpb[193] = 1024'd119656490562616398922074570885032875520740521943020578639169284942273872012344327074851988753620907865558982419195588912702857254400061894988523747200314070615072184060091907726742246520218074358423759821808931240944491208834289456730440376153450787299059412764343305471420197979340549461319192029730187577888;
            6'd48: xpb[193] = 1024'd103724354834398169329106104481869723314524597093294425229429844505836331685773696323889148120663826752781470431259272633354972368623711247182191893414909746872077236444625809564259918268720151684152533791236553630655001107925523755580984852501766630755044946569992750136540932052996722191989157205120634943581;
            6'd49: xpb[193] = 1024'd87792219106179939736137638078706571108308672243568271819690404069398791359203065572926307487706745640003958443322956354007087482847360599375860039629505423129082288829159711401777590017222229009881307760664176020365511007016758054431529328850082474211030480375642194801661666126652894922659122380511082309274;
            6'd50: xpb[193] = 1024'd71860083377961710143169171675543418902092747393842118409950963632961251032632434821963466854749664527226446455386640074659202597071009951569528185844101099386087341213693613239295261765724306335610081730091798410076020906107992353282073805198398317667016014181291639466782400200309067653329087555901529674967;
            6'd51: xpb[193] = 1024'd55927947649743480550200705272380266695876822544115965000211523196523710706061804071000626221792583414448934467450323795311317711294659303763196332058696775643092393598227515076812933514226383661338855699519420799786530805199226652132618281546714161123001547986941084131903134273965240383999052731291977040660;
            6'd52: xpb[193] = 1024'd39995811921525250957232238869217114489660897694389811590472082760086170379491173320037785588835502301671422479514007515963432825518308655956864478273292451900097445982761416914330605262728460987067629668947043189497040704290460950983162757895030004578987081792590528797023868347621413114669017906682424406353;
            6'd53: xpb[193] = 1024'd24063676193307021364263772466053962283444972844663658180732642323648630052920542569074944955878421188893910491577691236615547939741958008150532624487888128157102498367295318751848277011230538312796403638374665579207550603381695249833707234243345848034972615598239973462144602421277585845338983082072871772046;
            6'd54: xpb[193] = 1024'd8131540465088791771295306062890810077229047994937504770993201887211089726349911818112104322921340076116398503641374957267663053965607360344200770702483804414107550751829220589365948759732615638525177607802287968918060502472929548684251710591661691490958149403889418127265336494933758576008948257463319137739;
            6'd55: xpb[193] = 1024'd116266100420995303577125767064542090615711550270947035489385616515750444737088419977164334904621933272782035923162552112498842009030477047093029041933410521604803277705934339764513859699751898685564149185617150204992931251785060620499774756623206984213763586623655920822492598642518564323797603259479360987763;
            6'd56: xpb[193] = 1024'd100333964692777073984157300661378938409495625421220882079646176079312904410517789226201494271664852160004523935226235833150957123254126399286697188148006197861808330090468241602031531448253976011292923155044772594703441150876294919350319232971522827669749120429305365487613332716174737054467568434869808353456;
            6'd57: xpb[193] = 1024'd84401828964558844391188834258215786203279700571494728669906735642875364083947158475238653638707771047227011947289919553803072237477775751480365334362601874118813382475002143439549203196756053337021697124472394984413951049967529218200863709319838671125734654234954810152734066789830909785137533610260255719149;
            6'd58: xpb[193] = 1024'd68469693236340614798220367855052633997063775721768575260167295206437823757376527724275813005750689934449499959353603274455187351701425103674033480577197550375818434859536045277066874945258130662750471093900017374124460949058763517051408185668154514581720188040604254817854800863487082515807498785650703084842;
            6'd59: xpb[193] = 1024'd52537557508122385205251901451889481790847850872042421850427854770000283430805896973312972372793608821671987971417286995107302465925074455867701626791793226632823487244069947114584546693760207988479245063327639763834970848149997815901952662016470358037705721846253699482975534937143255246477463961041150450535;
            6'd60: xpb[193] = 1024'd36605421779904155612283435048726329584631926022316268440688414333562743104235266222350131739836527708894475983480970715759417580148723808061369773006388902889828539628603848952102218442262285314208019032755262153545480747241232114752497138364786201493691255651903144148096269010799427977147429136431597816228;
            6'd61: xpb[193] = 1024'd20673286051685926019314968645563177378416001172590115030948973897125202777664635471387291106879446596116963995544654436411532694372373160255037919220984579146833592013137750789619890190764362639936793002182884543255990646332466413603041614713102044949676789457552588813217003084455600707817394311822045181921;
            6'd62: xpb[193] = 1024'd4741150323467696426346502242400025172200076322863961621209533460687662451094004720424450473922365483339452007608338157063647808596022512448706065435580255403838644397671652627137561939266439965665566971610506932966500545423700712453586091061417888405662323263202033478337737158111773438487359487212492547614;
            6'd63: xpb[193] = 1024'd112875710279374208232176963244051305710682578598873492339601948089227017461832512879476681055622958680005089427129515312294826763660892199197534336666506972594534371351776771802285472879285723012704538549425369169041371294735831784269109137092963181128467760482968536173564999305696579186276014489228534397638;
        endcase
    end

    always_comb begin
        case(flag[64][16:12])
            5'd0: xpb[194] = 1024'd0;
            5'd1: xpb[194] = 1024'd96943574551155978639208496840888153504466653749147338929862507652789477135261882128513840422665877567227577439193199032946941877884541551391202482881102648851539423736310673639803144627787800338433312518852991558751881193827066083119653613441279024584453294288617980838685733379352751916945979664618981763331;
            5'd2: xpb[194] = 1024'd69820453418187215879618066276961874264234880372558993731593160240602058933214625347012609630674080825012005470928904631314819914927862768227244840745874256769388172903050129941976050064058394955556427429318743271139401537433235393274328657199328599902086685163118903647264938684776870816773269502612369042331;
            5'd3: xpb[194] = 1024'd42697332285218453120027635713035595024003106995970648533323812828414640731167368565511378838682284082796433502664610229682697951971183985063287198610645864687236922069789586244148955500328989572679542339784494983526921881039404703429003700957378175219720076037619826455844143990200989716600559340605756321331;
            5'd4: xpb[194] = 1024'd15574211152249690360437205149109315783771333619382303335054465416227222529120111784010148046690487340580861534400315828050575989014505201899329556475417472605085671236529042546321860936599584189802657250250246695914442224645574013583678744715427750537353466912120749264423349295625108616427849178599143600331;
            5'd5: xpb[194] = 1024'd112517785703405668999645701989997469288237987368529642264916973069016699664381993912523988469356364907808438973593514860997517866899046753290532039356520121456625094972839716186125005564387384528235969769103238254666323418472640096703332358156706775121806761200738730103109082674977860533373828843218125363662;
            5'd6: xpb[194] = 1024'd85394664570436906240055271426071190048006213991941297066647625656829281462334737131022757677364568165592867005329220459365395903942367970126574397221291729374473844139579172488297911000657979145359084679568989967053843762078809406858007401914756350439440152075239652911688287980401979433201118681211512642662;
            5'd7: xpb[194] = 1024'd58271543437468143480464840862144910807774440615352951868378278244641863260287480349521526885372771423377295037064926057733273940985689186962616755086063337292322593306318628790470816436928573762482199590034741679441364105684978717012682445672805925757073542949740575720267493285826098333028408519204899921662;
            5'd8: xpb[194] = 1024'd31148422304499380720874410298218631567542667238764606670108930832454445058240223568020296093380974681161723068800631656101151978029010403798659112950834945210171342473058085092643721873199168379605314500500493391828884449291148027167357489430855501074706933824241498528846698591250217232855698357198287200662;
            5'd9: xpb[194] = 1024'd4025301171530617961283979734292352327310893862176261471839583420267026856192966786519065301389177938946151100536337254469030015072331620634701470815606553128020091639797541394816627309469762996728429410966245104216404792897317337322032533188905076392340324698742421337425903896674336132682988195191674479662;
            5'd10: xpb[194] = 1024'd100968875722686596600492476575180505831777547611323600401702091073056503991454848915032905724055055506173728539729536287415971892956873172025903953696709201979559515376108215034619771937257563335161741929819236662968285986724383420441686146630184100976793618987360402176111637276027088049628967859810656242993;
            5'd11: xpb[194] = 1024'd73845754589717833840902046011254226591545774234735255203432743660869085789407592133531674932063258763958156571465241885783849930000194388861946311561480809897408264542847671336792677373528157952284856840284988375355806330330552730596361190388233676294427009861861324984690842581451206949456257697804043521993;
            5'd12: xpb[194] = 1024'd46722633456749071081311615447327947351314000858146910005163396248681667587360335352030444140071462021742584603200947484151727967043515605697988669426252417815257013709587127638965582809798752569407971750750740087743326673936722040751036234146283251612060400736362247793270047886875325849283547535797430800993;
            5'd13: xpb[194] = 1024'd19599512323780308321721184883401668111082227481558564806894048836494249385313078570529213348079665279527012634936653082519606004086836822534031027291024025733105762876326583941138488246069347186531086661216491800130847017542891350905711277904332826929693791610863170601849253192299444749110837373790818079993;
            5'd14: xpb[194] = 1024'd116543086874936286960929681724289821615548881230705903736756556489283726520574960699043053770745542846754590074129852115466547881971378373925233510172126674584645186612637257580941632873857147524964399180069483358882728211369957434025364891345611851514147085899481151440534986571652196666056817038409799843324;
            5'd15: xpb[194] = 1024'd89419965741967524201339251160363542375317107854117558538487209077096308318527703917541822978753746104539018105865557713834425919014699590761275868036898282502493935779376713883114538310127742142087514090535235071270248554976126744180039935103661426831780476773982074249114191877076315565884106876403187122324;
            5'd16: xpb[194] = 1024'd62296844608998761441748820596437263135085334477529213340217861664908890116480447136040592186761949362323446137601263312202303956058020807597318225901669890420342684946116170185287443746398336759210629001000986783657768898582296054334714978861711002149413867648482997057693397182500434465711396714396574401324;
            5'd17: xpb[194] = 1024'd35173723476029998682158390032510983894853561100940868141948514252721471914433190354539361394770152620107874169336968910570181993101342024433360583766441498338191434112855626487460349182668931376333743911466738496045289242188465364489390022619760577467047258522983919866272602487924553365538686552389961680324;
            5'd18: xpb[194] = 1024'd8050602343061235922567959468584704654621787724352522943679166840534053712385933573038130602778355877892302201072674508938060030144663241269402941631213106256040183279595082789633254618939525993456858821932490208432809585794634674644065066377810152784680649397484842674851807793348672265365976390383348959324;
            5'd19: xpb[194] = 1024'd104994176894217214561776456309472858159088441473499861873541674493323530847647815701551971025444233445119879640265873541885001908029204792660605424512315755107579607015905756429436399246727326331890171340785481767184690779621700757763718679819089177369133943686102823513537541172701424182311956055002330722655;
            5'd20: xpb[194] = 1024'd77871055761248451802186025745546578918856668096911516675272327081136112645600558920050740233452436702904307672001579140252879945072526009496647782377087363025428356182645212731609304682997920949013286251251233479572211123227870067918393723577138752686767334560603746322116746478125543082139245892995718001655;
            5'd21: xpb[194] = 1024'd50747934628279689042595595181620299678624894720323171477002979668948694443553302138549509441460639960688735703737284738620757982115847226332690140241858970943277105349384669033782210119268515566136401161716985191959731466834039378073068767335188328004400725435104669130695951783549661981966535730989105280655;
            5'd22: xpb[194] = 1024'd23624813495310926283005164617694020438393121343734826278733632256761276241506045357048278649468843218473163735472990336988636019159168443168732498106630578861125854516124125335955115555539110183259516072182736904347251810440208688227743811093237903322034116309605591939275157088973780881793825568982492559655;
            5'd23: xpb[194] = 1024'd120568388046466904922213661458582173942859775092882165208596139909550753376767927485562119072134720785700741174666189369935577897043709994559934980987733227712665278252434798975758260183326910521692828591035728463099133004267274771347397424534516927906487410598223572777960890468326532798739805233601474322986;
            5'd24: xpb[194] = 1024'd93445266913498142162623230894655894702628001716293820010326792497363335174720670704060888280142924043485169206401894968303455934087031211395977338852504835630514027419174255277931165619597505138815943501501480175486653347873444081502072468292566503224120801472724495586540095773750651698567095071594861601986;
            5'd25: xpb[194] = 1024'd66322145780529379403032800330729615462396228339705474812057445085175916972673413922559657488151127301269597238137600566671333971130352428232019696717276443548362776585913711580104071055868099755939058411967231887874173691479613391656747512050616078541754192347225418395119301079174770598394384909588248880986;
            5'd26: xpb[194] = 1024'd39199024647560616643442369766803336222164454963117129613788097672988498770626157141058426696159330559054025269873306165039212008173673645068062054582048051466211525752653167882276976492138694373062173322432983600261694035085782701811422555808665653859387583221726341203698506384598889498221674747581636159986;
            5'd27: xpb[194] = 1024'd12075903514591853883851939202877056981932681586528784415518750260801080568578900359557195904167533816838453301609011763407090045216994861904104412446819659384060274919392624184449881928409288990185288232898735312649214378691952011966097599566715229177020974096227264012277711690023008398048964585575023438986;
            5'd28: xpb[194] = 1024'd109019478065747832523060436043765210486399335335676123345381257913590557703840782488071036326833411384066030740802210796354031923101536413295306895327922308235599698655703297824253026556197089328618600751751726871401095572519018095085751213007994253761474268384845244850963445069375760314994944250194005202317;
            5'd29: xpb[194] = 1024'd81896356932779069763470005479838931246167561959087778147111910501403139501793525706569805534841614641850458772537916394721909960144857630131349253192693916153448447822442754126425931992467683945741715662217478583788615916125187405240426256766043829079107659259346167659542650374799879214822234088187392481317;
            5'd30: xpb[194] = 1024'd54773235799810307003879574915912652005935788582499432948842563089215721299746268925068574742849817899634886804273621993089787997188178846967391611057465524071297196989182210428598837428738278562864830572683230296176136259731356715395101300524093404396741050133847090468121855680223998114649523926180779760317;
            5'd31: xpb[194] = 1024'd27650114666841544244289144351986372765704015205911087750573215677028303097699012143567343950858021157419314836009327591457666034231500063803433968922237131989145946155921666730771742865008873179987945483148982008563656603337526025549776344282142979714374441008348013276701060985648117014476813764174167039317;
        endcase
    end

    always_comb begin
        case(flag[65][5:0])
            6'd0: xpb[195] = 1024'd0;
            6'd1: xpb[195] = 1024'd62296844608998761441748820596437263135085334477529213340217861664908890116480447136040592186761949362323446137601263312202303956058020807597318225901669890420342684946116170185287443746398336759210629001000986783657768898582296054334714978861711002149413867648482997057693397182500434465711396714396574401324;
            6'd2: xpb[195] = 1024'd526993533872781484698713788060093525472241829322742552303868264840884895651755362066113158866224415203742867745033189825544071274821280639476326787008739906994695322661123032944648301279467797111060393614733720951176946943695335704451388040192555032007831882848936085280266291072235914304103602167554318317;
            6'd3: xpb[195] = 1024'd62823838142871542926447534384497356660557576306851955892521729929749775012132202498106705345628173777527189005346296502027848027332842088236794552688678630327337380268777293218232092047677804556321689394615720504608945845525991390039166366901903557181421699531331933142973663473572670380015500316564128719641;
            6'd4: xpb[195] = 1024'd1053987067745562969397427576120187050944483658645485104607736529681769791303510724132226317732448830407485735490066379651088142549642561278952653574017479813989390645322246065889296602558935594222120787229467441902353893887390671408902776080385110064015663765697872170560532582144471828608207204335108636634;
            6'd5: xpb[195] = 1024'd63350831676744324411146248172557450186029818136174698444825598194590659907783957860172818504494398192730931873091329691853392098607663368876270879475687370234332075591438416251176740348957272353432749788230454225560122792469686725743617754942096112213429531414180869228253929764644906294319603918731683037958;
            6'd6: xpb[195] = 1024'd1580980601618344454096141364180280576416725487968227656911604794522654686955266086198339476598673245611228603235099569476632213824463841918428980361026219720984085967983369098833944903838403391333181180844201162853530840831086007113354164120577665096023495648546808255840798873216707742912310806502662954951;
            6'd7: xpb[195] = 1024'd63877825210617105895844961960617543711502059965497440997129466459431544803435713222238931663360622607934674740836362881678936169882484649515747206262696110141326770914099539284121388650236740150543810181845187946511299739413382061448069142982288667245437363297029805313534196055717142208623707520899237356275;
            6'd8: xpb[195] = 1024'd2107974135491125938794855152240374101888967317290970209215473059363539582607021448264452635464897660814971470980132759302176285099285122557905307148034959627978781290644492131778593205117871188444241574458934883804707787774781342817805552160770220128031327531395744341121065164288943657216414408670217273268;
            6'd9: xpb[195] = 1024'd64404818744489887380543675748677637236974301794820183549433334724272429699087468584305044822226847023138417608581396071504480241157305930155223533049704850048321466236760662317066036951516207947654870575459921667462476686357077397152520531022481222277445195179878741398814462346789378122927811123066791674592;
            6'd10: xpb[195] = 1024'd2634967669363907423493568940300467627361209146613712761519341324204424478258776810330565794331122076018714338725165949127720356374106403197381633935043699534973476613305615164723241506397338985555301968073668604755884734718476678522256940200962775160039159414244680426401331455361179571520518010837771591585;
            6'd11: xpb[195] = 1024'd64931812278362668865242389536737730762446543624142926101737202989113314594739223946371157981093071438342160476326429261330024312432127210794699859836713589955316161559421785350010685252795675744765930969074655388413653633300772732856971919062673777309453027062727677484094728637861614037231914725234345992909;
            6'd12: xpb[195] = 1024'd3161961203236688908192282728360561152833450975936455313823209589045309373910532172396678953197346491222457206470199138953264427648927683836857960722052439441968171935966738197667889807676806782666362361688402325707061681662172014226708328241155330192046991297093616511681597746433415485824621613005325909902;
            6'd13: xpb[195] = 1024'd65458805812235450349941103324797824287918785453465668654041071253954199490390979308437271139959295853545903344071462451155568383706948491434176186623722329862310856882082908382955333554075143541876991362689389109364830580244468068561423307102866332341460858945576613569374994928933849951536018327401900311226;
            6'd14: xpb[195] = 1024'd3688954737109470392890996516420654678305692805259197866127077853886194269562287534462792112063570906426200074215232328778808498923748964476334287509061179348962867258627861230612538108956274579777422755303136046658238628605867349931159716281347885224054823179942552596961864037505651400128725215172880228219;
            6'd15: xpb[195] = 1024'd65985799346108231834639817112857917813391027282788411206344939518795084386042734670503384298825520268749646211816495640981112454981769772073652513410731069769305552204744031415899981855354611338988051756304122830316007527188163404265874695143058887373468690828425549654655261220006085865840121929569454629543;
            6'd16: xpb[195] = 1024'd4215948270982251877589710304480748203777934634581940418430946118727079165214042896528905270929795321629942941960265518604352570198570245115810614296069919255957562581288984263557186410235742376888483148917869767609415575549562685635611104321540440256062655062791488682242130328577887314432828817340434546536;
            6'd17: xpb[195] = 1024'd66512792879981013319338530900918011338863269112111153758648807783635969281694490032569497457691744683953389079561528830806656526256591052713128840197739809676300247527405154448844630156634079136099112149918856551267184474131858739970326083183251442405476522711274485739935527511078321780144225531737008947860;
            6'd18: xpb[195] = 1024'd4742941804855033362288424092540841729250176463904682970734814383567964060865798258595018429796019736833685809705298708429896641473391525755286941083078659162952257903950107296501834711515210173999543542532603488560592522493258021340062492361732995288070486945640424767522396619650123228736932419507988864853;
            6'd19: xpb[195] = 1024'd67039786413853794804037244688978104864335510941433896310952676048476854177346245394635610616557969099157131947306562020632200597531412333352605166984748549583294942850066277481789278457913546933210172543533590272218361421075554075674777471223443997437484354594123421825215793802150557694448329133904563266177;
            6'd20: xpb[195] = 1024'd5269935338727814846987137880600935254722418293227425523038682648408848956517553620661131588662244152037428677450331898255440712748212806394763267870087399069946953226611230329446483012794677971110603936147337209511769469436953357044513880401925550320078318828489360852802662910722359143041036021675543183170;
            6'd21: xpb[195] = 1024'd67566779947726576288735958477038198389807752770756638863256544313317739072998000756701723775424193514360874815051595210457744668806233613992081493771757289490289638172727400514733926759193014730321232937148323993169538368019249411379228859263636552469492186476972357910496060093222793608752432736072117584494;
            6'd22: xpb[195] = 1024'd5796928872600596331685851668661028780194660122550168075342550913249733852169308982727244747528468567241171545195365088080984784023034087034239594657096138976941648549272353362391131314074145768221664329762070930462946416380648692748965268442118105352086150711338296938082929201794595057345139623843097501487;
            6'd23: xpb[195] = 1024'd68093773481599357773434672265098291915279994600079381415560412578158623968649756118767836934290417929564617682796628400283288740081054894631557820558766029397284333495388523547678575060472482527432293330763057714120715314962944747083680247303829107501500018359821293995776326384295029523056536338239671902811;
            6'd24: xpb[195] = 1024'd6323922406473377816384565456721122305666901951872910627646419178090618747821064344793357906394692982444914412940398277906528855297855367673715921444104878883936343871933476395335779615353613565332724723376804651414123363324344028453416656482310660384093982594187233023363195492866830971649243226010651819804;
            6'd25: xpb[195] = 1024'd68620767015472139258133386053158385440752236429402123967864280842999508864301511480833950093156642344768360550541661590108832811355876175271034147345774769304279028818049646580623223361751950324543353724377791435071892261906640082788131635344021662533507850242670230081056592675367265437360639940407226221128;
            6'd26: xpb[195] = 1024'd6850915940346159301083279244781215831139143781195653179950287442931503643472819706859471065260917397648657280685431467732072926572676648313192248231113618790931039194594599428280427916633081362443785116991538372365300310268039364157868044522503215416101814477036169108643461783939066885953346828178206138121;
            6'd27: xpb[195] = 1024'd69147760549344920742832099841218478966224478258724866520168149107840393759953266842900063252022866759972103418286694779934376882630697455910510474132783509211273724140710769613567871663031418121654414117992525156023069208850335418492583023384214217565515682125519166166336858966439501351664743542574780539445;
            6'd28: xpb[195] = 1024'd7377909474218940785781993032841309356611385610518395732254155707772388539124575068925584224127141812852400148430464657557616997847497928952668575018122358697925734517255722461225076217912549159554845510606272093316477257211734699862319432562695770448109646359885105193923728075011302800257450430345760456438;
            6'd29: xpb[195] = 1024'd69674754083217702227530813629278572491696720088047609072472017372681278655605022204966176410889091175175846286031727969759920953905518736549986800919792249118268419463371892646512519964310885918765474511607258876974246155794030754197034411424406772597523514008368102251617125257511737265968847144742334857762;
            6'd30: xpb[195] = 1024'd7904903008091722270480706820901402882083627439841138284558023972613273434776330430991697382993366228056143016175497847383161069122319209592144901805131098604920429839916845494169724519192016956665905904221005814267654204155430035566770820602888325480117478242734041279203994366083538714561554032513314774755;
            6'd31: xpb[195] = 1024'd70201747617090483712229527417338666017168961917370351624775885637522163551256777567032289569755315590379589153776761159585465025180340017189463127706800989025263114786033015679457168265590353715876534905221992597925423102737726089901485799464599327629531345891217038336897391548583973180272950746909889176079;
            6'd32: xpb[195] = 1024'd8431896541964503755179420608961496407555869269163880836861892237454158330428085793057810541859590643259885883920531037208705140397140490231621228592139838511915125162577968527114372820471484753776966297835739535218831151099125371271222208643080880512125310125582977364484260657155774628865657634680869093072;
            6'd33: xpb[195] = 1024'd70728741150963265196928241205398759542641203746693094177079753902363048446908532929098402728621540005583332021521794349411009096455161297828939454493809728932257810108694138712401816566869821512987595298836726318876600049681421425605937187504791882661539177774065974422177657839656209094577054349077443494396;
            6'd34: xpb[195] = 1024'd8958890075837285239878134397021589933028111098486623389165760502295043226079841155123923700725815058463628751665564227034249211671961770871097555379148578418909820485239091560059021121750952550888026691450473256170008098042820706975673596683273435544133142008431913449764526948228010543169761236848423411389;
            6'd35: xpb[195] = 1024'd71255734684836046681626954993458853068113445576015836729383622167203933342560288291164515887487764420787074889266827539236553167729982578468415781280818468839252505431355261745346464868149289310098655692451460039827776996625116761310388575544984437693547009656914910507457924130728445008881157951244997812713;
            6'd36: xpb[195] = 1024'd9485883609710066724576848185081683458500352927809365941469628767135928121731596517190036859592039473667371619410597416859793282946783051510573882166157318325904515807900214593003669423030420347999087085065206977121185044986516042680124984723465990576140973891280849535044793239300246457473864839015977729706;
            6'd37: xpb[195] = 1024'd71782728218708828166325668781518946593585687405338579281687490432044818238212043653230629046353988835990817757011860729062097239004803859107892108067827208746247200754016384778291113169428757107209716086066193760778953943568812097014839963585176992725554841539763846592738190421800680923185261553412552131030;
            6'd38: xpb[195] = 1024'd10012877143582848209275561973141776983972594757132108493773497031976813017383351879256150018458263888871114487155630606685337354221604332150050208953166058232899211130561337625948317724309888145110147478679940698072361991930211378384576372763658545608148805774129785620325059530372482371777968441183532048023;
            6'd39: xpb[195] = 1024'd72309721752581609651024382569579040119057929234661321833991358696885703133863799015296742205220213251194560624756893918887641310279625139747368434854835948653241896076677507811235761470708224904320776479680927481730130890512507432719291351625369547757562673422612782678018456712872916837489365155580106449347;
            6'd40: xpb[195] = 1024'd10539870677455629693974275761201870509444836586454851046077365296817697913035107241322263177324488304074857354900663796510881425496425612789526535740174798139893906453222460658892966025589355942221207872294674419023538938873906714089027760803851100640156637656978721705605325821444718286082072043351086366340;
            6'd41: xpb[195] = 1024'd72836715286454391135723096357639133644530171063984064386295226961726588029515554377362855364086437666398303492501927108713185381554446420386844761641844688560236591399338630844180409771987692701431836873295661202681307837456202768423742739665562102789570505305461718763298723003945152751793468757747660767664;
            6'd42: xpb[195] = 1024'd11066864211328411178672989549261964034917078415777593598381233561658582808686862603388376336190712719278600222645696986336425496771246893429002862527183538046888601775883583691837614326868823739332268265909408139974715885817602049793479148844043655672164469539827657790885592112516954200386175645518640684657;
            6'd43: xpb[195] = 1024'd73363708820327172620421810145699227170002412893306806938599095226567472925167309739428968522952662081602046360246960298538729452829267701026321088428853428467231286721999753877125058073267160498542897266910394923632484784399898104128194127705754657821578337188310654848578989295017388666097572359915215085981;
            6'd44: xpb[195] = 1024'd11593857745201192663371703337322057560389320245100336150685101826499467704338617965454489495056937134482343090390730176161969568046068174068479189314192277953883297098544706724782262628148291536443328659524141860925892832761297385497930536884236210704172301422676593876165858403589190114690279247686195002974;
            6'd45: xpb[195] = 1024'd73890702354199954105120523933759320695474654722629549490902963491408357820819065101495081681818886496805789227991993488364273524104088981665797415215862168374225982044660876910069706374546628295653957660525128644583661731343593439832645515745947212853586169071159590933859255586089624580401675962082769404298;
            6'd46: xpb[195] = 1024'd12120851279073974148070417125382151085861562074423078702988970091340352599990373327520602653923161549686085958135763365987513639320889454707955516101201017860877992421205829757726910929427759333554389053138875581877069779704992721202381924924428765736180133305525529961446124694661426028994382849853749321291;
            6'd47: xpb[195] = 1024'd74417695888072735589819237721819414220946896551952292043206831756249242716470820463561194840685110912009532095737026678189817595378910262305273742002870908281220677367321999943014354675826096092765018054139862365534838678287288775537096903786139767885594000954008527019139521877161860494705779564250323722615;
            6'd48: xpb[195] = 1024'd12647844812946755632769130913442244611333803903745821255292838356181237495642128689586715812789385964889828825880796555813057710595710735347431842888209757767872687743866952790671559230707227130665449446753609302828246726648688056906833312964621320768187965188374466046726390985733661943298486452021303639608;
            6'd49: xpb[195] = 1024'd74944689421945517074517951509879507746419138381275034595510700021090127612122575825627307999551335327213274963482059868015361666653731542944750068789879648188215372689983122975959002977105563889876078447754596086486015625230984111241548291826332322917601832836857463104419788168234096409009883166417878040932;
            6'd50: xpb[195] = 1024'd13174838346819537117467844701502338136806045733068563807596706621022122391293884051652828971655610380093571693625829745638601781870532015986908169675218497674867383066528075823616207531986694927776509840368343023779423673592383392611284701004813875800195797071223402132006657276805897857602590054188857957925;
            6'd51: xpb[195] = 1024'd75471682955818298559216665297939601271891380210597777147814568285931012507774331187693421158417559742417017831227093057840905737928552823584226395576888388095210068012644246008903651278385031686987138841369329807437192572174679446945999679866524877949609664719706399189700054459306332323313986768585432359249;
            6'd52: xpb[195] = 1024'd13701831880692318602166558489562431662278287562391306359900574885863007286945639413718942130521834795297314561370862935464145853145353296626384496462227237581862078389189198856560855833266162724887570233983076744730600620536078728315736089045006430832203628954072338217286923567878133771906693656356412276242;
            6'd53: xpb[195] = 1024'd75998676489691080043915379085999694797363622039920519700118436550771897403426086549759534317283784157620760698972126247666449809203374104223702722363897128002204763335305369041848299579664499484098199234984063528388369519118374782650451067906717432981617496602555335274980320750378568237618090370752986677566;
            6'd54: xpb[195] = 1024'd14228825414565100086865272277622525187750529391714048912204443150703892182597394775785055289388059210501057429115896125289689924420174577265860823249235977488856773711850321889505504134545630521998630627597810465681777567479774064020187477085198985864211460836921274302567189858950369686210797258523966594559;
            6'd55: xpb[195] = 1024'd76525670023563861528614092874059788322835863869243262252422304815612782299077841911825647476150008572824503566717159437491993880478195384863179049150905867909199458657966492074792947880943967281209259628598797249339546466062070118354902455946909988013625328485404271360260587041450804151922193972920540995883;
            6'd56: xpb[195] = 1024'd14755818948437881571563986065682618713222771221036791464508311415544777078249150137851168448254283625704800296860929315115233995694995857905337150036244717395851469034511444922450152435825098319109691021212544186632954514423469399724638865125391540896219292719770210387847456150022605600514900860691520912876;
            6'd57: xpb[195] = 1024'd77052663557436643013312806662119881848308105698566004804726173080453667194729597273891760635016232988028246434462192627317537951753016665502655375937914607816194153980627615107737596182223435078320320022213530970290723413005765454059353843987102543045633160368253207445540853332523040066226297575088095314200;
            6'd58: xpb[195] = 1024'd15282812482310663056262699853742712238695013050359534016812179680385661973900905499917281607120508040908543164605962504940778066969817138544813476823253457302846164357172567955394800737104566116220751414827277907584131461367164735429090253165584095928227124602619146473127722441094841514819004462859075231193;
            6'd59: xpb[195] = 1024'd77579657091309424498011520450179975373780347527888747357030041345294552090381352635957873793882457403231989302207225817143082023027837946142131702724923347723188849303288738140682244483502902875431380415828264691241900359949460789763805232027295098077640992251102143530821119623595275980530401177255649632517;
            6'd60: xpb[195] = 1024'd15809806016183444540961413641802805764167254879682276569116047945226546869552660861983394765986732456112286032350995694766322138244638419184289803610262197209840859679833690988339449038384033913331811808442011628535308408310860071133541641205776650960234956485468082558407988732167077429123108065026629549510;
            6'd61: xpb[195] = 1024'd78106650625182205982710234238240068899252589357211489909333909610135436986033107998023986952748681818435732169952259006968626094302659226781608029511932087630183544625949861173626892784782370672542440809442998412193077306893156125468256620067487653109648824133951079616101385914667511894834504779423203950834;
            6'd62: xpb[195] = 1024'd16336799550056226025660127429862899289639496709005019121419916210067431765204416224049507924852956871316028900096028884591866209519459699823766130397270937116835555002494814021284097339663501710442872202056745349486485355254555406837993029245969205992242788368317018643688255023239313343427211667194183867827;
            6'd63: xpb[195] = 1024'd78633644159054987467408948026300162424724831186534232461637777874976321881684863360090100111614906233639475037697292196794170165577480507421084356298940827537178239948610984206571541086061838469653501203057732133144254253836851461172708008107680208141656656016800015701381652205739747809138608381590758269151;
        endcase
    end

    always_comb begin
        case(flag[65][11:6])
            6'd0: xpb[196] = 1024'd0;
            6'd1: xpb[196] = 1024'd16863793083929007510358841217922992815111738538327761673723784474908316660856171586115621083719181286519771767841062074417410280794280980463242457184279677023830250325155937054228745640942969507553932595671479070437662302198250742542444417286161761024250620251165954728968521314311549257731315269361738186144;
            6'd2: xpb[196] = 1024'd33727586167858015020717682435845985630223477076655523347447568949816633321712343172231242167438362573039543535682124148834820561588561960926484914368559354047660500650311874108457491281885939015107865191342958140875324604396501485084888834572323522048501240502331909457937042628623098515462630538723476372288;
            6'd3: xpb[196] = 1024'd50591379251787022531076523653768978445335215614983285021171353424724949982568514758346863251157543859559315303523186223252230842382842941389727371552839031071490750975467811162686236922828908522661797787014437211312986906594752227627333251858485283072751860753497864186905563942934647773193945808085214558432;
            6'd4: xpb[196] = 1024'd67455172335716030041435364871691971260446954153311046694895137899633266643424686344462484334876725146079087071364248297669641123177123921852969828737118708095321001300623748216914982563771878030215730382685916281750649208793002970169777669144647044097002481004663818915874085257246197030925261077446952744576;
            6'd5: xpb[196] = 1024'd84318965419645037551794206089614964075558692691638808368618922374541583304280857930578105418595906432598858839205310372087051403971404902316212285921398385119151251625779685271143728204714847537769662978357395352188311510991253712712222086430808805121253101255829773644842606571557746288656576346808690930720;
            6'd6: xpb[196] = 1024'd101182758503574045062153047307537956890670431229966570042342706849449899965137029516693726502315087719118630607046372446504461684765685882779454743105678062142981501950935622325372473845657817045323595574028874422625973813189504455254666503716970566145503721506995728373811127885869295546387891616170429116864;
            6'd7: xpb[196] = 1024'd118046551587503052572511888525460949705782169768294331716066491324358216625993201102809347586034269005638402374887434520921871965559966863242697200289957739166811752276091559379601219486600786552877528169700353493063636115387755197797110921003132327169754341758161683102779649200180844804119206885532167303008;
            6'd8: xpb[196] = 1024'd10843648987307318684071802338569509776195481180886409261658420734289637949540233778909897455095775982715024735271003160760218405513027509150779532457906375256951328031676279096199725936026550339121263156984592717136937567365109167374576768606064638927185058595210579801641642440563761044731832328268311004821;
            6'd9: xpb[196] = 1024'd27707442071236326194430643556492502591307219719214170935382205209197954610396405365025518538814957269234796503112065235177628686307308489614021989642186052280781578356832216150428471576969519846675195752656071787574599869563359909917021185892226399951435678846376534530610163754875310302463147597630049190965;
            6'd10: xpb[196] = 1024'd44571235155165333704789484774415495406418958257541932609105989684106271271252576951141139622534138555754568270953127309595038967101589470077264446826465729304611828681988153204657217217912489354229128348327550858012262171761610652459465603178388160975686299097542489259578685069186859560194462866991787377109;
            6'd11: xpb[196] = 1024'd61435028239094341215148325992338488221530696795869694282829774159014587932108748537256760706253319842274340038794189384012449247895870450540506904010745406328442079007144090258885962858855458861783060943999029928449924473959861395001910020464549921999936919348708443988547206383498408817925778136353525563253;
            6'd12: xpb[196] = 1024'd78298821323023348725507167210261481036642435334197455956553558633922904592964920123372381789972501128794111806635251458429859528690151431003749361195025083352272329332300027313114708499798428369336993539670508998887586776158112137544354437750711683024187539599874398717515727697809958075657093405715263749397;
            6'd13: xpb[196] = 1024'd95162614406952356235866008428184473851754173872525217630277343108831221253821091709488002873691682415313883574476313532847269809484432411466991818379304760376102579657455964367343454140741397876890926135341988069325249078356362880086798855036873444048438159851040353446484249012121507333388408675077001935541;
            6'd14: xpb[196] = 1024'd112026407490881363746224849646107466666865912410852979304001127583739537914677263295603623957410863701833655342317375607264680090278713391930234275563584437399932829982611901421572199781684367384444858731013467139762911380554613622629243272323035205072688780102206308175452770326433056591119723944438740121685;
            6'd15: xpb[196] = 1024'd4823504890685629857784763459216026737279223823445056849593056993670959238224295971704173826472370678910277702700944247103026530231774037838316607731533073490072405738196621138170706231110131170688593718297706363836212832531967592206709119925967516830119496939255204874314763566815972831732349387174883823498;
            6'd16: xpb[196] = 1024'd21687297974614637368143604677139019552390962361772818523316841468579275899080467557819794910191551965430049470542006321520436811026055018301559064915812750513902656063352558192399451872053100678242526313969185434273875134730218334749153537212129277854370117190421159603283284881127522089463664656536622009642;
            6'd17: xpb[196] = 1024'd38551091058543644878502445895062012367502700900100580197040625943487592559936639143935415993910733251949821238383068395937847091820335998764801522100092427537732906388508495246628197512996070185796458909640664504711537436928469077291597954498291038878620737441587114332251806195439071347194979925898360195786;
            6'd18: xpb[196] = 1024'd55414884142472652388861287112985005182614439438428341870764410418395909220792810730051037077629914538469593006224130470355257372614616979228043979284372104561563156713664432300856943153939039693350391505312143575149199739126719819834042371784452799902871357692753069061220327509750620604926295195260098381930;
            6'd19: xpb[196] = 1024'd72278677226401659899220128330907997997726177976756103544488194893304225881648982316166658161349095824989364774065192544772667653408897959691286436468651781585393407038820369355085688794882009200904324100983622645586862041324970562376486789070614560927121977943919023790188848824062169862657610464621836568074;
            6'd20: xpb[196] = 1024'd89142470310330667409578969548830990812837916515083865218211979368212542542505153902282279245068277111509136541906254619190077934203178940154528893652931458609223657363976306409314434435824978708458256696655101716024524343523221304918931206356776321951372598195084978519157370138373719120388925733983574754218;
            6'd21: xpb[196] = 1024'd106006263394259674919937810766753983627949655053411626891935763843120859203361325488397900328787458398028908309747316693607488214997459920617771350837211135633053907689132243463543180076767948216012189292326580786462186645721472047461375623642938082975623218446250933248125891452685268378120241003345312940362;
            6'd22: xpb[196] = 1024'd122870056478188682430296651984676976443061393591739388565659548318029175864217497074513521412506639684548680077588378768024898495791740901081013808021490812656884158014288180517771925717710917723566121887998059856899848947919722790003820040929099843999873838697416887977094412766996817635851556272707051126506;
            6'd23: xpb[196] = 1024'd15667153877992948541856565797785536513474705004331466111251477727960597187764529750614071281568146661625302437971947407863244935744801546989096140189439448747023733769872900234370432167136681509809856875282299080973150399897076759581285888532032155757304555534465784675956406007379733876464181715443194828319;
            6'd24: xpb[196] = 1024'd32530946961921956052215407015708529328586443542659227784975262202868913848620701336729692365287327948145074205813009482280655216539082527452338597373719125770853984095028837288599177808079651017363789470953778151410812702095327502123730305818193916781555175785631739404924927321691283134195496984804933014463;
            6'd25: xpb[196] = 1024'd49394740045850963562574248233631522143698182080986989458699046677777230509476872922845313449006509234664845973654071556698065497333363507915581054557998802794684234420184774342827923449022620524917722066625257221848475004293578244666174723104355677805805796036797694133893448636002832391926812254166671200607;
            6'd26: xpb[196] = 1024'd66258533129779971072933089451554514958809920619314751132422831152685547170333044508960934532725690521184617741495133631115475778127644488378823511742278479818514484745340711397056669089965590032471654662296736292286137306491828987208619140390517438830056416287963648862861969950314381649658127523528409386751;
            6'd27: xpb[196] = 1024'd83122326213708978583291930669477507773921659157642512806146615627593863831189216095076555616444871807704389509336195705532886058921925468842065968926558156842344735070496648451285414730908559540025587257968215362723799608690079729751063557676679199854307036539129603591830491264625930907389442792890147572895;
            6'd28: xpb[196] = 1024'd99986119297637986093650771887400500589033397695970274479870400102502180492045387681192176700164053094224161277177257779950296339716206449305308426110837833866174985395652585505514160371851529047579519853639694433161461910888330472293507974962840960878557656790295558320799012578937480165120758062251885759039;
            6'd29: xpb[196] = 1024'd116849912381566993604009613105323493404145136234298036153594184577410497152901559267307797783883234380743933045018319854367706620510487429768550883295117510890005235720808522559742906012794498555133452449311173503599124213086581214835952392249002721902808277041461513049767533893249029422852073331613623945183;
            6'd30: xpb[196] = 1024'd9647009781371259715569526918432053474558447646890113699186113987341918476448591943408347652944741357820555405401888494206053060463548075676633215463066146980144811476393242276341412462220262341377187436595412727672425665063935184413418239851935033660238993878510409748629527133631945663464698774349767646996;
            6'd31: xpb[196] = 1024'd26510802865300267225928368136355046289670186185217875372909898462250235137304763529523968736663922644340327173242950568623463341257829056139875672647345824003975061801549179330570158103163231848931120032266891798110087967262185926955862657138096794684489614129676364477598048447943494921196014043711505833140;
            6'd32: xpb[196] = 1024'd43374595949229274736287209354278039104781924723545637046633682937158551798160935115639589820383103930860098941084012643040873622052110036603118129831625501027805312126705116384798903744106201356485052627938370868547750269460436669498307074424258555708740234380842319206566569762255044178927329313073244019284;
            6'd33: xpb[196] = 1024'd60238389033158282246646050572201031919893663261873398720357467412066868459017106701755210904102285217379870708925074717458283902846391017066360587015905178051635562451861053439027649385049170864038985223609849938985412571658687412040751491710420316732990854632008273935535091076566593436658644582434982205428;
            6'd34: xpb[196] = 1024'd77102182117087289757004891790124024735005401800201160394081251886975185119873278287870831987821466503899642476766136791875694183640671997529603044200184855075465812777016990493256395025992140371592917819281329009423074873856938154583195908996582077757241474883174228664503612390878142694389959851796720391572;
            6'd35: xpb[196] = 1024'd93965975201016297267363733008047017550117140338528922067805036361883501780729449873986453071540647790419414244607198866293104464434952977992845501384464532099296063102172927547485140666935109879146850414952808079860737176055188897125640326282743838781492095134340183393472133705189691952121275121158458577716;
            6'd36: xpb[196] = 1024'd110829768284945304777722574225970010365228878876856683741528820836791818441585621460102074155259829076939186012448260940710514745229233958456087958568744209123126313427328864601713886307878079386700783010624287150298399478253439639668084743568905599805742715385506138122440655019501241209852590390520196763860;
            6'd37: xpb[196] = 1024'd3626865684749570889282488039078570435642190289448761287120750246723239765132654136202624024321336054015808372831829580548861185182294604364170290736692845213265889182913584318312392757303843172944517997908526374371700930230793609245550591171837911563173432222555034821302648259884157450465215833256340465673;
            6'd38: xpb[196] = 1024'd20490658768678578399641329257001563250753928827776522960844534721631556425988825722318245108040517340535580140672891654966271465976575584827412747920972522237096139508069521372541138398246812680498450593580005444809363232429044351787995008457999672587424052473720989550271169574195706708196531102618078651817;
            6'd39: xpb[196] = 1024'd37354451852607585910000170474924556065865667366104284634568319196539873086844997308433866191759698627055351908513953729383681746770856565290655205105252199260926389833225458426769884039189782188052383189251484515247025534627295094330439425744161433611674672724886944279239690888507255965927846371979816837961;
            6'd40: xpb[196] = 1024'd54218244936536593420359011692847548880977405904432046308292103671448189747701168894549487275478879913575123676355015803801092027565137545753897662289531876284756640158381395480998629680132751695606315784922963585684687836825545836872883843030323194635925292976052899008208212202818805223659161641341555024105;
            6'd41: xpb[196] = 1024'd71082038020465600930717852910770541696089144442759807982015888146356506408557340480665108359198061200094895444196077878218502308359418526217140119473811553308586890483537332535227375321075721203160248380594442656122350139023796579415328260316484955660175913227218853737176733517130354481390476910703293210249;
            6'd42: xpb[196] = 1024'd87945831104394608441076694128693534511200882981087569655739672621264823069413512066780729442917242486614667212037139952635912589153699506680382576658091230332417140808693269589456120962018690710714180976265921726560012441222047321957772677602646716684426533478384808466145254831441903739121792180065031396393;
            6'd43: xpb[196] = 1024'd104809624188323615951435535346616527326312621519415331329463457096173139730269683652896350526636423773134438979878202027053322869947980487143625033842370907356247391133849206643684866602961660218268113571937400796997674743420298064500217094888808477708677153729550763195113776145753452996853107449426769582537;
            6'd44: xpb[196] = 1024'd121673417272252623461794376564539520141424360057743093003187241571081456391125855239011971610355605059654210747719264101470733150742261467606867491026650584380077641459005143697913612243904629725822046167608879867435337045618548807042661512174970238732927773980716717924082297460065002254584422718788507768681;
            6'd45: xpb[196] = 1024'd14470514672056889573354290377648080211837671470335170548779170981012877714672887915112521479417112036730833108102832741309079590695322113514949823194599220470217217214589863414512118693330393512065781154893119091508638497595902776620127359777902550490358490817765614622944290700447918495197048161524651470494;
            6'd46: xpb[196] = 1024'd31334307755985897083713131595571073026949410008662932222502955455921194375529059501228142563136293323250604875943894815726489871489603093978192280378878897494047467539745800468740864334273363019619713750564598161946300799794153519162571777064064311514609111068931569351912812014759467752928363430886389656638;
            6'd47: xpb[196] = 1024'd48198100839914904594071972813494065842061148546990693896226739930829511036385231087343763646855474609770376643784956890143900152283884074441434737563158574517877717864901737522969609975216332527173646346236077232383963101992404261705016194350226072538859731320097524080881333329071017010659678700248127842782;
            6'd48: xpb[196] = 1024'd65061893923843912104430814031417058657172887085318455569950524405737827697241402673459384730574655896290148411626018964561310433078165054904677194747438251541707968190057674577198355616159302034727578941907556302821625404190655004247460611636387833563110351571263478809849854643382566268390993969609866028926;
            6'd49: xpb[196] = 1024'd81925687007772919614789655249340051472284625623646217243674308880646144358097574259575005814293837182809920179467081038978720713872446035367919651931717928565538218515213611631427101257102271542281511537579035373259287706388905746789905028922549594587360971822429433538818375957694115526122309238971604215070;
            6'd50: xpb[196] = 1024'd98789480091701927125148496467263044287396364161973978917398093355554461018953745845690626898013018469329691947308143113396130994666727015831162109115997605589368468840369548685655846898045241049835444133250514443696950008587156489332349446208711355611611592073595388267786897272005664783853624508333342401214;
            6'd51: xpb[196] = 1024'd115653273175630934635507337685186037102508102700301740591121877830462777679809917431806247981732199755849463715149205187813541275461007996294404566300277282613198719165525485739884592538988210557389376728921993514134612310785407231874793863494873116635862212324761342996755418586317214041584939777695080587358;
            6'd52: xpb[196] = 1024'd8450370575435200747067251498294597172921414112893818136713807240394199003356950107906797850793706732926086075532773827651887715414068642202486898468225918703338294921110205456483098988413974343633111716206232738207913762762761201452259711097805428393292929161810239695617411826700130282197565220431224289171;
            6'd53: xpb[196] = 1024'd25314163659364208257426092716217589988033152651221579810437591715302515664213121694022418934512888019445857843373835902069297996208349622665729355652505595727168545246266142510711844629356943851187044311877711808645576064961011943994704128383967189417543549412976194424585933141011679539928880489792962475315;
            6'd54: xpb[196] = 1024'd42177956743293215767784933934140582803144891189549341484161376190210832325069293280138040018232069305965629611214897976486708277002630603128971812836785272750998795571422079564940590270299913358740976907549190879083238367159262686537148545670128950441794169664142149153554454455323228797660195759154700661459;
            6'd55: xpb[196] = 1024'd59041749827222223278143775152063575618256629727877103157885160665119148985925464866253661101951250592485401379055960050904118557796911583592214270021064949774829045896578016619169335911242882866294909503220669949520900669357513429079592962956290711466044789915308103882522975769634778055391511028516438847603;
            6'd56: xpb[196] = 1024'd75905542911151230788502616369986568433368368266204864831608945140027465646781636452369282185670431879005173146897022125321528838591192564055456727205344626798659296221733953673398081552185852373848842098892149019958562971555764171622037380242452472490295410166474058611491497083946327313122826297878177033747;
            6'd57: xpb[196] = 1024'd92769335995080238298861457587909561248480106804532626505332729614935782307637808038484903269389613165524944914738084199738939119385473544518699184389624303822489546546889890727626827193128821881402774694563628090396225273754014914164481797528614233514546030417640013340460018398257876570854141567239915219891;
            6'd58: xpb[196] = 1024'd109633129079009245809220298805832554063591845342860388179056514089844098968493979624600524353108794452044716682579146274156349400179754524981941641573903980846319796872045827781855572834071791388956707290235107160833887575952265656706926214814775994538796650668805968069428539712569425828585456836601653406035;
            6'd59: xpb[196] = 1024'd2430226478813511920780212618941114134005156755452465724648443499775520292041012300701074222170301429121339042962714913994695840132815170890023973741852616936459372627630547498454079283497555175200442277519346384907189027929619626284392062417708306296227367505854864768290532952952342069198082279337797107848;
            6'd60: xpb[196] = 1024'd19294019562742519431139053836864106949116895293780227398372227974683836952897183886816695305889482715641110810803776988412106120927096151353266430926132293960289622952786484552682824924440524682754374873190825455344851330127870368826836479703870067320477987757020819497259054267263891326929397548699535293992;
            6'd61: xpb[196] = 1024'd36157812646671526941497895054787099764228633832107989072096012449592153613753355472932316389608664002160882578644839062829516401721377131816508888110411970984119873277942421606911570565383494190308307468862304525782513632326121111369280896990031828344728608008186774226227575581575440584660712818061273480136;
            6'd62: xpb[196] = 1024'd53021605730600534451856736272710092579340372370435750745819796924500470274609527059047937473327845288680654346485901137246926682515658112279751345294691648007950123603098358661140316206326463697862240064533783596220175934524371853911725314276193589368979228259352728955196096895886989842392028087423011666280;
            6'd63: xpb[196] = 1024'd69885398814529541962215577490633085394452110908763512419543581399408786935465698645163558557047026575200426114326963211664336963309939092742993802478971325031780373928254295715369061847269433205416172660205262666657838236722622596454169731562355350393229848510518683684164618210198539100123343356784749852424;
        endcase
    end

    always_comb begin
        case(flag[65][16:12])
            5'd0: xpb[197] = 1024'd0;
            5'd1: xpb[197] = 1024'd86749191898458549472574418708556078209563849447091274093267365874317103596321870231279179640766207861720197882168025286081747244104220073206236259663251002055610624253410232769597807488212402712970105255876741737095500538920873338996614148848517111417480468761684638413133139524510088357854658626146488038568;
            5'd2: xpb[197] = 1024'd49431688112792357546349910012297723674429271768446864058402876683657311855334601552543288066874741413997246356878557137584430647367219811857312394310170963177530573937249248201565375784907599704630012903366243627826640227620849905028249728013804773568141034109252218796159750975091543698590627425667381592805;
            5'd3: xpb[197] = 1024'd12114184327126165620125401316039369139294694089802454023538387492997520114347332873807396492983274966274294831589088989087114050630219550508388528957090924299450523621088263633532944081602796696289920550855745518557779916320826471059885307179092435718801599456819799179186362425672999039326596225188275147042;
            5'd4: xpb[197] = 1024'd98863376225584715092699820024595447348858543536893728116805753367314623710669203105086576133749482827994492713757114275168861294734439623714624788620341926355061147874498496403130751569815199409260025806732487255653280455241699810056499456027609547136282068218504437592319501950183087397181254851334763185610;
            5'd5: xpb[197] = 1024'd61545872439918523166475311328337092813723965858249318081941264176654831969681934426350684559858016380271541188467646126671544697997439362365700923267261887476981097558337511835098319866510396400919933454221989146384420143941676376088135035192897209286942633566072017975346113400764542737917223650855656739847;
            5'd6: xpb[197] = 1024'd24228368654252331240250802632078738278589388179604908047076774985995040228694665747614792985966549932548589663178177978174228101260439101016777057914181848598901047242176527267065888163205593392579841101711491037115559832641652942119770614358184871437603198913639598358372724851345998078653192450376550294084;
            5'd7: xpb[197] = 1024'd110977560552710880712825221340634816488153237626696182140344140860312143825016535978893972626732757794268787545346203264255975345364659174223013317577432850654511671495586760036663695651417996105549946357588232774211060371562526281116384763206701982855083667675324236771505864375856086436507851076523038332652;
            5'd8: xpb[197] = 1024'd73660056767044688786600712644376461953018659948051772105479651669652352084029267300158081052841291346545836020056735115758658748627658912874089452224352811776431621179425775468631263948113193097209854005077734664942200060262502847148020342371989645005744233022891817154532475826437541777243819876043931886889;
            5'd9: xpb[197] = 1024'd36342552981378496860376203948118107417884082269407362070615162478992560343041998621422189478949824898822884494767266967261342151890658651525165586871272772898351570863264790900598832244808390088869761652567236555673339748962479413179655921537277307156404798370459397537559087277018997117979788675564825441126;
            5'd10: xpb[197] = 1024'd123091744879837046332950622656674185627447931716498636163882528353309663939363868852701369119716032760543082376935292253343089395994878724731401846534523774953962195116675023670196639733020792801839866908443978292768840287883352752176270070385794418573885267132144035950692226801529085475834447301711313479694;
            5'd11: xpb[197] = 1024'd85774241094170854406726113960415831092313354037854226129018039162649872198376600173965477545824566312820130851645824104845772799257878463382477981181443736075882144800514039102164208029715989793499774555933480183499979976583329318207905649551082080724545832479711616333718838252110540816570416101232207033931;
            5'd12: xpb[197] = 1024'd48456737308504662480501605264157476557178776359209816094153549971990080457389331495229585971933099865097179326356355956348456202520878202033554115828363697197802094484353054534131776326411186785159682203422982074231119665283305884239541228716369742875206397827279196716745449702691996157306384900753100588168;
            5'd13: xpb[197] = 1024'd11139233522838470554277096567899122022044198680565406059289060781330288716402062816493694398041633417374227801066887807851139605783877940684630250475283658319722044168192069966099344623106383776819589850912483964962259353983282450271176807881657405025866963174846777099772061153273451498042353700273994142405;
            5'd14: xpb[197] = 1024'd97888425421297020026851515276455200231608048127656680152556426655647392312723933047772874038807841279094425683234913093932886849888098013890866510138534660375332668421602302735697152111318786489789695106789225702057759892904155789267790956730174516443347431936531415512905200677783539855897012326420482180973;
            5'd15: xpb[197] = 1024'd60570921635630828100627006580196845696473470449012270117691937464987600571736664369036982464916374831371474157945444945435570253151097752541942644785454621497252618105441318167664720408013983481449602754278727592788899581604132355299426535895462178594007997284098995895931812128364995196632981125941375735210;
            5'd16: xpb[197] = 1024'd23253417849964636174402497883938491161338892770367860082827448274327808830749395690301090891024908383648522632655976796938253656414097491193018779432374582619172567789280333599632288704709180473109510401768229483520039270304108921331062115060749840744668562631666576278958423578946450537368949925462269289447;
            5'd17: xpb[197] = 1024'd110002609748423185646976916592494569370902742217459134176094814148644912427071265921580270531791116245368720514824002083020000900518317564399255039095625584674783192042690566369230096192921583186079615657644971220615539809224982260327676263909266952162149031393351214692091563103456538895223608551608757328015;
            5'd18: xpb[197] = 1024'd72685105962756993720752407896236214835768164538814724141230324957985120686083997242844378957899649797645768989534533934522684303781317303050331173742545545796703141726529581801197664489616780177739523305134473111346679497924958826359311843074554614312809596740918795075118174554037994235959577351129650882252;
            5'd19: xpb[197] = 1024'd35367602177090801794527899199977860300633586860170314106365835767325328945096728564108487384008183349922817464245065786025367707044317041701407308389465506918623091410368597233165232786311977169399430952623975002077819186624935392390947422239842276463470162088486375458144786004619449576695546150650544436489;
            5'd20: xpb[197] = 1024'd122116794075549351267102317908533938510197436307261588199633201641642432541418598795387667024774391211643015346413091072107114951148537114907643568052716508974233715663778830002763040274524379882369536208500716739173319725545808731387561571088359387880950630850171013871277925529129537934550204776797032475057;
            5'd21: xpb[197] = 1024'd84799290289883159340877809212275583975062858628617178164768712450982640800431330116651775450882924763920063821123622923609798354411536853558719702699636470096153665347617845434730608571219576874029443855990218629904459414245785297419197150253647050031611196197738594254304536979710993275286173576317926029294;
            5'd22: xpb[197] = 1024'd47481786504216967414653300516017229439928280949972768129904223260322849059444061437915883876991458316197112295834154775112481757674536592209795837346556431218073615031456860866698176867914773865689351503479720520635599102945761863450832729418934712182271761545306174637331148430292448616022142375838819583531;
            5'd23: xpb[197] = 1024'd10164282718550775488428791819758874904793703271328358095039734069663057318456792759179992303099991868474160770544686626615165160937536330860871971993476392339993564715295876298665745164609970857349259150969222411366738791645738429482468308584222374332932326892873755020357759880873903956758111175359713137768;
            5'd24: xpb[197] = 1024'd96913474617009324961003210528314953114357552718419632188307099943980160914778662990459171943866199730194358652712711912696912405041756404067108231656727394395604188968706109068263552652822373570319364406845964148462239330566611768479082457432739485750412795654558393433490899405383992314612769801506201176336;
            5'd25: xpb[197] = 1024'd59595970831343133034778701832056598579222975039775222153442610753320369173791394311723280369974733282471407127423243764199595808304756142718184366303647355517524138652545124500231120949517570561979272054335466039193379019266588334510718036598027147901073361002125973816517510855965447655348738601027094730573;
            5'd26: xpb[197] = 1024'd22278467045676941108554193135798244044088397361130812118578121562660577432804125632987388796083266834748455602133775615702279211567755881369260500950567316639444088336384139932198689246212767553639179701824967929924518707966564900542353615763314810051733926349693554199544122306546902996084707400547988284810;
            5'd27: xpb[197] = 1024'd109027658944135490581128611844354322253652246808222086211845487436977681029125995864266568436849474696468653484301800901784026455671975954575496760613818318695054712589794372701796496734425170266609284957701709667020019246887438239538967764611831921469214395111378192612677261831056991353939366026694476323378;
            5'd28: xpb[197] = 1024'd71710155158469298654904103148095967718517669129577676176980998246317889288138727185530676862958008248745701959012332753286709858934975693226572895260738279816974662273633388133764065031120367258269192605191211557751158935587414805570603343777119583619874960458945772995703873281638446694675334826215369877615;
            5'd29: xpb[197] = 1024'd34392651372803106728679594451837613183383091450933266142116509055658097547151458506794785289066541801022750433722864604789393262197975431877649029907658240938894611957472403565731633327815564249929100252680713448482298624287391371602238922942407245770535525806513353378730484732219902035411303625736263431852;
            5'd30: xpb[197] = 1024'd121141843271261656201254013160393691392946940898024540235383874929975201143473328738073964929832749662742948315890889890871140506302195505083885289570909242994505236210882636335329440816027966962899205508557455185577799163208264710598853071790924357188015994568197991791863624256729990393265962251882751470420;
            5'd31: xpb[197] = 1024'd83824339485595464275029504464135336857812363219380130200519385739315409402486060059338073355941283215019996790601421742373823909565195243734961424217829204116425185894721651767297009112723163954559113156046957076308938851908241276630488650956212019338676559915765572174890235707311445734001931051403645024657;
        endcase
    end



endmodule



module xpb_lut_final
(
    input logic [16:0] flag,
    output logic [1023:0] xpb[3]
);
        
        
    always_comb begin
        case(flag[5:0])
            6'd0: xpb[0] = 1024'd0;
            6'd1: xpb[0] = 1024'd55702617802106849374131591674088040617099270768494973145298226092755780468191824222693406107749861711676964472413899923079725927973196287937687305623143083444077218855294267938671980409728888398142885343697765922473789832121566108508934540857597787896530607270469240209840717864551083287716666502998629652885;
            6'd2: xpb[0] = 1024'd111405235604213698748263183348176081234198541536989946290596452185511560936383648445386812215499723423353928944827799846159451855946392575875374611246286166888154437710588535877343960819457776796285770687395531844947579664243132217017869081715195575793061214540938480419681435729102166575433333005997259305770;
            6'd3: xpb[0] = 1024'd43041157722195806723595847617449689106599385179749235307762823213290446067266333758065147108591910825587744009784206334660113943078368529257901791853098209398540981996311586478385702037669459473118458422706057921057008646143801552561825052889563914422771918397290662599415625519724616846031309682370294474324;
            6'd4: xpb[0] = 1024'd98743775524302656097727439291537729723698655948244208453061049306046226535458157980758553216341772537264708482198106257739839871051564817195589097476241292842618200851605854417057682447398347871261343766403823843530798478265367661070759593747161702319302525667759902809256343384275700133747976185368924127209;
            6'd5: xpb[0] = 1024'd30379697642284764073060103560811337596099499591003497470227420333825111666340843293436888109433959939498523547154512746240501958183540770578116278083053335353004745137328905018099423665610030548094031501714349919640227460166036996614715564921530040949013229524112084988990533174898150404345952861741959295763;
            6'd6: xpb[0] = 1024'd86082315444391613447191695234899378213198770359498470615525646426580892134532667516130294217183821651175488019568412669320227886156737058515803583706196418797081963992623172956771404075338918946236916845412115842114017292287603105123650105779127828845543836794581325198831251039449233692062619364740588948648;
            6'd7: xpb[0] = 1024'd17718237562373721422524359504172986085599614002257759632692017454359777265415352828808629110276009053409303084524819157820889973288713011898330764313008461307468508278346223557813145293550601623069604580722641918223446274188272440667606076953496167475254540650933507378565440830071683962660596041113624117202;
            6'd8: xpb[0] = 1024'd73420855364480570796655951178261026702698884770752732777990243547115557733607177051502035218025870765086267556938719080900615901261909299836018069936151544751545727133640491496485125703279490021212489924420407840697236106309838549176540617811093955371785147921402747588406158694622767250377262544112253770087;
            6'd9: xpb[0] = 1024'd5056777482462678771988615447534634575099728413512021795156614574894442864489862364180370111118058167320082621895125569401277988393885253218545250542963587261932271419363542097526866921491172698045177659730933916806665088210507884720496588985462294001495851777754929768140348485245217520975239220485288938641;
            6'd10: xpb[0] = 1024'd60759395284569528146120207121622675192198999182006994940454840667650223332681686586873776218867919878997047094309025492481003916367081541156232556166106670706009490274657810036198847331220061096188063003428699839280454920332073993229431129843060081898026459048224169977981066349796300808691905723483918591526;
            6'd11: xpb[0] = 1024'd116462013086676377520251798795710715809298269950501968085753066760406003800873510809567182326617781590674011566722925415560729844340277829093919861789249754150086709129952077974870827740948949494330948347126465761754244752453640101738365670700657869794557066318693410187821784214347384096408572226482548244411;
            6'd12: xpb[0] = 1024'd48097935204658485495584463064984323681699113593261257102919437788184888931756196122245517219709968992907826631679331904061391931472253782476447042396061796660473253415675128575912568959160632171163636082436991837863673734354309437282321641875026208424267770175045592367555974004969834367006548902855583412965;
            6'd13: xpb[0] = 1024'd103800553006765334869716054739072364298798384361756230248217663880940669399948020344938923327459830704584791104093231827141117859445450070414134348019204880104550472270969396514584549368889520569306521426134757760337463566475875545791256182732623996320798377445514832577396691869520917654723215405854213065850;
            6'd14: xpb[0] = 1024'd35436475124747442845048719008345972171199228004515519265384034908719554530830705657617258220552018106818606169049638315641779946577426023796661528626016922614937016556692447115626290587101203246139209161445283836446892548376544881335212153906992334950509081301867014757130881660143367925321192082227248234404;
            6'd15: xpb[0] = 1024'd91139092926854292219180310682434012788298498773010492410682261001475334999022529880310664328301879818495570641463538238721505874550622311734348834249160006059014235411986715054298270996830091644282094505143049758920682380498110989844146694764590122847039688572336254966971599524694451213037858585225877887289;
            6'd16: xpb[0] = 1024'd22775015044836400194512974951707620660699342415769781427848632029254220129905215192988999221394067220729385706419944727222167961682598265116876014855972048569400779697709765655340012215041774321114782240453575835030111362398780325388102665938958461476750392428688437146705789315316901483635835261598913055843;
            6'd17: xpb[0] = 1024'd78477632846943249568644566625795661277798613184264754573146858122010000598097039415682405329143928932406350178833844650301893889655794553054563320479115132013477998553004033594011992624770662719257667584151341757503901194520346433897037206796556249373280999699157677356546507179867984771352501764597542708728;
            6'd18: xpb[0] = 1024'd10113554964925357543977230895069269150199456827024043590313229149788885728979724728360740222236116334640165243790251138802555976787770506437090501085927174523864542838727084195053733842982345396090355319461867833613330176421015769440993177970924588002991703555509859536280696970490435041950478440970577877282;
            6'd19: xpb[0] = 1024'd65816172767032206918108822569157309767298727595519016735611455242544666197171548951054146329985978046317129716204151061882281904760966794374777806709070257967941761694021352133725714252711233794233240663159633756087120008542581877949927718828522375899522310825979099746121414835041518329667144943969207530167;
            6'd20: xpb[0] = 1024'd121518790569139056292240414243245350384397998364013989880909681335300446665363373173747552437735839757994094188618050984962007832734163082312465112332213341412018980549315620072397694662440122192376126006857399678560909840664147986458862259686120163796052918096448339955962132699592601617383811446967837183052;
            6'd21: xpb[0] = 1024'd53154712687121164267573078512518958256798842006773278898076052363079331796246058486425887330828027160227909253574457473462669919866139035694992292939025383922405524835038670673439435880651804869208813742167925754670338822564817322002818230860488502425763621952800522135696322490215051887981788123340872351606;
            6'd22: xpb[0] = 1024'd108857330489228013641704670186606998873898112775268252043374278455835112264437882709119293438577888871904873725988357396542395847839335323632679598562168467366482743690332938612111416290380693267351699085865691677144128654686383430511752771718086290322294229223269762345537040354766135175698454626339502004491;
            6'd23: xpb[0] = 1024'd40493252607210121617037334455880606746298956418027541060540649483613997395320568021797628331670076274138688790944763885043057934971311277015206779168980509876869287976055989213153157508592375944184386821176217753253557636587052766055708742892454628952004933079621944525271230145388585446296431302712537173045;
            6'd24: xpb[0] = 1024'd96195870409316970991168926129968647363398227186522514205838875576369777863512392244491034439419937985815653263358663808122783862944507564952894084792123593320946506831350257151825137918321264342327272164873983675727347468708618874564643283750052416848535540350091184735111948009939668734013097805711166825930;
            6'd25: xpb[0] = 1024'd27831792527299078966501590399242255235799070829281803223005246604148662994395077557169369332512125388049468328315070296623445950076483518335421265398935635831333051117073307752866879136532947019159959900184509751836776450609288210108599254924420755478246244206443366914846137800562119004611074482084201994484;
            6'd26: xpb[0] = 1024'd83534410329405928340633182073330295852898341597776776368303472696904443462586901779862775440261987099726432800728970219703171878049679806273108571022078719275410269972367575691538859546261835417302845243882275674310566282730854318617533795782018543374776851476912607124686855665113202292327740985082831647369;
            6'd27: xpb[0] = 1024'd15170332447388036315965846342603903725299185240536065385469843724683328593469587092541110333354174501960247865685376708203833965181655759655635751628890761785796814258090626292580600764473518094135532979192801750419995264631523654161489766956386882004487555333264789304421045455735652562925717661455866815923;
            6'd28: xpb[0] = 1024'd70872950249494885690097438016691944342398456009031038530768069817439109061661411315234516441104036213637212338099276631283559893154852047593323057252033845229874033113384894231252581174202406492278418322890567672893785096753089762670424307813984669901018162603734029514261763320286735850642384164454496468808;
            6'd29: xpb[0] = 1024'd2508872367476993665430102285965552214799299651790327547934440845217994192544096627912851334196223615871027403055683119784221980286828000975850237858845887740260577399107944832294322392414089169111106058201093749003214078653759098214380278988353008530728866460086211693995953110909186121240360840827531637362;
            6'd30: xpb[0] = 1024'd58211490169583843039561693960053592831898570420285300693232666937973774660735920850606257441946085327547991875469583042863947908260024288913537543481988971184337796254402212770966302802142977567253991401898859671477003910775325206723314819845950796427259473730555451903836670975460269408957027343826161290247;
            6'd31: xpb[0] = 1024'd113914107971690692413693285634141633448997841188780273838530893030729555128927745073299663549695947039224956347883482965943673836233220576851224849105132054628415015109696480709638283211871865965396876745596625593950793742896891315232249360703548584323790081001024692113677388840011352696673693846824790943132;
            6'd32: xpb[0] = 1024'd45550030089672800389025949903415241321398684831539562855697264058508440259810430385977998442788134441458771412839889454444335923365196530233752029711944097138801559395419531310680024430083548642229564480907151670060222724797560650776205331877916922953500784857376874293411578630633802967271670523197826111686;
            6'd33: xpb[0] = 1024'd101252647891779649763157541577503281938497955600034536000995490151264220728002254608671404550537996153135735885253789377524061851338392818171439335335087180582878778250713799249352004839812437040372449824604917592534012556919126759285139872735514710850031392127846114503252296495184886254988337026196455764571;
            6'd34: xpb[0] = 1024'd32888570009761757738490205846776889810898799242793825018161861179043105858884939921349739443630183555369550950210195866024723938470368771553966515941899223093265322536436849850393746058024119717205137559915443668643441538819796094829095843909883049479742095984198296682986486285807336525586313702569490933125;
            6'd35: xpb[0] = 1024'd88591187811868607112621797520864930427998070011288798163460087271798886327076764144043145551380045267046515422624095789104449866443565059491653821565042306537342541391731117789065726467753008115348022903613209591117231370941362203338030384767480837376272703254667536892827204150358419813302980205568120586010;
            6'd36: xpb[0] = 1024'd20227109929850715087954461790138538300398913654048087180626458299577771457959449456721480444472232669280330487580502277605111953575541012874181002171854349047729085677454168390107467685964690792180710638923735667226660352842031538881986355941849176005983407111019719072561393940980870083900956881941155754564;
            6'd37: xpb[0] = 1024'd75929727731957564462086053464226578917498184422543060325924684392333551926151273679414886552222094380957294959994402200684837881548737300811868307794997432491806304532748436328779448095693579190323595982621501589700450184963597647390920896799446963902514014381488959282402111805531953371617623384939785407449;
            6'd38: xpb[0] = 1024'd7565649849939672437418717733500186789899028065302349343091055420112437057033958992093221445314281783191110024950808689185499968680713254194395488401809475002192848818471486929821189313905261867156283717932027665809879166864266982934876867973815302532224718237841141462136301596154403642215600061312820576003;
            6'd39: xpb[0] = 1024'd63268267652046521811550309407588227406998298833797322488389281512868217525225783214786627553064143494868074497364708612265225896653909542132082794024952558446270067673765754868493169723634150265299169061629793588283668998985833091443811408831413090428755325508310381671977019460705486929932266564311450228888;
            6'd40: xpb[0] = 1024'd118970885454153371185681901081676268024097569602292295633687507605623997993417607437480033660814005206545038969778608535344951824627105830069770099648095641890347286529060022807165150133363038663442054405327559510757458831107399199952745949689010878325285932778779621881817737325256570217648933067310079881773;
            6'd41: xpb[0] = 1024'd50606807572135479161014565350949875896498413245051584650853878633402883124300292750158368553906192608778854034735015023845613911759081783452297280254907684400733830814783073408206891351574721340274742140638085586866887813008068535496701920863379216954996636635131804061551927115879020488246909743683115050327;
            6'd42: xpb[0] = 1024'd106309425374242328535146157025037916513597684013546557796152104726158663592492116972851774661656054320455818507148914946925339839732278071389984585878050767844811049670077341346878871761303609738417627484335851509340677645129634644005636461720977004851527243905601044271392644980430103775963576246681744703212;
            6'd43: xpb[0] = 1024'd37945347492224436510478821294311524385998527656305846813318475753937548723374802285530109554748241722689633572105321435426001926864254024772511766484862810355197593955800391947920612979515292415250315219646377585450106627030303979549592432895345343481237947761953226451126834771052554046561552923054779871766;
            6'd44: xpb[0] = 1024'd93647965294331285884610412968399565003097798424800819958616701846693329191566626508223515662498103434366598044519221358505727854837450312710199072108005893799274812811094659886592593389244180813393200563344143507923896459151870088058526973752943131377768555032422466660967552635603637334278219426053409524651;
            6'd45: xpb[0] = 1024'd25283887412313393859943077237673172875498642067560108975783072874472214322449311820901850555590290836600413109475627847006389941969426266092726252714817936309661357096817710487634334607455863490225888298654669584033325441052539423602482944927311470007479258888774648840701742426226087604876196102426444693205;
            6'd46: xpb[0] = 1024'd80986505214420243234074668911761213492597912836055082121081298967227994790641136043595256663340152548277377581889527770086115869942622554030413558337961019753738575952111978426306315017184751888368773642352435506507115273174105532111417485784909257904009866159243889050542460290777170892592862605425074346090;
            6'd47: xpb[0] = 1024'd12622427332402351209407333181034821364998756478814371138247669995006879921523821356273591556432339950511192646845934258586777957074598507412940738944773062264125120237835029027348056235396434565201461377662961582616544255074774867655373456959277596533720570015596071230276650081399621163190839281798109514644;
            6'd48: xpb[0] = 1024'd68325045134509200583538924855122861982098027247309344283545896087762660389715645578966997664182201662188157119259834181666503885047794795350628044567916145708202339093129296966020036645125322963344346721360727505090334087196340976164307997816875384430251177286065311440117367945950704450907505784796739167529;
            6'd49: xpb[0] = 1024'd124027662936616049957670516529210902599197298015804317428844122180518440857907469801660403771932063373865121591673734104746229813020991083288315350191059229152279557948423564904692017054854211361487232065058493427564123919317907084673242538674473172326781784556534551649958085810501787738624172287795368820414;
            6'd50: xpb[0] = 1024'd55663585054598157933003180798484510471598141658563606446010493208297325988790155114338738665024250776098936656630140593246891900152967036670842530797871271662666102234146615505733758273065894038319919800369019503673552901218576420217198509848841510956492488412886733829692275601124238009222148964168403988968;
            6'd51: xpb[0] = 1024'd111366202856705007307134772472572551088697412427058579591308719301053106456981979337032144772774112487775901129044040516326617828126163324608529836421014355106743321089440883444405738682794782436462805144066785426147342733340142528726133050706439298853023095683355974039532993465675321296938815467167033641853;
            6'd52: xpb[0] = 1024'd43002124974687115282467436741846158961098256069817868608475090328831991587864664649710479665866299890009716194000447004827279915258139277991057017027826397617129865375163934045447479901006465113295492879377311502256771715240811864270089021880807637482733799539708156219267183256297771567536792143540068810407;
            6'd53: xpb[0] = 1024'd98704742776793964656599028415934199578197526838312841753773316421587772056056488872403885773616161601686680666414346927907005843231335565928744322650969481061207084230458201984119460310735353511438378223075077424730561547362377972779023562738405425379264406810177396429107901120848854855253458646538698463292;
            6'd54: xpb[0] = 1024'd30340664894776072631931692685207807450598370481072130770939687449366657186939174185082220666708349003920495731370753416407667930363311519311271503257781523571593628516181252585161201528947036188271065958385603500839990529263047308322979533912773764008975110666529578608842090911471305125851435322911733631846;
            6'd55: xpb[0] = 1024'd86043282696882922006063284359295848067697641249567103916237913542122437655130998407775626774458210715597460203784653339487393858336507807248958808880924607015670847371475520523833181938675924586413951302083369423313780361384613416831914074770371551905505717936998818818682808776022388413568101825910363284731;
            6'd56: xpb[0] = 1024'd17679204814865029981395948628569455940098484892326392933404284569901322786013683720453961667550398117831275268741059827988055945468483760631485989487736649526057391657198571124874923156887607263246639037393895499423209343285282752375870045944739890535216421793351000998416998566644838684166078502283398453285;
            6'd57: xpb[0] = 1024'd73381822616971879355527540302657496557197755660821366078702510662657103254205507943147367775300259829508239741154959751067781873441680048569173295110879732970134610512492839063546903566616495661389524381091661421896999175406848860884804586802337678431747029063820241208257716431195921971882745005282028106170;
            6'd58: xpb[0] = 1024'd5017744734953987330860204571931104429598599303580655095868881690435988385088193255825702668392447231742054806111366239568443960573656001951700475717691775480521154798215889664588644784828178338222212116402187498006428157307518196428760557976706017061457732920172423387991906221818372242480721681655063274724;
            6'd59: xpb[0] = 1024'd60720362537060836704991796246019145046697870072075628241167107783191768853280017478519108776142308943419019278525266162648169888546852289889387781340834858924598373653510157603260625194557066736365097460099953420480217989429084304937695098834303804957988340190641663597832624086369455530197388184653692927609;
            6'd60: xpb[0] = 1024'd116422980339167686079123387920107185663797140840570601386465333875947549321471841701212514883892170655095983750939166085727895816520048577827075086963977942368675592508804425541932605604285955134507982803797719342954007821550650413446629639691901592854518947461110903807673341950920538817914054687652322580494;
            6'd61: xpb[0] = 1024'd48058902457149794054456052189380793536197984483329890403631704903726434452354527013890849776984358057329798815895572574228557903652024531209602267570789984879062136794527476142974346822497637811340670539108245419063436803451319748990585610866269931484229651317463085987407531741542989088512031364025357749048;
            6'd62: xpb[0] = 1024'd103761520259256643428587643863468834153297255251824863548929930996482214920546351236584255884734219769006763288309472497308283831625220819147289573193933068323139355649821744081646327232226526209483555882806011341537226635572885857499520151723867719380760258587932326197248249606094072376228697867023987401933;
            6'd63: xpb[0] = 1024'd35397442377238751403920308132742442025698098894584152566096302024261100051429036549262590777826407171240578353265878985808945918757196772529816753800745110833525899935544794682688068450438208886316243618116537417646655617473555193043476122898236058010470962444284508376982439396716522646826674543397022570487;
        endcase
    end

    always_comb begin
        case(flag[11:6])
            6'd0: xpb[1] = 1024'd0;
            6'd1: xpb[1] = 1024'd91100060179345600778051899806830482642797369663079125711394528117016880519620860771955996885576268882917542825679778908888671846730393060467504059423888194277603118790839062621360048860167097284459128961814303340120445449595121301552410663755833845907001569714753748586823157261267605934543341046395652223372;
            6'd2: xpb[1] = 1024'd58133424674566460157304872208846532540896312200422567294657201169056865701932582633896922556494863456391936243902064383198279852619565786379847993831445347621515563012106907905089858528816988847608060315241366833876530048969345830139842757828438242547183236015390439143539786448606578851967992266165709962413;
            6'd3: xpb[1] = 1024'd25166789169787319536557844610862582438995254737766008877919874221096850884244304495837848227413458029866329662124349857507887858508738512292191928239002500965428007233374753188819668197466880410756991668668430327632614648343570358727274851901042639187364902316027129700256415635945551769392643485935767701454;
            6'd4: xpb[1] = 1024'd116266849349132920314609744417693065081792624400845134589314402338113731403865165267793845112989726912783872487804128766396559705239131572759695987662890695243031126024213815810179717057633977695216120630482733667753060097938691660279685515656876485094366472030780878287079572897213157703935984532331419924826;
            6'd5: xpb[1] = 1024'd83300213844353779693862716819709114979891566938188576172577075390153716586176887129734770783908321486258265906026414240706167711128304298672039922070447848586943570245481661093909526726283869258365051983909797161509144697312916188867117609729480881734548138331417568843796202084552130621360635752101477663867;
            6'd6: xpb[1] = 1024'd50333578339574639073115689221725164877990509475532017755839748442193701768488608991675696454826916059732659324248699715015775717017477024584383856478005001930856014466749506377639336394933760821513983337336860655265229296687140717454549703802085278374729804632054259400512831271891103538785286971871535402908;
            6'd7: xpb[1] = 1024'd17366942834795498452368661623741214776089452012875459339102421494233686950800330853616622125745510633207052742470985189325383722906649750496727790885562155274768458688017351661369146063583652384662914690763924149021313896061365246041981797874689675014911470932690949957229460459230076456209938191641593141949;
            6'd8: xpb[1] = 1024'd108467003014141099230420561430571697418886821675954585050496949611250567470421191625572619011321779516124595568150764098214055569637042810964231850309450349552371577478856414282729194923750749669122043652578227489141759345656486547594392461630523520921913040647444698544052617720497682390753279238037245365321;
            6'd9: xpb[1] = 1024'd75500367509361958609673533832587747316985764213298026633759622663290552652732913487513544682240374089598988986373049572523663575526215536876575784717007502896284021700124259566459004592400641232270975006005290982897843945030711076181824555703127917562094706948081389100769246907836655308177930457807303104362;
            6'd10: xpb[1] = 1024'd42533732004582817988926506234603797215084706750641468217022295715330537835044635349454470353158968663073382404595335046833271581415388262788919719124564656240196465921392104850188814261050532795419906359432354476653928544404935604769256649775732314202276373248718079657485876095175628225602581677577360843403;
            6'd11: xpb[1] = 1024'd9567096499803677368179478636619847113183649287984909800284968767370523017356357211395396024077563236547775822817620521142879587304560988701263653532121809584108910142659950133918623929700424358568837712859417970410013143779160133356688743848336710842458039549354770214202505282514601143027232897347418582444;
            6'd12: xpb[1] = 1024'd100667156679149278146231378443450329755981018951064035511679496884387403536977217983351392909653832119465318648497399430031551434034954049168767712956010003861712028933499012755278672789867521643027966674673721310530458593374281434909099407604170556749459609264108518801025662543782207077570573943743070805816;
            6'd13: xpb[1] = 1024'd67700521174370137525484350845466379654079961488407477094942169936427388719288939845292318580572426692939712066719684904341159439924126775081111647363567157205624473154766858039008482458517413206176898028100784804286543192748505963496531501676774953389641275564745209357742291731121179994995225163513128544857;
            6'd14: xpb[1] = 1024'd34733885669590996904737323247482429552178904025750918678204842988467373901600661707233244251491021266414105484941970378650767445813299500993455581771124310549536917376034703322738292127167304769325829381527848298042627792122730492083963595749379350029822941865381899914458920918460152912419876383283186283898;
            6'd15: xpb[1] = 1024'd1767250164811856283990295649498479450277846563094360261467516040507359083912383569174169922409615839888498903164255852960375451702472226905799516178681463893449361597302548606468101795817196332474760734954911791798712391496955020671395689821983746670004608166018590471175550105799125829844527603053244022939;
            6'd16: xpb[1] = 1024'd92867310344157457062042195456328962093075216226173485972862044157524239603533244341130166807985884722806041728844034761849047298432865287373303575602569658171052480388141611227828150655984293616933889696769215131919157841092076322223806353577817592577006177880772339057998707367066731764387868649448896246311;
            6'd17: xpb[1] = 1024'd59900674839378316441295167858345011991174158763516927556124717209564224785844966203071092478904479296280435147066320236158655304322038013285647510010126811514964924609409456511557960324634185180082821050196278625675242440466300850811238447650421989217187844181409029614715336554405704681812519869218953985352;
            6'd18: xpb[1] = 1024'd26934039334599175820548140260361061889273101300860369139387390261604209968156688065012018149823073869754828565288605710468263310211210739197991444417683964858877368830677301795287769993284076743231752403623342119431327039840525379398670541723026385857369510482045720171431965741744677599237171088989011724393;
            6'd19: xpb[1] = 1024'd118034099513944776598600040067191544532070470963939494850781918378621090487777548836968015035399342752672371390968384619356935156941603799665495503841572159136480487621516364416647818853451174027690881365437645459551772489435646680951081205478860231764371080196799468758255123003012283533780512135384663947765;
            6'd20: xpb[1] = 1024'd85067464009165635977853012469207594430169413501282936434044591430661075670089270698908940706317937326146764809190670093666543162830776525577839438249129312480392931842784209700377628522101065590839812718864708953307857088809871209538513299551464628404552746497436159314971752190351256451205163355154721686806;
            6'd21: xpb[1] = 1024'd52100828504386495357105984871223644328268356038626378017307264482701060852400992560849866377236531899621158227412955567976151168719949251490183372656686465824305376064052054984107438190750957153988744072291772447063941688184095738125945393624069025044734412798072849871688381377690229368629814574924779425847;
            6'd22: xpb[1] = 1024'd19134192999607354736358957273239694226367298575969819600569937534741046034712714422790792048155126473095551645635241042285759174609121977402527307064243619168217820285319900267837247859400848717137675425718835940820026287558320266713377487696673421684916079098709540428405010565029202286054465794694837164888;
            6'd23: xpb[1] = 1024'd110234253178952955514410857080070176869164668239048945311964465651757926554333575194746788933731395356013094471315019951174431021339515037870031366488131813445820939076158962889197296719567946001596804387533139280940471737153441568265788151452507267591917648813463289015228167826296808220597806841090489388260;
            6'd24: xpb[1] = 1024'd77267617674173814893663829482086226767263610776392386895227138703797911736645297056687714604649989929487487889537305425484039027228687763782375300895688966789733383297426808172927106388217837564745735740960202774696556336527666096853220245525111664232099315114099979571944797013635781138022458060860547127301;
            6'd25: xpb[1] = 1024'd44300982169394674272916801884102276665362553313735828478489811755837896918957018918628640275568584502961881307759590899793647033117860489694719235303246120133645827518694653456656916056867729127894667094387266268452640935901890625440652339597716060872280981414736670128661426200974754055447109280630604866342;
            6'd26: xpb[1] = 1024'd11334346664615533652169774286118326563461495851079270061752484807877882101268740780569565946487179076436274725981876374103255039007033215607063169710803273477558271739962498740386725725517620691043598447814329762208725535276115154028084433670320457512462647715373360685378055388313726972871760500400662605383;
            6'd27: xpb[1] = 1024'd102434406843961134430221674092948809206258865514158395773147012924894762620889601552525562832063447959353817551661655282991926885737426276074567229134691467755161390530801561361746774585684717975502727409628633102329170984871236455580495097426154303419464217430127109272201212649581332907415101546796314828755;
            6'd28: xpb[1] = 1024'd69467771339181993809474646494964859104357808051501837356409685976934747803201323414466488502982042532828210969883940757301534891626599001986911163542248621099073834752069406645476584254334609538651658763055696596085255584245460984167927191498758700059645883730763799828917841836920305824839752766566372567796;
            6'd29: xpb[1] = 1024'd36501135834402853188727618896980909002456750588845278939672359028974732985513045276407414173900637106302604388106226231611142897515771727899255097949805774442986278973337251929206393922984501101800590116482760089841340183619685512755359285571363096699827550031400490385634471024259278742264403986336430306837;
            6'd30: xpb[1] = 1024'd3534500329623712567980591298996958900555693126188720522935032081014718167824767138348339844819231679776997806328511705920750903404944453811599032357362927786898723194605097212936203591634392664949521469909823583597424782993910041342791379643967493340009216332037180942351100211598251659689055206106488045878;
            6'd31: xpb[1] = 1024'd94634560508969313346032491105827441543353062789267846234329560198031598687445627910304336730395500562694540632008290614809422750135337514279103091781251122064501841985444159834296252451801489949408650431724126923717870232589031342895202043399801339247010786046790929529174257472865857594232396252502140269250;
            6'd32: xpb[1] = 1024'd61667925004190172725285463507843491441452005326611287817592233250071583869757349772245262401314095136168934050230576089119030756024510240191447026188808275408414286206712005118026062120451381512557581785151190417473954831963255871482634137472405735887192452347427620085890886660204830511657047472272198008291;
            6'd33: xpb[1] = 1024'd28701289499411032104538435909859541339550947863954729400854906302111569052069071634186188072232689709643327468452861563428638761913682966103790960596365428752326730427979850401755871789101273075706513138578253911230039431337480400070066231545010132527374118648064310642607515847543803429081698692042255747332;
            6'd34: xpb[1] = 1024'd119801349678756632882590335716690023982348317527033855112249434419128449571689932406142184957808958592560870294132640472317310608644076026571295020020253623029929849218818913023115920649268370360165642100392557251350484880932601701622476895300843978434375688362818059229430673108811409363625039738437907970704;
            6'd35: xpb[1] = 1024'd86834714173977492261843308118706073880447260064377296695512107471168434754001654268083110628727553166035263712354925946626918614533248752483638954427810776373842293440086758306845730317918261923314573453819620745106569480306826230209908989373448375074557354663454749786147302296150382281049690958207965709745;
            6'd36: xpb[1] = 1024'd53868078669198351641096280520722123778546202601720738278774780523208419936313376130024036299646147739509657130577211420936526620422421478395982888835367929717754737661354603590575539986568153486463504807246684238862654079681050758797341083446052771714739020964091440342863931483489355198474342177978023448786;
            6'd37: xpb[1] = 1024'd20901443164419211020349252922738173676645145139064179862037453575248405118625097991964961970564742312984050548799496895246134626311594204308326823242925083061667181882622448874305349655218045049612436160673747732618738679055275287384773177518657168354920687264728130899580560670828328115898993397748081187827;
            6'd38: xpb[1] = 1024'd112001503343764811798401152729568656319442514802143305573431981692265285638245958763920958856141011195901593374479275804134806473041987264775830882666813277339270300673461511495665398515385142334071565122488051072739184128650396588937183841274491014261922256979481879486403717932095934050442334444143733411199;
            6'd39: xpb[1] = 1024'd79034867838985671177654125131584706217541457339486747156694654744305270820557680625861884527059605769375986792701561278444414478931159990688174817074370430683182744894729356779395208184035033897220496475915114566495268728024621117524615935347095410902103923280118570043120347119434906967866985663913791150240;
            6'd40: xpb[1] = 1024'd46068232334206530556907097533600756115640399876830188739957327796345256002869402487802810197978200342850380210923846752754022484820332716600518751481927584027095189115997202063125017852684925460369427829342178060251353327398845646112048029419699807542285589580755260599836976306773879885291636883683848889281;
            6'd41: xpb[1] = 1024'd13101596829427389936160069935616806013739342414173630323220000848385241185181124349743735868896794916324773629146132227063630490709505442512862685889484737371007633337265047346854827521334817023518359182769241554007437926773070174699480123492304204182467255881391951156553605494112852802716288103453906628322;
            6'd42: xpb[1] = 1024'd104201657008772990714211969742447288656536712077252756034614528965402121704801985121699732754473063799242316454825911135952302337439898502980366745313372931648610752128104109968214876381501914307977488144583544894127883376368191476251890787248138050089468825596145699743376762755380458737259629149849558851694;
            6'd43: xpb[1] = 1024'd71235021503993850093464942144463338554635654614596197617877202017442106887113706983640658425391658372716709873048196610261910343329071228892710679720930084992523196349371955251944686050151805871126419498010608387883967975742416004839322881320742446729650491896782390300093391942719431654684280369619616590735;
            6'd44: xpb[1] = 1024'd38268385999214709472717914546479388452734597151939639201139875069482092069425428845581584096310252946191103291270482084571518349218243954805054614128487238336435640570639800535674495718801697434275350851437671881640052575116640533426754975393346843369832158197419080856810021130058404572108931589389674329776;
            6'd45: xpb[1] = 1024'd5301750494435568851970886948495438350833539689283080784402548121522077251737150707522509767228847519665496709492767558881126355107416680717398548536044391680348084791907645819404305387451588997424282204864735375396137174490865062014187069465951240010013824498055771413526650317397377489533582809159732068817;
            6'd46: xpb[1] = 1024'd96401810673781169630022786755325920993630909352362206495797076238538957771358011479478506652805116402583039535172546467769798201837809741184902607959932585957951203582746708440764354247618686281883411166679038715516582624085986363566597733221785085917015394212809520000349807578664983424076923855555384292189;
            6'd47: xpb[1] = 1024'd63435175169002029009275759157341970891729851889705648079059749290578942953669733341419432323723710976057432953394831942079406207726982467097246542367489739301863647804014553724494163916268577845032342520106102209272667223460210892154029827294389482557197060513446210557066436766003956341501575075325442031230;
            6'd48: xpb[1] = 1024'd30468539664222888388528731559358020789828794427049089662322422342618928135981455203360357994642305549531826371617117416389014213616155193009590476775046892645776092025282399008223973584918469408181273873533165703028751822834435420741461921366993879197378726814082901113783065953342929258926226295095499770271;
            6'd49: xpb[1] = 1024'd121568599843568489166580631366188503432626164090128215373716950459635808655602315975316354880218574432449369197296896325277686060346548253477094536198935086923379210816121461629584022445085566692640402835347469043149197272429556722293872585122827725104380296528836649700606223214610535193469567341491151993643;
            6'd50: xpb[1] = 1024'd88601964338789348545833603768204553330725106627471656956979623511675793837914037837257280551137169005923762615519181799587294066235720979389438470606492240267291655037389306913313832113735458255789334188774532536905281871803781250881304679195432121744561962829473340257322852401949508110894218561261209732684;
            6'd51: xpb[1] = 1024'd55635328834010207925086576170220603228824049164815098540242296563715779020225759699198206222055763579398156033741467273896902072124893705301782405014049393611204099258657152197043641782385349818938265542201596030661366471178005779468736773268036518384743629130110030814039481589288481028318869781031267471725;
            6'd52: xpb[1] = 1024'd22668693329231067304339548572236653126922991702158540123504969615755764202537481561139131892974358152872549451963752748206510078014066431214126339421606546955116543479924997480773451451035241382087196895628659524417451070552230308056168867340640915024925295430746721370756110776627453945743521000801325210766;
            6'd53: xpb[1] = 1024'd113768753508576668082391448379067135769720361365237665834899497732772644722158342333095128778550627035790092277643531657095181924744459491681630398845494741232719662270764060102133500311202338666546325857442962864537896520147351609608579531096474760931926865145500469957579268037895059880286862047196977434138;
            6'd54: xpb[1] = 1024'd80802118003797527461644420781083185667819303902581107418162170784812629904470064195036054449469221609264485695865817131404789930633632217593974333253051894576632106492031905385863309979852230229695257210870026358293981119521576138196011625169079157572108531446137160514295897225234032797711513266967035173179;
            6'd55: xpb[1] = 1024'd47835482499018386840897393183099235565918246439924549001424843836852615086781786056976980120387816182738879114088102605714397936522804943506318267660609047920544550713299750669593119648502121792844188564297089852050065718895800666783443719241683554212290197746773851071012526412573005715136164486737092912220;
            6'd56: xpb[1] = 1024'd14868846994239246220150365585115285464017188977267990584687516888892600269093507918917905791306410756213272532310388080024005942411977669418662202068166201264456994934567595953322929317152013355993119917724153345806150318270025195370875813314287950852471864047410541627729155599911978632560815706507150651261;
            6'd57: xpb[1] = 1024'd105968907173584846998202265391945768106814558640347116296082045005909480788714368690873902676882679639130815357990166988912677789142370729886166261492054395542060113725406658574682978177319110640452248879538456685926595767865146496923286477070121796759473433762164290214552312861179584567104156752902802874633;
            6'd58: xpb[1] = 1024'd73002271668805706377455237793961818004913501177690557879344718057949465971026090552814828347801274212605208776212452463222285795031543455798510195899611548885972557946674503858412787845969002203601180232965520179682680367239371025510718571142726193399655100062800980771268942048518557484528807972672860613674;
            6'd59: xpb[1] = 1024'd40035636164026565756708210195977867903012443715033999462607391109989451153337812414755754018719868786079602194434737937531893800920716181710854130307168702229885002167942349142142597514618893766750111586392583673438764966613595554098150665215330590039836766363437671327985571235857530401953459192442918352715;
            6'd60: xpb[1] = 1024'd7069000659247425135961182597993917801111386252377441045870064162029436335649534276696679689638463359553995612657023411841501806809888907623198064714725855573797446389210194425872407183268785329899042939819647167194849565987820082685582759287934986680018432664074361884702200423196503319378110412212976091756;
            6'd61: xpb[1] = 1024'd98169060838593025914013082404824400443908755915456566757264592279046316855270395048652676575214732242471538438336802320730173653540281968090702124138614049851400565180049257047232456043435882614358171901633950507315295015582941384237993423043768832587020002378828110471525357684464109253921451458608628315128;
            6'd62: xpb[1] = 1024'd65202425333813885293266054806840450342007698452800008340527265331086302037582116910593602246133326815945931856559087795039781659429454694003046058546171203195313009401317102330962265712085774177507103255061014001071379614957165912825425517116373229227201668679464801028241986871803082171346102678378686054169;
            6'd63: xpb[1] = 1024'd32235789829034744672519027208856500240106640990143449923789938383126287219893838772534527917051921389420325274781373269349389665318627419915389992953728356539225453622584947614692075380735665740656034608488077494827464214331390441412857611188977625867383334980101491584958616059142055088770753898148743793210;
        endcase
    end

    always_comb begin
        case(flag[16:12])
            5'd0: xpb[2] = 1024'd0;
            5'd1: xpb[2] = 1024'd123335850008380345450570927015686982882904010653222575635184466500143167739514699544490524802628190272337868100461152178238061512049020480382894052377616550816828572413424010236052124240902763025115163570302380834947909663926511742965268274944811471774384904694855240171781773320409661023314094944544396016582;
            5'd2: xpb[2] = 1024'd122605004332635949502342926626559533021109594180709467142237077935309440141720260178965978390598706235232586793464810921897059183256820626210627979738902060699966470257276803134474009290288320328920129532217521823531458477632126712965557980206393494281949905975593422313457018566890689029509500062463197548833;
            5'd3: xpb[2] = 1024'd121874158656891553554114926237432083159315177708196358649289689370475712543925820813441431978569222198127305486468469665556056854464620772038361907100187570583104368101129596032895894339673877632725095494132662812115007291337741682965847685467975516789514907256331604455132263813371717035704905180381999081084;
            5'd4: xpb[2] = 1024'd121143312981147157605886925848304633297520761235683250156342300805641984946131381447916885566539738161022024179472128409215054525672420917866095834461473080466242265944982388931317779389059434936530061456047803800698556105043356652966137390729557539297079908537069786596807509059852745041900310298300800613335;
            5'd5: xpb[2] = 1024'd120412467305402761657658925459177183435726344763170141663394912240808257348336942082392339154510254123916742872475787152874052196880221063693829761822758590349380163788835181829739664438444992240335027417962944789282104918748971622966427095991139561804644909817807968738482754306333773048095715416219602145586;
            5'd6: xpb[2] = 1024'd119681621629658365709430925070049733573931928290657033170447523675974529750542502716867792742480770086811461565479445896533049868088021209521563689184044100232518061632687974728161549487830549544139993379878085777865653732454586592966716801252721584312209911098546150880157999552814801054291120534138403677837;
            5'd7: xpb[2] = 1024'd118950775953913969761202924680922283712137511818143924677500135111140802152748063351343246330451286049706180258483104640192047539295821355349297616545329610115655959476540767626583434537216106847944959341793226766449202546160201562967006506514303606819774912379284333021833244799295829060486525652057205210088;
            5'd8: xpb[2] = 1024'd118219930278169573812974924291794833850343095345630816184552746546307074554953623985818699918421802012600898951486763383851045210503621501177031543906615119998793857320393560525005319586601664151749925303708367755032751359865816532967296211775885629327339913660022515163508490045776857066681930769976006742339;
            5'd9: xpb[2] = 1024'd117489084602425177864746923902667383988548678873117707691605357981473346957159184620294153506392317975495617644490422127510042881711421647004765471267900629881931755164246353423427204635987221455554891265623508743616300173571431502967585917037467651834904914940760697305183735292257885072877335887894808274590;
            5'd10: xpb[2] = 1024'd116758238926680781916518923513539934126754262400604599198657969416639619359364745254769607094362833938390336337494080871169040552919221792832499398629186139765069653008099146321849089685372778759359857227538649732199848987277046472967875622299049674342469916221498879446858980538738913079072741005813609806841;
            5'd11: xpb[2] = 1024'd116027393250936385968290923124412484264959845928091490705710580851805891761570305889245060682333349901285055030497739614828038224127021938660233325990471649648207550851951939220270974734758336063164823189453790720783397800982661442968165327560631696850034917502237061588534225785219941085268146123732411339092;
            5'd12: xpb[2] = 1024'd115296547575191990020062922735285034403165429455578382212763192286972164163775866523720514270303865864179773723501398358487035895334822084487967253351757159531345448695804732118692859784143893366969789151368931709366946614688276412968455032822213719357599918782975243730209471031700969091463551241651212871343;
            5'd13: xpb[2] = 1024'd114565701899447594071834922346157584541371012983065273719815803722138436565981427158195967858274381827074492416505057102146033566542622230315701180713042669414483346539657525017114744833529450670774755113284072697950495428393891382968744738083795741865164920063713425871884716278181997097658956359570014403594;
            5'd14: xpb[2] = 1024'd113834856223703198123606921957030134679576596510552165226868415157304708968186987792671421446244897789969211109508715845805031237750422376143435108074328179297621244383510317915536629882915007974579721075199213686534044242099506352969034443345377764372729921344451608013559961524663025103854361477488815935845;
            5'd15: xpb[2] = 1024'd113104010547958802175378921567902684817782180038039056733921026592470981370392548427146875034215413752863929802512374589464028908958222521971169035435613689180759142227363110813958514932300565278384687037114354675117593055805121322969324148606959786880294922625189790155235206771144053110049766595407617468096;
            5'd16: xpb[2] = 1024'd112373164872214406227150921178775234955987763565525948240973638027637253772598109061622328622185929715758648495516033333123026580166022667798902962796899199063897040071215903712380399981686122582189652999029495663701141869510736292969613853868541809387859923905927972296910452017625081116245171713326419000347;
            5'd17: xpb[2] = 1024'd111642319196470010278922920789647785094193347093012839748026249462803526174803669696097782210156445678653367188519692076782024251373822813626636890158184708947034937915068696610802285031071679885994618960944636652284690683216351262969903559130123831895424925186666154438585697264106109122440576831245220532598;
            5'd18: xpb[2] = 1024'd110911473520725614330694920400520335232398930620499731255078860897969798577009230330573235798126961641548085881523350820441021922581622959454370817519470218830172835758921489509224170080457237189799584922859777640868239496921966232970193264391705854402989926467404336580260942510587137128635981949164022064849;
            5'd19: xpb[2] = 1024'd110180627844981218382466920011392885370604514147986622762131472333136070979214790965048689386097477604442804574527009564100019593789423105282104744880755728713310733602774282407646055129842794493604550884774918629451788310627581202970482969653287876910554927748142518721936187757068165134831387067082823597100;
            5'd20: xpb[2] = 1024'd109449782169236822434238919622265435508810097675473514269184083768302343381420351599524142974067993567337523267530668307759017264997223251109838672242041238596448631446627075306067940179228351797409516846690059618035337124333196172970772674914869899418119929028880700863611433003549193141026792185001625129351;
            5'd21: xpb[2] = 1024'd108718936493492426486010919233137985647015681202960405776236695203468615783625912233999596562038509530232241960534327051418014936205023396937572599603326748479586529290479868204489825228613909101214482808605200606618885938038811142971062380176451921925684930309618883005286678250030221147222197302920426661602;
            5'd22: xpb[2] = 1024'd107988090817748030537782918844010535785221264730447297283289306638634888185831472868475050150009025493126960653537985795077012607412823542765306526964612258362724427134332661102911710277999466405019448770520341595202434751744426112971352085438033944433249931590357065146961923496511249153417602420839228193853;
            5'd23: xpb[2] = 1024'd107257245142003634589554918454883085923426848257934188790341918073801160588037033502950503737979541456021679346541644538736010278620623688593040454325897768245862324978185454001333595327385023708824414732435482583785983565450041082971641790699615966940814932871095247288637168742992277159613007538758029726104;
            5'd24: xpb[2] = 1024'd106526399466259238641326918065755636061632431785421080297394529508967432990242594137425957325950057418916398039545303282395007949828423834420774381687183278129000222822038246899755480376770581012629380694350623572369532379155656052971931495961197989448379934151833429430312413989473305165808412656676831258355;
            5'd25: xpb[2] = 1024'd105795553790514842693098917676628186199838015312907971804447140944133705392448154771901410913920573381811116732548962026054005621036223980248508309048468788012138120665891039798177365426156138316434346656265764560953081192861271022972221201222780011955944935432571611571987659235954333172003817774595632790606;
            5'd26: xpb[2] = 1024'd105064708114770446744870917287500736338043598840394863311499752379299977794653715406376864501891089344705835425552620769713003292244024126076242236409754297895276018509743832696599250475541695620239312618180905549536630006566885992972510906484362034463509936713309793713662904482435361178199222892514434322857;
            5'd27: xpb[2] = 1024'd104333862439026050796642916898373286476249182367881754818552363814466250196859276040852318089861605307600554118556279513372000963451824271903976163771039807778413916353596625595021135524927252924044278580096046538120178820272500962972800611745944056971074937994047975855338149728916389184394628010433235855108;
            5'd28: xpb[2] = 1024'd103603016763281654848414916509245836614454765895368646325604975249632522599064836675327771677832121270495272811559938257030998634659624417731710091132325317661551814197449418493443020574312810227849244542011187526703727633978115932973090317007526079478639939274786157997013394975397417190590033128352037387359;
            5'd29: xpb[2] = 1024'd102872171087537258900186916120118386752660349422855537832657586684798795001270397309803225265802637233389991504563597000689996305867424563559444018493610827544689712041302211391864905623698367531654210503926328515287276447683730902973380022269108101986204940555524340138688640221878445196785438246270838919610;
            5'd30: xpb[2] = 1024'd102141325411792862951958915730990936890865932950342429339710198119965067403475957944278678853773153196284710197567255744348993977075224709387177945854896337427827609885155004290286790673083924835459176465841469503870825261389345872973669727530690124493769941836262522280363885468359473202980843364189640451861;
            5'd31: xpb[2] = 1024'd101410479736048467003730915341863487029071516477829320846762809555131339805681518578754132441743669159179428890570914488007991648283024855214911873216181847310965507729007797188708675722469482139264142427756610492454374075094960842973959432792272147001334943117000704422039130714840501209176248482108441984112;
        endcase
    end



endmodule




module xpb_5_185
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h78d589ea10ce609e16a1e34b169f58c2f74e08cf6bf71b7bd02bc775570bc40026c9fdeeb2b883274cc25d3ea3da4f2123c6b1c6af4a438f275d620b6b7e4bdc54a88fa6895df379cec07c489d3a820a2b3807db01fffd63afa649e05db0d52ce6bc69d6a3fe4d444455fe0dcef9c81c1e82872d5dae3c6a3b078463bc22862d;
    5'b00010 : xpb = 1024'h40fdce7e5fae8c73623e4ebf1ce46a347d260e6e02769680227ad594fb14daf84a4b7e649b4a87bffa267b3664568d77e3733ba73be1b6d29e1b84b89c2a23073501ea9e632ae9ae8ae6f5eea1993fe3626b161d7779cdb6a9c001c6013707c79e7141839733a1fb01ec153ca6236a0eee2b2f786b111ba42f9f8dc2ef62a5ef;
    5'b00011 : xpb = 1024'h9261312ae8eb848addaba3323297ba602fe140c98f6118474c9e3b49f1df1f06dccfeda83dc8c58a78a992e24d2cbcea31fc587c8792a1614d9a765ccd5fa32155b45963cf7dfe3470d6f94a5f7fdbc999e245fecf39e09a3d9b9aba4bd3a62562619308a68f6b1bf822c6b7d4d0c01bdd3d7c37873fade2437972222a2c5b1;
    5'b00100 : xpb = 1024'h81fb9cfcbf5d18e6c47c9d7e39c8d468fa4c1cdc04ed2d0044f5ab29f629b5f09496fcc936950f7ff44cf66cc8ad1aefc6e6774e77c36da53c3709713854460e6a03d53cc655d35d15cdebdd43327fc6c4d62c3aeef39b6d5380038c026e0f8f3ce283072e6743f603d82a794c46d41ddc565ef0d62237485f3f1b85dec54bde;
    5'b00101 : xpb = 1024'h4a23e1910e3d44bc101908f2400de5da8024227a9b6ca8049744b9499a32cce8b8187d3f1f271418a1b11464892959468693012f045ae0e8b2f52c1e69001d394a5d3034a022c991d1f4658347913d9ffc093a7d646d6bc04d99bb71a5f44229f4975ab4219c98acc16e41a823707610abff073be385168253d724e512056ba0;
    5'b00110 : xpb = 1024'h124c26255d1d70915bb574664652f74c05fc281931ec2308e993c7693e3be3e0db99fdb507b918b14f15325c49a5979d463f8b0f90f2542c29b34ecb99abf4642ab68b2c79efbfc68e1adf294beffb79333c48bfd9e73c1347b37357497a74c4ac4c326114d1ed637f0458d6fa9a18037ba7af86f0e7f5bc486f2e4445458b62;
    5'b00111 : xpb = 1024'h8b21b00f6debd12f725757b15cf2500efd4a30e89de33e84b9bf8ede9547a7e10263fba3ba719bd89bd78f9aed7fe6be6a063cd6403c97bb5110b0d7052a40407f5f1ad3034db3405cdb5b71e92a7d835e74509adbe73976f759bd37a72b49f193089c37b8d03aa7c35a56e4c993e01f9a2a36b44e9632268376b2a80168118f;
    5'b01000 : xpb = 1024'h5349f4a3bccbfd04bdf3c32563376180832236873462b9890c0e9cfe3950bed925e57c19a303a071493bad92adfc251529b2c6b6ccd40afec7ced38435d6176b5fb875cadd1aa9751901d517ed893b5c95a75edd516109c9f173751d4ab17c8c4abd73e4ac058f5e80f06e13a0bd821269d2deff5bf91160780ebc0734a83151;
    5'b01001 : xpb = 1024'h1b7239380bac28da09902e99697c72f208fa3c25cae2348d5e5dab1ddd59d5d14966fc8f8b95a509f69fcb8a6e78636be95f5097596b7e423e8cf6316681ee964011d0c2b6e79fa9d5284ebdf1e7f935ccda6d1fc6dada1ceb8d2d02ee37af2702724b919f3ae4153e86854277e72405397b874a695bf09a6ca6c56667e85113;
    5'b01010 : xpb = 1024'h9447c3221c7a8978203211e4801bcbb5004844f536d950092e897293346599d17030fa7e3e4e2831436228c91252b28d0d26025e08b5c1d165ea583cd2003a7294ba606940459323a3e8cb068f227b3ff81274fac8dad7809b3376e34be88453e92eb5684339315982dc835046e0ec2157fe0e77c70a2d04a7ae49ca240ad740;
    5'b01011 : xpb = 1024'h5c7007b66b5ab54d6bce7d588660dd2686204a93cd58cb0d80d880b2d86eb0c993b27af426e02cc9f0c646c0d2cef0e3ccd28c3e954d3514dca87aea02ac119d7513bb611a128958600f44ac938139192f45833d3e54a7d3954d2ec8ef6eb6eea0e38d15366e861040729a7f1e0a8e1427a6b6c2d46d0c3e9c465329574af702;
    5'b01100 : xpb = 1024'h24984c4aba3ae122b76ae8cc8ca5ee980bf8503263d84611d3278ed27c77c7c1b733fb6a0f7231629e2a64b8934b2f3a8c7f161f21e4a85853669d973357e8c8556d1658f3df7f8d1c35be5297dff6f26678917fb3ce78268f66e6ae92f4e989589864c229a3dac6fe08b1adf5343006f74f5f0de1cfeb7890de5c888a8b16c4;
    5'b01101 : xpb = 1024'h9d6dd634cb0941c0ce0ccc17a345475b03465901cfcf618da3535647d3838bc1ddfdf958c22ab489eaecc1f737257e5bb045c7e5d12eebe77ac3ffa29ed634a4aa15a5ff7d3d7306eaf63a9b351a78fc91b0995ab5ce758a3f0d308ef0a5beb63f54ce98cda2280b425eafbbc42df82315d1e63b3f7e27e2cbe5e0ec46ad9cf1;
    5'b01110 : xpb = 1024'h65961ac919e96d9619a9378ba98a58cc891e5ea0664edc91f5a26467778ca2ba017f79ceaabcb9229850dfeef7a1bcb26ff251c65dc65f2af182224fcf820bcf8a6f00f7570a693ba71cb441397936d5c8e3a79d2b4845dd3926e874942bf150f709a645c0d77cc1fff4c6ea9b579a15e57a8e864ce1071cc07dea4b79edbcb3;
    5'b01111 : xpb = 1024'h2dbe5f5d68c9996b6545a2ffafcf6a3e0ef6643efcce579647f172871b95b9b22500fa44934ebdbb45b4fde6b81dfb092f9edba6ea5dd26e684044fd002de2fa6ac85bef30d75f7063432de73dd7f4af0016b5dfa0c216303340a05a37b223ebaebe7df2b40cd178bd8ade1972813c08b52336d15a43e656b515f3aaad2ddc75;
    5'b10000 : xpb = 1024'ha693e9477997fa097be7864ac66ec30106446d0e68c57312181d39fc72a17db24bcaf833460740e292775b255bf84a2a53658d6d99a815fd8f9da7086bac2ed6bf70eb95ba3552ea3203aa2fdb1276b92b4ebdbaa2c21393e2e6ea3a9562f918957ae7c9580b1ebd01e0dc27417b0424d3a5bdfeb7f222c0f01d780e695062a2;
    5'b10001 : xpb = 1024'h6ebc2ddbc87825dec783f1beccb3d4728c1c72acff44ee166a6c481c16aa94aa6f4c78a92e99457b3fdb791d1c7488811312174e263f8941065bc9b59c5806019fca468d9402491eee2a23d5df7134926281cbfd183be3e6dd00a22038e92bb34d2fbf764b407373bf76f35618a4a617a34e6649c55501fae4b5816d9c908264;
    5'b10010 : xpb = 1024'h36e47270175851b413205d32d2f8e5e411f4784b95c4691abcbb563bbab3aba292cdf91f172b4a13ed3f9714dcf0c6d7d2bea12eb2d6fc847d19ec62cd03dd2c8023a1856dcf3f53aa509d7be3cff26b99b4da3f8db5b439d71a5a05dc6f5e4e04e497233e75c82a7d0d0a84efce480a72f70e94d2b7e134d94d8acccfd0a226;
    5'b10011 : xpb = 1024'hafb9fc5a2826b25229c2407de9983ea70942811b01bb84968ce71db111bf6fa2b997f70dc9e3cd3b3a01f45380cb15f8f68552f562214013a4774e6e38822908d4cc312bf72d32cd791119c4810a7475c4ece21a8fb5b19d86c0a3e63a20337aeba100f9e274156ec1630892bec81026917995c230661d9f14550f308bf32853;
    5'b10100 : xpb = 1024'h77e240ee7706de27755eabf1efdd50188f1a86b9983aff9adf362bd0b5c8869add197783b275d1d3e766124b4147544fb631dcd5eeb8b3571b35711b692e0033b5258c23d0fa29023537936a8569324efc1ff05d052f81f080da5bcbdda66615a355d8a6d5a96a257ef91fc195f1b21961223e0d3dc8fcd908ed188fbf334815;
    5'b10101 : xpb = 1024'h400a8582c5e709fcc0fb1765f622618a14f28c582eba7a9f318539f059d19d93009af7f99b07d66c94ca304301c392a675de66b67b50269a91f393c899d9d75e957ee71baac71f36f15e0d1089c7f0283352fe9f7aa952437af413b1812c98b05b0ab053c8debedc3c8f36f06d1b540c30cae6584b2bdc12fd8521eef27367d7;
    5'b10110 : xpb = 1024'h832ca1714c735d20c9782d9fc6772fb9aca91f6c539f5a383d4480ffddab48b241c786f8399db05422e4e3ac23fd0fd358af09707e799de08b1b675ca85ae8975d842138494156bad8486b68e26ae016a860ce1f0232296750dcb9724b2cb4b12bf8800bc141392fa254e1f4444f5ff00738ea3588ebb4cf21d2b4e25b38799;
    5'b10111 : xpb = 1024'h8108540125959670233966251306cbbe92189ac63131111f54000f8554e6788b4ae6765e36525e2c8ef0ab79661a201e5951a25db731dd6d300f18813603fa65ca80d1ba0df208e57c4502ff2b61300b95be14bcf2231ffa24b415778263a077f97bf1d7601260d73e7b4c2d133ebe1b1ef615d0b63cf7b72d24afb1e1d60dc6;
    5'b11000 : xpb = 1024'h493098957475c2456ed5d199194bdd3017f0a064c7b08c23a64f1da4f8ef8f836e67f6d41ee462c53c54c97126965e7518fe2c3e43c950b0a6cd3b2e66afd190aada2cb1e7beff1a386b7ca52fbfede4ccf122ff679cf04d1ecdcd5d25e9d312b130c9845347b58dfc11635bea68600dee9ebe1bc39fd6f121bcb91115162d88;
    5'b11001 : xpb = 1024'h1158dd29c355ee1aba723d0d1f90eea19dc8a6035e300727f89e2bc49cf8a67b91e9774a0776675de9b8e768e7129ccbd8aab61ed060c3f41d8b5ddb975ba8bb8b3387a9c18bf54ef491f64b341eabbe04243141dd16c0a018e78542c97005ad68e5a131467d0a44b9a77a8ac1920200be476666d102b62b1654c27048564d4a;
    5'b11010 : xpb = 1024'h8a2e6713d4244eb8d1142058363047649516aed2ca2722a3c8c9f339f4046a7bb8b37538ba2eea85367b44a78aecebecfc7167e57fab078344e8bfe702d9f497dfdc17504ae9e8c8c3527293d1592dc82f5c391cdf16be03c88dcf232720dada4fa20b07ea7b5788fdfd7898908bca1cdcc9ed942eb0f295515c46d40478d377;
    5'b11011 : xpb = 1024'h5256aba823047a8e1cb08bcc3c7558d61aeeb47160a69da81b190159980d8173dc34f5aea2c0ef1de3df629f4b692a43bc1df1c60c427ac6bba6e2943385cbc2c035724824b6defd7f78ec39d5b7eba1668f475f54908e56c2a78708caa70d750756e2b4ddb0ac3fbb938fc767b56c0fac7295df3c13d1cf45f4503337b8f339;
    5'b11100 : xpb = 1024'h1a7ef03c71e4a663684cf74042ba6a47a0c6ba0ff72618ac6d680f793c16986bffb676248b52f3b6914380970be5689a7bca7ba698d9ee0a326505416431a2eda08ecd3ffe83d5323b9f65dfda16a97a9dc255a1ca0a5ea9bcc13eee6e2d400fbf0bba61d0e600f67929a6f63edf0e027c1b3e2a4976b1093a8c59926af912fb;
    5'b11101 : xpb = 1024'h93547a2682b307017eeeda8b5959c30a9814c2df631d34283d93d6ee93225c6c268074133e0b76ddde05ddd5afbfb7bb9f912d6d4824319959c2674ccfafeec9f5375ce687e1c8ac0a5fe22877512b84c8fa5d7ccc0a5c0d6c6788cecbde153ca5c8243874e44e3abd7fa5040dd8d61e9a9dc557a724ed737593ddf6271b9928;
    5'b11110 : xpb = 1024'h5b7cbebad19332d6ca8b45ff5f9ed47c1decc87df99caf2c8fe2e50e372b73644a01f489269d7b768b69fbcd703bf6125f3db74dd4bba4dcd08089fa005bc5f4d590b7de61aebee0c6865bce7bafe95e002d6bbf41842c60668140b46f6447d75d7cfbe56819a2f17b15bc32e50278116a466da2b487ccad6a2be7555a5bb8ea;
    5'b11111 : xpb = 1024'h23a5034f20735eac1627b17365e3e5eda3c4ce1c901c2a30e231f32ddb348a5c6d8374ff0f2f800f38ce19c530b834691eea412e61531820473eaca731079d1fb5ea12d63b7bb51582acd574800ea73737607a01b6fdfcb3609af89a12ea7a721531d3925b4ef7a838abd361bc2c1a0439ef15edc1eaabe75ec3f0b48d9bd8ac;
    endcase
end

endmodule

module xpb_5_925
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7aa6cb841adedf9dd229f6a7d46893cda81cfe52bc6fe0dee516393bfb62e8925a2224c120b57ee7ccdefb2158eb2456f76156449b799e7e90ed8361bb5fbe5e491637533e805a1b5e00d371f1e6665d88f4f3d0a9fd69310d7476e9e27ec9e3dbd182e5086051ebf81ed1c9d18c1f480ec709c44febeb3ea8c453901c2df200;
    5'b00010 : xpb = 1024'h44a051b273cf8a72d94e75789876e049dec3f974a36821464c4fb92243c3241cb0fbcc0977447f40fa5fb6fbce7837e38aa884a314406cb1713bc7653bed080b1ddd39f7cd6fb6f1a967a4414af1088a1de4ee08c774a551655c5bd90ad2f135889b73a05ff7ab4a697dbcb4ab481866ceb434a64f8c794d0b192c1baf797d95;
    5'b00011 : xpb = 1024'he99d7e0ccc03547e072f4495c852cc6156af4968a6061adb38939088c235fa707d57351cdd37f9a27e072d644054b701defb3018d073ae4518a0b68bc7a51b7f2a43c9c5c5f13c7f4ce7510a3fbaab6b2d4e840e4ebe171bd4440c8332718873565645bb78f04a8dadca79f850411858ea15f884f2d075b6d6e04a742c5092a;
    5'b00100 : xpb = 1024'h8940a364e79f14e5b29ceaf130edc093bd87f2e946d0428c989f72448786483961f79812ee88fe81f4bf6df79cf06fc7155109462880d962e2778eca77da10163bba73ef9adf6de352cf488295e211143bc9dc118ee94aa2cab8b7b215a5e26b1136e740bfef5694d2fb7969569030cd9d68694c9f18f29a163258375ef2fb2a;
    5'b00101 : xpb = 1024'h533a2993408fbfbab9c169c1f4fc0d0ff42eee0b2dc882f3ffd8f22acfe683c3b8d13f5b4517fedb224029d2127d8353a89837a4a147a795c2c5d2cdf86759c31081769429cecab99e361951eeecb340d0b9d649ac6086c322a09ca13dfa09bcbe00d7fc1786aff3445a6454304c29ec5d55942e9eb980a8788730c2f23e86bf;
    5'b00110 : xpb = 1024'h1d33afc199806a8fc0e5e892b90a598c2ad5e92d14c0c35b671272111846bf4e0faae6a39ba6ff344fc0e5ac880a96e03bdf66031a0e75c8a31416d178f4a36fe5487938b8be278fe99cea2147f7556d65a9d081c9d7c2e37a888190664e310e6acac8b76f1e0951b5b94f3f0a08230b1d42bf109e5a0eb6dadc094e858a1254;
    5'b00111 : xpb = 1024'h97da7b45b45f4a2d930fdf3a8d72ed59d2f2e77fd130a43a4c28ab4d13a9a7e069cd0b64bc5c7e1c1c9fe0cde0f5bb373340bc47b588144734019a33345461ce2e5eb08bf73e81ab479dbd9339ddbbcaee9ec45273d52c1487fcf87a48ccfaf2469c4b9c777e5b3dadd82108db9442532c09c8d4ee45f9f583a05cdea1b80454;
    5'b01000 : xpb = 1024'h61d401740d4ff5029a345e0b518139d60999e2a1b828e4a1b3622b335c09e36ac0a6b2ad12eb7e754a209ca85682cec3c687eaa62e4ee27a144fde36b4e1ab7b0325b330862dde8193048e6292e85df7838ebe8a914c6834dfe4dd6971212243f3663c57cf15b49c1f370bf3b5503b71ebf6f3b6ede68803e5f5356a35038fe9;
    5'b01001 : xpb = 1024'h2bcd87a266409fd7a158dcdc158f86524040ddc39f2125091a9bab19a46a1ef5178059f5697a7ece77a15882cc0fe25059cf1904a715b0acf49e223a356ef527d7ecb5d5151d3b57de6b5f31ebf30024187eb8c2aec3a45537ccc25899754995a0302d1326ad0dfa9095f6de8f0c3490abe41e98ed871612484a0df5c84f1b7e;
    5'b01010 : xpb = 1024'ha6745326811f7f757382d383e9f81a1fe85ddc165b9105e7ffb1e4559fcd078771a27eb68a2ffdb6448053a424fb06a751306f49428f4f2b858ba59bf0ceb3862102ed28539d95733c6c32a3ddd96681a173ac9358c10d86454139427bf413797c01aff82f0d5fe688b4c8a8609853d8baab285d3d730150f10e6185e47d0d7e;
    5'b01011 : xpb = 1024'h706dd954da102a4a7aa75254ae06669c1f04d7384289464f66eb643be82d4311c87c25fee0befe0f72010f7e9a881a33e4779da7bb561d5e65d9e99f715bfd32f5c9efcce28cf24987d3037336e408ae3663a6cb763849a69d291e31a4483acb28cba0b386a4b944fa13b3933a544cf77a98533f3d138f5f53633a1177c89913;
    5'b01100 : xpb = 1024'h3a675f833300d51f81cbd1257214b31855abd25a298186b6ce24e422308d7e9c1f55cd47374dfe689f81cb5910152dc077becc06341ceb9146282da2f1e946dfca90f271717c4f1fd339d4428feeaadacb53a10393af85c6f5110320cc9c621cd595916ede3c12a36b729e7e141046163a857e213cb41d6db5b8129d0b1424a8;
    5'b01101 : xpb = 1024'h460e5b18bf17ff488f04ff63622ff948c52cd7c1079c71e355e640878edba26762f748f8ddcfec1cd02873385a2414d0b05fa64ace3b9c4267671a67276908c9f57f516006babf61ea0a511e8f94d0760439b3bb126c1e74cf8e80ff4f0896e825f822a35d36c01dcd18968edcc3f34fa72a9033c54ab7c180ceb289e5fb03d;
    5'b01110 : xpb = 1024'h7f07b135a6d05f925b1a469e0a8b9362346fcbcecce9a7fd1a749d447450a2b8d0519950ae927da999e18254de8d65a4026750a9485d5842b763f5082dd64eeae86e2c693eec06117ca17883dadfb364e9388f0c5b242b185a6d5ef9d76f53525e31050f3e33bdedd4f05b32bf585e7d0939b2c78c4096bac0d13eb8ba8da23d;
    5'b01111 : xpb = 1024'h49013763ffc10a67623ec56ece99dfde6b16c6f0b3e1e86481ae1d2abcb0de43272b409905217e02c7623e2f541a793095ae7f07c124267597b2390bae639897bd352f0dcddb62e7c808495333ea55917e288944789b6738b25543e8ffc37aa40afaf5ca95cb174c464f461d9914579bc926dda98be124c9232617444dd92dd2;
    5'b10000 : xpb = 1024'h12fabd9258b1b53c6963443f92a82c5aa1bdc2129ada28cbe8e79d11051119cd7e04e7e15bb07e5bf4e2fa09c9a78cbd28f5ad6639eaf4a878007d0f2ef0e24491fc31b25ccabfbe136f1a228cf4f7be1318837c9612a3590a3d28d82817a1f5b7c4e685ed6270aab7ae310872d050ba8914088b8b81b2d7857aefcfe124b967;
    5'b10001 : xpb = 1024'h8da18916739094da3b8d3ae76710c02849dac065574a09aacdfdd64d0074025fd8270ca27c65fd43c1c1f52b2292b114205703aad564932708ee0070ea50a0a2db1269059b4b19d9716fed947edb5e1b9c0d774d40100c8a17b19fc20a966bd99396696af5c2c296afcd02d2445c700297db124fdb6d9e162e3f435ffd52ab67;
    5'b10010 : xpb = 1024'h579b0f44cc813faf42b1b9b82b1f0ca48081bb873e424a123537563348d43dea2f00b3ead2f4fd9cef42b105981fc4a0b39e32094e2b6159e93c44746addea4fafd96baa2a3a76afbcd6be63d7e6004830fd71855d8748aa6f9984b132ea932b40605a264d5a1bf5212bedbd1e18692157c83d31db0e2c2490941beb909e36fc;
    5'b10011 : xpb = 1024'h219495732571ea8449d63888ef2d5920b728b6a9253a8a799c70d6199134797485da5b332983fdf61cc36ce00dacd82d46e56067c6f22f8cc98a8877eb6b33fc84a06e4eb929d386083d8f3330f0a274c5ed6bbd7afe84cac78169a05b3eba7ced2a4ae1a4f17553928ad8a7f7d4624017b56813daaeba32f2e8f47723e9c291;
    5'b10100 : xpb = 1024'h9c3b60f74050ca221c002f30c395ecee5f45b4fbe1aa6b5881870f558c976206dffc7ff44a397cdde9a268016697fc843e46b6ac626bce0b5a780bd9a6caf25acdb6a5a1f7aa2da1663e62a522d708d24ee25f8e24fbedfbd4f5e08a3dbd8460c8fbcdc6ad51c73f8aa9aa71c9608188267c71d82a9aa5719bad48074017b491;
    5'b10101 : xpb = 1024'h6634e725994174f72324ae0187a4396a95ecb01dc8a2abbfe8c08f3bd4f79d9136d6273ca0c87d37172323dbdc251010d18de50adb329c3e3ac64fdd27583c07a27da84686998a77b1a533747be1aafee3d259c642732a1c2cddc5796611abb275c5be8204e9209dfc08955ca31c7aa6e6699cba2a3b337ffe022092d3634026;
    5'b10110 : xpb = 1024'h302e6d53f2321fcc2a492cd24bb285e6cc93ab3faf9aec274ffa0f221d57d91b8dafce84f7577d9044a3dfb651b2239d64d5136953f96a711b1493e0a7e585b47744aaeb1588e74dfd0c0443d4ec4d2b78c253fe5fea663c84c5aa688e65d304228faf3d5c8079fc6d6780477cd873c5a656c79c29dbc18e6056f91e66aecbbb;
    5'b10111 : xpb = 1024'haad538d80d10ff69fc73237a201b19b474b0a9926c0acd063510485e18bac1ade7d1f346180cfc781182dad7aa9d47f45c3669adef7308efac02174263454412c05ae23e540941695b0cd7b5c6d2b38901b747cf09e7cf6d923a215270e49ce7fe61322264e0cbe8658652114e64930db51dd16079c7accd091b4cae82dcbdbb;
    5'b11000 : xpb = 1024'h74cebf066601aa3f0397a24ae4296630ab57a4b453030d6d9c49c844611afd383eab9a8e6e9bfcd13f0396b2202a5b80ef7d980c6839d7228c505b45e3d28dbf9521e4e2e2f89e3fa673a8851fdd55b596a74207275f0b8dea2206419938c439ab2b22ddbc782546d6e53cfc28208c2c750afc4279683adb6b70253a16284950;
    5'b11001 : xpb = 1024'h3ec84534bef255140abc211ba837b2ace1fe9fd639fb4dd50383482aa97b38c2958541d6c52afd2a6c84528c95b76f0d82c4c66ae100a5556c9e9f49645fd76c69e8e78771e7fb15f1da795478e7f7e22b973c3f44d647ae4209eb30c18ceb8b57f51399140f7ea5484427e701dc854b34f827247908c8e9cdc4fdc5a973d4e5;
    5'b11010 : xpb = 1024'h8c1cb6317e2ffe911e09fec6c45ff2918a59af820f38e3c6abcc810f1db744cec5ee91f1bb9fd839a050e670b44829a160bf4c959c773884cece34ce4ed21193eafea2c00d757ec3d414a23d1f29a0ec0873677624d83ce99f1d01fe9e112dd04bf04546ba6d803b9a312d1db987e69f4e5520678a956f83019d6513cbf607a;
    5'b11011 : xpb = 1024'h836896e732c1df86e40a969440ae92f6c0c2994add636f1b4fd3014ced3e5cdf46810de03c6f7c6b66e40988642fa6f10d6d4b0df5411206ddda66aea04cdf7787c6217f3f57b2079b421d95c3d9006c497c2a480c4aecffa7664709cc5fdcc0e0908739740729efb1c1e49bad249db203ac5bcac8954236d8de29e158ed527a;
    5'b11100 : xpb = 1024'h4d621d158bb28a5beb2f156504bcdf72f769946cc45baf82b70c8133359e98699d5ab52892fe7cc49464c562d9bcba7da0b4796c6e07e039be28aab220da29245c8d2423ce470edde6a8ee651ce3a298de6c248029c2291fff4e2bf8f4b404128d5a77f4cb9e834e2320cf8686e096d0c39986acc835d0453b33026cec38de0f;
    5'b11101 : xpb = 1024'h175ba343e4a33530f2539435c8cb2bef2e108f8eab53efea1e4601197dfed3f3f4345c70e98d7d1dc1e5813d4f49ce0a33fba7cae6ceae6c9e76eeb5a16772d1315426c85d366bb4320fbf3475ee44c5735c1eb847396540573610e81d082b643a2468b02335dcac947fba71609c8fef8386b18ec7d65e539d87daf87f8469a4;
    5'b11110 : xpb = 1024'h92026ec7ff8214cec47d8add9d33bfbcd62d8de167c3d0c9035c3a557961bc864e5681320a42fc058ec47c5ea834f2612b5cfe0f82484ceb2f6472175cc7312f7a6a5e1b9bb6c5cf901092a667d4ab22fc511288f136ce7164aa87d1ff86f54815f5eb952b962e988c9e8c3b3228af37924dbb5317c24992464c2e889bb25ba4;
    5'b11111 : xpb = 1024'h5bfbf4f65872bfa3cba209ae61420c390cd489034ebc11306a95ba3bc1c1f810a530287a60d1fc5ebc4538391dc205edbea42c6dfb0f1b1e0fb2b61add547adc4f3160c02aa622a5db776375c0df4d4f91410cc10eae0a91bc926cc127db1c99c2bfdc50832d87f6fdfd77260be4a856523ae6351762d7a0a8a107142efde739;
    endcase
end

endmodule

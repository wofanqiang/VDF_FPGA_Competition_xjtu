module xpb_5_865
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h16fffc8d537e2aa0b0dc88f2d2411cc3fa32fca207234c2ed79d7cf233b8467f50f81331ccdafee921d305b1d8cace8225e99d760db9c2b741e078cb1c940ba8dc46bbe4ffacdfb105f5a21a3d01f157422c39f13331afa17504361b205895c6769473309e9b1e533ead4c4aeca9700f2858a038af96884666587bf56bb580a3;
    5'b00010 : xpb = 1024'h2dfff91aa6fc554161b911e5a4823987f465f9440e46985daf3af9e467708cfea1f0266399b5fdd243a60b63b1959d044bd33aec1b73856e83c0f19639281751b88d77c9ff59bf620beb44347a03e2ae845873e266635f42ea086c3640b12b8ced28e6613d363ca67d5a9895d952e01e50b140715f2d108cccb0f7ead76b0146;
    5'b00011 : xpb = 1024'h44fff5a7fa7a7fe212959ad876c3564bee98f5e61569e48c86d876d69b28d37df2e839956690fcbb657911158a606b8671bcd862292d4825c5a16a6155bc22fa94d433aeff069f1311e0e64eb705d405c684add399950ee45f0ca2516109c15363bd5991dbd15af9bc07e4e0c5fc502d7909e0aa0ec398d3330973e0432081e9;
    5'b00100 : xpb = 1024'h5bfff2354df8aa82c37223cb4904730fe8cbf2881c8d30bb5e75f3c8cee119fd43e04cc7336bfba4874c16c7632b3a0897a675d836e70add0781e32c72502ea3711aef93feb37ec417d68868f407c55d08b0e7c4ccc6be85d410d86c81625719da51ccc27a6c794cfab5312bb2a5c03ca16280e2be5a21199961efd5aed6028c;
    5'b00101 : xpb = 1024'h72ffeec2a176d523744eacbe1b458fd3e2feef2a23b07cea361370bb0299607c94d85ff90046fa8da91f1c793bf6088abd90134e44a0cd9449625bf78ee43a4c4d61ab78fe605e751dcc2a833109b6b44add21b5fff86e2749150e87a1baece050e63ff3190797a039627d769f4f304bc9bb211b6df0a95fffba6bcb1a8b832f;
    5'b00110 : xpb = 1024'h89ffeb4ff4f4ffc4252b35b0ed86ac97dd31ebcc2ad3c9190db0edad3651a6fbe5d0732acd21f976caf2222b14c0d70ce379b0c4525a904b8b42d4c2ab7845f529a8675dfe0d3e2623c1cc9d6e0ba80b8d095ba7332a1dc8be1944a2c21382a6c77ab323b7a2b5f3780fc9c18bf8a05af213c1541d8731a66612e7c0864103d2;
    5'b00111 : xpb = 1024'ha0ffe7dd48732a64d607bea3bfc7c95bd764e86e31f71547e54e6a9f6a09ed7b36c8865c99fcf85fecc527dced8ba58f09634e3a60145302cd234d8dc80c519e05ef2342fdba1dd729b76eb7ab0d9962cf359598665bcd6a331d7abde26c186d3e0f2654563dd446b6bd160c78a2106a1a6c618ccd1db9eccc6b63b5f1f68475;
    5'b01000 : xpb = 1024'h7529f14da03203cbbdecfbf81ae9ece6021e1df63a2c0ff3f0f2e3beabf86f284781c159cb178ba6f39ee47e2f86346cb32c3ca4b1b456e5e6486faa9cde8956de6aa794dd600431d130e2f4f33c6891d5cd5f10d074ffaf2951ede489a0ba1859c075b440ffa0c6eaa7b786d7b5a4ff3eb22e32c68e502ec5464a6d4c99ead;
    5'b01001 : xpb = 1024'h1e529ba22d814add6cbb58b253efbb925a54de816ac60d2e16acab2e1e77cd71d5702f47698c77a3910cf3f9bbc331c8f11c614058d50825a044ffc5c661f43e4a2d665e4d82dff42308b0498c35b7e05f890fe24038ff9c679954f968f2a167fc307a8be2ab185fad57c7c35a24ca5f1c43c31bdbff6d4952ace09c407f1f50;
    5'b01010 : xpb = 1024'h3552982f80ff757e1d97e1a52630d8565487db2371e9595cee4a2820523013f1266842793667768cb2dff9ab948e004b1705feb6668ecadce2257890e2f5ffe7267422434d2fbfa528fe5263c937a937a1b549d3736aaf3ddc9d8b14894b372e72c4edbc814636b2ec05140e46ce3a6e449c63548b95f58fb9055c91ac349ff3;
    5'b01011 : xpb = 1024'h4c5294bcd47da01ece746a97f871f51a4ebad7c5790ca58bc5e7a51285e85a70776055ab03427575d4b2ff5d6d58cecd3cef9c2c74488d942405f15bff8a0b9002bade284cdc9f562ef3f47e06399a8ee3e183c4a69c5edf51a1c12fa9a3ccf4e95960ed1fe155062ab260593377aa7d6cf5038d3b2c7dd61f5dd88717ea2096;
    5'b01100 : xpb = 1024'h6352914a27fbcabf7f50f38acab311de48edd467802ff1ba9d852204b9a0a0efc85868dcd01d745ef686050f46239d4f62d939a28202504b65e66a271c1e1738df019a0d4c897f0734e99698433b8be6260dbdb5d9ce0e80c6a5f74ac9fc62bb5fedd41dbe7c7359695faca420211a8c954da3c5eac3061c85b6547c839fa139;
    5'b01101 : xpb = 1024'h7a528dd77b79f560302d7c7d9cf42ea24320d10987533de975229ef6ed58e76f19507c0e9cf8734818590ac11eee6bd188c2d7188fbc1302a7c6e2f238b222e1bb4855f24c365eb83adf38b2803d7d3d6839f7a70cffbe223baa2d65ea54f881d682474e5d1791aca80cf8ef0cca8a9bbda643fe9a598e62ec0ed071ef5521dc;
    5'b01110 : xpb = 1024'h91528a64cef82000e10a05706f354b663d53cdab8e768a184cc01be921112dee6a488f4069d372313a2c1072f7b93a53aeac748e9d75d5b9e9a75bbd55462e8a978f11d74be33e6940d4daccbd3f6e94aa66319840316dc3b0ae63810aad8e484d16ba7efbb2afffe6ba4539f973faaae5fee43749f016a952674c675b0aa27f;
    5'b01111 : xpb = 1024'ha85286f222764aa191e68e634176682a3786ca4d9599d647245d98db54c9746dbb40a27236ae711a5bff1624d08408d5d4961204ab2f98712b87d48871da3a3373d5cdbc4b901e1a46ca7ce6fa415febec926b8973631d6525b2999c2b06240ec3ab2daf9a4dce5325679184e61d6aba0e57846ff9869eefb8bfc85cc6c02322;
    5'b10000 : xpb = 1024'hea53e29b406407977bd9f7f035d3d9cc043c3bec74581fe7e1e5c77d57f0de508f0382b3962f174de73dc8fc5f0c68d9665879496368adcbcc90df5539bd12adbcd54f29bac00863a261c5e9e678d123ab9abe21a0e9ff5e52a3dbc913417430b380eb6881ff418dd54f6f0daf6b49fe7d645c658d1ca05d8a8c94da9933d5a;
    5'b10001 : xpb = 1024'h25a53ab707846b1a289a2871d59e5a60ba76c060ce68ce2d55bbd96a0937546459e84b5d063df05e0046e2419ebb950fbc4f250aa3f04d93fea986c0702fdcd3b81410d79b58e037401bbe78db697e697ce5e5d34d404f975a2e73d7b18cad0981cc81e726bb126c1c02433bc7a024af102ee5ff0868524c3f0145431548bdfd;
    5'b10010 : xpb = 1024'h3ca537445b0295bad976b164a7df7724b4a9bd02d58c1a5c2d59565c3cef9ae3aae05e8ed318ef472219e7f377866391e238c280b1aa104b4089ff8b8cc3e87c945accbc9b05bfe846116093186b6fc0bf121fc48071ff38cf32a9f2d1e542cff860f517c55630bf5aaf8f86b44994be38878637b7feda92a559c13880fe3ea0;
    5'b10011 : xpb = 1024'h53a533d1ae80c05b8a533a577a2093e8aedcb9a4dcaf668b04f6d34e70a7e162fbd871c09ff3ee3043eceda55051321408225ff6bf63d302826a7856a957f42570a188a19ab29f994c0702ad556d6118013e59b5b3a3aeda4436e00df23dd8966ef5684863f14f12995cdbd1a0f304cd60e02670679562d90bb23d2decb3bf43;
    5'b10100 : xpb = 1024'h6aa5305f01feeafc3b2fc34a4c61b0aca90fb646e3d2b2b9dc945040a46027e24cd084f26cceed1965bff357291c00962e0bfd6ccd1d95b9c44af121c5ebffce4ce844869a5f7f4a51fca4c7926f526f436a93a6e6d55e7bb93b162912966e5ce589db79028c6d65d80a281c8d9c74dc8938c6a9172beb1f720ab92358693fe6;
    5'b10101 : xpb = 1024'h81a52cec557d159cec0c4c3d1ea2cd70a342b2e8eaf5fee8b431cd32d8186e619dc8982439a9ec028792f90901e6cf1853f59ae2dad75871062b69ece2800b77292f006b9a0c5efb57f246e1cf7143c68596cd981a070e1d2e3f4c4432ef04235c1e4ea9a1278bb916b774677a45e4ebb19166e1c6c27365d8633518c41ec089;
    5'b10110 : xpb = 1024'h98a52979a8fb403d9ce8d52ff0e3ea349d75af8af2194b178bcf4a250bd0b4e0eec0ab560684eaeba965febadab19d9a79df3858e8911b28480be2b7ff1417200575bc5099b93eac5de7e8fc0c73351dc7c307894d38bdbea343825f534799e9d2b2c1da3fc2aa0c5564c0b266ef54fad9ea071a7658fbac3ebbb10e2fd4412c;
    5'b10111 : xpb = 1024'hafa52606fc796ade4dc55e22c32506f897a8ac2cf93c9746636cc7173f88fb603fb8be87d35fe9d4cb39046cb37c6c1c9fc8d5cef64adddf89ec5b831ba822c8e1bc783599661e5d63dd8b164975267509ef417a806a6d601847b87a73a02fb04947350ade5dc85f94120cfd5398c50a0242a75325ef83f2a5142d039b89c1cf;
    5'b11000 : xpb = 1024'h15f7dd3e8e0960b6339c6f3e850bdc6b2065a59e2ae842fdbd2d8ab3c03e94d78d685440d6146a2f4dadcad7a8e929d461984b5ee151d04b1b2d94effd69b9c049b3ff6be98200c957392a8ded9b539b581681d32715eff0d7bf5c9ad9ce22e490d41611cc2fee254bff726948720eefdbc168a9853aaf08c4fd2df47e5cdc07;
    5'b11001 : xpb = 1024'h2cf7d9cbe1878b56e478f831574cf92f1a98a240320b8f2c94cb07a5f3f6db56de606772a2ef69186f80d08981b3f8568781e8d4ef0b93025d0e0dbb19fdc56925fabb50e92ee07a5d2ecca82a9d44f29a42bbc45a479f924cc392b5fa26b8ab076889426acb0c788aacbeb4351b7eff041a08e234d1374f2b55a9e9ea125caa;
    5'b11010 : xpb = 1024'h43f7d6593505b5f795558124298e15f314cb9ee2392edb5b6c68849827af21d62f587aa46fca68019153d63b5a7ec6d8ad6b864afcc555b99eee86863691d11202417735e8dbc02b63246ec2679f3649dc6ef5b58d794f33c1c7c8d11a7f4e717dfcfc7309662acbc95a0aff21c4ef0e2c72a91ae467bf9591ae25df55c7dd4d;
    5'b11011 : xpb = 1024'h5af7d2e68883e09846320a16fbcf32b70efe9b844052278a4406018a5b67685580508dd63ca566eab326dbed3349955ad35523c10a7f1870e0ceff515325dcbade88331ae8889fdc691a10dca4a127a11e9b2fa6c0aafed536cbfeec3ad7e437f4916fa3a801491f0807574a0e6e5f1d54cb495393fe47dbf806a1d4c17d5df0;
    5'b11100 : xpb = 1024'h71f7cf73dc020b38f70e9309ce104f7b09319826477573b91ba37e7c8f1faed4d148a108098065d3d4f9e19f0c1463dcf93ec1371838db2822af781c6fb9e863baceeeffe8357f8d6f0fb2f6e1a318f860c76997f3dcae76abd035075b3079fe6b25e2d4469c677246b4a394fb17cf2c7d23e98c4394d0225e5f1dca2d32de93;
    5'b11101 : xpb = 1024'h88f7cc012f8035d9a7eb1bfca0516c3f036494c84e98bfe7f340fb6ec2d7f5542240b439d65b64bcf6cce750e4df325f1f285ead25f29ddf648ff0e78c4df40c9715aae4e7e25f3e750555111ea50a4fa2f3a389270e5e1820d46b227b890fc4e1ba5604e53785c58561efdfe7c13f3ba57c89c4f32b5868c4b799bf98e85f36;
    5'b11110 : xpb = 1024'h9ff7c88e82fe607a58c7a4ef72928902fd97916a55bc0c16cade7860f6903bd37338c76ba33663a6189fed02bdaa00e14511fc2333ac6096a67069b2a8e1ffb5735c66c9e78f3eef7afaf72b5ba6fba6e51fdd7a5a400db995d8a13d9be1a58b584ec93583d2a418c40f3c2ad46aaf4acdd529fda2c1e0af2b1015b5049ddfd9;
    5'b11111 : xpb = 1024'h64a7fc6148e56523e9eb60b34795e7586548adb8767b7ce249f3bfd7745d54ac0e85d24a5eae4009b14b36db316be9906e171b31eb3530237b1a31f8aa396acdb53ee0037ab215b6e5696a2ffcd28cd33471dd300eb904a5550455e020f98bf9fdbaa3c71a4c9de7bfca196c943f930a753eb54020d0bc54af916a5e770fa11;
    endcase
end

endmodule

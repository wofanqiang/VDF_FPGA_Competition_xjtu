module xpb_5_485
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha2faf86643bd35390cfcdd6e6ad8b53c38c2bee7714c48b8bc406c26462e5eeb6fb5d8b73d6801c442688eed6e94b678a59a1428db8dccb5bcfcd7724ab34ba85751be2722b106299aefdeac7d507446b05e6c81d94206e22d42b371d69ab01506679c78461754470042e165f33ab7e1a268aab6dca74d50a64ee464aa5f6e46;
    5'b00010 : xpb = 1024'h9548ab76c58c35a94ef44305c5572327000f7a9e0d20f0f9faa41ef6d95a10cedc2333f5b0a984f9e572de93f9cb5c26e71a006b9468c91fc95a6f865a94229f3a54479f95d10f0e2345bab661c5245c6cb7df6b25fde0b3a4f8d4e8f30abd97ddc7a6c6db65b00079c5dbeceea54999f5f7768b69033d71062e4dc4cbdc7621;
    5'b00011 : xpb = 1024'h87965e87475b361990eba89d1fd59111c75c3654a8f5993b3907d1c76c85c2b248908f3423eb082f887d2e3a850201d52899ecae4d43c589d5b8079a6a74f9961d56d11808f117f2ab9b96c04639d4722911525472b9ba851caef6600f7acb1ab527b11570b40bb9f348d673ea0fdb524986425ff55f2d91660db724ed597dfc;
    5'b00100 : xpb = 1024'h79e41197c92a3689d2e30e347a53fefc8ea8f20b44ca417c776b8497ffb17495b4fdea72972c8b652b877de11038a7836a19d8f1061ec1f3e2159fae7a55d08d00595a907c1120d733f172ca2aae8487e56ac53dbf759456946517d72bead89d8c87bb64060267736ccbd0fae57a6d0a9d150e3481bb1db1c5ed20850ed685d7;
    5'b00101 : xpb = 1024'h6c31c4a84af936fa14da73cbd4d26ce755f5adc1e09ee9bdb5cf376892dd2679216b45b10a6e0e9ace91cd879b6f4d31ab99c533bef9be5dee7337c28a36a783e35be408ef3129bbbc474ed40f23349da1c438270c316e280c1b394e485ae62063e7c5b29b50c32ce64ecb81e0e4fec2f0a3da090e170dd225cc89e530538db2;
    5'b00110 : xpb = 1024'h5e7f77b8ccc8376a56d1d9632f50dad21d4269787c7391fef432ea392608d85c8dd8a0ef7daf91d0719c1d2e26a5f2dfed19b17677d4bac7fad0cfd69a177e7ac65e6d81625132a0449d2addf397e4b35e1dab1058ed47f983d15ac564caf3a33b47d001309f1ee65fd1c608dc4f907b4432a5dd9a72fdf285abf34551d0958d;
    5'b00111 : xpb = 1024'h50cd2ac94e9737da98c93efa89cf48bce48f252f18483a4032969d09b9348a3ffa45fc2df0f1150614a66cd4b1dc988e2e999db930afb732072e67eaa9f85571a960f6f9d5713b84ccf306e7d80c94c91a771df9a5a921cafb877c3c813b012612a7da4fc5ed7a9fd954c08fd7ba223397c171b226ceee12e58b5ca5734d9d68;
    5'b01000 : xpb = 1024'h431addd9d066384adac0a491e44db6a7abdbe0e5b41ce28170fa4fda4c603c2366b3576c6432983bb7b0bc7b3d133e3c701989fbe98ab39c138bfffeb9d92c688c638072489144695548e2f1bc8144ded6d090e2f264fb9c733d9db39dab0ea8ea07e49e5b3bd65952d7bb16d324b3ebeb503d86b32ade33456ac60594caa543;
    5'b01001 : xpb = 1024'h356890ea523538bb1cb80a293ecc249273289c9c4ff18ac2af5e02aadf8bee06d320b2aad7741b715abb0c21c849e3eab199763ea265b0061fe99812c9ba035f6f6609eabbb14d4ddd9ebefba0f5f4f4932a03cc3f20d56deaf3bf2aba1b1c2bc167eeecf08a3212cc5ab59dce8f45a43edf095b3f86ce53a54a2f65b647ad1e;
    5'b01010 : xpb = 1024'h27b643fad404392b5eaf6fc0994a927d3a755852ebc63303edc1b57b72b79fea3f8e0de94ab59ea6fdc55bc853808998f31962815b40ac702c473026d99ada56526893632ed1563265f49b05856aa50a4f8376b58bdcaf3f62a9e0a1d68b29ae98c7f93b85d88dcc45ddb024c9f9d75c926dd52fcbe2be74052998c5d7c4b4f9;
    5'b01011 : xpb = 1024'h1a03f70b55d3399ba0a6d557f3c9006801c21409879adb452c25684c05e351cdabfb6927bdf721dca0cfab6edeb72f4734994ec4141ba8da38a4c83ae97bb14d356b1cdba1f15f16ee4a770f69df55200bdce99ed8988910da600218f2fb37317028038a1b26e985bf60aaabc5646914e5fca104583eae9465090225f941bcd4;
    5'b01100 : xpb = 1024'hc51aa1bd7a23a0be29e3aef4e476e52c90ecfc0236f83866a891b1c990f03b11868c4663138a51243d9fb1569edd4f576193b06ccf6a5444502604ef95c8844186da654151167fb76a053194e540535c8365c88255462e2521623900f6b44b447880dd8b075453f38e3a532c0cefacd398b6cd8e49a9eb4c4e86b861abec4af;
    5'b01101 : xpb = 1024'haf4ca2821b5f6f44ef9b185db920238f01d18ea794bbcc3f26c98742df3d629c881e9d1d6ea0a6d686428a02d8828b6e1bb34f2fa88471fa01ff37c1440fd3ec6fbf647b37c26e25119031c5cba4797c7894c909fe9669c47f58d701e605f4c94defaa50f68c998639268698b409b2aedbf4178fc141ec056b374feac51e32f5;
    5'b01110 : xpb = 1024'ha19a55929d2e6fb531927df5139e9179c91e4a5e30907480652d3a137269147ff48bf85be1e22a0c294cd9a963b9311c5d333b72615f6e640e5ccfd553f0aae352c1edf3aae2770999e60dcfb019299234ee3bf34b524395f70ef8790276024c254fb49f8bdaf53fb2a9811faf7444672f82e3644d9ddc25cb16b94ae69b3ad0;
    5'b01111 : xpb = 1024'h93e808a31efd70257389e38c6e1cff64906b0614cc651cc1a390ece40594c66360f9539a5523ad41cc57294feeefd6ca9eb327b51a3a6ace1aba67e963d181da35c4776c1e027fee223be9d9948dd9a7f147aedc980e1d676ec519f01ee60fcefcafbeee212950f92c2c7ba6aaded61f8311af38d9f9cc462af622ab081842ab;
    5'b10000 : xpb = 1024'h8635bbb3a0cc7095b5814923c89b6d4f57b7c1cb6839c502e1f49fb498c07846cd66aed8c86530776f6178f67a267c78e03313f7d31567382717fffd73b258d118c700e4912288d2aa91c5e3790289bdada121c5e4c9f738e67b3b673b561d51d40fc93cb677acb2a5af762da64967d7d6a07b0d6655bc668ad58c0b29954a86;
    5'b10001 : xpb = 1024'h78836ec4229b7105f778aebb2319db3a1f047d82040e6d44205852852bec2a2a39d40a173ba6b3ad126bc89d055d222721b3003a8bf063a23375981183932fc7fbc98a5d044291b732e7a1ed5d7739d369fa94af3185d10a5e315cde57c62ad4ab6fd38b4bc6086c1f3270b4a1b3f9902a2f46e1f2b1ac86eab4f56b4b125261;
    5'b10010 : xpb = 1024'h6ad121d4a46a7176397014527d984924e65139389fe315855ebc0555bf17dc0da6416555aee836e2b57618439093c7d56332ec7d44cb600c3fd33025937406bedecc13d577629a9bbb3d7df741ebe9e9265407987e41aadbd5e77e557436385782cfddd9e114642598b56b3b9d1e8b487dbe12b67f0d9ca74a945ecb6c8f5a3c;
    5'b10011 : xpb = 1024'h5d1ed4e5263971e67b6779e9d816b70fad9df4ef3bb7bdc69d1fb82652438df112aec0942229ba18588067ea1bca6d83a4b2d8bffda65c764c30c839a354ddb5c1ce9d4dea82a38043935a01266099fee2ad7a81cafd84ad4d9d9fcc90a645da5a2fe8287662bfdf123865c298891d00d14cde8b0b698cc7aa73c82b8e0c6217;
    5'b10100 : xpb = 1024'h4f6c87f5a8087256bd5edf81329524fa74eab0a5d78c6607db836af6e56f3fd47f1c1bd2956b3d4dfb8ab790a7011331e632c502b68158e0588e604db335b4aca4d126c65da2ac64cbe9360b0ad54a149f06ed6b17b95e7ec553c143ad16535d318ff2770bb11b988bbb604993f3aeb924dbaa5f97c57ce80a53318baf8969f2;
    5'b10101 : xpb = 1024'h41ba3b0629d772c6ff5645188d1392e53c376c5c73610e4919e71dc7789af1b7eb89771108acc0839e9507373237b8e027b2b1456f5c554a64ebf861c3168ba387d3b03ed0c2b549543f1214ef49fa2a5b606054647538503d09e2bac98660e008effcc5a0ff7752053e5ad08f5e4071786a763424216d086a329aebd10671cd;
    5'b10110 : xpb = 1024'h3407ee16aba67337414daaafe79200d0038428130f35b68a584ad0980bc6a39b57f6d24f7bee43b9419f56ddbd6e5e8e69329d88283751b471499075d2f7629a6ad639b743e2be2ddc94ee1ed3beaa4017b9d33db1311221b4c00431e5f66e62e0500714364dd30b7ec155578ac8d229cbf94208b07d5d28ca12044bf28379a8;
    5'b10111 : xpb = 1024'h2655a1272d7573a78345104742106ebacad0e3c9ab0a5ecb96ae83689ef2557ec4642d8def2fc6eee4a9a68448a5043caab289cae1124e1e7da72889e2d839914dd8c32fb702c71264eaca28b8335a55d4134626fdecebf32c7625a902667be5b7b01162cb9c2ec4f8444fde863363e21f880ddd3cd94d4929f16dac14008183;
    5'b11000 : xpb = 1024'h18a35437af447417c53c75de9c8edca5921d9f8046df070cd5123639321e076230d188cc62714a2487b3f62ad3dba9eaec32760d99ed4a888a04c09df2b9108830db4ca82a22cff6ed40a6329ca80a6b906cb9104aa8c5c4a42c47201ed689688f101bb160ea8a7e71c74a65819df59a7316d9b1c9353d6989d0d70c357d895e;
    5'b11001 : xpb = 1024'haf10748311374880733db75f70d4a90596a5b36e2b3af4e1375e909c549b9459d3ee40ad5b2cd5a2abe45d15f124f992db2625052c846f2966258b20299e77f13ddd6209d42d8db7596823c811cba814cc62bf997649f961be268973b4696eb667025fff638e637eb4a44ec7d088752c6a5a58655912d89e9b0406c56fa9139;
    5'b11010 : xpb = 1024'hadebffae74d0a9c11430b8e461e5ffcc922d1a1e53fff806cfb655300b7818310cf4bcc2131acf1e6d26d4becda70611d34c76792e5613a8535f30244d4d33276b2f9447bff3df05108660e8fe6d2ec7fd24987b70a6a67849251c0911e147006cd7c2783c503a7eeb8d265270433f34690e503d32387ada8fff24d10159ff7f;
    5'b11011 : xpb = 1024'ha039b2bef69faa3156281e7bbc646db75979d5d4efd4a0480e1a08009ea3ca1479621800865c52541031246558ddabc014cc62bbe73110125fbcc8385d2e0a1e4e321dc03313e7e998dc3cf2e2e1deddb97e0b64bd628049c0db3d802e5154834437ccc6d19e9638651020d96badd0ecbc9d1c11be946afaefde8e3122d7075a;
    5'b11100 : xpb = 1024'h928765cf786eaaa1981f841316e2dba220c6918b8ba948894c7dbad131cf7bf7e5cf733ef99dd589b33b740be414516e564c4efea00c0c7c6c1a604c6d0ee1153134a738a633f0ce213218fcc7568ef375d77e4e0a1e5a1b38915ef74ac162061b97d71566ecf1f1de931b60671862a5102be7e64af05b1b4fbdf79144540f35;
    5'b11101 : xpb = 1024'h84d518dffa3dab11da16e9aa7161498ce8134d42277df0ca8ae16da1c4fb2ddb523cce7d6cdf58bf5645c3b26f4af71c97cc3b4158e708e67877f8607cefb80c143730b11953f9b2a987f506abcb3f093230f13756da33ecb047806e67316f88f2f7e163fc3b4dab581615e76282f45d63bab3bad74c4b3baf9d60f165d11710;
    5'b11110 : xpb = 1024'h7722cbf07c0cab821c0e4f41cbdfb777af6008f8c352990bc94520725826dfbebeaa29bbe020dbf4f9501358fa819ccad94c278411c2055084d590748cd08f02f739ba298c74029731ddd110903fef1eee8a6420a3960dbe27fda1e583a17d0bca57ebb29189a964d199106e5ded8615b7497f8f63a83b5c0f7cca51874e1eeb;
    5'b11111 : xpb = 1024'h69707f00fddbabf25e05b4d9265e256276acc4af5f27414d07a8d342eb5291a22b1784fa53625f2a9c5a62ff85b842791acc13c6ca9d01ba913328889cb165f9da3c43a1ff940b7bba33ad1a74b49f34aae3d709f051e78f9fb3c35ca0118a8ea1b7f60126d8051e4b1c0af5595817ce0ad84b63f0042b7c6f5c33b1a8cb26c6;
    endcase
end

endmodule

module compressor_array_512_16_1024
(
    input  [511:0] col_in_0,
    input  [511:0] col_in_1,
    input  [511:0] col_in_2,
    input  [511:0] col_in_3,
    input  [511:0] col_in_4,
    input  [511:0] col_in_5,
    input  [511:0] col_in_6,
    input  [511:0] col_in_7,
    input  [511:0] col_in_8,
    input  [511:0] col_in_9,
    input  [511:0] col_in_10,
    input  [511:0] col_in_11,
    input  [511:0] col_in_12,
    input  [511:0] col_in_13,
    input  [511:0] col_in_14,
    input  [511:0] col_in_15,
    input  [511:0] col_in_16,
    input  [511:0] col_in_17,
    input  [511:0] col_in_18,
    input  [511:0] col_in_19,
    input  [511:0] col_in_20,
    input  [511:0] col_in_21,
    input  [511:0] col_in_22,
    input  [511:0] col_in_23,
    input  [511:0] col_in_24,
    input  [511:0] col_in_25,
    input  [511:0] col_in_26,
    input  [511:0] col_in_27,
    input  [511:0] col_in_28,
    input  [511:0] col_in_29,
    input  [511:0] col_in_30,
    input  [511:0] col_in_31,
    input  [511:0] col_in_32,
    input  [511:0] col_in_33,
    input  [511:0] col_in_34,
    input  [511:0] col_in_35,
    input  [511:0] col_in_36,
    input  [511:0] col_in_37,
    input  [511:0] col_in_38,
    input  [511:0] col_in_39,
    input  [511:0] col_in_40,
    input  [511:0] col_in_41,
    input  [511:0] col_in_42,
    input  [511:0] col_in_43,
    input  [511:0] col_in_44,
    input  [511:0] col_in_45,
    input  [511:0] col_in_46,
    input  [511:0] col_in_47,
    input  [511:0] col_in_48,
    input  [511:0] col_in_49,
    input  [511:0] col_in_50,
    input  [511:0] col_in_51,
    input  [511:0] col_in_52,
    input  [511:0] col_in_53,
    input  [511:0] col_in_54,
    input  [511:0] col_in_55,
    input  [511:0] col_in_56,
    input  [511:0] col_in_57,
    input  [511:0] col_in_58,
    input  [511:0] col_in_59,
    input  [511:0] col_in_60,
    input  [511:0] col_in_61,
    input  [511:0] col_in_62,
    input  [511:0] col_in_63,
    input  [511:0] col_in_64,
    input  [511:0] col_in_65,
    input  [511:0] col_in_66,
    input  [511:0] col_in_67,
    input  [511:0] col_in_68,
    input  [511:0] col_in_69,
    input  [511:0] col_in_70,
    input  [511:0] col_in_71,
    input  [511:0] col_in_72,
    input  [511:0] col_in_73,
    input  [511:0] col_in_74,
    input  [511:0] col_in_75,
    input  [511:0] col_in_76,
    input  [511:0] col_in_77,
    input  [511:0] col_in_78,
    input  [511:0] col_in_79,
    input  [511:0] col_in_80,
    input  [511:0] col_in_81,
    input  [511:0] col_in_82,
    input  [511:0] col_in_83,
    input  [511:0] col_in_84,
    input  [511:0] col_in_85,
    input  [511:0] col_in_86,
    input  [511:0] col_in_87,
    input  [511:0] col_in_88,
    input  [511:0] col_in_89,
    input  [511:0] col_in_90,
    input  [511:0] col_in_91,
    input  [511:0] col_in_92,
    input  [511:0] col_in_93,
    input  [511:0] col_in_94,
    input  [511:0] col_in_95,
    input  [511:0] col_in_96,
    input  [511:0] col_in_97,
    input  [511:0] col_in_98,
    input  [511:0] col_in_99,
    input  [511:0] col_in_100,
    input  [511:0] col_in_101,
    input  [511:0] col_in_102,
    input  [511:0] col_in_103,
    input  [511:0] col_in_104,
    input  [511:0] col_in_105,
    input  [511:0] col_in_106,
    input  [511:0] col_in_107,
    input  [511:0] col_in_108,
    input  [511:0] col_in_109,
    input  [511:0] col_in_110,
    input  [511:0] col_in_111,
    input  [511:0] col_in_112,
    input  [511:0] col_in_113,
    input  [511:0] col_in_114,
    input  [511:0] col_in_115,
    input  [511:0] col_in_116,
    input  [511:0] col_in_117,
    input  [511:0] col_in_118,
    input  [511:0] col_in_119,
    input  [511:0] col_in_120,
    input  [511:0] col_in_121,
    input  [511:0] col_in_122,
    input  [511:0] col_in_123,
    input  [511:0] col_in_124,
    input  [511:0] col_in_125,
    input  [511:0] col_in_126,
    input  [511:0] col_in_127,
    input  [511:0] col_in_128,
    input  [511:0] col_in_129,
    input  [511:0] col_in_130,
    input  [511:0] col_in_131,
    input  [511:0] col_in_132,
    input  [511:0] col_in_133,
    input  [511:0] col_in_134,
    input  [511:0] col_in_135,
    input  [511:0] col_in_136,
    input  [511:0] col_in_137,
    input  [511:0] col_in_138,
    input  [511:0] col_in_139,
    input  [511:0] col_in_140,
    input  [511:0] col_in_141,
    input  [511:0] col_in_142,
    input  [511:0] col_in_143,
    input  [511:0] col_in_144,
    input  [511:0] col_in_145,
    input  [511:0] col_in_146,
    input  [511:0] col_in_147,
    input  [511:0] col_in_148,
    input  [511:0] col_in_149,
    input  [511:0] col_in_150,
    input  [511:0] col_in_151,
    input  [511:0] col_in_152,
    input  [511:0] col_in_153,
    input  [511:0] col_in_154,
    input  [511:0] col_in_155,
    input  [511:0] col_in_156,
    input  [511:0] col_in_157,
    input  [511:0] col_in_158,
    input  [511:0] col_in_159,
    input  [511:0] col_in_160,
    input  [511:0] col_in_161,
    input  [511:0] col_in_162,
    input  [511:0] col_in_163,
    input  [511:0] col_in_164,
    input  [511:0] col_in_165,
    input  [511:0] col_in_166,
    input  [511:0] col_in_167,
    input  [511:0] col_in_168,
    input  [511:0] col_in_169,
    input  [511:0] col_in_170,
    input  [511:0] col_in_171,
    input  [511:0] col_in_172,
    input  [511:0] col_in_173,
    input  [511:0] col_in_174,
    input  [511:0] col_in_175,
    input  [511:0] col_in_176,
    input  [511:0] col_in_177,
    input  [511:0] col_in_178,
    input  [511:0] col_in_179,
    input  [511:0] col_in_180,
    input  [511:0] col_in_181,
    input  [511:0] col_in_182,
    input  [511:0] col_in_183,
    input  [511:0] col_in_184,
    input  [511:0] col_in_185,
    input  [511:0] col_in_186,
    input  [511:0] col_in_187,
    input  [511:0] col_in_188,
    input  [511:0] col_in_189,
    input  [511:0] col_in_190,
    input  [511:0] col_in_191,
    input  [511:0] col_in_192,
    input  [511:0] col_in_193,
    input  [511:0] col_in_194,
    input  [511:0] col_in_195,
    input  [511:0] col_in_196,
    input  [511:0] col_in_197,
    input  [511:0] col_in_198,
    input  [511:0] col_in_199,
    input  [511:0] col_in_200,
    input  [511:0] col_in_201,
    input  [511:0] col_in_202,
    input  [511:0] col_in_203,
    input  [511:0] col_in_204,
    input  [511:0] col_in_205,
    input  [511:0] col_in_206,
    input  [511:0] col_in_207,
    input  [511:0] col_in_208,
    input  [511:0] col_in_209,
    input  [511:0] col_in_210,
    input  [511:0] col_in_211,
    input  [511:0] col_in_212,
    input  [511:0] col_in_213,
    input  [511:0] col_in_214,
    input  [511:0] col_in_215,
    input  [511:0] col_in_216,
    input  [511:0] col_in_217,
    input  [511:0] col_in_218,
    input  [511:0] col_in_219,
    input  [511:0] col_in_220,
    input  [511:0] col_in_221,
    input  [511:0] col_in_222,
    input  [511:0] col_in_223,
    input  [511:0] col_in_224,
    input  [511:0] col_in_225,
    input  [511:0] col_in_226,
    input  [511:0] col_in_227,
    input  [511:0] col_in_228,
    input  [511:0] col_in_229,
    input  [511:0] col_in_230,
    input  [511:0] col_in_231,
    input  [511:0] col_in_232,
    input  [511:0] col_in_233,
    input  [511:0] col_in_234,
    input  [511:0] col_in_235,
    input  [511:0] col_in_236,
    input  [511:0] col_in_237,
    input  [511:0] col_in_238,
    input  [511:0] col_in_239,
    input  [511:0] col_in_240,
    input  [511:0] col_in_241,
    input  [511:0] col_in_242,
    input  [511:0] col_in_243,
    input  [511:0] col_in_244,
    input  [511:0] col_in_245,
    input  [511:0] col_in_246,
    input  [511:0] col_in_247,
    input  [511:0] col_in_248,
    input  [511:0] col_in_249,
    input  [511:0] col_in_250,
    input  [511:0] col_in_251,
    input  [511:0] col_in_252,
    input  [511:0] col_in_253,
    input  [511:0] col_in_254,
    input  [511:0] col_in_255,
    input  [511:0] col_in_256,
    input  [511:0] col_in_257,
    input  [511:0] col_in_258,
    input  [511:0] col_in_259,
    input  [511:0] col_in_260,
    input  [511:0] col_in_261,
    input  [511:0] col_in_262,
    input  [511:0] col_in_263,
    input  [511:0] col_in_264,
    input  [511:0] col_in_265,
    input  [511:0] col_in_266,
    input  [511:0] col_in_267,
    input  [511:0] col_in_268,
    input  [511:0] col_in_269,
    input  [511:0] col_in_270,
    input  [511:0] col_in_271,
    input  [511:0] col_in_272,
    input  [511:0] col_in_273,
    input  [511:0] col_in_274,
    input  [511:0] col_in_275,
    input  [511:0] col_in_276,
    input  [511:0] col_in_277,
    input  [511:0] col_in_278,
    input  [511:0] col_in_279,
    input  [511:0] col_in_280,
    input  [511:0] col_in_281,
    input  [511:0] col_in_282,
    input  [511:0] col_in_283,
    input  [511:0] col_in_284,
    input  [511:0] col_in_285,
    input  [511:0] col_in_286,
    input  [511:0] col_in_287,
    input  [511:0] col_in_288,
    input  [511:0] col_in_289,
    input  [511:0] col_in_290,
    input  [511:0] col_in_291,
    input  [511:0] col_in_292,
    input  [511:0] col_in_293,
    input  [511:0] col_in_294,
    input  [511:0] col_in_295,
    input  [511:0] col_in_296,
    input  [511:0] col_in_297,
    input  [511:0] col_in_298,
    input  [511:0] col_in_299,
    input  [511:0] col_in_300,
    input  [511:0] col_in_301,
    input  [511:0] col_in_302,
    input  [511:0] col_in_303,
    input  [511:0] col_in_304,
    input  [511:0] col_in_305,
    input  [511:0] col_in_306,
    input  [511:0] col_in_307,
    input  [511:0] col_in_308,
    input  [511:0] col_in_309,
    input  [511:0] col_in_310,
    input  [511:0] col_in_311,
    input  [511:0] col_in_312,
    input  [511:0] col_in_313,
    input  [511:0] col_in_314,
    input  [511:0] col_in_315,
    input  [511:0] col_in_316,
    input  [511:0] col_in_317,
    input  [511:0] col_in_318,
    input  [511:0] col_in_319,
    input  [511:0] col_in_320,
    input  [511:0] col_in_321,
    input  [511:0] col_in_322,
    input  [511:0] col_in_323,
    input  [511:0] col_in_324,
    input  [511:0] col_in_325,
    input  [511:0] col_in_326,
    input  [511:0] col_in_327,
    input  [511:0] col_in_328,
    input  [511:0] col_in_329,
    input  [511:0] col_in_330,
    input  [511:0] col_in_331,
    input  [511:0] col_in_332,
    input  [511:0] col_in_333,
    input  [511:0] col_in_334,
    input  [511:0] col_in_335,
    input  [511:0] col_in_336,
    input  [511:0] col_in_337,
    input  [511:0] col_in_338,
    input  [511:0] col_in_339,
    input  [511:0] col_in_340,
    input  [511:0] col_in_341,
    input  [511:0] col_in_342,
    input  [511:0] col_in_343,
    input  [511:0] col_in_344,
    input  [511:0] col_in_345,
    input  [511:0] col_in_346,
    input  [511:0] col_in_347,
    input  [511:0] col_in_348,
    input  [511:0] col_in_349,
    input  [511:0] col_in_350,
    input  [511:0] col_in_351,
    input  [511:0] col_in_352,
    input  [511:0] col_in_353,
    input  [511:0] col_in_354,
    input  [511:0] col_in_355,
    input  [511:0] col_in_356,
    input  [511:0] col_in_357,
    input  [511:0] col_in_358,
    input  [511:0] col_in_359,
    input  [511:0] col_in_360,
    input  [511:0] col_in_361,
    input  [511:0] col_in_362,
    input  [511:0] col_in_363,
    input  [511:0] col_in_364,
    input  [511:0] col_in_365,
    input  [511:0] col_in_366,
    input  [511:0] col_in_367,
    input  [511:0] col_in_368,
    input  [511:0] col_in_369,
    input  [511:0] col_in_370,
    input  [511:0] col_in_371,
    input  [511:0] col_in_372,
    input  [511:0] col_in_373,
    input  [511:0] col_in_374,
    input  [511:0] col_in_375,
    input  [511:0] col_in_376,
    input  [511:0] col_in_377,
    input  [511:0] col_in_378,
    input  [511:0] col_in_379,
    input  [511:0] col_in_380,
    input  [511:0] col_in_381,
    input  [511:0] col_in_382,
    input  [511:0] col_in_383,
    input  [511:0] col_in_384,
    input  [511:0] col_in_385,
    input  [511:0] col_in_386,
    input  [511:0] col_in_387,
    input  [511:0] col_in_388,
    input  [511:0] col_in_389,
    input  [511:0] col_in_390,
    input  [511:0] col_in_391,
    input  [511:0] col_in_392,
    input  [511:0] col_in_393,
    input  [511:0] col_in_394,
    input  [511:0] col_in_395,
    input  [511:0] col_in_396,
    input  [511:0] col_in_397,
    input  [511:0] col_in_398,
    input  [511:0] col_in_399,
    input  [511:0] col_in_400,
    input  [511:0] col_in_401,
    input  [511:0] col_in_402,
    input  [511:0] col_in_403,
    input  [511:0] col_in_404,
    input  [511:0] col_in_405,
    input  [511:0] col_in_406,
    input  [511:0] col_in_407,
    input  [511:0] col_in_408,
    input  [511:0] col_in_409,
    input  [511:0] col_in_410,
    input  [511:0] col_in_411,
    input  [511:0] col_in_412,
    input  [511:0] col_in_413,
    input  [511:0] col_in_414,
    input  [511:0] col_in_415,
    input  [511:0] col_in_416,
    input  [511:0] col_in_417,
    input  [511:0] col_in_418,
    input  [511:0] col_in_419,
    input  [511:0] col_in_420,
    input  [511:0] col_in_421,
    input  [511:0] col_in_422,
    input  [511:0] col_in_423,
    input  [511:0] col_in_424,
    input  [511:0] col_in_425,
    input  [511:0] col_in_426,
    input  [511:0] col_in_427,
    input  [511:0] col_in_428,
    input  [511:0] col_in_429,
    input  [511:0] col_in_430,
    input  [511:0] col_in_431,
    input  [511:0] col_in_432,
    input  [511:0] col_in_433,
    input  [511:0] col_in_434,
    input  [511:0] col_in_435,
    input  [511:0] col_in_436,
    input  [511:0] col_in_437,
    input  [511:0] col_in_438,
    input  [511:0] col_in_439,
    input  [511:0] col_in_440,
    input  [511:0] col_in_441,
    input  [511:0] col_in_442,
    input  [511:0] col_in_443,
    input  [511:0] col_in_444,
    input  [511:0] col_in_445,
    input  [511:0] col_in_446,
    input  [511:0] col_in_447,
    input  [511:0] col_in_448,
    input  [511:0] col_in_449,
    input  [511:0] col_in_450,
    input  [511:0] col_in_451,
    input  [511:0] col_in_452,
    input  [511:0] col_in_453,
    input  [511:0] col_in_454,
    input  [511:0] col_in_455,
    input  [511:0] col_in_456,
    input  [511:0] col_in_457,
    input  [511:0] col_in_458,
    input  [511:0] col_in_459,
    input  [511:0] col_in_460,
    input  [511:0] col_in_461,
    input  [511:0] col_in_462,
    input  [511:0] col_in_463,
    input  [511:0] col_in_464,
    input  [511:0] col_in_465,
    input  [511:0] col_in_466,
    input  [511:0] col_in_467,
    input  [511:0] col_in_468,
    input  [511:0] col_in_469,
    input  [511:0] col_in_470,
    input  [511:0] col_in_471,
    input  [511:0] col_in_472,
    input  [511:0] col_in_473,
    input  [511:0] col_in_474,
    input  [511:0] col_in_475,
    input  [511:0] col_in_476,
    input  [511:0] col_in_477,
    input  [511:0] col_in_478,
    input  [511:0] col_in_479,
    input  [511:0] col_in_480,
    input  [511:0] col_in_481,
    input  [511:0] col_in_482,
    input  [511:0] col_in_483,
    input  [511:0] col_in_484,
    input  [511:0] col_in_485,
    input  [511:0] col_in_486,
    input  [511:0] col_in_487,
    input  [511:0] col_in_488,
    input  [511:0] col_in_489,
    input  [511:0] col_in_490,
    input  [511:0] col_in_491,
    input  [511:0] col_in_492,
    input  [511:0] col_in_493,
    input  [511:0] col_in_494,
    input  [511:0] col_in_495,
    input  [511:0] col_in_496,
    input  [511:0] col_in_497,
    input  [511:0] col_in_498,
    input  [511:0] col_in_499,
    input  [511:0] col_in_500,
    input  [511:0] col_in_501,
    input  [511:0] col_in_502,
    input  [511:0] col_in_503,
    input  [511:0] col_in_504,
    input  [511:0] col_in_505,
    input  [511:0] col_in_506,
    input  [511:0] col_in_507,
    input  [511:0] col_in_508,
    input  [511:0] col_in_509,
    input  [511:0] col_in_510,
    input  [511:0] col_in_511,
    input  [511:0] col_in_512,
    input  [511:0] col_in_513,
    input  [511:0] col_in_514,
    input  [511:0] col_in_515,
    input  [511:0] col_in_516,
    input  [511:0] col_in_517,
    input  [511:0] col_in_518,
    input  [511:0] col_in_519,
    input  [511:0] col_in_520,
    input  [511:0] col_in_521,
    input  [511:0] col_in_522,
    input  [511:0] col_in_523,
    input  [511:0] col_in_524,
    input  [511:0] col_in_525,
    input  [511:0] col_in_526,
    input  [511:0] col_in_527,
    input  [511:0] col_in_528,
    input  [511:0] col_in_529,
    input  [511:0] col_in_530,
    input  [511:0] col_in_531,
    input  [511:0] col_in_532,
    input  [511:0] col_in_533,
    input  [511:0] col_in_534,
    input  [511:0] col_in_535,
    input  [511:0] col_in_536,
    input  [511:0] col_in_537,
    input  [511:0] col_in_538,
    input  [511:0] col_in_539,
    input  [511:0] col_in_540,
    input  [511:0] col_in_541,
    input  [511:0] col_in_542,
    input  [511:0] col_in_543,
    input  [511:0] col_in_544,
    input  [511:0] col_in_545,
    input  [511:0] col_in_546,
    input  [511:0] col_in_547,
    input  [511:0] col_in_548,
    input  [511:0] col_in_549,
    input  [511:0] col_in_550,
    input  [511:0] col_in_551,
    input  [511:0] col_in_552,
    input  [511:0] col_in_553,
    input  [511:0] col_in_554,
    input  [511:0] col_in_555,
    input  [511:0] col_in_556,
    input  [511:0] col_in_557,
    input  [511:0] col_in_558,
    input  [511:0] col_in_559,
    input  [511:0] col_in_560,
    input  [511:0] col_in_561,
    input  [511:0] col_in_562,
    input  [511:0] col_in_563,
    input  [511:0] col_in_564,
    input  [511:0] col_in_565,
    input  [511:0] col_in_566,
    input  [511:0] col_in_567,
    input  [511:0] col_in_568,
    input  [511:0] col_in_569,
    input  [511:0] col_in_570,
    input  [511:0] col_in_571,
    input  [511:0] col_in_572,
    input  [511:0] col_in_573,
    input  [511:0] col_in_574,
    input  [511:0] col_in_575,
    input  [511:0] col_in_576,
    input  [511:0] col_in_577,
    input  [511:0] col_in_578,
    input  [511:0] col_in_579,
    input  [511:0] col_in_580,
    input  [511:0] col_in_581,
    input  [511:0] col_in_582,
    input  [511:0] col_in_583,
    input  [511:0] col_in_584,
    input  [511:0] col_in_585,
    input  [511:0] col_in_586,
    input  [511:0] col_in_587,
    input  [511:0] col_in_588,
    input  [511:0] col_in_589,
    input  [511:0] col_in_590,
    input  [511:0] col_in_591,
    input  [511:0] col_in_592,
    input  [511:0] col_in_593,
    input  [511:0] col_in_594,
    input  [511:0] col_in_595,
    input  [511:0] col_in_596,
    input  [511:0] col_in_597,
    input  [511:0] col_in_598,
    input  [511:0] col_in_599,
    input  [511:0] col_in_600,
    input  [511:0] col_in_601,
    input  [511:0] col_in_602,
    input  [511:0] col_in_603,
    input  [511:0] col_in_604,
    input  [511:0] col_in_605,
    input  [511:0] col_in_606,
    input  [511:0] col_in_607,
    input  [511:0] col_in_608,
    input  [511:0] col_in_609,
    input  [511:0] col_in_610,
    input  [511:0] col_in_611,
    input  [511:0] col_in_612,
    input  [511:0] col_in_613,
    input  [511:0] col_in_614,
    input  [511:0] col_in_615,
    input  [511:0] col_in_616,
    input  [511:0] col_in_617,
    input  [511:0] col_in_618,
    input  [511:0] col_in_619,
    input  [511:0] col_in_620,
    input  [511:0] col_in_621,
    input  [511:0] col_in_622,
    input  [511:0] col_in_623,
    input  [511:0] col_in_624,
    input  [511:0] col_in_625,
    input  [511:0] col_in_626,
    input  [511:0] col_in_627,
    input  [511:0] col_in_628,
    input  [511:0] col_in_629,
    input  [511:0] col_in_630,
    input  [511:0] col_in_631,
    input  [511:0] col_in_632,
    input  [511:0] col_in_633,
    input  [511:0] col_in_634,
    input  [511:0] col_in_635,
    input  [511:0] col_in_636,
    input  [511:0] col_in_637,
    input  [511:0] col_in_638,
    input  [511:0] col_in_639,
    input  [511:0] col_in_640,
    input  [511:0] col_in_641,
    input  [511:0] col_in_642,
    input  [511:0] col_in_643,
    input  [511:0] col_in_644,
    input  [511:0] col_in_645,
    input  [511:0] col_in_646,
    input  [511:0] col_in_647,
    input  [511:0] col_in_648,
    input  [511:0] col_in_649,
    input  [511:0] col_in_650,
    input  [511:0] col_in_651,
    input  [511:0] col_in_652,
    input  [511:0] col_in_653,
    input  [511:0] col_in_654,
    input  [511:0] col_in_655,
    input  [511:0] col_in_656,
    input  [511:0] col_in_657,
    input  [511:0] col_in_658,
    input  [511:0] col_in_659,
    input  [511:0] col_in_660,
    input  [511:0] col_in_661,
    input  [511:0] col_in_662,
    input  [511:0] col_in_663,
    input  [511:0] col_in_664,
    input  [511:0] col_in_665,
    input  [511:0] col_in_666,
    input  [511:0] col_in_667,
    input  [511:0] col_in_668,
    input  [511:0] col_in_669,
    input  [511:0] col_in_670,
    input  [511:0] col_in_671,
    input  [511:0] col_in_672,
    input  [511:0] col_in_673,
    input  [511:0] col_in_674,
    input  [511:0] col_in_675,
    input  [511:0] col_in_676,
    input  [511:0] col_in_677,
    input  [511:0] col_in_678,
    input  [511:0] col_in_679,
    input  [511:0] col_in_680,
    input  [511:0] col_in_681,
    input  [511:0] col_in_682,
    input  [511:0] col_in_683,
    input  [511:0] col_in_684,
    input  [511:0] col_in_685,
    input  [511:0] col_in_686,
    input  [511:0] col_in_687,
    input  [511:0] col_in_688,
    input  [511:0] col_in_689,
    input  [511:0] col_in_690,
    input  [511:0] col_in_691,
    input  [511:0] col_in_692,
    input  [511:0] col_in_693,
    input  [511:0] col_in_694,
    input  [511:0] col_in_695,
    input  [511:0] col_in_696,
    input  [511:0] col_in_697,
    input  [511:0] col_in_698,
    input  [511:0] col_in_699,
    input  [511:0] col_in_700,
    input  [511:0] col_in_701,
    input  [511:0] col_in_702,
    input  [511:0] col_in_703,
    input  [511:0] col_in_704,
    input  [511:0] col_in_705,
    input  [511:0] col_in_706,
    input  [511:0] col_in_707,
    input  [511:0] col_in_708,
    input  [511:0] col_in_709,
    input  [511:0] col_in_710,
    input  [511:0] col_in_711,
    input  [511:0] col_in_712,
    input  [511:0] col_in_713,
    input  [511:0] col_in_714,
    input  [511:0] col_in_715,
    input  [511:0] col_in_716,
    input  [511:0] col_in_717,
    input  [511:0] col_in_718,
    input  [511:0] col_in_719,
    input  [511:0] col_in_720,
    input  [511:0] col_in_721,
    input  [511:0] col_in_722,
    input  [511:0] col_in_723,
    input  [511:0] col_in_724,
    input  [511:0] col_in_725,
    input  [511:0] col_in_726,
    input  [511:0] col_in_727,
    input  [511:0] col_in_728,
    input  [511:0] col_in_729,
    input  [511:0] col_in_730,
    input  [511:0] col_in_731,
    input  [511:0] col_in_732,
    input  [511:0] col_in_733,
    input  [511:0] col_in_734,
    input  [511:0] col_in_735,
    input  [511:0] col_in_736,
    input  [511:0] col_in_737,
    input  [511:0] col_in_738,
    input  [511:0] col_in_739,
    input  [511:0] col_in_740,
    input  [511:0] col_in_741,
    input  [511:0] col_in_742,
    input  [511:0] col_in_743,
    input  [511:0] col_in_744,
    input  [511:0] col_in_745,
    input  [511:0] col_in_746,
    input  [511:0] col_in_747,
    input  [511:0] col_in_748,
    input  [511:0] col_in_749,
    input  [511:0] col_in_750,
    input  [511:0] col_in_751,
    input  [511:0] col_in_752,
    input  [511:0] col_in_753,
    input  [511:0] col_in_754,
    input  [511:0] col_in_755,
    input  [511:0] col_in_756,
    input  [511:0] col_in_757,
    input  [511:0] col_in_758,
    input  [511:0] col_in_759,
    input  [511:0] col_in_760,
    input  [511:0] col_in_761,
    input  [511:0] col_in_762,
    input  [511:0] col_in_763,
    input  [511:0] col_in_764,
    input  [511:0] col_in_765,
    input  [511:0] col_in_766,
    input  [511:0] col_in_767,
    input  [511:0] col_in_768,
    input  [511:0] col_in_769,
    input  [511:0] col_in_770,
    input  [511:0] col_in_771,
    input  [511:0] col_in_772,
    input  [511:0] col_in_773,
    input  [511:0] col_in_774,
    input  [511:0] col_in_775,
    input  [511:0] col_in_776,
    input  [511:0] col_in_777,
    input  [511:0] col_in_778,
    input  [511:0] col_in_779,
    input  [511:0] col_in_780,
    input  [511:0] col_in_781,
    input  [511:0] col_in_782,
    input  [511:0] col_in_783,
    input  [511:0] col_in_784,
    input  [511:0] col_in_785,
    input  [511:0] col_in_786,
    input  [511:0] col_in_787,
    input  [511:0] col_in_788,
    input  [511:0] col_in_789,
    input  [511:0] col_in_790,
    input  [511:0] col_in_791,
    input  [511:0] col_in_792,
    input  [511:0] col_in_793,
    input  [511:0] col_in_794,
    input  [511:0] col_in_795,
    input  [511:0] col_in_796,
    input  [511:0] col_in_797,
    input  [511:0] col_in_798,
    input  [511:0] col_in_799,
    input  [511:0] col_in_800,
    input  [511:0] col_in_801,
    input  [511:0] col_in_802,
    input  [511:0] col_in_803,
    input  [511:0] col_in_804,
    input  [511:0] col_in_805,
    input  [511:0] col_in_806,
    input  [511:0] col_in_807,
    input  [511:0] col_in_808,
    input  [511:0] col_in_809,
    input  [511:0] col_in_810,
    input  [511:0] col_in_811,
    input  [511:0] col_in_812,
    input  [511:0] col_in_813,
    input  [511:0] col_in_814,
    input  [511:0] col_in_815,
    input  [511:0] col_in_816,
    input  [511:0] col_in_817,
    input  [511:0] col_in_818,
    input  [511:0] col_in_819,
    input  [511:0] col_in_820,
    input  [511:0] col_in_821,
    input  [511:0] col_in_822,
    input  [511:0] col_in_823,
    input  [511:0] col_in_824,
    input  [511:0] col_in_825,
    input  [511:0] col_in_826,
    input  [511:0] col_in_827,
    input  [511:0] col_in_828,
    input  [511:0] col_in_829,
    input  [511:0] col_in_830,
    input  [511:0] col_in_831,
    input  [511:0] col_in_832,
    input  [511:0] col_in_833,
    input  [511:0] col_in_834,
    input  [511:0] col_in_835,
    input  [511:0] col_in_836,
    input  [511:0] col_in_837,
    input  [511:0] col_in_838,
    input  [511:0] col_in_839,
    input  [511:0] col_in_840,
    input  [511:0] col_in_841,
    input  [511:0] col_in_842,
    input  [511:0] col_in_843,
    input  [511:0] col_in_844,
    input  [511:0] col_in_845,
    input  [511:0] col_in_846,
    input  [511:0] col_in_847,
    input  [511:0] col_in_848,
    input  [511:0] col_in_849,
    input  [511:0] col_in_850,
    input  [511:0] col_in_851,
    input  [511:0] col_in_852,
    input  [511:0] col_in_853,
    input  [511:0] col_in_854,
    input  [511:0] col_in_855,
    input  [511:0] col_in_856,
    input  [511:0] col_in_857,
    input  [511:0] col_in_858,
    input  [511:0] col_in_859,
    input  [511:0] col_in_860,
    input  [511:0] col_in_861,
    input  [511:0] col_in_862,
    input  [511:0] col_in_863,
    input  [511:0] col_in_864,
    input  [511:0] col_in_865,
    input  [511:0] col_in_866,
    input  [511:0] col_in_867,
    input  [511:0] col_in_868,
    input  [511:0] col_in_869,
    input  [511:0] col_in_870,
    input  [511:0] col_in_871,
    input  [511:0] col_in_872,
    input  [511:0] col_in_873,
    input  [511:0] col_in_874,
    input  [511:0] col_in_875,
    input  [511:0] col_in_876,
    input  [511:0] col_in_877,
    input  [511:0] col_in_878,
    input  [511:0] col_in_879,
    input  [511:0] col_in_880,
    input  [511:0] col_in_881,
    input  [511:0] col_in_882,
    input  [511:0] col_in_883,
    input  [511:0] col_in_884,
    input  [511:0] col_in_885,
    input  [511:0] col_in_886,
    input  [511:0] col_in_887,
    input  [511:0] col_in_888,
    input  [511:0] col_in_889,
    input  [511:0] col_in_890,
    input  [511:0] col_in_891,
    input  [511:0] col_in_892,
    input  [511:0] col_in_893,
    input  [511:0] col_in_894,
    input  [511:0] col_in_895,
    input  [511:0] col_in_896,
    input  [511:0] col_in_897,
    input  [511:0] col_in_898,
    input  [511:0] col_in_899,
    input  [511:0] col_in_900,
    input  [511:0] col_in_901,
    input  [511:0] col_in_902,
    input  [511:0] col_in_903,
    input  [511:0] col_in_904,
    input  [511:0] col_in_905,
    input  [511:0] col_in_906,
    input  [511:0] col_in_907,
    input  [511:0] col_in_908,
    input  [511:0] col_in_909,
    input  [511:0] col_in_910,
    input  [511:0] col_in_911,
    input  [511:0] col_in_912,
    input  [511:0] col_in_913,
    input  [511:0] col_in_914,
    input  [511:0] col_in_915,
    input  [511:0] col_in_916,
    input  [511:0] col_in_917,
    input  [511:0] col_in_918,
    input  [511:0] col_in_919,
    input  [511:0] col_in_920,
    input  [511:0] col_in_921,
    input  [511:0] col_in_922,
    input  [511:0] col_in_923,
    input  [511:0] col_in_924,
    input  [511:0] col_in_925,
    input  [511:0] col_in_926,
    input  [511:0] col_in_927,
    input  [511:0] col_in_928,
    input  [511:0] col_in_929,
    input  [511:0] col_in_930,
    input  [511:0] col_in_931,
    input  [511:0] col_in_932,
    input  [511:0] col_in_933,
    input  [511:0] col_in_934,
    input  [511:0] col_in_935,
    input  [511:0] col_in_936,
    input  [511:0] col_in_937,
    input  [511:0] col_in_938,
    input  [511:0] col_in_939,
    input  [511:0] col_in_940,
    input  [511:0] col_in_941,
    input  [511:0] col_in_942,
    input  [511:0] col_in_943,
    input  [511:0] col_in_944,
    input  [511:0] col_in_945,
    input  [511:0] col_in_946,
    input  [511:0] col_in_947,
    input  [511:0] col_in_948,
    input  [511:0] col_in_949,
    input  [511:0] col_in_950,
    input  [511:0] col_in_951,
    input  [511:0] col_in_952,
    input  [511:0] col_in_953,
    input  [511:0] col_in_954,
    input  [511:0] col_in_955,
    input  [511:0] col_in_956,
    input  [511:0] col_in_957,
    input  [511:0] col_in_958,
    input  [511:0] col_in_959,
    input  [511:0] col_in_960,
    input  [511:0] col_in_961,
    input  [511:0] col_in_962,
    input  [511:0] col_in_963,
    input  [511:0] col_in_964,
    input  [511:0] col_in_965,
    input  [511:0] col_in_966,
    input  [511:0] col_in_967,
    input  [511:0] col_in_968,
    input  [511:0] col_in_969,
    input  [511:0] col_in_970,
    input  [511:0] col_in_971,
    input  [511:0] col_in_972,
    input  [511:0] col_in_973,
    input  [511:0] col_in_974,
    input  [511:0] col_in_975,
    input  [511:0] col_in_976,
    input  [511:0] col_in_977,
    input  [511:0] col_in_978,
    input  [511:0] col_in_979,
    input  [511:0] col_in_980,
    input  [511:0] col_in_981,
    input  [511:0] col_in_982,
    input  [511:0] col_in_983,
    input  [511:0] col_in_984,
    input  [511:0] col_in_985,
    input  [511:0] col_in_986,
    input  [511:0] col_in_987,
    input  [511:0] col_in_988,
    input  [511:0] col_in_989,
    input  [511:0] col_in_990,
    input  [511:0] col_in_991,
    input  [511:0] col_in_992,
    input  [511:0] col_in_993,
    input  [511:0] col_in_994,
    input  [511:0] col_in_995,
    input  [511:0] col_in_996,
    input  [511:0] col_in_997,
    input  [511:0] col_in_998,
    input  [511:0] col_in_999,
    input  [511:0] col_in_1000,
    input  [511:0] col_in_1001,
    input  [511:0] col_in_1002,
    input  [511:0] col_in_1003,
    input  [511:0] col_in_1004,
    input  [511:0] col_in_1005,
    input  [511:0] col_in_1006,
    input  [511:0] col_in_1007,
    input  [511:0] col_in_1008,
    input  [511:0] col_in_1009,
    input  [511:0] col_in_1010,
    input  [511:0] col_in_1011,
    input  [511:0] col_in_1012,
    input  [511:0] col_in_1013,
    input  [511:0] col_in_1014,
    input  [511:0] col_in_1015,
    input  [511:0] col_in_1016,
    input  [511:0] col_in_1017,
    input  [511:0] col_in_1018,
    input  [511:0] col_in_1019,
    input  [511:0] col_in_1020,
    input  [511:0] col_in_1021,
    input  [511:0] col_in_1022,
    input  [511:0] col_in_1023,




    output [15:0] col_out_0,
    output [15:0] col_out_1,
    output [15:0] col_out_2,
    output [15:0] col_out_3,
    output [15:0] col_out_4,
    output [15:0] col_out_5,
    output [15:0] col_out_6,
    output [15:0] col_out_7,
    output [15:0] col_out_8,
    output [15:0] col_out_9,
    output [15:0] col_out_10,
    output [15:0] col_out_11,
    output [15:0] col_out_12,
    output [15:0] col_out_13,
    output [15:0] col_out_14,
    output [15:0] col_out_15,
    output [15:0] col_out_16,
    output [15:0] col_out_17,
    output [15:0] col_out_18,
    output [15:0] col_out_19,
    output [15:0] col_out_20,
    output [15:0] col_out_21,
    output [15:0] col_out_22,
    output [15:0] col_out_23,
    output [15:0] col_out_24,
    output [15:0] col_out_25,
    output [15:0] col_out_26,
    output [15:0] col_out_27,
    output [15:0] col_out_28,
    output [15:0] col_out_29,
    output [15:0] col_out_30,
    output [15:0] col_out_31,
    output [15:0] col_out_32,
    output [15:0] col_out_33,
    output [15:0] col_out_34,
    output [15:0] col_out_35,
    output [15:0] col_out_36,
    output [15:0] col_out_37,
    output [15:0] col_out_38,
    output [15:0] col_out_39,
    output [15:0] col_out_40,
    output [15:0] col_out_41,
    output [15:0] col_out_42,
    output [15:0] col_out_43,
    output [15:0] col_out_44,
    output [15:0] col_out_45,
    output [15:0] col_out_46,
    output [15:0] col_out_47,
    output [15:0] col_out_48,
    output [15:0] col_out_49,
    output [15:0] col_out_50,
    output [15:0] col_out_51,
    output [15:0] col_out_52,
    output [15:0] col_out_53,
    output [15:0] col_out_54,
    output [15:0] col_out_55,
    output [15:0] col_out_56,
    output [15:0] col_out_57,
    output [15:0] col_out_58,
    output [15:0] col_out_59,
    output [15:0] col_out_60,
    output [15:0] col_out_61,
    output [15:0] col_out_62,
    output [15:0] col_out_63,
    output [15:0] col_out_64,
    output [15:0] col_out_65,
    output [15:0] col_out_66,
    output [15:0] col_out_67,
    output [15:0] col_out_68,
    output [15:0] col_out_69,
    output [15:0] col_out_70,
    output [15:0] col_out_71,
    output [15:0] col_out_72,
    output [15:0] col_out_73,
    output [15:0] col_out_74,
    output [15:0] col_out_75,
    output [15:0] col_out_76,
    output [15:0] col_out_77,
    output [15:0] col_out_78,
    output [15:0] col_out_79,
    output [15:0] col_out_80,
    output [15:0] col_out_81,
    output [15:0] col_out_82,
    output [15:0] col_out_83,
    output [15:0] col_out_84,
    output [15:0] col_out_85,
    output [15:0] col_out_86,
    output [15:0] col_out_87,
    output [15:0] col_out_88,
    output [15:0] col_out_89,
    output [15:0] col_out_90,
    output [15:0] col_out_91,
    output [15:0] col_out_92,
    output [15:0] col_out_93,
    output [15:0] col_out_94,
    output [15:0] col_out_95,
    output [15:0] col_out_96,
    output [15:0] col_out_97,
    output [15:0] col_out_98,
    output [15:0] col_out_99,
    output [15:0] col_out_100,
    output [15:0] col_out_101,
    output [15:0] col_out_102,
    output [15:0] col_out_103,
    output [15:0] col_out_104,
    output [15:0] col_out_105,
    output [15:0] col_out_106,
    output [15:0] col_out_107,
    output [15:0] col_out_108,
    output [15:0] col_out_109,
    output [15:0] col_out_110,
    output [15:0] col_out_111,
    output [15:0] col_out_112,
    output [15:0] col_out_113,
    output [15:0] col_out_114,
    output [15:0] col_out_115,
    output [15:0] col_out_116,
    output [15:0] col_out_117,
    output [15:0] col_out_118,
    output [15:0] col_out_119,
    output [15:0] col_out_120,
    output [15:0] col_out_121,
    output [15:0] col_out_122,
    output [15:0] col_out_123,
    output [15:0] col_out_124,
    output [15:0] col_out_125,
    output [15:0] col_out_126,
    output [15:0] col_out_127,
    output [15:0] col_out_128,
    output [15:0] col_out_129,
    output [15:0] col_out_130,
    output [15:0] col_out_131,
    output [15:0] col_out_132,
    output [15:0] col_out_133,
    output [15:0] col_out_134,
    output [15:0] col_out_135,
    output [15:0] col_out_136,
    output [15:0] col_out_137,
    output [15:0] col_out_138,
    output [15:0] col_out_139,
    output [15:0] col_out_140,
    output [15:0] col_out_141,
    output [15:0] col_out_142,
    output [15:0] col_out_143,
    output [15:0] col_out_144,
    output [15:0] col_out_145,
    output [15:0] col_out_146,
    output [15:0] col_out_147,
    output [15:0] col_out_148,
    output [15:0] col_out_149,
    output [15:0] col_out_150,
    output [15:0] col_out_151,
    output [15:0] col_out_152,
    output [15:0] col_out_153,
    output [15:0] col_out_154,
    output [15:0] col_out_155,
    output [15:0] col_out_156,
    output [15:0] col_out_157,
    output [15:0] col_out_158,
    output [15:0] col_out_159,
    output [15:0] col_out_160,
    output [15:0] col_out_161,
    output [15:0] col_out_162,
    output [15:0] col_out_163,
    output [15:0] col_out_164,
    output [15:0] col_out_165,
    output [15:0] col_out_166,
    output [15:0] col_out_167,
    output [15:0] col_out_168,
    output [15:0] col_out_169,
    output [15:0] col_out_170,
    output [15:0] col_out_171,
    output [15:0] col_out_172,
    output [15:0] col_out_173,
    output [15:0] col_out_174,
    output [15:0] col_out_175,
    output [15:0] col_out_176,
    output [15:0] col_out_177,
    output [15:0] col_out_178,
    output [15:0] col_out_179,
    output [15:0] col_out_180,
    output [15:0] col_out_181,
    output [15:0] col_out_182,
    output [15:0] col_out_183,
    output [15:0] col_out_184,
    output [15:0] col_out_185,
    output [15:0] col_out_186,
    output [15:0] col_out_187,
    output [15:0] col_out_188,
    output [15:0] col_out_189,
    output [15:0] col_out_190,
    output [15:0] col_out_191,
    output [15:0] col_out_192,
    output [15:0] col_out_193,
    output [15:0] col_out_194,
    output [15:0] col_out_195,
    output [15:0] col_out_196,
    output [15:0] col_out_197,
    output [15:0] col_out_198,
    output [15:0] col_out_199,
    output [15:0] col_out_200,
    output [15:0] col_out_201,
    output [15:0] col_out_202,
    output [15:0] col_out_203,
    output [15:0] col_out_204,
    output [15:0] col_out_205,
    output [15:0] col_out_206,
    output [15:0] col_out_207,
    output [15:0] col_out_208,
    output [15:0] col_out_209,
    output [15:0] col_out_210,
    output [15:0] col_out_211,
    output [15:0] col_out_212,
    output [15:0] col_out_213,
    output [15:0] col_out_214,
    output [15:0] col_out_215,
    output [15:0] col_out_216,
    output [15:0] col_out_217,
    output [15:0] col_out_218,
    output [15:0] col_out_219,
    output [15:0] col_out_220,
    output [15:0] col_out_221,
    output [15:0] col_out_222,
    output [15:0] col_out_223,
    output [15:0] col_out_224,
    output [15:0] col_out_225,
    output [15:0] col_out_226,
    output [15:0] col_out_227,
    output [15:0] col_out_228,
    output [15:0] col_out_229,
    output [15:0] col_out_230,
    output [15:0] col_out_231,
    output [15:0] col_out_232,
    output [15:0] col_out_233,
    output [15:0] col_out_234,
    output [15:0] col_out_235,
    output [15:0] col_out_236,
    output [15:0] col_out_237,
    output [15:0] col_out_238,
    output [15:0] col_out_239,
    output [15:0] col_out_240,
    output [15:0] col_out_241,
    output [15:0] col_out_242,
    output [15:0] col_out_243,
    output [15:0] col_out_244,
    output [15:0] col_out_245,
    output [15:0] col_out_246,
    output [15:0] col_out_247,
    output [15:0] col_out_248,
    output [15:0] col_out_249,
    output [15:0] col_out_250,
    output [15:0] col_out_251,
    output [15:0] col_out_252,
    output [15:0] col_out_253,
    output [15:0] col_out_254,
    output [15:0] col_out_255,
    output [15:0] col_out_256,
    output [15:0] col_out_257,
    output [15:0] col_out_258,
    output [15:0] col_out_259,
    output [15:0] col_out_260,
    output [15:0] col_out_261,
    output [15:0] col_out_262,
    output [15:0] col_out_263,
    output [15:0] col_out_264,
    output [15:0] col_out_265,
    output [15:0] col_out_266,
    output [15:0] col_out_267,
    output [15:0] col_out_268,
    output [15:0] col_out_269,
    output [15:0] col_out_270,
    output [15:0] col_out_271,
    output [15:0] col_out_272,
    output [15:0] col_out_273,
    output [15:0] col_out_274,
    output [15:0] col_out_275,
    output [15:0] col_out_276,
    output [15:0] col_out_277,
    output [15:0] col_out_278,
    output [15:0] col_out_279,
    output [15:0] col_out_280,
    output [15:0] col_out_281,
    output [15:0] col_out_282,
    output [15:0] col_out_283,
    output [15:0] col_out_284,
    output [15:0] col_out_285,
    output [15:0] col_out_286,
    output [15:0] col_out_287,
    output [15:0] col_out_288,
    output [15:0] col_out_289,
    output [15:0] col_out_290,
    output [15:0] col_out_291,
    output [15:0] col_out_292,
    output [15:0] col_out_293,
    output [15:0] col_out_294,
    output [15:0] col_out_295,
    output [15:0] col_out_296,
    output [15:0] col_out_297,
    output [15:0] col_out_298,
    output [15:0] col_out_299,
    output [15:0] col_out_300,
    output [15:0] col_out_301,
    output [15:0] col_out_302,
    output [15:0] col_out_303,
    output [15:0] col_out_304,
    output [15:0] col_out_305,
    output [15:0] col_out_306,
    output [15:0] col_out_307,
    output [15:0] col_out_308,
    output [15:0] col_out_309,
    output [15:0] col_out_310,
    output [15:0] col_out_311,
    output [15:0] col_out_312,
    output [15:0] col_out_313,
    output [15:0] col_out_314,
    output [15:0] col_out_315,
    output [15:0] col_out_316,
    output [15:0] col_out_317,
    output [15:0] col_out_318,
    output [15:0] col_out_319,
    output [15:0] col_out_320,
    output [15:0] col_out_321,
    output [15:0] col_out_322,
    output [15:0] col_out_323,
    output [15:0] col_out_324,
    output [15:0] col_out_325,
    output [15:0] col_out_326,
    output [15:0] col_out_327,
    output [15:0] col_out_328,
    output [15:0] col_out_329,
    output [15:0] col_out_330,
    output [15:0] col_out_331,
    output [15:0] col_out_332,
    output [15:0] col_out_333,
    output [15:0] col_out_334,
    output [15:0] col_out_335,
    output [15:0] col_out_336,
    output [15:0] col_out_337,
    output [15:0] col_out_338,
    output [15:0] col_out_339,
    output [15:0] col_out_340,
    output [15:0] col_out_341,
    output [15:0] col_out_342,
    output [15:0] col_out_343,
    output [15:0] col_out_344,
    output [15:0] col_out_345,
    output [15:0] col_out_346,
    output [15:0] col_out_347,
    output [15:0] col_out_348,
    output [15:0] col_out_349,
    output [15:0] col_out_350,
    output [15:0] col_out_351,
    output [15:0] col_out_352,
    output [15:0] col_out_353,
    output [15:0] col_out_354,
    output [15:0] col_out_355,
    output [15:0] col_out_356,
    output [15:0] col_out_357,
    output [15:0] col_out_358,
    output [15:0] col_out_359,
    output [15:0] col_out_360,
    output [15:0] col_out_361,
    output [15:0] col_out_362,
    output [15:0] col_out_363,
    output [15:0] col_out_364,
    output [15:0] col_out_365,
    output [15:0] col_out_366,
    output [15:0] col_out_367,
    output [15:0] col_out_368,
    output [15:0] col_out_369,
    output [15:0] col_out_370,
    output [15:0] col_out_371,
    output [15:0] col_out_372,
    output [15:0] col_out_373,
    output [15:0] col_out_374,
    output [15:0] col_out_375,
    output [15:0] col_out_376,
    output [15:0] col_out_377,
    output [15:0] col_out_378,
    output [15:0] col_out_379,
    output [15:0] col_out_380,
    output [15:0] col_out_381,
    output [15:0] col_out_382,
    output [15:0] col_out_383,
    output [15:0] col_out_384,
    output [15:0] col_out_385,
    output [15:0] col_out_386,
    output [15:0] col_out_387,
    output [15:0] col_out_388,
    output [15:0] col_out_389,
    output [15:0] col_out_390,
    output [15:0] col_out_391,
    output [15:0] col_out_392,
    output [15:0] col_out_393,
    output [15:0] col_out_394,
    output [15:0] col_out_395,
    output [15:0] col_out_396,
    output [15:0] col_out_397,
    output [15:0] col_out_398,
    output [15:0] col_out_399,
    output [15:0] col_out_400,
    output [15:0] col_out_401,
    output [15:0] col_out_402,
    output [15:0] col_out_403,
    output [15:0] col_out_404,
    output [15:0] col_out_405,
    output [15:0] col_out_406,
    output [15:0] col_out_407,
    output [15:0] col_out_408,
    output [15:0] col_out_409,
    output [15:0] col_out_410,
    output [15:0] col_out_411,
    output [15:0] col_out_412,
    output [15:0] col_out_413,
    output [15:0] col_out_414,
    output [15:0] col_out_415,
    output [15:0] col_out_416,
    output [15:0] col_out_417,
    output [15:0] col_out_418,
    output [15:0] col_out_419,
    output [15:0] col_out_420,
    output [15:0] col_out_421,
    output [15:0] col_out_422,
    output [15:0] col_out_423,
    output [15:0] col_out_424,
    output [15:0] col_out_425,
    output [15:0] col_out_426,
    output [15:0] col_out_427,
    output [15:0] col_out_428,
    output [15:0] col_out_429,
    output [15:0] col_out_430,
    output [15:0] col_out_431,
    output [15:0] col_out_432,
    output [15:0] col_out_433,
    output [15:0] col_out_434,
    output [15:0] col_out_435,
    output [15:0] col_out_436,
    output [15:0] col_out_437,
    output [15:0] col_out_438,
    output [15:0] col_out_439,
    output [15:0] col_out_440,
    output [15:0] col_out_441,
    output [15:0] col_out_442,
    output [15:0] col_out_443,
    output [15:0] col_out_444,
    output [15:0] col_out_445,
    output [15:0] col_out_446,
    output [15:0] col_out_447,
    output [15:0] col_out_448,
    output [15:0] col_out_449,
    output [15:0] col_out_450,
    output [15:0] col_out_451,
    output [15:0] col_out_452,
    output [15:0] col_out_453,
    output [15:0] col_out_454,
    output [15:0] col_out_455,
    output [15:0] col_out_456,
    output [15:0] col_out_457,
    output [15:0] col_out_458,
    output [15:0] col_out_459,
    output [15:0] col_out_460,
    output [15:0] col_out_461,
    output [15:0] col_out_462,
    output [15:0] col_out_463,
    output [15:0] col_out_464,
    output [15:0] col_out_465,
    output [15:0] col_out_466,
    output [15:0] col_out_467,
    output [15:0] col_out_468,
    output [15:0] col_out_469,
    output [15:0] col_out_470,
    output [15:0] col_out_471,
    output [15:0] col_out_472,
    output [15:0] col_out_473,
    output [15:0] col_out_474,
    output [15:0] col_out_475,
    output [15:0] col_out_476,
    output [15:0] col_out_477,
    output [15:0] col_out_478,
    output [15:0] col_out_479,
    output [15:0] col_out_480,
    output [15:0] col_out_481,
    output [15:0] col_out_482,
    output [15:0] col_out_483,
    output [15:0] col_out_484,
    output [15:0] col_out_485,
    output [15:0] col_out_486,
    output [15:0] col_out_487,
    output [15:0] col_out_488,
    output [15:0] col_out_489,
    output [15:0] col_out_490,
    output [15:0] col_out_491,
    output [15:0] col_out_492,
    output [15:0] col_out_493,
    output [15:0] col_out_494,
    output [15:0] col_out_495,
    output [15:0] col_out_496,
    output [15:0] col_out_497,
    output [15:0] col_out_498,
    output [15:0] col_out_499,
    output [15:0] col_out_500,
    output [15:0] col_out_501,
    output [15:0] col_out_502,
    output [15:0] col_out_503,
    output [15:0] col_out_504,
    output [15:0] col_out_505,
    output [15:0] col_out_506,
    output [15:0] col_out_507,
    output [15:0] col_out_508,
    output [15:0] col_out_509,
    output [15:0] col_out_510,
    output [15:0] col_out_511,
    output [15:0] col_out_512,
    output [15:0] col_out_513,
    output [15:0] col_out_514,
    output [15:0] col_out_515,
    output [15:0] col_out_516,
    output [15:0] col_out_517,
    output [15:0] col_out_518,
    output [15:0] col_out_519,
    output [15:0] col_out_520,
    output [15:0] col_out_521,
    output [15:0] col_out_522,
    output [15:0] col_out_523,
    output [15:0] col_out_524,
    output [15:0] col_out_525,
    output [15:0] col_out_526,
    output [15:0] col_out_527,
    output [15:0] col_out_528,
    output [15:0] col_out_529,
    output [15:0] col_out_530,
    output [15:0] col_out_531,
    output [15:0] col_out_532,
    output [15:0] col_out_533,
    output [15:0] col_out_534,
    output [15:0] col_out_535,
    output [15:0] col_out_536,
    output [15:0] col_out_537,
    output [15:0] col_out_538,
    output [15:0] col_out_539,
    output [15:0] col_out_540,
    output [15:0] col_out_541,
    output [15:0] col_out_542,
    output [15:0] col_out_543,
    output [15:0] col_out_544,
    output [15:0] col_out_545,
    output [15:0] col_out_546,
    output [15:0] col_out_547,
    output [15:0] col_out_548,
    output [15:0] col_out_549,
    output [15:0] col_out_550,
    output [15:0] col_out_551,
    output [15:0] col_out_552,
    output [15:0] col_out_553,
    output [15:0] col_out_554,
    output [15:0] col_out_555,
    output [15:0] col_out_556,
    output [15:0] col_out_557,
    output [15:0] col_out_558,
    output [15:0] col_out_559,
    output [15:0] col_out_560,
    output [15:0] col_out_561,
    output [15:0] col_out_562,
    output [15:0] col_out_563,
    output [15:0] col_out_564,
    output [15:0] col_out_565,
    output [15:0] col_out_566,
    output [15:0] col_out_567,
    output [15:0] col_out_568,
    output [15:0] col_out_569,
    output [15:0] col_out_570,
    output [15:0] col_out_571,
    output [15:0] col_out_572,
    output [15:0] col_out_573,
    output [15:0] col_out_574,
    output [15:0] col_out_575,
    output [15:0] col_out_576,
    output [15:0] col_out_577,
    output [15:0] col_out_578,
    output [15:0] col_out_579,
    output [15:0] col_out_580,
    output [15:0] col_out_581,
    output [15:0] col_out_582,
    output [15:0] col_out_583,
    output [15:0] col_out_584,
    output [15:0] col_out_585,
    output [15:0] col_out_586,
    output [15:0] col_out_587,
    output [15:0] col_out_588,
    output [15:0] col_out_589,
    output [15:0] col_out_590,
    output [15:0] col_out_591,
    output [15:0] col_out_592,
    output [15:0] col_out_593,
    output [15:0] col_out_594,
    output [15:0] col_out_595,
    output [15:0] col_out_596,
    output [15:0] col_out_597,
    output [15:0] col_out_598,
    output [15:0] col_out_599,
    output [15:0] col_out_600,
    output [15:0] col_out_601,
    output [15:0] col_out_602,
    output [15:0] col_out_603,
    output [15:0] col_out_604,
    output [15:0] col_out_605,
    output [15:0] col_out_606,
    output [15:0] col_out_607,
    output [15:0] col_out_608,
    output [15:0] col_out_609,
    output [15:0] col_out_610,
    output [15:0] col_out_611,
    output [15:0] col_out_612,
    output [15:0] col_out_613,
    output [15:0] col_out_614,
    output [15:0] col_out_615,
    output [15:0] col_out_616,
    output [15:0] col_out_617,
    output [15:0] col_out_618,
    output [15:0] col_out_619,
    output [15:0] col_out_620,
    output [15:0] col_out_621,
    output [15:0] col_out_622,
    output [15:0] col_out_623,
    output [15:0] col_out_624,
    output [15:0] col_out_625,
    output [15:0] col_out_626,
    output [15:0] col_out_627,
    output [15:0] col_out_628,
    output [15:0] col_out_629,
    output [15:0] col_out_630,
    output [15:0] col_out_631,
    output [15:0] col_out_632,
    output [15:0] col_out_633,
    output [15:0] col_out_634,
    output [15:0] col_out_635,
    output [15:0] col_out_636,
    output [15:0] col_out_637,
    output [15:0] col_out_638,
    output [15:0] col_out_639,
    output [15:0] col_out_640,
    output [15:0] col_out_641,
    output [15:0] col_out_642,
    output [15:0] col_out_643,
    output [15:0] col_out_644,
    output [15:0] col_out_645,
    output [15:0] col_out_646,
    output [15:0] col_out_647,
    output [15:0] col_out_648,
    output [15:0] col_out_649,
    output [15:0] col_out_650,
    output [15:0] col_out_651,
    output [15:0] col_out_652,
    output [15:0] col_out_653,
    output [15:0] col_out_654,
    output [15:0] col_out_655,
    output [15:0] col_out_656,
    output [15:0] col_out_657,
    output [15:0] col_out_658,
    output [15:0] col_out_659,
    output [15:0] col_out_660,
    output [15:0] col_out_661,
    output [15:0] col_out_662,
    output [15:0] col_out_663,
    output [15:0] col_out_664,
    output [15:0] col_out_665,
    output [15:0] col_out_666,
    output [15:0] col_out_667,
    output [15:0] col_out_668,
    output [15:0] col_out_669,
    output [15:0] col_out_670,
    output [15:0] col_out_671,
    output [15:0] col_out_672,
    output [15:0] col_out_673,
    output [15:0] col_out_674,
    output [15:0] col_out_675,
    output [15:0] col_out_676,
    output [15:0] col_out_677,
    output [15:0] col_out_678,
    output [15:0] col_out_679,
    output [15:0] col_out_680,
    output [15:0] col_out_681,
    output [15:0] col_out_682,
    output [15:0] col_out_683,
    output [15:0] col_out_684,
    output [15:0] col_out_685,
    output [15:0] col_out_686,
    output [15:0] col_out_687,
    output [15:0] col_out_688,
    output [15:0] col_out_689,
    output [15:0] col_out_690,
    output [15:0] col_out_691,
    output [15:0] col_out_692,
    output [15:0] col_out_693,
    output [15:0] col_out_694,
    output [15:0] col_out_695,
    output [15:0] col_out_696,
    output [15:0] col_out_697,
    output [15:0] col_out_698,
    output [15:0] col_out_699,
    output [15:0] col_out_700,
    output [15:0] col_out_701,
    output [15:0] col_out_702,
    output [15:0] col_out_703,
    output [15:0] col_out_704,
    output [15:0] col_out_705,
    output [15:0] col_out_706,
    output [15:0] col_out_707,
    output [15:0] col_out_708,
    output [15:0] col_out_709,
    output [15:0] col_out_710,
    output [15:0] col_out_711,
    output [15:0] col_out_712,
    output [15:0] col_out_713,
    output [15:0] col_out_714,
    output [15:0] col_out_715,
    output [15:0] col_out_716,
    output [15:0] col_out_717,
    output [15:0] col_out_718,
    output [15:0] col_out_719,
    output [15:0] col_out_720,
    output [15:0] col_out_721,
    output [15:0] col_out_722,
    output [15:0] col_out_723,
    output [15:0] col_out_724,
    output [15:0] col_out_725,
    output [15:0] col_out_726,
    output [15:0] col_out_727,
    output [15:0] col_out_728,
    output [15:0] col_out_729,
    output [15:0] col_out_730,
    output [15:0] col_out_731,
    output [15:0] col_out_732,
    output [15:0] col_out_733,
    output [15:0] col_out_734,
    output [15:0] col_out_735,
    output [15:0] col_out_736,
    output [15:0] col_out_737,
    output [15:0] col_out_738,
    output [15:0] col_out_739,
    output [15:0] col_out_740,
    output [15:0] col_out_741,
    output [15:0] col_out_742,
    output [15:0] col_out_743,
    output [15:0] col_out_744,
    output [15:0] col_out_745,
    output [15:0] col_out_746,
    output [15:0] col_out_747,
    output [15:0] col_out_748,
    output [15:0] col_out_749,
    output [15:0] col_out_750,
    output [15:0] col_out_751,
    output [15:0] col_out_752,
    output [15:0] col_out_753,
    output [15:0] col_out_754,
    output [15:0] col_out_755,
    output [15:0] col_out_756,
    output [15:0] col_out_757,
    output [15:0] col_out_758,
    output [15:0] col_out_759,
    output [15:0] col_out_760,
    output [15:0] col_out_761,
    output [15:0] col_out_762,
    output [15:0] col_out_763,
    output [15:0] col_out_764,
    output [15:0] col_out_765,
    output [15:0] col_out_766,
    output [15:0] col_out_767,
    output [15:0] col_out_768,
    output [15:0] col_out_769,
    output [15:0] col_out_770,
    output [15:0] col_out_771,
    output [15:0] col_out_772,
    output [15:0] col_out_773,
    output [15:0] col_out_774,
    output [15:0] col_out_775,
    output [15:0] col_out_776,
    output [15:0] col_out_777,
    output [15:0] col_out_778,
    output [15:0] col_out_779,
    output [15:0] col_out_780,
    output [15:0] col_out_781,
    output [15:0] col_out_782,
    output [15:0] col_out_783,
    output [15:0] col_out_784,
    output [15:0] col_out_785,
    output [15:0] col_out_786,
    output [15:0] col_out_787,
    output [15:0] col_out_788,
    output [15:0] col_out_789,
    output [15:0] col_out_790,
    output [15:0] col_out_791,
    output [15:0] col_out_792,
    output [15:0] col_out_793,
    output [15:0] col_out_794,
    output [15:0] col_out_795,
    output [15:0] col_out_796,
    output [15:0] col_out_797,
    output [15:0] col_out_798,
    output [15:0] col_out_799,
    output [15:0] col_out_800,
    output [15:0] col_out_801,
    output [15:0] col_out_802,
    output [15:0] col_out_803,
    output [15:0] col_out_804,
    output [15:0] col_out_805,
    output [15:0] col_out_806,
    output [15:0] col_out_807,
    output [15:0] col_out_808,
    output [15:0] col_out_809,
    output [15:0] col_out_810,
    output [15:0] col_out_811,
    output [15:0] col_out_812,
    output [15:0] col_out_813,
    output [15:0] col_out_814,
    output [15:0] col_out_815,
    output [15:0] col_out_816,
    output [15:0] col_out_817,
    output [15:0] col_out_818,
    output [15:0] col_out_819,
    output [15:0] col_out_820,
    output [15:0] col_out_821,
    output [15:0] col_out_822,
    output [15:0] col_out_823,
    output [15:0] col_out_824,
    output [15:0] col_out_825,
    output [15:0] col_out_826,
    output [15:0] col_out_827,
    output [15:0] col_out_828,
    output [15:0] col_out_829,
    output [15:0] col_out_830,
    output [15:0] col_out_831,
    output [15:0] col_out_832,
    output [15:0] col_out_833,
    output [15:0] col_out_834,
    output [15:0] col_out_835,
    output [15:0] col_out_836,
    output [15:0] col_out_837,
    output [15:0] col_out_838,
    output [15:0] col_out_839,
    output [15:0] col_out_840,
    output [15:0] col_out_841,
    output [15:0] col_out_842,
    output [15:0] col_out_843,
    output [15:0] col_out_844,
    output [15:0] col_out_845,
    output [15:0] col_out_846,
    output [15:0] col_out_847,
    output [15:0] col_out_848,
    output [15:0] col_out_849,
    output [15:0] col_out_850,
    output [15:0] col_out_851,
    output [15:0] col_out_852,
    output [15:0] col_out_853,
    output [15:0] col_out_854,
    output [15:0] col_out_855,
    output [15:0] col_out_856,
    output [15:0] col_out_857,
    output [15:0] col_out_858,
    output [15:0] col_out_859,
    output [15:0] col_out_860,
    output [15:0] col_out_861,
    output [15:0] col_out_862,
    output [15:0] col_out_863,
    output [15:0] col_out_864,
    output [15:0] col_out_865,
    output [15:0] col_out_866,
    output [15:0] col_out_867,
    output [15:0] col_out_868,
    output [15:0] col_out_869,
    output [15:0] col_out_870,
    output [15:0] col_out_871,
    output [15:0] col_out_872,
    output [15:0] col_out_873,
    output [15:0] col_out_874,
    output [15:0] col_out_875,
    output [15:0] col_out_876,
    output [15:0] col_out_877,
    output [15:0] col_out_878,
    output [15:0] col_out_879,
    output [15:0] col_out_880,
    output [15:0] col_out_881,
    output [15:0] col_out_882,
    output [15:0] col_out_883,
    output [15:0] col_out_884,
    output [15:0] col_out_885,
    output [15:0] col_out_886,
    output [15:0] col_out_887,
    output [15:0] col_out_888,
    output [15:0] col_out_889,
    output [15:0] col_out_890,
    output [15:0] col_out_891,
    output [15:0] col_out_892,
    output [15:0] col_out_893,
    output [15:0] col_out_894,
    output [15:0] col_out_895,
    output [15:0] col_out_896,
    output [15:0] col_out_897,
    output [15:0] col_out_898,
    output [15:0] col_out_899,
    output [15:0] col_out_900,
    output [15:0] col_out_901,
    output [15:0] col_out_902,
    output [15:0] col_out_903,
    output [15:0] col_out_904,
    output [15:0] col_out_905,
    output [15:0] col_out_906,
    output [15:0] col_out_907,
    output [15:0] col_out_908,
    output [15:0] col_out_909,
    output [15:0] col_out_910,
    output [15:0] col_out_911,
    output [15:0] col_out_912,
    output [15:0] col_out_913,
    output [15:0] col_out_914,
    output [15:0] col_out_915,
    output [15:0] col_out_916,
    output [15:0] col_out_917,
    output [15:0] col_out_918,
    output [15:0] col_out_919,
    output [15:0] col_out_920,
    output [15:0] col_out_921,
    output [15:0] col_out_922,
    output [15:0] col_out_923,
    output [15:0] col_out_924,
    output [15:0] col_out_925,
    output [15:0] col_out_926,
    output [15:0] col_out_927,
    output [15:0] col_out_928,
    output [15:0] col_out_929,
    output [15:0] col_out_930,
    output [15:0] col_out_931,
    output [15:0] col_out_932,
    output [15:0] col_out_933,
    output [15:0] col_out_934,
    output [15:0] col_out_935,
    output [15:0] col_out_936,
    output [15:0] col_out_937,
    output [15:0] col_out_938,
    output [15:0] col_out_939,
    output [15:0] col_out_940,
    output [15:0] col_out_941,
    output [15:0] col_out_942,
    output [15:0] col_out_943,
    output [15:0] col_out_944,
    output [15:0] col_out_945,
    output [15:0] col_out_946,
    output [15:0] col_out_947,
    output [15:0] col_out_948,
    output [15:0] col_out_949,
    output [15:0] col_out_950,
    output [15:0] col_out_951,
    output [15:0] col_out_952,
    output [15:0] col_out_953,
    output [15:0] col_out_954,
    output [15:0] col_out_955,
    output [15:0] col_out_956,
    output [15:0] col_out_957,
    output [15:0] col_out_958,
    output [15:0] col_out_959,
    output [15:0] col_out_960,
    output [15:0] col_out_961,
    output [15:0] col_out_962,
    output [15:0] col_out_963,
    output [15:0] col_out_964,
    output [15:0] col_out_965,
    output [15:0] col_out_966,
    output [15:0] col_out_967,
    output [15:0] col_out_968,
    output [15:0] col_out_969,
    output [15:0] col_out_970,
    output [15:0] col_out_971,
    output [15:0] col_out_972,
    output [15:0] col_out_973,
    output [15:0] col_out_974,
    output [15:0] col_out_975,
    output [15:0] col_out_976,
    output [15:0] col_out_977,
    output [15:0] col_out_978,
    output [15:0] col_out_979,
    output [15:0] col_out_980,
    output [15:0] col_out_981,
    output [15:0] col_out_982,
    output [15:0] col_out_983,
    output [15:0] col_out_984,
    output [15:0] col_out_985,
    output [15:0] col_out_986,
    output [15:0] col_out_987,
    output [15:0] col_out_988,
    output [15:0] col_out_989,
    output [15:0] col_out_990,
    output [15:0] col_out_991,
    output [15:0] col_out_992,
    output [15:0] col_out_993,
    output [15:0] col_out_994,
    output [15:0] col_out_995,
    output [15:0] col_out_996,
    output [15:0] col_out_997,
    output [15:0] col_out_998,
    output [15:0] col_out_999,
    output [15:0] col_out_1000,
    output [15:0] col_out_1001,
    output [15:0] col_out_1002,
    output [15:0] col_out_1003,
    output [15:0] col_out_1004,
    output [15:0] col_out_1005,
    output [15:0] col_out_1006,
    output [15:0] col_out_1007,
    output [15:0] col_out_1008,
    output [15:0] col_out_1009,
    output [15:0] col_out_1010,
    output [15:0] col_out_1011,
    output [15:0] col_out_1012,
    output [15:0] col_out_1013,
    output [15:0] col_out_1014,
    output [15:0] col_out_1015,
    output [15:0] col_out_1016,
    output [15:0] col_out_1017,
    output [15:0] col_out_1018,
    output [15:0] col_out_1019,
    output [15:0] col_out_1020,
    output [15:0] col_out_1021,
    output [15:0] col_out_1022,
    output [15:0] col_out_1023,
    output [15:0] col_out_1024,
    output [15:0] col_out_1025,
    output [15:0] col_out_1026,
    output [15:0] col_out_1027,
    output [15:0] col_out_1028,
    output [15:0] col_out_1029,
    output [15:0] col_out_1030,
    output [15:0] col_out_1031,
    output [15:0] col_out_1032


);


//*****************************************************
//**************u0输入定义******************************
//*****************************************************
wire [511:0] u0_col_in_0;
wire [511:0] u0_col_in_1;
wire [511:0] u0_col_in_2;
wire [511:0] u0_col_in_3;
wire [511:0] u0_col_in_4;
wire [511:0] u0_col_in_5;
wire [511:0] u0_col_in_6;
wire [511:0] u0_col_in_7;
wire [511:0] u0_col_in_8;
wire [511:0] u0_col_in_9;
wire [511:0] u0_col_in_10;
wire [511:0] u0_col_in_11;
wire [511:0] u0_col_in_12;
wire [511:0] u0_col_in_13;
wire [511:0] u0_col_in_14;
wire [511:0] u0_col_in_15;
wire [511:0] u0_col_in_16;
wire [511:0] u0_col_in_17;
wire [511:0] u0_col_in_18;
wire [511:0] u0_col_in_19;
wire [511:0] u0_col_in_20;
wire [511:0] u0_col_in_21;
wire [511:0] u0_col_in_22;
wire [511:0] u0_col_in_23;
wire [511:0] u0_col_in_24;
wire [511:0] u0_col_in_25;
wire [511:0] u0_col_in_26;
wire [511:0] u0_col_in_27;
wire [511:0] u0_col_in_28;
wire [511:0] u0_col_in_29;
wire [511:0] u0_col_in_30;
wire [511:0] u0_col_in_31;
wire [511:0] u0_col_in_32;
wire [511:0] u0_col_in_33;
wire [511:0] u0_col_in_34;
wire [511:0] u0_col_in_35;
wire [511:0] u0_col_in_36;
wire [511:0] u0_col_in_37;
wire [511:0] u0_col_in_38;
wire [511:0] u0_col_in_39;
wire [511:0] u0_col_in_40;
wire [511:0] u0_col_in_41;
wire [511:0] u0_col_in_42;
wire [511:0] u0_col_in_43;
wire [511:0] u0_col_in_44;
wire [511:0] u0_col_in_45;
wire [511:0] u0_col_in_46;
wire [511:0] u0_col_in_47;
wire [511:0] u0_col_in_48;
wire [511:0] u0_col_in_49;
wire [511:0] u0_col_in_50;
wire [511:0] u0_col_in_51;
wire [511:0] u0_col_in_52;
wire [511:0] u0_col_in_53;
wire [511:0] u0_col_in_54;
wire [511:0] u0_col_in_55;
wire [511:0] u0_col_in_56;
wire [511:0] u0_col_in_57;
wire [511:0] u0_col_in_58;
wire [511:0] u0_col_in_59;
wire [511:0] u0_col_in_60;
wire [511:0] u0_col_in_61;
wire [511:0] u0_col_in_62;
wire [511:0] u0_col_in_63;
wire [511:0] u0_col_in_64;
wire [511:0] u0_col_in_65;
wire [511:0] u0_col_in_66;
wire [511:0] u0_col_in_67;
wire [511:0] u0_col_in_68;
wire [511:0] u0_col_in_69;
wire [511:0] u0_col_in_70;
wire [511:0] u0_col_in_71;
wire [511:0] u0_col_in_72;
wire [511:0] u0_col_in_73;
wire [511:0] u0_col_in_74;
wire [511:0] u0_col_in_75;
wire [511:0] u0_col_in_76;
wire [511:0] u0_col_in_77;
wire [511:0] u0_col_in_78;
wire [511:0] u0_col_in_79;
wire [511:0] u0_col_in_80;
wire [511:0] u0_col_in_81;
wire [511:0] u0_col_in_82;
wire [511:0] u0_col_in_83;
wire [511:0] u0_col_in_84;
wire [511:0] u0_col_in_85;
wire [511:0] u0_col_in_86;
wire [511:0] u0_col_in_87;
wire [511:0] u0_col_in_88;
wire [511:0] u0_col_in_89;
wire [511:0] u0_col_in_90;
wire [511:0] u0_col_in_91;
wire [511:0] u0_col_in_92;
wire [511:0] u0_col_in_93;
wire [511:0] u0_col_in_94;
wire [511:0] u0_col_in_95;
wire [511:0] u0_col_in_96;
wire [511:0] u0_col_in_97;
wire [511:0] u0_col_in_98;
wire [511:0] u0_col_in_99;
wire [511:0] u0_col_in_100;
wire [511:0] u0_col_in_101;
wire [511:0] u0_col_in_102;
wire [511:0] u0_col_in_103;
wire [511:0] u0_col_in_104;
wire [511:0] u0_col_in_105;
wire [511:0] u0_col_in_106;
wire [511:0] u0_col_in_107;
wire [511:0] u0_col_in_108;
wire [511:0] u0_col_in_109;
wire [511:0] u0_col_in_110;
wire [511:0] u0_col_in_111;
wire [511:0] u0_col_in_112;
wire [511:0] u0_col_in_113;
wire [511:0] u0_col_in_114;
wire [511:0] u0_col_in_115;
wire [511:0] u0_col_in_116;
wire [511:0] u0_col_in_117;
wire [511:0] u0_col_in_118;
wire [511:0] u0_col_in_119;
wire [511:0] u0_col_in_120;
wire [511:0] u0_col_in_121;
wire [511:0] u0_col_in_122;
wire [511:0] u0_col_in_123;
wire [511:0] u0_col_in_124;
wire [511:0] u0_col_in_125;
wire [511:0] u0_col_in_126;
wire [511:0] u0_col_in_127;
wire [511:0] u0_col_in_128;
wire [511:0] u0_col_in_129;
wire [511:0] u0_col_in_130;
wire [511:0] u0_col_in_131;
wire [511:0] u0_col_in_132;
wire [511:0] u0_col_in_133;
wire [511:0] u0_col_in_134;
wire [511:0] u0_col_in_135;
wire [511:0] u0_col_in_136;
wire [511:0] u0_col_in_137;
wire [511:0] u0_col_in_138;
wire [511:0] u0_col_in_139;
wire [511:0] u0_col_in_140;
wire [511:0] u0_col_in_141;
wire [511:0] u0_col_in_142;
wire [511:0] u0_col_in_143;
wire [511:0] u0_col_in_144;
wire [511:0] u0_col_in_145;
wire [511:0] u0_col_in_146;
wire [511:0] u0_col_in_147;
wire [511:0] u0_col_in_148;
wire [511:0] u0_col_in_149;
wire [511:0] u0_col_in_150;
wire [511:0] u0_col_in_151;
wire [511:0] u0_col_in_152;
wire [511:0] u0_col_in_153;
wire [511:0] u0_col_in_154;
wire [511:0] u0_col_in_155;
wire [511:0] u0_col_in_156;
wire [511:0] u0_col_in_157;
wire [511:0] u0_col_in_158;
wire [511:0] u0_col_in_159;
wire [511:0] u0_col_in_160;
wire [511:0] u0_col_in_161;
wire [511:0] u0_col_in_162;
wire [511:0] u0_col_in_163;
wire [511:0] u0_col_in_164;
wire [511:0] u0_col_in_165;
wire [511:0] u0_col_in_166;
wire [511:0] u0_col_in_167;
wire [511:0] u0_col_in_168;
wire [511:0] u0_col_in_169;
wire [511:0] u0_col_in_170;
wire [511:0] u0_col_in_171;
wire [511:0] u0_col_in_172;
wire [511:0] u0_col_in_173;
wire [511:0] u0_col_in_174;
wire [511:0] u0_col_in_175;
wire [511:0] u0_col_in_176;
wire [511:0] u0_col_in_177;
wire [511:0] u0_col_in_178;
wire [511:0] u0_col_in_179;
wire [511:0] u0_col_in_180;
wire [511:0] u0_col_in_181;
wire [511:0] u0_col_in_182;
wire [511:0] u0_col_in_183;
wire [511:0] u0_col_in_184;
wire [511:0] u0_col_in_185;
wire [511:0] u0_col_in_186;
wire [511:0] u0_col_in_187;
wire [511:0] u0_col_in_188;
wire [511:0] u0_col_in_189;
wire [511:0] u0_col_in_190;
wire [511:0] u0_col_in_191;
wire [511:0] u0_col_in_192;
wire [511:0] u0_col_in_193;
wire [511:0] u0_col_in_194;
wire [511:0] u0_col_in_195;
wire [511:0] u0_col_in_196;
wire [511:0] u0_col_in_197;
wire [511:0] u0_col_in_198;
wire [511:0] u0_col_in_199;
wire [511:0] u0_col_in_200;
wire [511:0] u0_col_in_201;
wire [511:0] u0_col_in_202;
wire [511:0] u0_col_in_203;
wire [511:0] u0_col_in_204;
wire [511:0] u0_col_in_205;
wire [511:0] u0_col_in_206;
wire [511:0] u0_col_in_207;
wire [511:0] u0_col_in_208;
wire [511:0] u0_col_in_209;
wire [511:0] u0_col_in_210;
wire [511:0] u0_col_in_211;
wire [511:0] u0_col_in_212;
wire [511:0] u0_col_in_213;
wire [511:0] u0_col_in_214;
wire [511:0] u0_col_in_215;
wire [511:0] u0_col_in_216;
wire [511:0] u0_col_in_217;
wire [511:0] u0_col_in_218;
wire [511:0] u0_col_in_219;
wire [511:0] u0_col_in_220;
wire [511:0] u0_col_in_221;
wire [511:0] u0_col_in_222;
wire [511:0] u0_col_in_223;
wire [511:0] u0_col_in_224;
wire [511:0] u0_col_in_225;
wire [511:0] u0_col_in_226;
wire [511:0] u0_col_in_227;
wire [511:0] u0_col_in_228;
wire [511:0] u0_col_in_229;
wire [511:0] u0_col_in_230;
wire [511:0] u0_col_in_231;
wire [511:0] u0_col_in_232;
wire [511:0] u0_col_in_233;
wire [511:0] u0_col_in_234;
wire [511:0] u0_col_in_235;
wire [511:0] u0_col_in_236;
wire [511:0] u0_col_in_237;
wire [511:0] u0_col_in_238;
wire [511:0] u0_col_in_239;
wire [511:0] u0_col_in_240;
wire [511:0] u0_col_in_241;
wire [511:0] u0_col_in_242;
wire [511:0] u0_col_in_243;
wire [511:0] u0_col_in_244;
wire [511:0] u0_col_in_245;
wire [511:0] u0_col_in_246;
wire [511:0] u0_col_in_247;
wire [511:0] u0_col_in_248;
wire [511:0] u0_col_in_249;
wire [511:0] u0_col_in_250;
wire [511:0] u0_col_in_251;
wire [511:0] u0_col_in_252;
wire [511:0] u0_col_in_253;
wire [511:0] u0_col_in_254;
wire [511:0] u0_col_in_255;
wire [511:0] u0_col_in_256;
wire [511:0] u0_col_in_257;
wire [511:0] u0_col_in_258;
wire [511:0] u0_col_in_259;
wire [511:0] u0_col_in_260;
wire [511:0] u0_col_in_261;
wire [511:0] u0_col_in_262;
wire [511:0] u0_col_in_263;
wire [511:0] u0_col_in_264;
wire [511:0] u0_col_in_265;
wire [511:0] u0_col_in_266;
wire [511:0] u0_col_in_267;
wire [511:0] u0_col_in_268;
wire [511:0] u0_col_in_269;
wire [511:0] u0_col_in_270;
wire [511:0] u0_col_in_271;
wire [511:0] u0_col_in_272;
wire [511:0] u0_col_in_273;
wire [511:0] u0_col_in_274;
wire [511:0] u0_col_in_275;
wire [511:0] u0_col_in_276;
wire [511:0] u0_col_in_277;
wire [511:0] u0_col_in_278;
wire [511:0] u0_col_in_279;
wire [511:0] u0_col_in_280;
wire [511:0] u0_col_in_281;
wire [511:0] u0_col_in_282;
wire [511:0] u0_col_in_283;
wire [511:0] u0_col_in_284;
wire [511:0] u0_col_in_285;
wire [511:0] u0_col_in_286;
wire [511:0] u0_col_in_287;
wire [511:0] u0_col_in_288;
wire [511:0] u0_col_in_289;
wire [511:0] u0_col_in_290;
wire [511:0] u0_col_in_291;
wire [511:0] u0_col_in_292;
wire [511:0] u0_col_in_293;
wire [511:0] u0_col_in_294;
wire [511:0] u0_col_in_295;
wire [511:0] u0_col_in_296;
wire [511:0] u0_col_in_297;
wire [511:0] u0_col_in_298;
wire [511:0] u0_col_in_299;
wire [511:0] u0_col_in_300;
wire [511:0] u0_col_in_301;
wire [511:0] u0_col_in_302;
wire [511:0] u0_col_in_303;
wire [511:0] u0_col_in_304;
wire [511:0] u0_col_in_305;
wire [511:0] u0_col_in_306;
wire [511:0] u0_col_in_307;
wire [511:0] u0_col_in_308;
wire [511:0] u0_col_in_309;
wire [511:0] u0_col_in_310;
wire [511:0] u0_col_in_311;
wire [511:0] u0_col_in_312;
wire [511:0] u0_col_in_313;
wire [511:0] u0_col_in_314;
wire [511:0] u0_col_in_315;
wire [511:0] u0_col_in_316;
wire [511:0] u0_col_in_317;
wire [511:0] u0_col_in_318;
wire [511:0] u0_col_in_319;
wire [511:0] u0_col_in_320;
wire [511:0] u0_col_in_321;
wire [511:0] u0_col_in_322;
wire [511:0] u0_col_in_323;
wire [511:0] u0_col_in_324;
wire [511:0] u0_col_in_325;
wire [511:0] u0_col_in_326;
wire [511:0] u0_col_in_327;
wire [511:0] u0_col_in_328;
wire [511:0] u0_col_in_329;
wire [511:0] u0_col_in_330;
wire [511:0] u0_col_in_331;
wire [511:0] u0_col_in_332;
wire [511:0] u0_col_in_333;
wire [511:0] u0_col_in_334;
wire [511:0] u0_col_in_335;
wire [511:0] u0_col_in_336;
wire [511:0] u0_col_in_337;
wire [511:0] u0_col_in_338;
wire [511:0] u0_col_in_339;
wire [511:0] u0_col_in_340;
wire [511:0] u0_col_in_341;
wire [511:0] u0_col_in_342;
wire [511:0] u0_col_in_343;
wire [511:0] u0_col_in_344;
wire [511:0] u0_col_in_345;
wire [511:0] u0_col_in_346;
wire [511:0] u0_col_in_347;
wire [511:0] u0_col_in_348;
wire [511:0] u0_col_in_349;
wire [511:0] u0_col_in_350;
wire [511:0] u0_col_in_351;
wire [511:0] u0_col_in_352;
wire [511:0] u0_col_in_353;
wire [511:0] u0_col_in_354;
wire [511:0] u0_col_in_355;
wire [511:0] u0_col_in_356;
wire [511:0] u0_col_in_357;
wire [511:0] u0_col_in_358;
wire [511:0] u0_col_in_359;
wire [511:0] u0_col_in_360;
wire [511:0] u0_col_in_361;
wire [511:0] u0_col_in_362;
wire [511:0] u0_col_in_363;
wire [511:0] u0_col_in_364;
wire [511:0] u0_col_in_365;
wire [511:0] u0_col_in_366;
wire [511:0] u0_col_in_367;
wire [511:0] u0_col_in_368;
wire [511:0] u0_col_in_369;
wire [511:0] u0_col_in_370;
wire [511:0] u0_col_in_371;
wire [511:0] u0_col_in_372;
wire [511:0] u0_col_in_373;
wire [511:0] u0_col_in_374;
wire [511:0] u0_col_in_375;
wire [511:0] u0_col_in_376;
wire [511:0] u0_col_in_377;
wire [511:0] u0_col_in_378;
wire [511:0] u0_col_in_379;
wire [511:0] u0_col_in_380;
wire [511:0] u0_col_in_381;
wire [511:0] u0_col_in_382;
wire [511:0] u0_col_in_383;
wire [511:0] u0_col_in_384;
wire [511:0] u0_col_in_385;
wire [511:0] u0_col_in_386;
wire [511:0] u0_col_in_387;
wire [511:0] u0_col_in_388;
wire [511:0] u0_col_in_389;
wire [511:0] u0_col_in_390;
wire [511:0] u0_col_in_391;
wire [511:0] u0_col_in_392;
wire [511:0] u0_col_in_393;
wire [511:0] u0_col_in_394;
wire [511:0] u0_col_in_395;
wire [511:0] u0_col_in_396;
wire [511:0] u0_col_in_397;
wire [511:0] u0_col_in_398;
wire [511:0] u0_col_in_399;
wire [511:0] u0_col_in_400;
wire [511:0] u0_col_in_401;
wire [511:0] u0_col_in_402;
wire [511:0] u0_col_in_403;
wire [511:0] u0_col_in_404;
wire [511:0] u0_col_in_405;
wire [511:0] u0_col_in_406;
wire [511:0] u0_col_in_407;
wire [511:0] u0_col_in_408;
wire [511:0] u0_col_in_409;
wire [511:0] u0_col_in_410;
wire [511:0] u0_col_in_411;
wire [511:0] u0_col_in_412;
wire [511:0] u0_col_in_413;
wire [511:0] u0_col_in_414;
wire [511:0] u0_col_in_415;
wire [511:0] u0_col_in_416;
wire [511:0] u0_col_in_417;
wire [511:0] u0_col_in_418;
wire [511:0] u0_col_in_419;
wire [511:0] u0_col_in_420;
wire [511:0] u0_col_in_421;
wire [511:0] u0_col_in_422;
wire [511:0] u0_col_in_423;
wire [511:0] u0_col_in_424;
wire [511:0] u0_col_in_425;
wire [511:0] u0_col_in_426;
wire [511:0] u0_col_in_427;
wire [511:0] u0_col_in_428;
wire [511:0] u0_col_in_429;
wire [511:0] u0_col_in_430;
wire [511:0] u0_col_in_431;
wire [511:0] u0_col_in_432;
wire [511:0] u0_col_in_433;
wire [511:0] u0_col_in_434;
wire [511:0] u0_col_in_435;
wire [511:0] u0_col_in_436;
wire [511:0] u0_col_in_437;
wire [511:0] u0_col_in_438;
wire [511:0] u0_col_in_439;
wire [511:0] u0_col_in_440;
wire [511:0] u0_col_in_441;
wire [511:0] u0_col_in_442;
wire [511:0] u0_col_in_443;
wire [511:0] u0_col_in_444;
wire [511:0] u0_col_in_445;
wire [511:0] u0_col_in_446;
wire [511:0] u0_col_in_447;
wire [511:0] u0_col_in_448;
wire [511:0] u0_col_in_449;
wire [511:0] u0_col_in_450;
wire [511:0] u0_col_in_451;
wire [511:0] u0_col_in_452;
wire [511:0] u0_col_in_453;
wire [511:0] u0_col_in_454;
wire [511:0] u0_col_in_455;
wire [511:0] u0_col_in_456;
wire [511:0] u0_col_in_457;
wire [511:0] u0_col_in_458;
wire [511:0] u0_col_in_459;
wire [511:0] u0_col_in_460;
wire [511:0] u0_col_in_461;
wire [511:0] u0_col_in_462;
wire [511:0] u0_col_in_463;
wire [511:0] u0_col_in_464;
wire [511:0] u0_col_in_465;
wire [511:0] u0_col_in_466;
wire [511:0] u0_col_in_467;
wire [511:0] u0_col_in_468;
wire [511:0] u0_col_in_469;
wire [511:0] u0_col_in_470;
wire [511:0] u0_col_in_471;
wire [511:0] u0_col_in_472;
wire [511:0] u0_col_in_473;
wire [511:0] u0_col_in_474;
wire [511:0] u0_col_in_475;
wire [511:0] u0_col_in_476;
wire [511:0] u0_col_in_477;
wire [511:0] u0_col_in_478;
wire [511:0] u0_col_in_479;
wire [511:0] u0_col_in_480;
wire [511:0] u0_col_in_481;
wire [511:0] u0_col_in_482;
wire [511:0] u0_col_in_483;
wire [511:0] u0_col_in_484;
wire [511:0] u0_col_in_485;
wire [511:0] u0_col_in_486;
wire [511:0] u0_col_in_487;
wire [511:0] u0_col_in_488;
wire [511:0] u0_col_in_489;
wire [511:0] u0_col_in_490;
wire [511:0] u0_col_in_491;
wire [511:0] u0_col_in_492;
wire [511:0] u0_col_in_493;
wire [511:0] u0_col_in_494;
wire [511:0] u0_col_in_495;
wire [511:0] u0_col_in_496;
wire [511:0] u0_col_in_497;
wire [511:0] u0_col_in_498;
wire [511:0] u0_col_in_499;
wire [511:0] u0_col_in_500;
wire [511:0] u0_col_in_501;
wire [511:0] u0_col_in_502;
wire [511:0] u0_col_in_503;
wire [511:0] u0_col_in_504;
wire [511:0] u0_col_in_505;
wire [511:0] u0_col_in_506;
wire [511:0] u0_col_in_507;
wire [511:0] u0_col_in_508;
wire [511:0] u0_col_in_509;
wire [511:0] u0_col_in_510;
wire [511:0] u0_col_in_511;
wire [511:0] u0_col_in_512;
wire [511:0] u0_col_in_513;
wire [511:0] u0_col_in_514;
wire [511:0] u0_col_in_515;
wire [511:0] u0_col_in_516;
wire [511:0] u0_col_in_517;
wire [511:0] u0_col_in_518;
wire [511:0] u0_col_in_519;
wire [511:0] u0_col_in_520;
wire [511:0] u0_col_in_521;
wire [511:0] u0_col_in_522;
wire [511:0] u0_col_in_523;
wire [511:0] u0_col_in_524;
wire [511:0] u0_col_in_525;
wire [511:0] u0_col_in_526;
wire [511:0] u0_col_in_527;
wire [511:0] u0_col_in_528;
wire [511:0] u0_col_in_529;
wire [511:0] u0_col_in_530;
wire [511:0] u0_col_in_531;
wire [511:0] u0_col_in_532;
wire [511:0] u0_col_in_533;
wire [511:0] u0_col_in_534;
wire [511:0] u0_col_in_535;
wire [511:0] u0_col_in_536;
wire [511:0] u0_col_in_537;
wire [511:0] u0_col_in_538;
wire [511:0] u0_col_in_539;
wire [511:0] u0_col_in_540;
wire [511:0] u0_col_in_541;
wire [511:0] u0_col_in_542;
wire [511:0] u0_col_in_543;
wire [511:0] u0_col_in_544;
wire [511:0] u0_col_in_545;
wire [511:0] u0_col_in_546;
wire [511:0] u0_col_in_547;
wire [511:0] u0_col_in_548;
wire [511:0] u0_col_in_549;
wire [511:0] u0_col_in_550;
wire [511:0] u0_col_in_551;
wire [511:0] u0_col_in_552;
wire [511:0] u0_col_in_553;
wire [511:0] u0_col_in_554;
wire [511:0] u0_col_in_555;
wire [511:0] u0_col_in_556;
wire [511:0] u0_col_in_557;
wire [511:0] u0_col_in_558;
wire [511:0] u0_col_in_559;
wire [511:0] u0_col_in_560;
wire [511:0] u0_col_in_561;
wire [511:0] u0_col_in_562;
wire [511:0] u0_col_in_563;
wire [511:0] u0_col_in_564;
wire [511:0] u0_col_in_565;
wire [511:0] u0_col_in_566;
wire [511:0] u0_col_in_567;
wire [511:0] u0_col_in_568;
wire [511:0] u0_col_in_569;
wire [511:0] u0_col_in_570;
wire [511:0] u0_col_in_571;
wire [511:0] u0_col_in_572;
wire [511:0] u0_col_in_573;
wire [511:0] u0_col_in_574;
wire [511:0] u0_col_in_575;
wire [511:0] u0_col_in_576;
wire [511:0] u0_col_in_577;
wire [511:0] u0_col_in_578;
wire [511:0] u0_col_in_579;
wire [511:0] u0_col_in_580;
wire [511:0] u0_col_in_581;
wire [511:0] u0_col_in_582;
wire [511:0] u0_col_in_583;
wire [511:0] u0_col_in_584;
wire [511:0] u0_col_in_585;
wire [511:0] u0_col_in_586;
wire [511:0] u0_col_in_587;
wire [511:0] u0_col_in_588;
wire [511:0] u0_col_in_589;
wire [511:0] u0_col_in_590;
wire [511:0] u0_col_in_591;
wire [511:0] u0_col_in_592;
wire [511:0] u0_col_in_593;
wire [511:0] u0_col_in_594;
wire [511:0] u0_col_in_595;
wire [511:0] u0_col_in_596;
wire [511:0] u0_col_in_597;
wire [511:0] u0_col_in_598;
wire [511:0] u0_col_in_599;
wire [511:0] u0_col_in_600;
wire [511:0] u0_col_in_601;
wire [511:0] u0_col_in_602;
wire [511:0] u0_col_in_603;
wire [511:0] u0_col_in_604;
wire [511:0] u0_col_in_605;
wire [511:0] u0_col_in_606;
wire [511:0] u0_col_in_607;
wire [511:0] u0_col_in_608;
wire [511:0] u0_col_in_609;
wire [511:0] u0_col_in_610;
wire [511:0] u0_col_in_611;
wire [511:0] u0_col_in_612;
wire [511:0] u0_col_in_613;
wire [511:0] u0_col_in_614;
wire [511:0] u0_col_in_615;
wire [511:0] u0_col_in_616;
wire [511:0] u0_col_in_617;
wire [511:0] u0_col_in_618;
wire [511:0] u0_col_in_619;
wire [511:0] u0_col_in_620;
wire [511:0] u0_col_in_621;
wire [511:0] u0_col_in_622;
wire [511:0] u0_col_in_623;
wire [511:0] u0_col_in_624;
wire [511:0] u0_col_in_625;
wire [511:0] u0_col_in_626;
wire [511:0] u0_col_in_627;
wire [511:0] u0_col_in_628;
wire [511:0] u0_col_in_629;
wire [511:0] u0_col_in_630;
wire [511:0] u0_col_in_631;
wire [511:0] u0_col_in_632;
wire [511:0] u0_col_in_633;
wire [511:0] u0_col_in_634;
wire [511:0] u0_col_in_635;
wire [511:0] u0_col_in_636;
wire [511:0] u0_col_in_637;
wire [511:0] u0_col_in_638;
wire [511:0] u0_col_in_639;
wire [511:0] u0_col_in_640;
wire [511:0] u0_col_in_641;
wire [511:0] u0_col_in_642;
wire [511:0] u0_col_in_643;
wire [511:0] u0_col_in_644;
wire [511:0] u0_col_in_645;
wire [511:0] u0_col_in_646;
wire [511:0] u0_col_in_647;
wire [511:0] u0_col_in_648;
wire [511:0] u0_col_in_649;
wire [511:0] u0_col_in_650;
wire [511:0] u0_col_in_651;
wire [511:0] u0_col_in_652;
wire [511:0] u0_col_in_653;
wire [511:0] u0_col_in_654;
wire [511:0] u0_col_in_655;
wire [511:0] u0_col_in_656;
wire [511:0] u0_col_in_657;
wire [511:0] u0_col_in_658;
wire [511:0] u0_col_in_659;
wire [511:0] u0_col_in_660;
wire [511:0] u0_col_in_661;
wire [511:0] u0_col_in_662;
wire [511:0] u0_col_in_663;
wire [511:0] u0_col_in_664;
wire [511:0] u0_col_in_665;
wire [511:0] u0_col_in_666;
wire [511:0] u0_col_in_667;
wire [511:0] u0_col_in_668;
wire [511:0] u0_col_in_669;
wire [511:0] u0_col_in_670;
wire [511:0] u0_col_in_671;
wire [511:0] u0_col_in_672;
wire [511:0] u0_col_in_673;
wire [511:0] u0_col_in_674;
wire [511:0] u0_col_in_675;
wire [511:0] u0_col_in_676;
wire [511:0] u0_col_in_677;
wire [511:0] u0_col_in_678;
wire [511:0] u0_col_in_679;
wire [511:0] u0_col_in_680;
wire [511:0] u0_col_in_681;
wire [511:0] u0_col_in_682;
wire [511:0] u0_col_in_683;
wire [511:0] u0_col_in_684;
wire [511:0] u0_col_in_685;
wire [511:0] u0_col_in_686;
wire [511:0] u0_col_in_687;
wire [511:0] u0_col_in_688;
wire [511:0] u0_col_in_689;
wire [511:0] u0_col_in_690;
wire [511:0] u0_col_in_691;
wire [511:0] u0_col_in_692;
wire [511:0] u0_col_in_693;
wire [511:0] u0_col_in_694;
wire [511:0] u0_col_in_695;
wire [511:0] u0_col_in_696;
wire [511:0] u0_col_in_697;
wire [511:0] u0_col_in_698;
wire [511:0] u0_col_in_699;
wire [511:0] u0_col_in_700;
wire [511:0] u0_col_in_701;
wire [511:0] u0_col_in_702;
wire [511:0] u0_col_in_703;
wire [511:0] u0_col_in_704;
wire [511:0] u0_col_in_705;
wire [511:0] u0_col_in_706;
wire [511:0] u0_col_in_707;
wire [511:0] u0_col_in_708;
wire [511:0] u0_col_in_709;
wire [511:0] u0_col_in_710;
wire [511:0] u0_col_in_711;
wire [511:0] u0_col_in_712;
wire [511:0] u0_col_in_713;
wire [511:0] u0_col_in_714;
wire [511:0] u0_col_in_715;
wire [511:0] u0_col_in_716;
wire [511:0] u0_col_in_717;
wire [511:0] u0_col_in_718;
wire [511:0] u0_col_in_719;
wire [511:0] u0_col_in_720;
wire [511:0] u0_col_in_721;
wire [511:0] u0_col_in_722;
wire [511:0] u0_col_in_723;
wire [511:0] u0_col_in_724;
wire [511:0] u0_col_in_725;
wire [511:0] u0_col_in_726;
wire [511:0] u0_col_in_727;
wire [511:0] u0_col_in_728;
wire [511:0] u0_col_in_729;
wire [511:0] u0_col_in_730;
wire [511:0] u0_col_in_731;
wire [511:0] u0_col_in_732;
wire [511:0] u0_col_in_733;
wire [511:0] u0_col_in_734;
wire [511:0] u0_col_in_735;
wire [511:0] u0_col_in_736;
wire [511:0] u0_col_in_737;
wire [511:0] u0_col_in_738;
wire [511:0] u0_col_in_739;
wire [511:0] u0_col_in_740;
wire [511:0] u0_col_in_741;
wire [511:0] u0_col_in_742;
wire [511:0] u0_col_in_743;
wire [511:0] u0_col_in_744;
wire [511:0] u0_col_in_745;
wire [511:0] u0_col_in_746;
wire [511:0] u0_col_in_747;
wire [511:0] u0_col_in_748;
wire [511:0] u0_col_in_749;
wire [511:0] u0_col_in_750;
wire [511:0] u0_col_in_751;
wire [511:0] u0_col_in_752;
wire [511:0] u0_col_in_753;
wire [511:0] u0_col_in_754;
wire [511:0] u0_col_in_755;
wire [511:0] u0_col_in_756;
wire [511:0] u0_col_in_757;
wire [511:0] u0_col_in_758;
wire [511:0] u0_col_in_759;
wire [511:0] u0_col_in_760;
wire [511:0] u0_col_in_761;
wire [511:0] u0_col_in_762;
wire [511:0] u0_col_in_763;
wire [511:0] u0_col_in_764;
wire [511:0] u0_col_in_765;
wire [511:0] u0_col_in_766;
wire [511:0] u0_col_in_767;
wire [511:0] u0_col_in_768;
wire [511:0] u0_col_in_769;
wire [511:0] u0_col_in_770;
wire [511:0] u0_col_in_771;
wire [511:0] u0_col_in_772;
wire [511:0] u0_col_in_773;
wire [511:0] u0_col_in_774;
wire [511:0] u0_col_in_775;
wire [511:0] u0_col_in_776;
wire [511:0] u0_col_in_777;
wire [511:0] u0_col_in_778;
wire [511:0] u0_col_in_779;
wire [511:0] u0_col_in_780;
wire [511:0] u0_col_in_781;
wire [511:0] u0_col_in_782;
wire [511:0] u0_col_in_783;
wire [511:0] u0_col_in_784;
wire [511:0] u0_col_in_785;
wire [511:0] u0_col_in_786;
wire [511:0] u0_col_in_787;
wire [511:0] u0_col_in_788;
wire [511:0] u0_col_in_789;
wire [511:0] u0_col_in_790;
wire [511:0] u0_col_in_791;
wire [511:0] u0_col_in_792;
wire [511:0] u0_col_in_793;
wire [511:0] u0_col_in_794;
wire [511:0] u0_col_in_795;
wire [511:0] u0_col_in_796;
wire [511:0] u0_col_in_797;
wire [511:0] u0_col_in_798;
wire [511:0] u0_col_in_799;
wire [511:0] u0_col_in_800;
wire [511:0] u0_col_in_801;
wire [511:0] u0_col_in_802;
wire [511:0] u0_col_in_803;
wire [511:0] u0_col_in_804;
wire [511:0] u0_col_in_805;
wire [511:0] u0_col_in_806;
wire [511:0] u0_col_in_807;
wire [511:0] u0_col_in_808;
wire [511:0] u0_col_in_809;
wire [511:0] u0_col_in_810;
wire [511:0] u0_col_in_811;
wire [511:0] u0_col_in_812;
wire [511:0] u0_col_in_813;
wire [511:0] u0_col_in_814;
wire [511:0] u0_col_in_815;
wire [511:0] u0_col_in_816;
wire [511:0] u0_col_in_817;
wire [511:0] u0_col_in_818;
wire [511:0] u0_col_in_819;
wire [511:0] u0_col_in_820;
wire [511:0] u0_col_in_821;
wire [511:0] u0_col_in_822;
wire [511:0] u0_col_in_823;
wire [511:0] u0_col_in_824;
wire [511:0] u0_col_in_825;
wire [511:0] u0_col_in_826;
wire [511:0] u0_col_in_827;
wire [511:0] u0_col_in_828;
wire [511:0] u0_col_in_829;
wire [511:0] u0_col_in_830;
wire [511:0] u0_col_in_831;
wire [511:0] u0_col_in_832;
wire [511:0] u0_col_in_833;
wire [511:0] u0_col_in_834;
wire [511:0] u0_col_in_835;
wire [511:0] u0_col_in_836;
wire [511:0] u0_col_in_837;
wire [511:0] u0_col_in_838;
wire [511:0] u0_col_in_839;
wire [511:0] u0_col_in_840;
wire [511:0] u0_col_in_841;
wire [511:0] u0_col_in_842;
wire [511:0] u0_col_in_843;
wire [511:0] u0_col_in_844;
wire [511:0] u0_col_in_845;
wire [511:0] u0_col_in_846;
wire [511:0] u0_col_in_847;
wire [511:0] u0_col_in_848;
wire [511:0] u0_col_in_849;
wire [511:0] u0_col_in_850;
wire [511:0] u0_col_in_851;
wire [511:0] u0_col_in_852;
wire [511:0] u0_col_in_853;
wire [511:0] u0_col_in_854;
wire [511:0] u0_col_in_855;
wire [511:0] u0_col_in_856;
wire [511:0] u0_col_in_857;
wire [511:0] u0_col_in_858;
wire [511:0] u0_col_in_859;
wire [511:0] u0_col_in_860;
wire [511:0] u0_col_in_861;
wire [511:0] u0_col_in_862;
wire [511:0] u0_col_in_863;
wire [511:0] u0_col_in_864;
wire [511:0] u0_col_in_865;
wire [511:0] u0_col_in_866;
wire [511:0] u0_col_in_867;
wire [511:0] u0_col_in_868;
wire [511:0] u0_col_in_869;
wire [511:0] u0_col_in_870;
wire [511:0] u0_col_in_871;
wire [511:0] u0_col_in_872;
wire [511:0] u0_col_in_873;
wire [511:0] u0_col_in_874;
wire [511:0] u0_col_in_875;
wire [511:0] u0_col_in_876;
wire [511:0] u0_col_in_877;
wire [511:0] u0_col_in_878;
wire [511:0] u0_col_in_879;
wire [511:0] u0_col_in_880;
wire [511:0] u0_col_in_881;
wire [511:0] u0_col_in_882;
wire [511:0] u0_col_in_883;
wire [511:0] u0_col_in_884;
wire [511:0] u0_col_in_885;
wire [511:0] u0_col_in_886;
wire [511:0] u0_col_in_887;
wire [511:0] u0_col_in_888;
wire [511:0] u0_col_in_889;
wire [511:0] u0_col_in_890;
wire [511:0] u0_col_in_891;
wire [511:0] u0_col_in_892;
wire [511:0] u0_col_in_893;
wire [511:0] u0_col_in_894;
wire [511:0] u0_col_in_895;
wire [511:0] u0_col_in_896;
wire [511:0] u0_col_in_897;
wire [511:0] u0_col_in_898;
wire [511:0] u0_col_in_899;
wire [511:0] u0_col_in_900;
wire [511:0] u0_col_in_901;
wire [511:0] u0_col_in_902;
wire [511:0] u0_col_in_903;
wire [511:0] u0_col_in_904;
wire [511:0] u0_col_in_905;
wire [511:0] u0_col_in_906;
wire [511:0] u0_col_in_907;
wire [511:0] u0_col_in_908;
wire [511:0] u0_col_in_909;
wire [511:0] u0_col_in_910;
wire [511:0] u0_col_in_911;
wire [511:0] u0_col_in_912;
wire [511:0] u0_col_in_913;
wire [511:0] u0_col_in_914;
wire [511:0] u0_col_in_915;
wire [511:0] u0_col_in_916;
wire [511:0] u0_col_in_917;
wire [511:0] u0_col_in_918;
wire [511:0] u0_col_in_919;
wire [511:0] u0_col_in_920;
wire [511:0] u0_col_in_921;
wire [511:0] u0_col_in_922;
wire [511:0] u0_col_in_923;
wire [511:0] u0_col_in_924;
wire [511:0] u0_col_in_925;
wire [511:0] u0_col_in_926;
wire [511:0] u0_col_in_927;
wire [511:0] u0_col_in_928;
wire [511:0] u0_col_in_929;
wire [511:0] u0_col_in_930;
wire [511:0] u0_col_in_931;
wire [511:0] u0_col_in_932;
wire [511:0] u0_col_in_933;
wire [511:0] u0_col_in_934;
wire [511:0] u0_col_in_935;
wire [511:0] u0_col_in_936;
wire [511:0] u0_col_in_937;
wire [511:0] u0_col_in_938;
wire [511:0] u0_col_in_939;
wire [511:0] u0_col_in_940;
wire [511:0] u0_col_in_941;
wire [511:0] u0_col_in_942;
wire [511:0] u0_col_in_943;
wire [511:0] u0_col_in_944;
wire [511:0] u0_col_in_945;
wire [511:0] u0_col_in_946;
wire [511:0] u0_col_in_947;
wire [511:0] u0_col_in_948;
wire [511:0] u0_col_in_949;
wire [511:0] u0_col_in_950;
wire [511:0] u0_col_in_951;
wire [511:0] u0_col_in_952;
wire [511:0] u0_col_in_953;
wire [511:0] u0_col_in_954;
wire [511:0] u0_col_in_955;
wire [511:0] u0_col_in_956;
wire [511:0] u0_col_in_957;
wire [511:0] u0_col_in_958;
wire [511:0] u0_col_in_959;
wire [511:0] u0_col_in_960;
wire [511:0] u0_col_in_961;
wire [511:0] u0_col_in_962;
wire [511:0] u0_col_in_963;
wire [511:0] u0_col_in_964;
wire [511:0] u0_col_in_965;
wire [511:0] u0_col_in_966;
wire [511:0] u0_col_in_967;
wire [511:0] u0_col_in_968;
wire [511:0] u0_col_in_969;
wire [511:0] u0_col_in_970;
wire [511:0] u0_col_in_971;
wire [511:0] u0_col_in_972;
wire [511:0] u0_col_in_973;
wire [511:0] u0_col_in_974;
wire [511:0] u0_col_in_975;
wire [511:0] u0_col_in_976;
wire [511:0] u0_col_in_977;
wire [511:0] u0_col_in_978;
wire [511:0] u0_col_in_979;
wire [511:0] u0_col_in_980;
wire [511:0] u0_col_in_981;
wire [511:0] u0_col_in_982;
wire [511:0] u0_col_in_983;
wire [511:0] u0_col_in_984;
wire [511:0] u0_col_in_985;
wire [511:0] u0_col_in_986;
wire [511:0] u0_col_in_987;
wire [511:0] u0_col_in_988;
wire [511:0] u0_col_in_989;
wire [511:0] u0_col_in_990;
wire [511:0] u0_col_in_991;
wire [511:0] u0_col_in_992;
wire [511:0] u0_col_in_993;
wire [511:0] u0_col_in_994;
wire [511:0] u0_col_in_995;
wire [511:0] u0_col_in_996;
wire [511:0] u0_col_in_997;
wire [511:0] u0_col_in_998;
wire [511:0] u0_col_in_999;
wire [511:0] u0_col_in_1000;
wire [511:0] u0_col_in_1001;
wire [511:0] u0_col_in_1002;
wire [511:0] u0_col_in_1003;
wire [511:0] u0_col_in_1004;
wire [511:0] u0_col_in_1005;
wire [511:0] u0_col_in_1006;
wire [511:0] u0_col_in_1007;
wire [511:0] u0_col_in_1008;
wire [511:0] u0_col_in_1009;
wire [511:0] u0_col_in_1010;
wire [511:0] u0_col_in_1011;
wire [511:0] u0_col_in_1012;
wire [511:0] u0_col_in_1013;
wire [511:0] u0_col_in_1014;
wire [511:0] u0_col_in_1015;
wire [511:0] u0_col_in_1016;
wire [511:0] u0_col_in_1017;
wire [511:0] u0_col_in_1018;
wire [511:0] u0_col_in_1019;
wire [511:0] u0_col_in_1020;
wire [511:0] u0_col_in_1021;
wire [511:0] u0_col_in_1022;
wire [511:0] u0_col_in_1023;






//*****************************************************
//**************u0输出定义******************************
//*****************************************************
wire [151:0] u0_col_out_0;
wire [151:0] u0_col_out_1;
wire [151:0] u0_col_out_2;
wire [151:0] u0_col_out_3;
wire [151:0] u0_col_out_4;
wire [151:0] u0_col_out_5;
wire [151:0] u0_col_out_6;
wire [151:0] u0_col_out_7;
wire [151:0] u0_col_out_8;
wire [151:0] u0_col_out_9;
wire [151:0] u0_col_out_10;
wire [151:0] u0_col_out_11;
wire [151:0] u0_col_out_12;
wire [151:0] u0_col_out_13;
wire [151:0] u0_col_out_14;
wire [151:0] u0_col_out_15;
wire [151:0] u0_col_out_16;
wire [151:0] u0_col_out_17;
wire [151:0] u0_col_out_18;
wire [151:0] u0_col_out_19;
wire [151:0] u0_col_out_20;
wire [151:0] u0_col_out_21;
wire [151:0] u0_col_out_22;
wire [151:0] u0_col_out_23;
wire [151:0] u0_col_out_24;
wire [151:0] u0_col_out_25;
wire [151:0] u0_col_out_26;
wire [151:0] u0_col_out_27;
wire [151:0] u0_col_out_28;
wire [151:0] u0_col_out_29;
wire [151:0] u0_col_out_30;
wire [151:0] u0_col_out_31;
wire [151:0] u0_col_out_32;
wire [151:0] u0_col_out_33;
wire [151:0] u0_col_out_34;
wire [151:0] u0_col_out_35;
wire [151:0] u0_col_out_36;
wire [151:0] u0_col_out_37;
wire [151:0] u0_col_out_38;
wire [151:0] u0_col_out_39;
wire [151:0] u0_col_out_40;
wire [151:0] u0_col_out_41;
wire [151:0] u0_col_out_42;
wire [151:0] u0_col_out_43;
wire [151:0] u0_col_out_44;
wire [151:0] u0_col_out_45;
wire [151:0] u0_col_out_46;
wire [151:0] u0_col_out_47;
wire [151:0] u0_col_out_48;
wire [151:0] u0_col_out_49;
wire [151:0] u0_col_out_50;
wire [151:0] u0_col_out_51;
wire [151:0] u0_col_out_52;
wire [151:0] u0_col_out_53;
wire [151:0] u0_col_out_54;
wire [151:0] u0_col_out_55;
wire [151:0] u0_col_out_56;
wire [151:0] u0_col_out_57;
wire [151:0] u0_col_out_58;
wire [151:0] u0_col_out_59;
wire [151:0] u0_col_out_60;
wire [151:0] u0_col_out_61;
wire [151:0] u0_col_out_62;
wire [151:0] u0_col_out_63;
wire [151:0] u0_col_out_64;
wire [151:0] u0_col_out_65;
wire [151:0] u0_col_out_66;
wire [151:0] u0_col_out_67;
wire [151:0] u0_col_out_68;
wire [151:0] u0_col_out_69;
wire [151:0] u0_col_out_70;
wire [151:0] u0_col_out_71;
wire [151:0] u0_col_out_72;
wire [151:0] u0_col_out_73;
wire [151:0] u0_col_out_74;
wire [151:0] u0_col_out_75;
wire [151:0] u0_col_out_76;
wire [151:0] u0_col_out_77;
wire [151:0] u0_col_out_78;
wire [151:0] u0_col_out_79;
wire [151:0] u0_col_out_80;
wire [151:0] u0_col_out_81;
wire [151:0] u0_col_out_82;
wire [151:0] u0_col_out_83;
wire [151:0] u0_col_out_84;
wire [151:0] u0_col_out_85;
wire [151:0] u0_col_out_86;
wire [151:0] u0_col_out_87;
wire [151:0] u0_col_out_88;
wire [151:0] u0_col_out_89;
wire [151:0] u0_col_out_90;
wire [151:0] u0_col_out_91;
wire [151:0] u0_col_out_92;
wire [151:0] u0_col_out_93;
wire [151:0] u0_col_out_94;
wire [151:0] u0_col_out_95;
wire [151:0] u0_col_out_96;
wire [151:0] u0_col_out_97;
wire [151:0] u0_col_out_98;
wire [151:0] u0_col_out_99;
wire [151:0] u0_col_out_100;
wire [151:0] u0_col_out_101;
wire [151:0] u0_col_out_102;
wire [151:0] u0_col_out_103;
wire [151:0] u0_col_out_104;
wire [151:0] u0_col_out_105;
wire [151:0] u0_col_out_106;
wire [151:0] u0_col_out_107;
wire [151:0] u0_col_out_108;
wire [151:0] u0_col_out_109;
wire [151:0] u0_col_out_110;
wire [151:0] u0_col_out_111;
wire [151:0] u0_col_out_112;
wire [151:0] u0_col_out_113;
wire [151:0] u0_col_out_114;
wire [151:0] u0_col_out_115;
wire [151:0] u0_col_out_116;
wire [151:0] u0_col_out_117;
wire [151:0] u0_col_out_118;
wire [151:0] u0_col_out_119;
wire [151:0] u0_col_out_120;
wire [151:0] u0_col_out_121;
wire [151:0] u0_col_out_122;
wire [151:0] u0_col_out_123;
wire [151:0] u0_col_out_124;
wire [151:0] u0_col_out_125;
wire [151:0] u0_col_out_126;
wire [151:0] u0_col_out_127;
wire [151:0] u0_col_out_128;
wire [151:0] u0_col_out_129;
wire [151:0] u0_col_out_130;
wire [151:0] u0_col_out_131;
wire [151:0] u0_col_out_132;
wire [151:0] u0_col_out_133;
wire [151:0] u0_col_out_134;
wire [151:0] u0_col_out_135;
wire [151:0] u0_col_out_136;
wire [151:0] u0_col_out_137;
wire [151:0] u0_col_out_138;
wire [151:0] u0_col_out_139;
wire [151:0] u0_col_out_140;
wire [151:0] u0_col_out_141;
wire [151:0] u0_col_out_142;
wire [151:0] u0_col_out_143;
wire [151:0] u0_col_out_144;
wire [151:0] u0_col_out_145;
wire [151:0] u0_col_out_146;
wire [151:0] u0_col_out_147;
wire [151:0] u0_col_out_148;
wire [151:0] u0_col_out_149;
wire [151:0] u0_col_out_150;
wire [151:0] u0_col_out_151;
wire [151:0] u0_col_out_152;
wire [151:0] u0_col_out_153;
wire [151:0] u0_col_out_154;
wire [151:0] u0_col_out_155;
wire [151:0] u0_col_out_156;
wire [151:0] u0_col_out_157;
wire [151:0] u0_col_out_158;
wire [151:0] u0_col_out_159;
wire [151:0] u0_col_out_160;
wire [151:0] u0_col_out_161;
wire [151:0] u0_col_out_162;
wire [151:0] u0_col_out_163;
wire [151:0] u0_col_out_164;
wire [151:0] u0_col_out_165;
wire [151:0] u0_col_out_166;
wire [151:0] u0_col_out_167;
wire [151:0] u0_col_out_168;
wire [151:0] u0_col_out_169;
wire [151:0] u0_col_out_170;
wire [151:0] u0_col_out_171;
wire [151:0] u0_col_out_172;
wire [151:0] u0_col_out_173;
wire [151:0] u0_col_out_174;
wire [151:0] u0_col_out_175;
wire [151:0] u0_col_out_176;
wire [151:0] u0_col_out_177;
wire [151:0] u0_col_out_178;
wire [151:0] u0_col_out_179;
wire [151:0] u0_col_out_180;
wire [151:0] u0_col_out_181;
wire [151:0] u0_col_out_182;
wire [151:0] u0_col_out_183;
wire [151:0] u0_col_out_184;
wire [151:0] u0_col_out_185;
wire [151:0] u0_col_out_186;
wire [151:0] u0_col_out_187;
wire [151:0] u0_col_out_188;
wire [151:0] u0_col_out_189;
wire [151:0] u0_col_out_190;
wire [151:0] u0_col_out_191;
wire [151:0] u0_col_out_192;
wire [151:0] u0_col_out_193;
wire [151:0] u0_col_out_194;
wire [151:0] u0_col_out_195;
wire [151:0] u0_col_out_196;
wire [151:0] u0_col_out_197;
wire [151:0] u0_col_out_198;
wire [151:0] u0_col_out_199;
wire [151:0] u0_col_out_200;
wire [151:0] u0_col_out_201;
wire [151:0] u0_col_out_202;
wire [151:0] u0_col_out_203;
wire [151:0] u0_col_out_204;
wire [151:0] u0_col_out_205;
wire [151:0] u0_col_out_206;
wire [151:0] u0_col_out_207;
wire [151:0] u0_col_out_208;
wire [151:0] u0_col_out_209;
wire [151:0] u0_col_out_210;
wire [151:0] u0_col_out_211;
wire [151:0] u0_col_out_212;
wire [151:0] u0_col_out_213;
wire [151:0] u0_col_out_214;
wire [151:0] u0_col_out_215;
wire [151:0] u0_col_out_216;
wire [151:0] u0_col_out_217;
wire [151:0] u0_col_out_218;
wire [151:0] u0_col_out_219;
wire [151:0] u0_col_out_220;
wire [151:0] u0_col_out_221;
wire [151:0] u0_col_out_222;
wire [151:0] u0_col_out_223;
wire [151:0] u0_col_out_224;
wire [151:0] u0_col_out_225;
wire [151:0] u0_col_out_226;
wire [151:0] u0_col_out_227;
wire [151:0] u0_col_out_228;
wire [151:0] u0_col_out_229;
wire [151:0] u0_col_out_230;
wire [151:0] u0_col_out_231;
wire [151:0] u0_col_out_232;
wire [151:0] u0_col_out_233;
wire [151:0] u0_col_out_234;
wire [151:0] u0_col_out_235;
wire [151:0] u0_col_out_236;
wire [151:0] u0_col_out_237;
wire [151:0] u0_col_out_238;
wire [151:0] u0_col_out_239;
wire [151:0] u0_col_out_240;
wire [151:0] u0_col_out_241;
wire [151:0] u0_col_out_242;
wire [151:0] u0_col_out_243;
wire [151:0] u0_col_out_244;
wire [151:0] u0_col_out_245;
wire [151:0] u0_col_out_246;
wire [151:0] u0_col_out_247;
wire [151:0] u0_col_out_248;
wire [151:0] u0_col_out_249;
wire [151:0] u0_col_out_250;
wire [151:0] u0_col_out_251;
wire [151:0] u0_col_out_252;
wire [151:0] u0_col_out_253;
wire [151:0] u0_col_out_254;
wire [151:0] u0_col_out_255;
wire [151:0] u0_col_out_256;
wire [151:0] u0_col_out_257;
wire [151:0] u0_col_out_258;
wire [151:0] u0_col_out_259;
wire [151:0] u0_col_out_260;
wire [151:0] u0_col_out_261;
wire [151:0] u0_col_out_262;
wire [151:0] u0_col_out_263;
wire [151:0] u0_col_out_264;
wire [151:0] u0_col_out_265;
wire [151:0] u0_col_out_266;
wire [151:0] u0_col_out_267;
wire [151:0] u0_col_out_268;
wire [151:0] u0_col_out_269;
wire [151:0] u0_col_out_270;
wire [151:0] u0_col_out_271;
wire [151:0] u0_col_out_272;
wire [151:0] u0_col_out_273;
wire [151:0] u0_col_out_274;
wire [151:0] u0_col_out_275;
wire [151:0] u0_col_out_276;
wire [151:0] u0_col_out_277;
wire [151:0] u0_col_out_278;
wire [151:0] u0_col_out_279;
wire [151:0] u0_col_out_280;
wire [151:0] u0_col_out_281;
wire [151:0] u0_col_out_282;
wire [151:0] u0_col_out_283;
wire [151:0] u0_col_out_284;
wire [151:0] u0_col_out_285;
wire [151:0] u0_col_out_286;
wire [151:0] u0_col_out_287;
wire [151:0] u0_col_out_288;
wire [151:0] u0_col_out_289;
wire [151:0] u0_col_out_290;
wire [151:0] u0_col_out_291;
wire [151:0] u0_col_out_292;
wire [151:0] u0_col_out_293;
wire [151:0] u0_col_out_294;
wire [151:0] u0_col_out_295;
wire [151:0] u0_col_out_296;
wire [151:0] u0_col_out_297;
wire [151:0] u0_col_out_298;
wire [151:0] u0_col_out_299;
wire [151:0] u0_col_out_300;
wire [151:0] u0_col_out_301;
wire [151:0] u0_col_out_302;
wire [151:0] u0_col_out_303;
wire [151:0] u0_col_out_304;
wire [151:0] u0_col_out_305;
wire [151:0] u0_col_out_306;
wire [151:0] u0_col_out_307;
wire [151:0] u0_col_out_308;
wire [151:0] u0_col_out_309;
wire [151:0] u0_col_out_310;
wire [151:0] u0_col_out_311;
wire [151:0] u0_col_out_312;
wire [151:0] u0_col_out_313;
wire [151:0] u0_col_out_314;
wire [151:0] u0_col_out_315;
wire [151:0] u0_col_out_316;
wire [151:0] u0_col_out_317;
wire [151:0] u0_col_out_318;
wire [151:0] u0_col_out_319;
wire [151:0] u0_col_out_320;
wire [151:0] u0_col_out_321;
wire [151:0] u0_col_out_322;
wire [151:0] u0_col_out_323;
wire [151:0] u0_col_out_324;
wire [151:0] u0_col_out_325;
wire [151:0] u0_col_out_326;
wire [151:0] u0_col_out_327;
wire [151:0] u0_col_out_328;
wire [151:0] u0_col_out_329;
wire [151:0] u0_col_out_330;
wire [151:0] u0_col_out_331;
wire [151:0] u0_col_out_332;
wire [151:0] u0_col_out_333;
wire [151:0] u0_col_out_334;
wire [151:0] u0_col_out_335;
wire [151:0] u0_col_out_336;
wire [151:0] u0_col_out_337;
wire [151:0] u0_col_out_338;
wire [151:0] u0_col_out_339;
wire [151:0] u0_col_out_340;
wire [151:0] u0_col_out_341;
wire [151:0] u0_col_out_342;
wire [151:0] u0_col_out_343;
wire [151:0] u0_col_out_344;
wire [151:0] u0_col_out_345;
wire [151:0] u0_col_out_346;
wire [151:0] u0_col_out_347;
wire [151:0] u0_col_out_348;
wire [151:0] u0_col_out_349;
wire [151:0] u0_col_out_350;
wire [151:0] u0_col_out_351;
wire [151:0] u0_col_out_352;
wire [151:0] u0_col_out_353;
wire [151:0] u0_col_out_354;
wire [151:0] u0_col_out_355;
wire [151:0] u0_col_out_356;
wire [151:0] u0_col_out_357;
wire [151:0] u0_col_out_358;
wire [151:0] u0_col_out_359;
wire [151:0] u0_col_out_360;
wire [151:0] u0_col_out_361;
wire [151:0] u0_col_out_362;
wire [151:0] u0_col_out_363;
wire [151:0] u0_col_out_364;
wire [151:0] u0_col_out_365;
wire [151:0] u0_col_out_366;
wire [151:0] u0_col_out_367;
wire [151:0] u0_col_out_368;
wire [151:0] u0_col_out_369;
wire [151:0] u0_col_out_370;
wire [151:0] u0_col_out_371;
wire [151:0] u0_col_out_372;
wire [151:0] u0_col_out_373;
wire [151:0] u0_col_out_374;
wire [151:0] u0_col_out_375;
wire [151:0] u0_col_out_376;
wire [151:0] u0_col_out_377;
wire [151:0] u0_col_out_378;
wire [151:0] u0_col_out_379;
wire [151:0] u0_col_out_380;
wire [151:0] u0_col_out_381;
wire [151:0] u0_col_out_382;
wire [151:0] u0_col_out_383;
wire [151:0] u0_col_out_384;
wire [151:0] u0_col_out_385;
wire [151:0] u0_col_out_386;
wire [151:0] u0_col_out_387;
wire [151:0] u0_col_out_388;
wire [151:0] u0_col_out_389;
wire [151:0] u0_col_out_390;
wire [151:0] u0_col_out_391;
wire [151:0] u0_col_out_392;
wire [151:0] u0_col_out_393;
wire [151:0] u0_col_out_394;
wire [151:0] u0_col_out_395;
wire [151:0] u0_col_out_396;
wire [151:0] u0_col_out_397;
wire [151:0] u0_col_out_398;
wire [151:0] u0_col_out_399;
wire [151:0] u0_col_out_400;
wire [151:0] u0_col_out_401;
wire [151:0] u0_col_out_402;
wire [151:0] u0_col_out_403;
wire [151:0] u0_col_out_404;
wire [151:0] u0_col_out_405;
wire [151:0] u0_col_out_406;
wire [151:0] u0_col_out_407;
wire [151:0] u0_col_out_408;
wire [151:0] u0_col_out_409;
wire [151:0] u0_col_out_410;
wire [151:0] u0_col_out_411;
wire [151:0] u0_col_out_412;
wire [151:0] u0_col_out_413;
wire [151:0] u0_col_out_414;
wire [151:0] u0_col_out_415;
wire [151:0] u0_col_out_416;
wire [151:0] u0_col_out_417;
wire [151:0] u0_col_out_418;
wire [151:0] u0_col_out_419;
wire [151:0] u0_col_out_420;
wire [151:0] u0_col_out_421;
wire [151:0] u0_col_out_422;
wire [151:0] u0_col_out_423;
wire [151:0] u0_col_out_424;
wire [151:0] u0_col_out_425;
wire [151:0] u0_col_out_426;
wire [151:0] u0_col_out_427;
wire [151:0] u0_col_out_428;
wire [151:0] u0_col_out_429;
wire [151:0] u0_col_out_430;
wire [151:0] u0_col_out_431;
wire [151:0] u0_col_out_432;
wire [151:0] u0_col_out_433;
wire [151:0] u0_col_out_434;
wire [151:0] u0_col_out_435;
wire [151:0] u0_col_out_436;
wire [151:0] u0_col_out_437;
wire [151:0] u0_col_out_438;
wire [151:0] u0_col_out_439;
wire [151:0] u0_col_out_440;
wire [151:0] u0_col_out_441;
wire [151:0] u0_col_out_442;
wire [151:0] u0_col_out_443;
wire [151:0] u0_col_out_444;
wire [151:0] u0_col_out_445;
wire [151:0] u0_col_out_446;
wire [151:0] u0_col_out_447;
wire [151:0] u0_col_out_448;
wire [151:0] u0_col_out_449;
wire [151:0] u0_col_out_450;
wire [151:0] u0_col_out_451;
wire [151:0] u0_col_out_452;
wire [151:0] u0_col_out_453;
wire [151:0] u0_col_out_454;
wire [151:0] u0_col_out_455;
wire [151:0] u0_col_out_456;
wire [151:0] u0_col_out_457;
wire [151:0] u0_col_out_458;
wire [151:0] u0_col_out_459;
wire [151:0] u0_col_out_460;
wire [151:0] u0_col_out_461;
wire [151:0] u0_col_out_462;
wire [151:0] u0_col_out_463;
wire [151:0] u0_col_out_464;
wire [151:0] u0_col_out_465;
wire [151:0] u0_col_out_466;
wire [151:0] u0_col_out_467;
wire [151:0] u0_col_out_468;
wire [151:0] u0_col_out_469;
wire [151:0] u0_col_out_470;
wire [151:0] u0_col_out_471;
wire [151:0] u0_col_out_472;
wire [151:0] u0_col_out_473;
wire [151:0] u0_col_out_474;
wire [151:0] u0_col_out_475;
wire [151:0] u0_col_out_476;
wire [151:0] u0_col_out_477;
wire [151:0] u0_col_out_478;
wire [151:0] u0_col_out_479;
wire [151:0] u0_col_out_480;
wire [151:0] u0_col_out_481;
wire [151:0] u0_col_out_482;
wire [151:0] u0_col_out_483;
wire [151:0] u0_col_out_484;
wire [151:0] u0_col_out_485;
wire [151:0] u0_col_out_486;
wire [151:0] u0_col_out_487;
wire [151:0] u0_col_out_488;
wire [151:0] u0_col_out_489;
wire [151:0] u0_col_out_490;
wire [151:0] u0_col_out_491;
wire [151:0] u0_col_out_492;
wire [151:0] u0_col_out_493;
wire [151:0] u0_col_out_494;
wire [151:0] u0_col_out_495;
wire [151:0] u0_col_out_496;
wire [151:0] u0_col_out_497;
wire [151:0] u0_col_out_498;
wire [151:0] u0_col_out_499;
wire [151:0] u0_col_out_500;
wire [151:0] u0_col_out_501;
wire [151:0] u0_col_out_502;
wire [151:0] u0_col_out_503;
wire [151:0] u0_col_out_504;
wire [151:0] u0_col_out_505;
wire [151:0] u0_col_out_506;
wire [151:0] u0_col_out_507;
wire [151:0] u0_col_out_508;
wire [151:0] u0_col_out_509;
wire [151:0] u0_col_out_510;
wire [151:0] u0_col_out_511;
wire [151:0] u0_col_out_512;
wire [151:0] u0_col_out_513;
wire [151:0] u0_col_out_514;
wire [151:0] u0_col_out_515;
wire [151:0] u0_col_out_516;
wire [151:0] u0_col_out_517;
wire [151:0] u0_col_out_518;
wire [151:0] u0_col_out_519;
wire [151:0] u0_col_out_520;
wire [151:0] u0_col_out_521;
wire [151:0] u0_col_out_522;
wire [151:0] u0_col_out_523;
wire [151:0] u0_col_out_524;
wire [151:0] u0_col_out_525;
wire [151:0] u0_col_out_526;
wire [151:0] u0_col_out_527;
wire [151:0] u0_col_out_528;
wire [151:0] u0_col_out_529;
wire [151:0] u0_col_out_530;
wire [151:0] u0_col_out_531;
wire [151:0] u0_col_out_532;
wire [151:0] u0_col_out_533;
wire [151:0] u0_col_out_534;
wire [151:0] u0_col_out_535;
wire [151:0] u0_col_out_536;
wire [151:0] u0_col_out_537;
wire [151:0] u0_col_out_538;
wire [151:0] u0_col_out_539;
wire [151:0] u0_col_out_540;
wire [151:0] u0_col_out_541;
wire [151:0] u0_col_out_542;
wire [151:0] u0_col_out_543;
wire [151:0] u0_col_out_544;
wire [151:0] u0_col_out_545;
wire [151:0] u0_col_out_546;
wire [151:0] u0_col_out_547;
wire [151:0] u0_col_out_548;
wire [151:0] u0_col_out_549;
wire [151:0] u0_col_out_550;
wire [151:0] u0_col_out_551;
wire [151:0] u0_col_out_552;
wire [151:0] u0_col_out_553;
wire [151:0] u0_col_out_554;
wire [151:0] u0_col_out_555;
wire [151:0] u0_col_out_556;
wire [151:0] u0_col_out_557;
wire [151:0] u0_col_out_558;
wire [151:0] u0_col_out_559;
wire [151:0] u0_col_out_560;
wire [151:0] u0_col_out_561;
wire [151:0] u0_col_out_562;
wire [151:0] u0_col_out_563;
wire [151:0] u0_col_out_564;
wire [151:0] u0_col_out_565;
wire [151:0] u0_col_out_566;
wire [151:0] u0_col_out_567;
wire [151:0] u0_col_out_568;
wire [151:0] u0_col_out_569;
wire [151:0] u0_col_out_570;
wire [151:0] u0_col_out_571;
wire [151:0] u0_col_out_572;
wire [151:0] u0_col_out_573;
wire [151:0] u0_col_out_574;
wire [151:0] u0_col_out_575;
wire [151:0] u0_col_out_576;
wire [151:0] u0_col_out_577;
wire [151:0] u0_col_out_578;
wire [151:0] u0_col_out_579;
wire [151:0] u0_col_out_580;
wire [151:0] u0_col_out_581;
wire [151:0] u0_col_out_582;
wire [151:0] u0_col_out_583;
wire [151:0] u0_col_out_584;
wire [151:0] u0_col_out_585;
wire [151:0] u0_col_out_586;
wire [151:0] u0_col_out_587;
wire [151:0] u0_col_out_588;
wire [151:0] u0_col_out_589;
wire [151:0] u0_col_out_590;
wire [151:0] u0_col_out_591;
wire [151:0] u0_col_out_592;
wire [151:0] u0_col_out_593;
wire [151:0] u0_col_out_594;
wire [151:0] u0_col_out_595;
wire [151:0] u0_col_out_596;
wire [151:0] u0_col_out_597;
wire [151:0] u0_col_out_598;
wire [151:0] u0_col_out_599;
wire [151:0] u0_col_out_600;
wire [151:0] u0_col_out_601;
wire [151:0] u0_col_out_602;
wire [151:0] u0_col_out_603;
wire [151:0] u0_col_out_604;
wire [151:0] u0_col_out_605;
wire [151:0] u0_col_out_606;
wire [151:0] u0_col_out_607;
wire [151:0] u0_col_out_608;
wire [151:0] u0_col_out_609;
wire [151:0] u0_col_out_610;
wire [151:0] u0_col_out_611;
wire [151:0] u0_col_out_612;
wire [151:0] u0_col_out_613;
wire [151:0] u0_col_out_614;
wire [151:0] u0_col_out_615;
wire [151:0] u0_col_out_616;
wire [151:0] u0_col_out_617;
wire [151:0] u0_col_out_618;
wire [151:0] u0_col_out_619;
wire [151:0] u0_col_out_620;
wire [151:0] u0_col_out_621;
wire [151:0] u0_col_out_622;
wire [151:0] u0_col_out_623;
wire [151:0] u0_col_out_624;
wire [151:0] u0_col_out_625;
wire [151:0] u0_col_out_626;
wire [151:0] u0_col_out_627;
wire [151:0] u0_col_out_628;
wire [151:0] u0_col_out_629;
wire [151:0] u0_col_out_630;
wire [151:0] u0_col_out_631;
wire [151:0] u0_col_out_632;
wire [151:0] u0_col_out_633;
wire [151:0] u0_col_out_634;
wire [151:0] u0_col_out_635;
wire [151:0] u0_col_out_636;
wire [151:0] u0_col_out_637;
wire [151:0] u0_col_out_638;
wire [151:0] u0_col_out_639;
wire [151:0] u0_col_out_640;
wire [151:0] u0_col_out_641;
wire [151:0] u0_col_out_642;
wire [151:0] u0_col_out_643;
wire [151:0] u0_col_out_644;
wire [151:0] u0_col_out_645;
wire [151:0] u0_col_out_646;
wire [151:0] u0_col_out_647;
wire [151:0] u0_col_out_648;
wire [151:0] u0_col_out_649;
wire [151:0] u0_col_out_650;
wire [151:0] u0_col_out_651;
wire [151:0] u0_col_out_652;
wire [151:0] u0_col_out_653;
wire [151:0] u0_col_out_654;
wire [151:0] u0_col_out_655;
wire [151:0] u0_col_out_656;
wire [151:0] u0_col_out_657;
wire [151:0] u0_col_out_658;
wire [151:0] u0_col_out_659;
wire [151:0] u0_col_out_660;
wire [151:0] u0_col_out_661;
wire [151:0] u0_col_out_662;
wire [151:0] u0_col_out_663;
wire [151:0] u0_col_out_664;
wire [151:0] u0_col_out_665;
wire [151:0] u0_col_out_666;
wire [151:0] u0_col_out_667;
wire [151:0] u0_col_out_668;
wire [151:0] u0_col_out_669;
wire [151:0] u0_col_out_670;
wire [151:0] u0_col_out_671;
wire [151:0] u0_col_out_672;
wire [151:0] u0_col_out_673;
wire [151:0] u0_col_out_674;
wire [151:0] u0_col_out_675;
wire [151:0] u0_col_out_676;
wire [151:0] u0_col_out_677;
wire [151:0] u0_col_out_678;
wire [151:0] u0_col_out_679;
wire [151:0] u0_col_out_680;
wire [151:0] u0_col_out_681;
wire [151:0] u0_col_out_682;
wire [151:0] u0_col_out_683;
wire [151:0] u0_col_out_684;
wire [151:0] u0_col_out_685;
wire [151:0] u0_col_out_686;
wire [151:0] u0_col_out_687;
wire [151:0] u0_col_out_688;
wire [151:0] u0_col_out_689;
wire [151:0] u0_col_out_690;
wire [151:0] u0_col_out_691;
wire [151:0] u0_col_out_692;
wire [151:0] u0_col_out_693;
wire [151:0] u0_col_out_694;
wire [151:0] u0_col_out_695;
wire [151:0] u0_col_out_696;
wire [151:0] u0_col_out_697;
wire [151:0] u0_col_out_698;
wire [151:0] u0_col_out_699;
wire [151:0] u0_col_out_700;
wire [151:0] u0_col_out_701;
wire [151:0] u0_col_out_702;
wire [151:0] u0_col_out_703;
wire [151:0] u0_col_out_704;
wire [151:0] u0_col_out_705;
wire [151:0] u0_col_out_706;
wire [151:0] u0_col_out_707;
wire [151:0] u0_col_out_708;
wire [151:0] u0_col_out_709;
wire [151:0] u0_col_out_710;
wire [151:0] u0_col_out_711;
wire [151:0] u0_col_out_712;
wire [151:0] u0_col_out_713;
wire [151:0] u0_col_out_714;
wire [151:0] u0_col_out_715;
wire [151:0] u0_col_out_716;
wire [151:0] u0_col_out_717;
wire [151:0] u0_col_out_718;
wire [151:0] u0_col_out_719;
wire [151:0] u0_col_out_720;
wire [151:0] u0_col_out_721;
wire [151:0] u0_col_out_722;
wire [151:0] u0_col_out_723;
wire [151:0] u0_col_out_724;
wire [151:0] u0_col_out_725;
wire [151:0] u0_col_out_726;
wire [151:0] u0_col_out_727;
wire [151:0] u0_col_out_728;
wire [151:0] u0_col_out_729;
wire [151:0] u0_col_out_730;
wire [151:0] u0_col_out_731;
wire [151:0] u0_col_out_732;
wire [151:0] u0_col_out_733;
wire [151:0] u0_col_out_734;
wire [151:0] u0_col_out_735;
wire [151:0] u0_col_out_736;
wire [151:0] u0_col_out_737;
wire [151:0] u0_col_out_738;
wire [151:0] u0_col_out_739;
wire [151:0] u0_col_out_740;
wire [151:0] u0_col_out_741;
wire [151:0] u0_col_out_742;
wire [151:0] u0_col_out_743;
wire [151:0] u0_col_out_744;
wire [151:0] u0_col_out_745;
wire [151:0] u0_col_out_746;
wire [151:0] u0_col_out_747;
wire [151:0] u0_col_out_748;
wire [151:0] u0_col_out_749;
wire [151:0] u0_col_out_750;
wire [151:0] u0_col_out_751;
wire [151:0] u0_col_out_752;
wire [151:0] u0_col_out_753;
wire [151:0] u0_col_out_754;
wire [151:0] u0_col_out_755;
wire [151:0] u0_col_out_756;
wire [151:0] u0_col_out_757;
wire [151:0] u0_col_out_758;
wire [151:0] u0_col_out_759;
wire [151:0] u0_col_out_760;
wire [151:0] u0_col_out_761;
wire [151:0] u0_col_out_762;
wire [151:0] u0_col_out_763;
wire [151:0] u0_col_out_764;
wire [151:0] u0_col_out_765;
wire [151:0] u0_col_out_766;
wire [151:0] u0_col_out_767;
wire [151:0] u0_col_out_768;
wire [151:0] u0_col_out_769;
wire [151:0] u0_col_out_770;
wire [151:0] u0_col_out_771;
wire [151:0] u0_col_out_772;
wire [151:0] u0_col_out_773;
wire [151:0] u0_col_out_774;
wire [151:0] u0_col_out_775;
wire [151:0] u0_col_out_776;
wire [151:0] u0_col_out_777;
wire [151:0] u0_col_out_778;
wire [151:0] u0_col_out_779;
wire [151:0] u0_col_out_780;
wire [151:0] u0_col_out_781;
wire [151:0] u0_col_out_782;
wire [151:0] u0_col_out_783;
wire [151:0] u0_col_out_784;
wire [151:0] u0_col_out_785;
wire [151:0] u0_col_out_786;
wire [151:0] u0_col_out_787;
wire [151:0] u0_col_out_788;
wire [151:0] u0_col_out_789;
wire [151:0] u0_col_out_790;
wire [151:0] u0_col_out_791;
wire [151:0] u0_col_out_792;
wire [151:0] u0_col_out_793;
wire [151:0] u0_col_out_794;
wire [151:0] u0_col_out_795;
wire [151:0] u0_col_out_796;
wire [151:0] u0_col_out_797;
wire [151:0] u0_col_out_798;
wire [151:0] u0_col_out_799;
wire [151:0] u0_col_out_800;
wire [151:0] u0_col_out_801;
wire [151:0] u0_col_out_802;
wire [151:0] u0_col_out_803;
wire [151:0] u0_col_out_804;
wire [151:0] u0_col_out_805;
wire [151:0] u0_col_out_806;
wire [151:0] u0_col_out_807;
wire [151:0] u0_col_out_808;
wire [151:0] u0_col_out_809;
wire [151:0] u0_col_out_810;
wire [151:0] u0_col_out_811;
wire [151:0] u0_col_out_812;
wire [151:0] u0_col_out_813;
wire [151:0] u0_col_out_814;
wire [151:0] u0_col_out_815;
wire [151:0] u0_col_out_816;
wire [151:0] u0_col_out_817;
wire [151:0] u0_col_out_818;
wire [151:0] u0_col_out_819;
wire [151:0] u0_col_out_820;
wire [151:0] u0_col_out_821;
wire [151:0] u0_col_out_822;
wire [151:0] u0_col_out_823;
wire [151:0] u0_col_out_824;
wire [151:0] u0_col_out_825;
wire [151:0] u0_col_out_826;
wire [151:0] u0_col_out_827;
wire [151:0] u0_col_out_828;
wire [151:0] u0_col_out_829;
wire [151:0] u0_col_out_830;
wire [151:0] u0_col_out_831;
wire [151:0] u0_col_out_832;
wire [151:0] u0_col_out_833;
wire [151:0] u0_col_out_834;
wire [151:0] u0_col_out_835;
wire [151:0] u0_col_out_836;
wire [151:0] u0_col_out_837;
wire [151:0] u0_col_out_838;
wire [151:0] u0_col_out_839;
wire [151:0] u0_col_out_840;
wire [151:0] u0_col_out_841;
wire [151:0] u0_col_out_842;
wire [151:0] u0_col_out_843;
wire [151:0] u0_col_out_844;
wire [151:0] u0_col_out_845;
wire [151:0] u0_col_out_846;
wire [151:0] u0_col_out_847;
wire [151:0] u0_col_out_848;
wire [151:0] u0_col_out_849;
wire [151:0] u0_col_out_850;
wire [151:0] u0_col_out_851;
wire [151:0] u0_col_out_852;
wire [151:0] u0_col_out_853;
wire [151:0] u0_col_out_854;
wire [151:0] u0_col_out_855;
wire [151:0] u0_col_out_856;
wire [151:0] u0_col_out_857;
wire [151:0] u0_col_out_858;
wire [151:0] u0_col_out_859;
wire [151:0] u0_col_out_860;
wire [151:0] u0_col_out_861;
wire [151:0] u0_col_out_862;
wire [151:0] u0_col_out_863;
wire [151:0] u0_col_out_864;
wire [151:0] u0_col_out_865;
wire [151:0] u0_col_out_866;
wire [151:0] u0_col_out_867;
wire [151:0] u0_col_out_868;
wire [151:0] u0_col_out_869;
wire [151:0] u0_col_out_870;
wire [151:0] u0_col_out_871;
wire [151:0] u0_col_out_872;
wire [151:0] u0_col_out_873;
wire [151:0] u0_col_out_874;
wire [151:0] u0_col_out_875;
wire [151:0] u0_col_out_876;
wire [151:0] u0_col_out_877;
wire [151:0] u0_col_out_878;
wire [151:0] u0_col_out_879;
wire [151:0] u0_col_out_880;
wire [151:0] u0_col_out_881;
wire [151:0] u0_col_out_882;
wire [151:0] u0_col_out_883;
wire [151:0] u0_col_out_884;
wire [151:0] u0_col_out_885;
wire [151:0] u0_col_out_886;
wire [151:0] u0_col_out_887;
wire [151:0] u0_col_out_888;
wire [151:0] u0_col_out_889;
wire [151:0] u0_col_out_890;
wire [151:0] u0_col_out_891;
wire [151:0] u0_col_out_892;
wire [151:0] u0_col_out_893;
wire [151:0] u0_col_out_894;
wire [151:0] u0_col_out_895;
wire [151:0] u0_col_out_896;
wire [151:0] u0_col_out_897;
wire [151:0] u0_col_out_898;
wire [151:0] u0_col_out_899;
wire [151:0] u0_col_out_900;
wire [151:0] u0_col_out_901;
wire [151:0] u0_col_out_902;
wire [151:0] u0_col_out_903;
wire [151:0] u0_col_out_904;
wire [151:0] u0_col_out_905;
wire [151:0] u0_col_out_906;
wire [151:0] u0_col_out_907;
wire [151:0] u0_col_out_908;
wire [151:0] u0_col_out_909;
wire [151:0] u0_col_out_910;
wire [151:0] u0_col_out_911;
wire [151:0] u0_col_out_912;
wire [151:0] u0_col_out_913;
wire [151:0] u0_col_out_914;
wire [151:0] u0_col_out_915;
wire [151:0] u0_col_out_916;
wire [151:0] u0_col_out_917;
wire [151:0] u0_col_out_918;
wire [151:0] u0_col_out_919;
wire [151:0] u0_col_out_920;
wire [151:0] u0_col_out_921;
wire [151:0] u0_col_out_922;
wire [151:0] u0_col_out_923;
wire [151:0] u0_col_out_924;
wire [151:0] u0_col_out_925;
wire [151:0] u0_col_out_926;
wire [151:0] u0_col_out_927;
wire [151:0] u0_col_out_928;
wire [151:0] u0_col_out_929;
wire [151:0] u0_col_out_930;
wire [151:0] u0_col_out_931;
wire [151:0] u0_col_out_932;
wire [151:0] u0_col_out_933;
wire [151:0] u0_col_out_934;
wire [151:0] u0_col_out_935;
wire [151:0] u0_col_out_936;
wire [151:0] u0_col_out_937;
wire [151:0] u0_col_out_938;
wire [151:0] u0_col_out_939;
wire [151:0] u0_col_out_940;
wire [151:0] u0_col_out_941;
wire [151:0] u0_col_out_942;
wire [151:0] u0_col_out_943;
wire [151:0] u0_col_out_944;
wire [151:0] u0_col_out_945;
wire [151:0] u0_col_out_946;
wire [151:0] u0_col_out_947;
wire [151:0] u0_col_out_948;
wire [151:0] u0_col_out_949;
wire [151:0] u0_col_out_950;
wire [151:0] u0_col_out_951;
wire [151:0] u0_col_out_952;
wire [151:0] u0_col_out_953;
wire [151:0] u0_col_out_954;
wire [151:0] u0_col_out_955;
wire [151:0] u0_col_out_956;
wire [151:0] u0_col_out_957;
wire [151:0] u0_col_out_958;
wire [151:0] u0_col_out_959;
wire [151:0] u0_col_out_960;
wire [151:0] u0_col_out_961;
wire [151:0] u0_col_out_962;
wire [151:0] u0_col_out_963;
wire [151:0] u0_col_out_964;
wire [151:0] u0_col_out_965;
wire [151:0] u0_col_out_966;
wire [151:0] u0_col_out_967;
wire [151:0] u0_col_out_968;
wire [151:0] u0_col_out_969;
wire [151:0] u0_col_out_970;
wire [151:0] u0_col_out_971;
wire [151:0] u0_col_out_972;
wire [151:0] u0_col_out_973;
wire [151:0] u0_col_out_974;
wire [151:0] u0_col_out_975;
wire [151:0] u0_col_out_976;
wire [151:0] u0_col_out_977;
wire [151:0] u0_col_out_978;
wire [151:0] u0_col_out_979;
wire [151:0] u0_col_out_980;
wire [151:0] u0_col_out_981;
wire [151:0] u0_col_out_982;
wire [151:0] u0_col_out_983;
wire [151:0] u0_col_out_984;
wire [151:0] u0_col_out_985;
wire [151:0] u0_col_out_986;
wire [151:0] u0_col_out_987;
wire [151:0] u0_col_out_988;
wire [151:0] u0_col_out_989;
wire [151:0] u0_col_out_990;
wire [151:0] u0_col_out_991;
wire [151:0] u0_col_out_992;
wire [151:0] u0_col_out_993;
wire [151:0] u0_col_out_994;
wire [151:0] u0_col_out_995;
wire [151:0] u0_col_out_996;
wire [151:0] u0_col_out_997;
wire [151:0] u0_col_out_998;
wire [151:0] u0_col_out_999;
wire [151:0] u0_col_out_1000;
wire [151:0] u0_col_out_1001;
wire [151:0] u0_col_out_1002;
wire [151:0] u0_col_out_1003;
wire [151:0] u0_col_out_1004;
wire [151:0] u0_col_out_1005;
wire [151:0] u0_col_out_1006;
wire [151:0] u0_col_out_1007;
wire [151:0] u0_col_out_1008;
wire [151:0] u0_col_out_1009;
wire [151:0] u0_col_out_1010;
wire [151:0] u0_col_out_1011;
wire [151:0] u0_col_out_1012;
wire [151:0] u0_col_out_1013;
wire [151:0] u0_col_out_1014;
wire [151:0] u0_col_out_1015;
wire [151:0] u0_col_out_1016;
wire [151:0] u0_col_out_1017;
wire [151:0] u0_col_out_1018;
wire [151:0] u0_col_out_1019;
wire [151:0] u0_col_out_1020;
wire [151:0] u0_col_out_1021;
wire [151:0] u0_col_out_1022;
wire [151:0] u0_col_out_1023;
wire [151:0] u0_col_out_1024;
wire [151:0] u0_col_out_1025;
wire [151:0] u0_col_out_1026;






//*****************************************************
//**************u0输入赋值******************************
//*****************************************************
assign u0_col_in_0 = col_in_0;
assign u0_col_in_1 = col_in_1;
assign u0_col_in_2 = col_in_2;
assign u0_col_in_3 = col_in_3;
assign u0_col_in_4 = col_in_4;
assign u0_col_in_5 = col_in_5;
assign u0_col_in_6 = col_in_6;
assign u0_col_in_7 = col_in_7;
assign u0_col_in_8 = col_in_8;
assign u0_col_in_9 = col_in_9;
assign u0_col_in_10 = col_in_10;
assign u0_col_in_11 = col_in_11;
assign u0_col_in_12 = col_in_12;
assign u0_col_in_13 = col_in_13;
assign u0_col_in_14 = col_in_14;
assign u0_col_in_15 = col_in_15;
assign u0_col_in_16 = col_in_16;
assign u0_col_in_17 = col_in_17;
assign u0_col_in_18 = col_in_18;
assign u0_col_in_19 = col_in_19;
assign u0_col_in_20 = col_in_20;
assign u0_col_in_21 = col_in_21;
assign u0_col_in_22 = col_in_22;
assign u0_col_in_23 = col_in_23;
assign u0_col_in_24 = col_in_24;
assign u0_col_in_25 = col_in_25;
assign u0_col_in_26 = col_in_26;
assign u0_col_in_27 = col_in_27;
assign u0_col_in_28 = col_in_28;
assign u0_col_in_29 = col_in_29;
assign u0_col_in_30 = col_in_30;
assign u0_col_in_31 = col_in_31;
assign u0_col_in_32 = col_in_32;
assign u0_col_in_33 = col_in_33;
assign u0_col_in_34 = col_in_34;
assign u0_col_in_35 = col_in_35;
assign u0_col_in_36 = col_in_36;
assign u0_col_in_37 = col_in_37;
assign u0_col_in_38 = col_in_38;
assign u0_col_in_39 = col_in_39;
assign u0_col_in_40 = col_in_40;
assign u0_col_in_41 = col_in_41;
assign u0_col_in_42 = col_in_42;
assign u0_col_in_43 = col_in_43;
assign u0_col_in_44 = col_in_44;
assign u0_col_in_45 = col_in_45;
assign u0_col_in_46 = col_in_46;
assign u0_col_in_47 = col_in_47;
assign u0_col_in_48 = col_in_48;
assign u0_col_in_49 = col_in_49;
assign u0_col_in_50 = col_in_50;
assign u0_col_in_51 = col_in_51;
assign u0_col_in_52 = col_in_52;
assign u0_col_in_53 = col_in_53;
assign u0_col_in_54 = col_in_54;
assign u0_col_in_55 = col_in_55;
assign u0_col_in_56 = col_in_56;
assign u0_col_in_57 = col_in_57;
assign u0_col_in_58 = col_in_58;
assign u0_col_in_59 = col_in_59;
assign u0_col_in_60 = col_in_60;
assign u0_col_in_61 = col_in_61;
assign u0_col_in_62 = col_in_62;
assign u0_col_in_63 = col_in_63;
assign u0_col_in_64 = col_in_64;
assign u0_col_in_65 = col_in_65;
assign u0_col_in_66 = col_in_66;
assign u0_col_in_67 = col_in_67;
assign u0_col_in_68 = col_in_68;
assign u0_col_in_69 = col_in_69;
assign u0_col_in_70 = col_in_70;
assign u0_col_in_71 = col_in_71;
assign u0_col_in_72 = col_in_72;
assign u0_col_in_73 = col_in_73;
assign u0_col_in_74 = col_in_74;
assign u0_col_in_75 = col_in_75;
assign u0_col_in_76 = col_in_76;
assign u0_col_in_77 = col_in_77;
assign u0_col_in_78 = col_in_78;
assign u0_col_in_79 = col_in_79;
assign u0_col_in_80 = col_in_80;
assign u0_col_in_81 = col_in_81;
assign u0_col_in_82 = col_in_82;
assign u0_col_in_83 = col_in_83;
assign u0_col_in_84 = col_in_84;
assign u0_col_in_85 = col_in_85;
assign u0_col_in_86 = col_in_86;
assign u0_col_in_87 = col_in_87;
assign u0_col_in_88 = col_in_88;
assign u0_col_in_89 = col_in_89;
assign u0_col_in_90 = col_in_90;
assign u0_col_in_91 = col_in_91;
assign u0_col_in_92 = col_in_92;
assign u0_col_in_93 = col_in_93;
assign u0_col_in_94 = col_in_94;
assign u0_col_in_95 = col_in_95;
assign u0_col_in_96 = col_in_96;
assign u0_col_in_97 = col_in_97;
assign u0_col_in_98 = col_in_98;
assign u0_col_in_99 = col_in_99;
assign u0_col_in_100 = col_in_100;
assign u0_col_in_101 = col_in_101;
assign u0_col_in_102 = col_in_102;
assign u0_col_in_103 = col_in_103;
assign u0_col_in_104 = col_in_104;
assign u0_col_in_105 = col_in_105;
assign u0_col_in_106 = col_in_106;
assign u0_col_in_107 = col_in_107;
assign u0_col_in_108 = col_in_108;
assign u0_col_in_109 = col_in_109;
assign u0_col_in_110 = col_in_110;
assign u0_col_in_111 = col_in_111;
assign u0_col_in_112 = col_in_112;
assign u0_col_in_113 = col_in_113;
assign u0_col_in_114 = col_in_114;
assign u0_col_in_115 = col_in_115;
assign u0_col_in_116 = col_in_116;
assign u0_col_in_117 = col_in_117;
assign u0_col_in_118 = col_in_118;
assign u0_col_in_119 = col_in_119;
assign u0_col_in_120 = col_in_120;
assign u0_col_in_121 = col_in_121;
assign u0_col_in_122 = col_in_122;
assign u0_col_in_123 = col_in_123;
assign u0_col_in_124 = col_in_124;
assign u0_col_in_125 = col_in_125;
assign u0_col_in_126 = col_in_126;
assign u0_col_in_127 = col_in_127;
assign u0_col_in_128 = col_in_128;
assign u0_col_in_129 = col_in_129;
assign u0_col_in_130 = col_in_130;
assign u0_col_in_131 = col_in_131;
assign u0_col_in_132 = col_in_132;
assign u0_col_in_133 = col_in_133;
assign u0_col_in_134 = col_in_134;
assign u0_col_in_135 = col_in_135;
assign u0_col_in_136 = col_in_136;
assign u0_col_in_137 = col_in_137;
assign u0_col_in_138 = col_in_138;
assign u0_col_in_139 = col_in_139;
assign u0_col_in_140 = col_in_140;
assign u0_col_in_141 = col_in_141;
assign u0_col_in_142 = col_in_142;
assign u0_col_in_143 = col_in_143;
assign u0_col_in_144 = col_in_144;
assign u0_col_in_145 = col_in_145;
assign u0_col_in_146 = col_in_146;
assign u0_col_in_147 = col_in_147;
assign u0_col_in_148 = col_in_148;
assign u0_col_in_149 = col_in_149;
assign u0_col_in_150 = col_in_150;
assign u0_col_in_151 = col_in_151;
assign u0_col_in_152 = col_in_152;
assign u0_col_in_153 = col_in_153;
assign u0_col_in_154 = col_in_154;
assign u0_col_in_155 = col_in_155;
assign u0_col_in_156 = col_in_156;
assign u0_col_in_157 = col_in_157;
assign u0_col_in_158 = col_in_158;
assign u0_col_in_159 = col_in_159;
assign u0_col_in_160 = col_in_160;
assign u0_col_in_161 = col_in_161;
assign u0_col_in_162 = col_in_162;
assign u0_col_in_163 = col_in_163;
assign u0_col_in_164 = col_in_164;
assign u0_col_in_165 = col_in_165;
assign u0_col_in_166 = col_in_166;
assign u0_col_in_167 = col_in_167;
assign u0_col_in_168 = col_in_168;
assign u0_col_in_169 = col_in_169;
assign u0_col_in_170 = col_in_170;
assign u0_col_in_171 = col_in_171;
assign u0_col_in_172 = col_in_172;
assign u0_col_in_173 = col_in_173;
assign u0_col_in_174 = col_in_174;
assign u0_col_in_175 = col_in_175;
assign u0_col_in_176 = col_in_176;
assign u0_col_in_177 = col_in_177;
assign u0_col_in_178 = col_in_178;
assign u0_col_in_179 = col_in_179;
assign u0_col_in_180 = col_in_180;
assign u0_col_in_181 = col_in_181;
assign u0_col_in_182 = col_in_182;
assign u0_col_in_183 = col_in_183;
assign u0_col_in_184 = col_in_184;
assign u0_col_in_185 = col_in_185;
assign u0_col_in_186 = col_in_186;
assign u0_col_in_187 = col_in_187;
assign u0_col_in_188 = col_in_188;
assign u0_col_in_189 = col_in_189;
assign u0_col_in_190 = col_in_190;
assign u0_col_in_191 = col_in_191;
assign u0_col_in_192 = col_in_192;
assign u0_col_in_193 = col_in_193;
assign u0_col_in_194 = col_in_194;
assign u0_col_in_195 = col_in_195;
assign u0_col_in_196 = col_in_196;
assign u0_col_in_197 = col_in_197;
assign u0_col_in_198 = col_in_198;
assign u0_col_in_199 = col_in_199;
assign u0_col_in_200 = col_in_200;
assign u0_col_in_201 = col_in_201;
assign u0_col_in_202 = col_in_202;
assign u0_col_in_203 = col_in_203;
assign u0_col_in_204 = col_in_204;
assign u0_col_in_205 = col_in_205;
assign u0_col_in_206 = col_in_206;
assign u0_col_in_207 = col_in_207;
assign u0_col_in_208 = col_in_208;
assign u0_col_in_209 = col_in_209;
assign u0_col_in_210 = col_in_210;
assign u0_col_in_211 = col_in_211;
assign u0_col_in_212 = col_in_212;
assign u0_col_in_213 = col_in_213;
assign u0_col_in_214 = col_in_214;
assign u0_col_in_215 = col_in_215;
assign u0_col_in_216 = col_in_216;
assign u0_col_in_217 = col_in_217;
assign u0_col_in_218 = col_in_218;
assign u0_col_in_219 = col_in_219;
assign u0_col_in_220 = col_in_220;
assign u0_col_in_221 = col_in_221;
assign u0_col_in_222 = col_in_222;
assign u0_col_in_223 = col_in_223;
assign u0_col_in_224 = col_in_224;
assign u0_col_in_225 = col_in_225;
assign u0_col_in_226 = col_in_226;
assign u0_col_in_227 = col_in_227;
assign u0_col_in_228 = col_in_228;
assign u0_col_in_229 = col_in_229;
assign u0_col_in_230 = col_in_230;
assign u0_col_in_231 = col_in_231;
assign u0_col_in_232 = col_in_232;
assign u0_col_in_233 = col_in_233;
assign u0_col_in_234 = col_in_234;
assign u0_col_in_235 = col_in_235;
assign u0_col_in_236 = col_in_236;
assign u0_col_in_237 = col_in_237;
assign u0_col_in_238 = col_in_238;
assign u0_col_in_239 = col_in_239;
assign u0_col_in_240 = col_in_240;
assign u0_col_in_241 = col_in_241;
assign u0_col_in_242 = col_in_242;
assign u0_col_in_243 = col_in_243;
assign u0_col_in_244 = col_in_244;
assign u0_col_in_245 = col_in_245;
assign u0_col_in_246 = col_in_246;
assign u0_col_in_247 = col_in_247;
assign u0_col_in_248 = col_in_248;
assign u0_col_in_249 = col_in_249;
assign u0_col_in_250 = col_in_250;
assign u0_col_in_251 = col_in_251;
assign u0_col_in_252 = col_in_252;
assign u0_col_in_253 = col_in_253;
assign u0_col_in_254 = col_in_254;
assign u0_col_in_255 = col_in_255;
assign u0_col_in_256 = col_in_256;
assign u0_col_in_257 = col_in_257;
assign u0_col_in_258 = col_in_258;
assign u0_col_in_259 = col_in_259;
assign u0_col_in_260 = col_in_260;
assign u0_col_in_261 = col_in_261;
assign u0_col_in_262 = col_in_262;
assign u0_col_in_263 = col_in_263;
assign u0_col_in_264 = col_in_264;
assign u0_col_in_265 = col_in_265;
assign u0_col_in_266 = col_in_266;
assign u0_col_in_267 = col_in_267;
assign u0_col_in_268 = col_in_268;
assign u0_col_in_269 = col_in_269;
assign u0_col_in_270 = col_in_270;
assign u0_col_in_271 = col_in_271;
assign u0_col_in_272 = col_in_272;
assign u0_col_in_273 = col_in_273;
assign u0_col_in_274 = col_in_274;
assign u0_col_in_275 = col_in_275;
assign u0_col_in_276 = col_in_276;
assign u0_col_in_277 = col_in_277;
assign u0_col_in_278 = col_in_278;
assign u0_col_in_279 = col_in_279;
assign u0_col_in_280 = col_in_280;
assign u0_col_in_281 = col_in_281;
assign u0_col_in_282 = col_in_282;
assign u0_col_in_283 = col_in_283;
assign u0_col_in_284 = col_in_284;
assign u0_col_in_285 = col_in_285;
assign u0_col_in_286 = col_in_286;
assign u0_col_in_287 = col_in_287;
assign u0_col_in_288 = col_in_288;
assign u0_col_in_289 = col_in_289;
assign u0_col_in_290 = col_in_290;
assign u0_col_in_291 = col_in_291;
assign u0_col_in_292 = col_in_292;
assign u0_col_in_293 = col_in_293;
assign u0_col_in_294 = col_in_294;
assign u0_col_in_295 = col_in_295;
assign u0_col_in_296 = col_in_296;
assign u0_col_in_297 = col_in_297;
assign u0_col_in_298 = col_in_298;
assign u0_col_in_299 = col_in_299;
assign u0_col_in_300 = col_in_300;
assign u0_col_in_301 = col_in_301;
assign u0_col_in_302 = col_in_302;
assign u0_col_in_303 = col_in_303;
assign u0_col_in_304 = col_in_304;
assign u0_col_in_305 = col_in_305;
assign u0_col_in_306 = col_in_306;
assign u0_col_in_307 = col_in_307;
assign u0_col_in_308 = col_in_308;
assign u0_col_in_309 = col_in_309;
assign u0_col_in_310 = col_in_310;
assign u0_col_in_311 = col_in_311;
assign u0_col_in_312 = col_in_312;
assign u0_col_in_313 = col_in_313;
assign u0_col_in_314 = col_in_314;
assign u0_col_in_315 = col_in_315;
assign u0_col_in_316 = col_in_316;
assign u0_col_in_317 = col_in_317;
assign u0_col_in_318 = col_in_318;
assign u0_col_in_319 = col_in_319;
assign u0_col_in_320 = col_in_320;
assign u0_col_in_321 = col_in_321;
assign u0_col_in_322 = col_in_322;
assign u0_col_in_323 = col_in_323;
assign u0_col_in_324 = col_in_324;
assign u0_col_in_325 = col_in_325;
assign u0_col_in_326 = col_in_326;
assign u0_col_in_327 = col_in_327;
assign u0_col_in_328 = col_in_328;
assign u0_col_in_329 = col_in_329;
assign u0_col_in_330 = col_in_330;
assign u0_col_in_331 = col_in_331;
assign u0_col_in_332 = col_in_332;
assign u0_col_in_333 = col_in_333;
assign u0_col_in_334 = col_in_334;
assign u0_col_in_335 = col_in_335;
assign u0_col_in_336 = col_in_336;
assign u0_col_in_337 = col_in_337;
assign u0_col_in_338 = col_in_338;
assign u0_col_in_339 = col_in_339;
assign u0_col_in_340 = col_in_340;
assign u0_col_in_341 = col_in_341;
assign u0_col_in_342 = col_in_342;
assign u0_col_in_343 = col_in_343;
assign u0_col_in_344 = col_in_344;
assign u0_col_in_345 = col_in_345;
assign u0_col_in_346 = col_in_346;
assign u0_col_in_347 = col_in_347;
assign u0_col_in_348 = col_in_348;
assign u0_col_in_349 = col_in_349;
assign u0_col_in_350 = col_in_350;
assign u0_col_in_351 = col_in_351;
assign u0_col_in_352 = col_in_352;
assign u0_col_in_353 = col_in_353;
assign u0_col_in_354 = col_in_354;
assign u0_col_in_355 = col_in_355;
assign u0_col_in_356 = col_in_356;
assign u0_col_in_357 = col_in_357;
assign u0_col_in_358 = col_in_358;
assign u0_col_in_359 = col_in_359;
assign u0_col_in_360 = col_in_360;
assign u0_col_in_361 = col_in_361;
assign u0_col_in_362 = col_in_362;
assign u0_col_in_363 = col_in_363;
assign u0_col_in_364 = col_in_364;
assign u0_col_in_365 = col_in_365;
assign u0_col_in_366 = col_in_366;
assign u0_col_in_367 = col_in_367;
assign u0_col_in_368 = col_in_368;
assign u0_col_in_369 = col_in_369;
assign u0_col_in_370 = col_in_370;
assign u0_col_in_371 = col_in_371;
assign u0_col_in_372 = col_in_372;
assign u0_col_in_373 = col_in_373;
assign u0_col_in_374 = col_in_374;
assign u0_col_in_375 = col_in_375;
assign u0_col_in_376 = col_in_376;
assign u0_col_in_377 = col_in_377;
assign u0_col_in_378 = col_in_378;
assign u0_col_in_379 = col_in_379;
assign u0_col_in_380 = col_in_380;
assign u0_col_in_381 = col_in_381;
assign u0_col_in_382 = col_in_382;
assign u0_col_in_383 = col_in_383;
assign u0_col_in_384 = col_in_384;
assign u0_col_in_385 = col_in_385;
assign u0_col_in_386 = col_in_386;
assign u0_col_in_387 = col_in_387;
assign u0_col_in_388 = col_in_388;
assign u0_col_in_389 = col_in_389;
assign u0_col_in_390 = col_in_390;
assign u0_col_in_391 = col_in_391;
assign u0_col_in_392 = col_in_392;
assign u0_col_in_393 = col_in_393;
assign u0_col_in_394 = col_in_394;
assign u0_col_in_395 = col_in_395;
assign u0_col_in_396 = col_in_396;
assign u0_col_in_397 = col_in_397;
assign u0_col_in_398 = col_in_398;
assign u0_col_in_399 = col_in_399;
assign u0_col_in_400 = col_in_400;
assign u0_col_in_401 = col_in_401;
assign u0_col_in_402 = col_in_402;
assign u0_col_in_403 = col_in_403;
assign u0_col_in_404 = col_in_404;
assign u0_col_in_405 = col_in_405;
assign u0_col_in_406 = col_in_406;
assign u0_col_in_407 = col_in_407;
assign u0_col_in_408 = col_in_408;
assign u0_col_in_409 = col_in_409;
assign u0_col_in_410 = col_in_410;
assign u0_col_in_411 = col_in_411;
assign u0_col_in_412 = col_in_412;
assign u0_col_in_413 = col_in_413;
assign u0_col_in_414 = col_in_414;
assign u0_col_in_415 = col_in_415;
assign u0_col_in_416 = col_in_416;
assign u0_col_in_417 = col_in_417;
assign u0_col_in_418 = col_in_418;
assign u0_col_in_419 = col_in_419;
assign u0_col_in_420 = col_in_420;
assign u0_col_in_421 = col_in_421;
assign u0_col_in_422 = col_in_422;
assign u0_col_in_423 = col_in_423;
assign u0_col_in_424 = col_in_424;
assign u0_col_in_425 = col_in_425;
assign u0_col_in_426 = col_in_426;
assign u0_col_in_427 = col_in_427;
assign u0_col_in_428 = col_in_428;
assign u0_col_in_429 = col_in_429;
assign u0_col_in_430 = col_in_430;
assign u0_col_in_431 = col_in_431;
assign u0_col_in_432 = col_in_432;
assign u0_col_in_433 = col_in_433;
assign u0_col_in_434 = col_in_434;
assign u0_col_in_435 = col_in_435;
assign u0_col_in_436 = col_in_436;
assign u0_col_in_437 = col_in_437;
assign u0_col_in_438 = col_in_438;
assign u0_col_in_439 = col_in_439;
assign u0_col_in_440 = col_in_440;
assign u0_col_in_441 = col_in_441;
assign u0_col_in_442 = col_in_442;
assign u0_col_in_443 = col_in_443;
assign u0_col_in_444 = col_in_444;
assign u0_col_in_445 = col_in_445;
assign u0_col_in_446 = col_in_446;
assign u0_col_in_447 = col_in_447;
assign u0_col_in_448 = col_in_448;
assign u0_col_in_449 = col_in_449;
assign u0_col_in_450 = col_in_450;
assign u0_col_in_451 = col_in_451;
assign u0_col_in_452 = col_in_452;
assign u0_col_in_453 = col_in_453;
assign u0_col_in_454 = col_in_454;
assign u0_col_in_455 = col_in_455;
assign u0_col_in_456 = col_in_456;
assign u0_col_in_457 = col_in_457;
assign u0_col_in_458 = col_in_458;
assign u0_col_in_459 = col_in_459;
assign u0_col_in_460 = col_in_460;
assign u0_col_in_461 = col_in_461;
assign u0_col_in_462 = col_in_462;
assign u0_col_in_463 = col_in_463;
assign u0_col_in_464 = col_in_464;
assign u0_col_in_465 = col_in_465;
assign u0_col_in_466 = col_in_466;
assign u0_col_in_467 = col_in_467;
assign u0_col_in_468 = col_in_468;
assign u0_col_in_469 = col_in_469;
assign u0_col_in_470 = col_in_470;
assign u0_col_in_471 = col_in_471;
assign u0_col_in_472 = col_in_472;
assign u0_col_in_473 = col_in_473;
assign u0_col_in_474 = col_in_474;
assign u0_col_in_475 = col_in_475;
assign u0_col_in_476 = col_in_476;
assign u0_col_in_477 = col_in_477;
assign u0_col_in_478 = col_in_478;
assign u0_col_in_479 = col_in_479;
assign u0_col_in_480 = col_in_480;
assign u0_col_in_481 = col_in_481;
assign u0_col_in_482 = col_in_482;
assign u0_col_in_483 = col_in_483;
assign u0_col_in_484 = col_in_484;
assign u0_col_in_485 = col_in_485;
assign u0_col_in_486 = col_in_486;
assign u0_col_in_487 = col_in_487;
assign u0_col_in_488 = col_in_488;
assign u0_col_in_489 = col_in_489;
assign u0_col_in_490 = col_in_490;
assign u0_col_in_491 = col_in_491;
assign u0_col_in_492 = col_in_492;
assign u0_col_in_493 = col_in_493;
assign u0_col_in_494 = col_in_494;
assign u0_col_in_495 = col_in_495;
assign u0_col_in_496 = col_in_496;
assign u0_col_in_497 = col_in_497;
assign u0_col_in_498 = col_in_498;
assign u0_col_in_499 = col_in_499;
assign u0_col_in_500 = col_in_500;
assign u0_col_in_501 = col_in_501;
assign u0_col_in_502 = col_in_502;
assign u0_col_in_503 = col_in_503;
assign u0_col_in_504 = col_in_504;
assign u0_col_in_505 = col_in_505;
assign u0_col_in_506 = col_in_506;
assign u0_col_in_507 = col_in_507;
assign u0_col_in_508 = col_in_508;
assign u0_col_in_509 = col_in_509;
assign u0_col_in_510 = col_in_510;
assign u0_col_in_511 = col_in_511;
assign u0_col_in_512 = col_in_512;
assign u0_col_in_513 = col_in_513;
assign u0_col_in_514 = col_in_514;
assign u0_col_in_515 = col_in_515;
assign u0_col_in_516 = col_in_516;
assign u0_col_in_517 = col_in_517;
assign u0_col_in_518 = col_in_518;
assign u0_col_in_519 = col_in_519;
assign u0_col_in_520 = col_in_520;
assign u0_col_in_521 = col_in_521;
assign u0_col_in_522 = col_in_522;
assign u0_col_in_523 = col_in_523;
assign u0_col_in_524 = col_in_524;
assign u0_col_in_525 = col_in_525;
assign u0_col_in_526 = col_in_526;
assign u0_col_in_527 = col_in_527;
assign u0_col_in_528 = col_in_528;
assign u0_col_in_529 = col_in_529;
assign u0_col_in_530 = col_in_530;
assign u0_col_in_531 = col_in_531;
assign u0_col_in_532 = col_in_532;
assign u0_col_in_533 = col_in_533;
assign u0_col_in_534 = col_in_534;
assign u0_col_in_535 = col_in_535;
assign u0_col_in_536 = col_in_536;
assign u0_col_in_537 = col_in_537;
assign u0_col_in_538 = col_in_538;
assign u0_col_in_539 = col_in_539;
assign u0_col_in_540 = col_in_540;
assign u0_col_in_541 = col_in_541;
assign u0_col_in_542 = col_in_542;
assign u0_col_in_543 = col_in_543;
assign u0_col_in_544 = col_in_544;
assign u0_col_in_545 = col_in_545;
assign u0_col_in_546 = col_in_546;
assign u0_col_in_547 = col_in_547;
assign u0_col_in_548 = col_in_548;
assign u0_col_in_549 = col_in_549;
assign u0_col_in_550 = col_in_550;
assign u0_col_in_551 = col_in_551;
assign u0_col_in_552 = col_in_552;
assign u0_col_in_553 = col_in_553;
assign u0_col_in_554 = col_in_554;
assign u0_col_in_555 = col_in_555;
assign u0_col_in_556 = col_in_556;
assign u0_col_in_557 = col_in_557;
assign u0_col_in_558 = col_in_558;
assign u0_col_in_559 = col_in_559;
assign u0_col_in_560 = col_in_560;
assign u0_col_in_561 = col_in_561;
assign u0_col_in_562 = col_in_562;
assign u0_col_in_563 = col_in_563;
assign u0_col_in_564 = col_in_564;
assign u0_col_in_565 = col_in_565;
assign u0_col_in_566 = col_in_566;
assign u0_col_in_567 = col_in_567;
assign u0_col_in_568 = col_in_568;
assign u0_col_in_569 = col_in_569;
assign u0_col_in_570 = col_in_570;
assign u0_col_in_571 = col_in_571;
assign u0_col_in_572 = col_in_572;
assign u0_col_in_573 = col_in_573;
assign u0_col_in_574 = col_in_574;
assign u0_col_in_575 = col_in_575;
assign u0_col_in_576 = col_in_576;
assign u0_col_in_577 = col_in_577;
assign u0_col_in_578 = col_in_578;
assign u0_col_in_579 = col_in_579;
assign u0_col_in_580 = col_in_580;
assign u0_col_in_581 = col_in_581;
assign u0_col_in_582 = col_in_582;
assign u0_col_in_583 = col_in_583;
assign u0_col_in_584 = col_in_584;
assign u0_col_in_585 = col_in_585;
assign u0_col_in_586 = col_in_586;
assign u0_col_in_587 = col_in_587;
assign u0_col_in_588 = col_in_588;
assign u0_col_in_589 = col_in_589;
assign u0_col_in_590 = col_in_590;
assign u0_col_in_591 = col_in_591;
assign u0_col_in_592 = col_in_592;
assign u0_col_in_593 = col_in_593;
assign u0_col_in_594 = col_in_594;
assign u0_col_in_595 = col_in_595;
assign u0_col_in_596 = col_in_596;
assign u0_col_in_597 = col_in_597;
assign u0_col_in_598 = col_in_598;
assign u0_col_in_599 = col_in_599;
assign u0_col_in_600 = col_in_600;
assign u0_col_in_601 = col_in_601;
assign u0_col_in_602 = col_in_602;
assign u0_col_in_603 = col_in_603;
assign u0_col_in_604 = col_in_604;
assign u0_col_in_605 = col_in_605;
assign u0_col_in_606 = col_in_606;
assign u0_col_in_607 = col_in_607;
assign u0_col_in_608 = col_in_608;
assign u0_col_in_609 = col_in_609;
assign u0_col_in_610 = col_in_610;
assign u0_col_in_611 = col_in_611;
assign u0_col_in_612 = col_in_612;
assign u0_col_in_613 = col_in_613;
assign u0_col_in_614 = col_in_614;
assign u0_col_in_615 = col_in_615;
assign u0_col_in_616 = col_in_616;
assign u0_col_in_617 = col_in_617;
assign u0_col_in_618 = col_in_618;
assign u0_col_in_619 = col_in_619;
assign u0_col_in_620 = col_in_620;
assign u0_col_in_621 = col_in_621;
assign u0_col_in_622 = col_in_622;
assign u0_col_in_623 = col_in_623;
assign u0_col_in_624 = col_in_624;
assign u0_col_in_625 = col_in_625;
assign u0_col_in_626 = col_in_626;
assign u0_col_in_627 = col_in_627;
assign u0_col_in_628 = col_in_628;
assign u0_col_in_629 = col_in_629;
assign u0_col_in_630 = col_in_630;
assign u0_col_in_631 = col_in_631;
assign u0_col_in_632 = col_in_632;
assign u0_col_in_633 = col_in_633;
assign u0_col_in_634 = col_in_634;
assign u0_col_in_635 = col_in_635;
assign u0_col_in_636 = col_in_636;
assign u0_col_in_637 = col_in_637;
assign u0_col_in_638 = col_in_638;
assign u0_col_in_639 = col_in_639;
assign u0_col_in_640 = col_in_640;
assign u0_col_in_641 = col_in_641;
assign u0_col_in_642 = col_in_642;
assign u0_col_in_643 = col_in_643;
assign u0_col_in_644 = col_in_644;
assign u0_col_in_645 = col_in_645;
assign u0_col_in_646 = col_in_646;
assign u0_col_in_647 = col_in_647;
assign u0_col_in_648 = col_in_648;
assign u0_col_in_649 = col_in_649;
assign u0_col_in_650 = col_in_650;
assign u0_col_in_651 = col_in_651;
assign u0_col_in_652 = col_in_652;
assign u0_col_in_653 = col_in_653;
assign u0_col_in_654 = col_in_654;
assign u0_col_in_655 = col_in_655;
assign u0_col_in_656 = col_in_656;
assign u0_col_in_657 = col_in_657;
assign u0_col_in_658 = col_in_658;
assign u0_col_in_659 = col_in_659;
assign u0_col_in_660 = col_in_660;
assign u0_col_in_661 = col_in_661;
assign u0_col_in_662 = col_in_662;
assign u0_col_in_663 = col_in_663;
assign u0_col_in_664 = col_in_664;
assign u0_col_in_665 = col_in_665;
assign u0_col_in_666 = col_in_666;
assign u0_col_in_667 = col_in_667;
assign u0_col_in_668 = col_in_668;
assign u0_col_in_669 = col_in_669;
assign u0_col_in_670 = col_in_670;
assign u0_col_in_671 = col_in_671;
assign u0_col_in_672 = col_in_672;
assign u0_col_in_673 = col_in_673;
assign u0_col_in_674 = col_in_674;
assign u0_col_in_675 = col_in_675;
assign u0_col_in_676 = col_in_676;
assign u0_col_in_677 = col_in_677;
assign u0_col_in_678 = col_in_678;
assign u0_col_in_679 = col_in_679;
assign u0_col_in_680 = col_in_680;
assign u0_col_in_681 = col_in_681;
assign u0_col_in_682 = col_in_682;
assign u0_col_in_683 = col_in_683;
assign u0_col_in_684 = col_in_684;
assign u0_col_in_685 = col_in_685;
assign u0_col_in_686 = col_in_686;
assign u0_col_in_687 = col_in_687;
assign u0_col_in_688 = col_in_688;
assign u0_col_in_689 = col_in_689;
assign u0_col_in_690 = col_in_690;
assign u0_col_in_691 = col_in_691;
assign u0_col_in_692 = col_in_692;
assign u0_col_in_693 = col_in_693;
assign u0_col_in_694 = col_in_694;
assign u0_col_in_695 = col_in_695;
assign u0_col_in_696 = col_in_696;
assign u0_col_in_697 = col_in_697;
assign u0_col_in_698 = col_in_698;
assign u0_col_in_699 = col_in_699;
assign u0_col_in_700 = col_in_700;
assign u0_col_in_701 = col_in_701;
assign u0_col_in_702 = col_in_702;
assign u0_col_in_703 = col_in_703;
assign u0_col_in_704 = col_in_704;
assign u0_col_in_705 = col_in_705;
assign u0_col_in_706 = col_in_706;
assign u0_col_in_707 = col_in_707;
assign u0_col_in_708 = col_in_708;
assign u0_col_in_709 = col_in_709;
assign u0_col_in_710 = col_in_710;
assign u0_col_in_711 = col_in_711;
assign u0_col_in_712 = col_in_712;
assign u0_col_in_713 = col_in_713;
assign u0_col_in_714 = col_in_714;
assign u0_col_in_715 = col_in_715;
assign u0_col_in_716 = col_in_716;
assign u0_col_in_717 = col_in_717;
assign u0_col_in_718 = col_in_718;
assign u0_col_in_719 = col_in_719;
assign u0_col_in_720 = col_in_720;
assign u0_col_in_721 = col_in_721;
assign u0_col_in_722 = col_in_722;
assign u0_col_in_723 = col_in_723;
assign u0_col_in_724 = col_in_724;
assign u0_col_in_725 = col_in_725;
assign u0_col_in_726 = col_in_726;
assign u0_col_in_727 = col_in_727;
assign u0_col_in_728 = col_in_728;
assign u0_col_in_729 = col_in_729;
assign u0_col_in_730 = col_in_730;
assign u0_col_in_731 = col_in_731;
assign u0_col_in_732 = col_in_732;
assign u0_col_in_733 = col_in_733;
assign u0_col_in_734 = col_in_734;
assign u0_col_in_735 = col_in_735;
assign u0_col_in_736 = col_in_736;
assign u0_col_in_737 = col_in_737;
assign u0_col_in_738 = col_in_738;
assign u0_col_in_739 = col_in_739;
assign u0_col_in_740 = col_in_740;
assign u0_col_in_741 = col_in_741;
assign u0_col_in_742 = col_in_742;
assign u0_col_in_743 = col_in_743;
assign u0_col_in_744 = col_in_744;
assign u0_col_in_745 = col_in_745;
assign u0_col_in_746 = col_in_746;
assign u0_col_in_747 = col_in_747;
assign u0_col_in_748 = col_in_748;
assign u0_col_in_749 = col_in_749;
assign u0_col_in_750 = col_in_750;
assign u0_col_in_751 = col_in_751;
assign u0_col_in_752 = col_in_752;
assign u0_col_in_753 = col_in_753;
assign u0_col_in_754 = col_in_754;
assign u0_col_in_755 = col_in_755;
assign u0_col_in_756 = col_in_756;
assign u0_col_in_757 = col_in_757;
assign u0_col_in_758 = col_in_758;
assign u0_col_in_759 = col_in_759;
assign u0_col_in_760 = col_in_760;
assign u0_col_in_761 = col_in_761;
assign u0_col_in_762 = col_in_762;
assign u0_col_in_763 = col_in_763;
assign u0_col_in_764 = col_in_764;
assign u0_col_in_765 = col_in_765;
assign u0_col_in_766 = col_in_766;
assign u0_col_in_767 = col_in_767;
assign u0_col_in_768 = col_in_768;
assign u0_col_in_769 = col_in_769;
assign u0_col_in_770 = col_in_770;
assign u0_col_in_771 = col_in_771;
assign u0_col_in_772 = col_in_772;
assign u0_col_in_773 = col_in_773;
assign u0_col_in_774 = col_in_774;
assign u0_col_in_775 = col_in_775;
assign u0_col_in_776 = col_in_776;
assign u0_col_in_777 = col_in_777;
assign u0_col_in_778 = col_in_778;
assign u0_col_in_779 = col_in_779;
assign u0_col_in_780 = col_in_780;
assign u0_col_in_781 = col_in_781;
assign u0_col_in_782 = col_in_782;
assign u0_col_in_783 = col_in_783;
assign u0_col_in_784 = col_in_784;
assign u0_col_in_785 = col_in_785;
assign u0_col_in_786 = col_in_786;
assign u0_col_in_787 = col_in_787;
assign u0_col_in_788 = col_in_788;
assign u0_col_in_789 = col_in_789;
assign u0_col_in_790 = col_in_790;
assign u0_col_in_791 = col_in_791;
assign u0_col_in_792 = col_in_792;
assign u0_col_in_793 = col_in_793;
assign u0_col_in_794 = col_in_794;
assign u0_col_in_795 = col_in_795;
assign u0_col_in_796 = col_in_796;
assign u0_col_in_797 = col_in_797;
assign u0_col_in_798 = col_in_798;
assign u0_col_in_799 = col_in_799;
assign u0_col_in_800 = col_in_800;
assign u0_col_in_801 = col_in_801;
assign u0_col_in_802 = col_in_802;
assign u0_col_in_803 = col_in_803;
assign u0_col_in_804 = col_in_804;
assign u0_col_in_805 = col_in_805;
assign u0_col_in_806 = col_in_806;
assign u0_col_in_807 = col_in_807;
assign u0_col_in_808 = col_in_808;
assign u0_col_in_809 = col_in_809;
assign u0_col_in_810 = col_in_810;
assign u0_col_in_811 = col_in_811;
assign u0_col_in_812 = col_in_812;
assign u0_col_in_813 = col_in_813;
assign u0_col_in_814 = col_in_814;
assign u0_col_in_815 = col_in_815;
assign u0_col_in_816 = col_in_816;
assign u0_col_in_817 = col_in_817;
assign u0_col_in_818 = col_in_818;
assign u0_col_in_819 = col_in_819;
assign u0_col_in_820 = col_in_820;
assign u0_col_in_821 = col_in_821;
assign u0_col_in_822 = col_in_822;
assign u0_col_in_823 = col_in_823;
assign u0_col_in_824 = col_in_824;
assign u0_col_in_825 = col_in_825;
assign u0_col_in_826 = col_in_826;
assign u0_col_in_827 = col_in_827;
assign u0_col_in_828 = col_in_828;
assign u0_col_in_829 = col_in_829;
assign u0_col_in_830 = col_in_830;
assign u0_col_in_831 = col_in_831;
assign u0_col_in_832 = col_in_832;
assign u0_col_in_833 = col_in_833;
assign u0_col_in_834 = col_in_834;
assign u0_col_in_835 = col_in_835;
assign u0_col_in_836 = col_in_836;
assign u0_col_in_837 = col_in_837;
assign u0_col_in_838 = col_in_838;
assign u0_col_in_839 = col_in_839;
assign u0_col_in_840 = col_in_840;
assign u0_col_in_841 = col_in_841;
assign u0_col_in_842 = col_in_842;
assign u0_col_in_843 = col_in_843;
assign u0_col_in_844 = col_in_844;
assign u0_col_in_845 = col_in_845;
assign u0_col_in_846 = col_in_846;
assign u0_col_in_847 = col_in_847;
assign u0_col_in_848 = col_in_848;
assign u0_col_in_849 = col_in_849;
assign u0_col_in_850 = col_in_850;
assign u0_col_in_851 = col_in_851;
assign u0_col_in_852 = col_in_852;
assign u0_col_in_853 = col_in_853;
assign u0_col_in_854 = col_in_854;
assign u0_col_in_855 = col_in_855;
assign u0_col_in_856 = col_in_856;
assign u0_col_in_857 = col_in_857;
assign u0_col_in_858 = col_in_858;
assign u0_col_in_859 = col_in_859;
assign u0_col_in_860 = col_in_860;
assign u0_col_in_861 = col_in_861;
assign u0_col_in_862 = col_in_862;
assign u0_col_in_863 = col_in_863;
assign u0_col_in_864 = col_in_864;
assign u0_col_in_865 = col_in_865;
assign u0_col_in_866 = col_in_866;
assign u0_col_in_867 = col_in_867;
assign u0_col_in_868 = col_in_868;
assign u0_col_in_869 = col_in_869;
assign u0_col_in_870 = col_in_870;
assign u0_col_in_871 = col_in_871;
assign u0_col_in_872 = col_in_872;
assign u0_col_in_873 = col_in_873;
assign u0_col_in_874 = col_in_874;
assign u0_col_in_875 = col_in_875;
assign u0_col_in_876 = col_in_876;
assign u0_col_in_877 = col_in_877;
assign u0_col_in_878 = col_in_878;
assign u0_col_in_879 = col_in_879;
assign u0_col_in_880 = col_in_880;
assign u0_col_in_881 = col_in_881;
assign u0_col_in_882 = col_in_882;
assign u0_col_in_883 = col_in_883;
assign u0_col_in_884 = col_in_884;
assign u0_col_in_885 = col_in_885;
assign u0_col_in_886 = col_in_886;
assign u0_col_in_887 = col_in_887;
assign u0_col_in_888 = col_in_888;
assign u0_col_in_889 = col_in_889;
assign u0_col_in_890 = col_in_890;
assign u0_col_in_891 = col_in_891;
assign u0_col_in_892 = col_in_892;
assign u0_col_in_893 = col_in_893;
assign u0_col_in_894 = col_in_894;
assign u0_col_in_895 = col_in_895;
assign u0_col_in_896 = col_in_896;
assign u0_col_in_897 = col_in_897;
assign u0_col_in_898 = col_in_898;
assign u0_col_in_899 = col_in_899;
assign u0_col_in_900 = col_in_900;
assign u0_col_in_901 = col_in_901;
assign u0_col_in_902 = col_in_902;
assign u0_col_in_903 = col_in_903;
assign u0_col_in_904 = col_in_904;
assign u0_col_in_905 = col_in_905;
assign u0_col_in_906 = col_in_906;
assign u0_col_in_907 = col_in_907;
assign u0_col_in_908 = col_in_908;
assign u0_col_in_909 = col_in_909;
assign u0_col_in_910 = col_in_910;
assign u0_col_in_911 = col_in_911;
assign u0_col_in_912 = col_in_912;
assign u0_col_in_913 = col_in_913;
assign u0_col_in_914 = col_in_914;
assign u0_col_in_915 = col_in_915;
assign u0_col_in_916 = col_in_916;
assign u0_col_in_917 = col_in_917;
assign u0_col_in_918 = col_in_918;
assign u0_col_in_919 = col_in_919;
assign u0_col_in_920 = col_in_920;
assign u0_col_in_921 = col_in_921;
assign u0_col_in_922 = col_in_922;
assign u0_col_in_923 = col_in_923;
assign u0_col_in_924 = col_in_924;
assign u0_col_in_925 = col_in_925;
assign u0_col_in_926 = col_in_926;
assign u0_col_in_927 = col_in_927;
assign u0_col_in_928 = col_in_928;
assign u0_col_in_929 = col_in_929;
assign u0_col_in_930 = col_in_930;
assign u0_col_in_931 = col_in_931;
assign u0_col_in_932 = col_in_932;
assign u0_col_in_933 = col_in_933;
assign u0_col_in_934 = col_in_934;
assign u0_col_in_935 = col_in_935;
assign u0_col_in_936 = col_in_936;
assign u0_col_in_937 = col_in_937;
assign u0_col_in_938 = col_in_938;
assign u0_col_in_939 = col_in_939;
assign u0_col_in_940 = col_in_940;
assign u0_col_in_941 = col_in_941;
assign u0_col_in_942 = col_in_942;
assign u0_col_in_943 = col_in_943;
assign u0_col_in_944 = col_in_944;
assign u0_col_in_945 = col_in_945;
assign u0_col_in_946 = col_in_946;
assign u0_col_in_947 = col_in_947;
assign u0_col_in_948 = col_in_948;
assign u0_col_in_949 = col_in_949;
assign u0_col_in_950 = col_in_950;
assign u0_col_in_951 = col_in_951;
assign u0_col_in_952 = col_in_952;
assign u0_col_in_953 = col_in_953;
assign u0_col_in_954 = col_in_954;
assign u0_col_in_955 = col_in_955;
assign u0_col_in_956 = col_in_956;
assign u0_col_in_957 = col_in_957;
assign u0_col_in_958 = col_in_958;
assign u0_col_in_959 = col_in_959;
assign u0_col_in_960 = col_in_960;
assign u0_col_in_961 = col_in_961;
assign u0_col_in_962 = col_in_962;
assign u0_col_in_963 = col_in_963;
assign u0_col_in_964 = col_in_964;
assign u0_col_in_965 = col_in_965;
assign u0_col_in_966 = col_in_966;
assign u0_col_in_967 = col_in_967;
assign u0_col_in_968 = col_in_968;
assign u0_col_in_969 = col_in_969;
assign u0_col_in_970 = col_in_970;
assign u0_col_in_971 = col_in_971;
assign u0_col_in_972 = col_in_972;
assign u0_col_in_973 = col_in_973;
assign u0_col_in_974 = col_in_974;
assign u0_col_in_975 = col_in_975;
assign u0_col_in_976 = col_in_976;
assign u0_col_in_977 = col_in_977;
assign u0_col_in_978 = col_in_978;
assign u0_col_in_979 = col_in_979;
assign u0_col_in_980 = col_in_980;
assign u0_col_in_981 = col_in_981;
assign u0_col_in_982 = col_in_982;
assign u0_col_in_983 = col_in_983;
assign u0_col_in_984 = col_in_984;
assign u0_col_in_985 = col_in_985;
assign u0_col_in_986 = col_in_986;
assign u0_col_in_987 = col_in_987;
assign u0_col_in_988 = col_in_988;
assign u0_col_in_989 = col_in_989;
assign u0_col_in_990 = col_in_990;
assign u0_col_in_991 = col_in_991;
assign u0_col_in_992 = col_in_992;
assign u0_col_in_993 = col_in_993;
assign u0_col_in_994 = col_in_994;
assign u0_col_in_995 = col_in_995;
assign u0_col_in_996 = col_in_996;
assign u0_col_in_997 = col_in_997;
assign u0_col_in_998 = col_in_998;
assign u0_col_in_999 = col_in_999;
assign u0_col_in_1000 = col_in_1000;
assign u0_col_in_1001 = col_in_1001;
assign u0_col_in_1002 = col_in_1002;
assign u0_col_in_1003 = col_in_1003;
assign u0_col_in_1004 = col_in_1004;
assign u0_col_in_1005 = col_in_1005;
assign u0_col_in_1006 = col_in_1006;
assign u0_col_in_1007 = col_in_1007;
assign u0_col_in_1008 = col_in_1008;
assign u0_col_in_1009 = col_in_1009;
assign u0_col_in_1010 = col_in_1010;
assign u0_col_in_1011 = col_in_1011;
assign u0_col_in_1012 = col_in_1012;
assign u0_col_in_1013 = col_in_1013;
assign u0_col_in_1014 = col_in_1014;
assign u0_col_in_1015 = col_in_1015;
assign u0_col_in_1016 = col_in_1016;
assign u0_col_in_1017 = col_in_1017;
assign u0_col_in_1018 = col_in_1018;
assign u0_col_in_1019 = col_in_1019;
assign u0_col_in_1020 = col_in_1020;
assign u0_col_in_1021 = col_in_1021;
assign u0_col_in_1022 = col_in_1022;
assign u0_col_in_1023 = col_in_1023;


//*****************************************************
//**************u0压缩阵列******************************
//*****************************************************
compressor_array_512_152_1024 u0_ca_512_152_1024
(
    .col_in_0(u0_col_in_0),
    .col_in_1(u0_col_in_1),
    .col_in_2(u0_col_in_2),
    .col_in_3(u0_col_in_3),
    .col_in_4(u0_col_in_4),
    .col_in_5(u0_col_in_5),
    .col_in_6(u0_col_in_6),
    .col_in_7(u0_col_in_7),
    .col_in_8(u0_col_in_8),
    .col_in_9(u0_col_in_9),
    .col_in_10(u0_col_in_10),
    .col_in_11(u0_col_in_11),
    .col_in_12(u0_col_in_12),
    .col_in_13(u0_col_in_13),
    .col_in_14(u0_col_in_14),
    .col_in_15(u0_col_in_15),
    .col_in_16(u0_col_in_16),
    .col_in_17(u0_col_in_17),
    .col_in_18(u0_col_in_18),
    .col_in_19(u0_col_in_19),
    .col_in_20(u0_col_in_20),
    .col_in_21(u0_col_in_21),
    .col_in_22(u0_col_in_22),
    .col_in_23(u0_col_in_23),
    .col_in_24(u0_col_in_24),
    .col_in_25(u0_col_in_25),
    .col_in_26(u0_col_in_26),
    .col_in_27(u0_col_in_27),
    .col_in_28(u0_col_in_28),
    .col_in_29(u0_col_in_29),
    .col_in_30(u0_col_in_30),
    .col_in_31(u0_col_in_31),
    .col_in_32(u0_col_in_32),
    .col_in_33(u0_col_in_33),
    .col_in_34(u0_col_in_34),
    .col_in_35(u0_col_in_35),
    .col_in_36(u0_col_in_36),
    .col_in_37(u0_col_in_37),
    .col_in_38(u0_col_in_38),
    .col_in_39(u0_col_in_39),
    .col_in_40(u0_col_in_40),
    .col_in_41(u0_col_in_41),
    .col_in_42(u0_col_in_42),
    .col_in_43(u0_col_in_43),
    .col_in_44(u0_col_in_44),
    .col_in_45(u0_col_in_45),
    .col_in_46(u0_col_in_46),
    .col_in_47(u0_col_in_47),
    .col_in_48(u0_col_in_48),
    .col_in_49(u0_col_in_49),
    .col_in_50(u0_col_in_50),
    .col_in_51(u0_col_in_51),
    .col_in_52(u0_col_in_52),
    .col_in_53(u0_col_in_53),
    .col_in_54(u0_col_in_54),
    .col_in_55(u0_col_in_55),
    .col_in_56(u0_col_in_56),
    .col_in_57(u0_col_in_57),
    .col_in_58(u0_col_in_58),
    .col_in_59(u0_col_in_59),
    .col_in_60(u0_col_in_60),
    .col_in_61(u0_col_in_61),
    .col_in_62(u0_col_in_62),
    .col_in_63(u0_col_in_63),
    .col_in_64(u0_col_in_64),
    .col_in_65(u0_col_in_65),
    .col_in_66(u0_col_in_66),
    .col_in_67(u0_col_in_67),
    .col_in_68(u0_col_in_68),
    .col_in_69(u0_col_in_69),
    .col_in_70(u0_col_in_70),
    .col_in_71(u0_col_in_71),
    .col_in_72(u0_col_in_72),
    .col_in_73(u0_col_in_73),
    .col_in_74(u0_col_in_74),
    .col_in_75(u0_col_in_75),
    .col_in_76(u0_col_in_76),
    .col_in_77(u0_col_in_77),
    .col_in_78(u0_col_in_78),
    .col_in_79(u0_col_in_79),
    .col_in_80(u0_col_in_80),
    .col_in_81(u0_col_in_81),
    .col_in_82(u0_col_in_82),
    .col_in_83(u0_col_in_83),
    .col_in_84(u0_col_in_84),
    .col_in_85(u0_col_in_85),
    .col_in_86(u0_col_in_86),
    .col_in_87(u0_col_in_87),
    .col_in_88(u0_col_in_88),
    .col_in_89(u0_col_in_89),
    .col_in_90(u0_col_in_90),
    .col_in_91(u0_col_in_91),
    .col_in_92(u0_col_in_92),
    .col_in_93(u0_col_in_93),
    .col_in_94(u0_col_in_94),
    .col_in_95(u0_col_in_95),
    .col_in_96(u0_col_in_96),
    .col_in_97(u0_col_in_97),
    .col_in_98(u0_col_in_98),
    .col_in_99(u0_col_in_99),
    .col_in_100(u0_col_in_100),
    .col_in_101(u0_col_in_101),
    .col_in_102(u0_col_in_102),
    .col_in_103(u0_col_in_103),
    .col_in_104(u0_col_in_104),
    .col_in_105(u0_col_in_105),
    .col_in_106(u0_col_in_106),
    .col_in_107(u0_col_in_107),
    .col_in_108(u0_col_in_108),
    .col_in_109(u0_col_in_109),
    .col_in_110(u0_col_in_110),
    .col_in_111(u0_col_in_111),
    .col_in_112(u0_col_in_112),
    .col_in_113(u0_col_in_113),
    .col_in_114(u0_col_in_114),
    .col_in_115(u0_col_in_115),
    .col_in_116(u0_col_in_116),
    .col_in_117(u0_col_in_117),
    .col_in_118(u0_col_in_118),
    .col_in_119(u0_col_in_119),
    .col_in_120(u0_col_in_120),
    .col_in_121(u0_col_in_121),
    .col_in_122(u0_col_in_122),
    .col_in_123(u0_col_in_123),
    .col_in_124(u0_col_in_124),
    .col_in_125(u0_col_in_125),
    .col_in_126(u0_col_in_126),
    .col_in_127(u0_col_in_127),
    .col_in_128(u0_col_in_128),
    .col_in_129(u0_col_in_129),
    .col_in_130(u0_col_in_130),
    .col_in_131(u0_col_in_131),
    .col_in_132(u0_col_in_132),
    .col_in_133(u0_col_in_133),
    .col_in_134(u0_col_in_134),
    .col_in_135(u0_col_in_135),
    .col_in_136(u0_col_in_136),
    .col_in_137(u0_col_in_137),
    .col_in_138(u0_col_in_138),
    .col_in_139(u0_col_in_139),
    .col_in_140(u0_col_in_140),
    .col_in_141(u0_col_in_141),
    .col_in_142(u0_col_in_142),
    .col_in_143(u0_col_in_143),
    .col_in_144(u0_col_in_144),
    .col_in_145(u0_col_in_145),
    .col_in_146(u0_col_in_146),
    .col_in_147(u0_col_in_147),
    .col_in_148(u0_col_in_148),
    .col_in_149(u0_col_in_149),
    .col_in_150(u0_col_in_150),
    .col_in_151(u0_col_in_151),
    .col_in_152(u0_col_in_152),
    .col_in_153(u0_col_in_153),
    .col_in_154(u0_col_in_154),
    .col_in_155(u0_col_in_155),
    .col_in_156(u0_col_in_156),
    .col_in_157(u0_col_in_157),
    .col_in_158(u0_col_in_158),
    .col_in_159(u0_col_in_159),
    .col_in_160(u0_col_in_160),
    .col_in_161(u0_col_in_161),
    .col_in_162(u0_col_in_162),
    .col_in_163(u0_col_in_163),
    .col_in_164(u0_col_in_164),
    .col_in_165(u0_col_in_165),
    .col_in_166(u0_col_in_166),
    .col_in_167(u0_col_in_167),
    .col_in_168(u0_col_in_168),
    .col_in_169(u0_col_in_169),
    .col_in_170(u0_col_in_170),
    .col_in_171(u0_col_in_171),
    .col_in_172(u0_col_in_172),
    .col_in_173(u0_col_in_173),
    .col_in_174(u0_col_in_174),
    .col_in_175(u0_col_in_175),
    .col_in_176(u0_col_in_176),
    .col_in_177(u0_col_in_177),
    .col_in_178(u0_col_in_178),
    .col_in_179(u0_col_in_179),
    .col_in_180(u0_col_in_180),
    .col_in_181(u0_col_in_181),
    .col_in_182(u0_col_in_182),
    .col_in_183(u0_col_in_183),
    .col_in_184(u0_col_in_184),
    .col_in_185(u0_col_in_185),
    .col_in_186(u0_col_in_186),
    .col_in_187(u0_col_in_187),
    .col_in_188(u0_col_in_188),
    .col_in_189(u0_col_in_189),
    .col_in_190(u0_col_in_190),
    .col_in_191(u0_col_in_191),
    .col_in_192(u0_col_in_192),
    .col_in_193(u0_col_in_193),
    .col_in_194(u0_col_in_194),
    .col_in_195(u0_col_in_195),
    .col_in_196(u0_col_in_196),
    .col_in_197(u0_col_in_197),
    .col_in_198(u0_col_in_198),
    .col_in_199(u0_col_in_199),
    .col_in_200(u0_col_in_200),
    .col_in_201(u0_col_in_201),
    .col_in_202(u0_col_in_202),
    .col_in_203(u0_col_in_203),
    .col_in_204(u0_col_in_204),
    .col_in_205(u0_col_in_205),
    .col_in_206(u0_col_in_206),
    .col_in_207(u0_col_in_207),
    .col_in_208(u0_col_in_208),
    .col_in_209(u0_col_in_209),
    .col_in_210(u0_col_in_210),
    .col_in_211(u0_col_in_211),
    .col_in_212(u0_col_in_212),
    .col_in_213(u0_col_in_213),
    .col_in_214(u0_col_in_214),
    .col_in_215(u0_col_in_215),
    .col_in_216(u0_col_in_216),
    .col_in_217(u0_col_in_217),
    .col_in_218(u0_col_in_218),
    .col_in_219(u0_col_in_219),
    .col_in_220(u0_col_in_220),
    .col_in_221(u0_col_in_221),
    .col_in_222(u0_col_in_222),
    .col_in_223(u0_col_in_223),
    .col_in_224(u0_col_in_224),
    .col_in_225(u0_col_in_225),
    .col_in_226(u0_col_in_226),
    .col_in_227(u0_col_in_227),
    .col_in_228(u0_col_in_228),
    .col_in_229(u0_col_in_229),
    .col_in_230(u0_col_in_230),
    .col_in_231(u0_col_in_231),
    .col_in_232(u0_col_in_232),
    .col_in_233(u0_col_in_233),
    .col_in_234(u0_col_in_234),
    .col_in_235(u0_col_in_235),
    .col_in_236(u0_col_in_236),
    .col_in_237(u0_col_in_237),
    .col_in_238(u0_col_in_238),
    .col_in_239(u0_col_in_239),
    .col_in_240(u0_col_in_240),
    .col_in_241(u0_col_in_241),
    .col_in_242(u0_col_in_242),
    .col_in_243(u0_col_in_243),
    .col_in_244(u0_col_in_244),
    .col_in_245(u0_col_in_245),
    .col_in_246(u0_col_in_246),
    .col_in_247(u0_col_in_247),
    .col_in_248(u0_col_in_248),
    .col_in_249(u0_col_in_249),
    .col_in_250(u0_col_in_250),
    .col_in_251(u0_col_in_251),
    .col_in_252(u0_col_in_252),
    .col_in_253(u0_col_in_253),
    .col_in_254(u0_col_in_254),
    .col_in_255(u0_col_in_255),
    .col_in_256(u0_col_in_256),
    .col_in_257(u0_col_in_257),
    .col_in_258(u0_col_in_258),
    .col_in_259(u0_col_in_259),
    .col_in_260(u0_col_in_260),
    .col_in_261(u0_col_in_261),
    .col_in_262(u0_col_in_262),
    .col_in_263(u0_col_in_263),
    .col_in_264(u0_col_in_264),
    .col_in_265(u0_col_in_265),
    .col_in_266(u0_col_in_266),
    .col_in_267(u0_col_in_267),
    .col_in_268(u0_col_in_268),
    .col_in_269(u0_col_in_269),
    .col_in_270(u0_col_in_270),
    .col_in_271(u0_col_in_271),
    .col_in_272(u0_col_in_272),
    .col_in_273(u0_col_in_273),
    .col_in_274(u0_col_in_274),
    .col_in_275(u0_col_in_275),
    .col_in_276(u0_col_in_276),
    .col_in_277(u0_col_in_277),
    .col_in_278(u0_col_in_278),
    .col_in_279(u0_col_in_279),
    .col_in_280(u0_col_in_280),
    .col_in_281(u0_col_in_281),
    .col_in_282(u0_col_in_282),
    .col_in_283(u0_col_in_283),
    .col_in_284(u0_col_in_284),
    .col_in_285(u0_col_in_285),
    .col_in_286(u0_col_in_286),
    .col_in_287(u0_col_in_287),
    .col_in_288(u0_col_in_288),
    .col_in_289(u0_col_in_289),
    .col_in_290(u0_col_in_290),
    .col_in_291(u0_col_in_291),
    .col_in_292(u0_col_in_292),
    .col_in_293(u0_col_in_293),
    .col_in_294(u0_col_in_294),
    .col_in_295(u0_col_in_295),
    .col_in_296(u0_col_in_296),
    .col_in_297(u0_col_in_297),
    .col_in_298(u0_col_in_298),
    .col_in_299(u0_col_in_299),
    .col_in_300(u0_col_in_300),
    .col_in_301(u0_col_in_301),
    .col_in_302(u0_col_in_302),
    .col_in_303(u0_col_in_303),
    .col_in_304(u0_col_in_304),
    .col_in_305(u0_col_in_305),
    .col_in_306(u0_col_in_306),
    .col_in_307(u0_col_in_307),
    .col_in_308(u0_col_in_308),
    .col_in_309(u0_col_in_309),
    .col_in_310(u0_col_in_310),
    .col_in_311(u0_col_in_311),
    .col_in_312(u0_col_in_312),
    .col_in_313(u0_col_in_313),
    .col_in_314(u0_col_in_314),
    .col_in_315(u0_col_in_315),
    .col_in_316(u0_col_in_316),
    .col_in_317(u0_col_in_317),
    .col_in_318(u0_col_in_318),
    .col_in_319(u0_col_in_319),
    .col_in_320(u0_col_in_320),
    .col_in_321(u0_col_in_321),
    .col_in_322(u0_col_in_322),
    .col_in_323(u0_col_in_323),
    .col_in_324(u0_col_in_324),
    .col_in_325(u0_col_in_325),
    .col_in_326(u0_col_in_326),
    .col_in_327(u0_col_in_327),
    .col_in_328(u0_col_in_328),
    .col_in_329(u0_col_in_329),
    .col_in_330(u0_col_in_330),
    .col_in_331(u0_col_in_331),
    .col_in_332(u0_col_in_332),
    .col_in_333(u0_col_in_333),
    .col_in_334(u0_col_in_334),
    .col_in_335(u0_col_in_335),
    .col_in_336(u0_col_in_336),
    .col_in_337(u0_col_in_337),
    .col_in_338(u0_col_in_338),
    .col_in_339(u0_col_in_339),
    .col_in_340(u0_col_in_340),
    .col_in_341(u0_col_in_341),
    .col_in_342(u0_col_in_342),
    .col_in_343(u0_col_in_343),
    .col_in_344(u0_col_in_344),
    .col_in_345(u0_col_in_345),
    .col_in_346(u0_col_in_346),
    .col_in_347(u0_col_in_347),
    .col_in_348(u0_col_in_348),
    .col_in_349(u0_col_in_349),
    .col_in_350(u0_col_in_350),
    .col_in_351(u0_col_in_351),
    .col_in_352(u0_col_in_352),
    .col_in_353(u0_col_in_353),
    .col_in_354(u0_col_in_354),
    .col_in_355(u0_col_in_355),
    .col_in_356(u0_col_in_356),
    .col_in_357(u0_col_in_357),
    .col_in_358(u0_col_in_358),
    .col_in_359(u0_col_in_359),
    .col_in_360(u0_col_in_360),
    .col_in_361(u0_col_in_361),
    .col_in_362(u0_col_in_362),
    .col_in_363(u0_col_in_363),
    .col_in_364(u0_col_in_364),
    .col_in_365(u0_col_in_365),
    .col_in_366(u0_col_in_366),
    .col_in_367(u0_col_in_367),
    .col_in_368(u0_col_in_368),
    .col_in_369(u0_col_in_369),
    .col_in_370(u0_col_in_370),
    .col_in_371(u0_col_in_371),
    .col_in_372(u0_col_in_372),
    .col_in_373(u0_col_in_373),
    .col_in_374(u0_col_in_374),
    .col_in_375(u0_col_in_375),
    .col_in_376(u0_col_in_376),
    .col_in_377(u0_col_in_377),
    .col_in_378(u0_col_in_378),
    .col_in_379(u0_col_in_379),
    .col_in_380(u0_col_in_380),
    .col_in_381(u0_col_in_381),
    .col_in_382(u0_col_in_382),
    .col_in_383(u0_col_in_383),
    .col_in_384(u0_col_in_384),
    .col_in_385(u0_col_in_385),
    .col_in_386(u0_col_in_386),
    .col_in_387(u0_col_in_387),
    .col_in_388(u0_col_in_388),
    .col_in_389(u0_col_in_389),
    .col_in_390(u0_col_in_390),
    .col_in_391(u0_col_in_391),
    .col_in_392(u0_col_in_392),
    .col_in_393(u0_col_in_393),
    .col_in_394(u0_col_in_394),
    .col_in_395(u0_col_in_395),
    .col_in_396(u0_col_in_396),
    .col_in_397(u0_col_in_397),
    .col_in_398(u0_col_in_398),
    .col_in_399(u0_col_in_399),
    .col_in_400(u0_col_in_400),
    .col_in_401(u0_col_in_401),
    .col_in_402(u0_col_in_402),
    .col_in_403(u0_col_in_403),
    .col_in_404(u0_col_in_404),
    .col_in_405(u0_col_in_405),
    .col_in_406(u0_col_in_406),
    .col_in_407(u0_col_in_407),
    .col_in_408(u0_col_in_408),
    .col_in_409(u0_col_in_409),
    .col_in_410(u0_col_in_410),
    .col_in_411(u0_col_in_411),
    .col_in_412(u0_col_in_412),
    .col_in_413(u0_col_in_413),
    .col_in_414(u0_col_in_414),
    .col_in_415(u0_col_in_415),
    .col_in_416(u0_col_in_416),
    .col_in_417(u0_col_in_417),
    .col_in_418(u0_col_in_418),
    .col_in_419(u0_col_in_419),
    .col_in_420(u0_col_in_420),
    .col_in_421(u0_col_in_421),
    .col_in_422(u0_col_in_422),
    .col_in_423(u0_col_in_423),
    .col_in_424(u0_col_in_424),
    .col_in_425(u0_col_in_425),
    .col_in_426(u0_col_in_426),
    .col_in_427(u0_col_in_427),
    .col_in_428(u0_col_in_428),
    .col_in_429(u0_col_in_429),
    .col_in_430(u0_col_in_430),
    .col_in_431(u0_col_in_431),
    .col_in_432(u0_col_in_432),
    .col_in_433(u0_col_in_433),
    .col_in_434(u0_col_in_434),
    .col_in_435(u0_col_in_435),
    .col_in_436(u0_col_in_436),
    .col_in_437(u0_col_in_437),
    .col_in_438(u0_col_in_438),
    .col_in_439(u0_col_in_439),
    .col_in_440(u0_col_in_440),
    .col_in_441(u0_col_in_441),
    .col_in_442(u0_col_in_442),
    .col_in_443(u0_col_in_443),
    .col_in_444(u0_col_in_444),
    .col_in_445(u0_col_in_445),
    .col_in_446(u0_col_in_446),
    .col_in_447(u0_col_in_447),
    .col_in_448(u0_col_in_448),
    .col_in_449(u0_col_in_449),
    .col_in_450(u0_col_in_450),
    .col_in_451(u0_col_in_451),
    .col_in_452(u0_col_in_452),
    .col_in_453(u0_col_in_453),
    .col_in_454(u0_col_in_454),
    .col_in_455(u0_col_in_455),
    .col_in_456(u0_col_in_456),
    .col_in_457(u0_col_in_457),
    .col_in_458(u0_col_in_458),
    .col_in_459(u0_col_in_459),
    .col_in_460(u0_col_in_460),
    .col_in_461(u0_col_in_461),
    .col_in_462(u0_col_in_462),
    .col_in_463(u0_col_in_463),
    .col_in_464(u0_col_in_464),
    .col_in_465(u0_col_in_465),
    .col_in_466(u0_col_in_466),
    .col_in_467(u0_col_in_467),
    .col_in_468(u0_col_in_468),
    .col_in_469(u0_col_in_469),
    .col_in_470(u0_col_in_470),
    .col_in_471(u0_col_in_471),
    .col_in_472(u0_col_in_472),
    .col_in_473(u0_col_in_473),
    .col_in_474(u0_col_in_474),
    .col_in_475(u0_col_in_475),
    .col_in_476(u0_col_in_476),
    .col_in_477(u0_col_in_477),
    .col_in_478(u0_col_in_478),
    .col_in_479(u0_col_in_479),
    .col_in_480(u0_col_in_480),
    .col_in_481(u0_col_in_481),
    .col_in_482(u0_col_in_482),
    .col_in_483(u0_col_in_483),
    .col_in_484(u0_col_in_484),
    .col_in_485(u0_col_in_485),
    .col_in_486(u0_col_in_486),
    .col_in_487(u0_col_in_487),
    .col_in_488(u0_col_in_488),
    .col_in_489(u0_col_in_489),
    .col_in_490(u0_col_in_490),
    .col_in_491(u0_col_in_491),
    .col_in_492(u0_col_in_492),
    .col_in_493(u0_col_in_493),
    .col_in_494(u0_col_in_494),
    .col_in_495(u0_col_in_495),
    .col_in_496(u0_col_in_496),
    .col_in_497(u0_col_in_497),
    .col_in_498(u0_col_in_498),
    .col_in_499(u0_col_in_499),
    .col_in_500(u0_col_in_500),
    .col_in_501(u0_col_in_501),
    .col_in_502(u0_col_in_502),
    .col_in_503(u0_col_in_503),
    .col_in_504(u0_col_in_504),
    .col_in_505(u0_col_in_505),
    .col_in_506(u0_col_in_506),
    .col_in_507(u0_col_in_507),
    .col_in_508(u0_col_in_508),
    .col_in_509(u0_col_in_509),
    .col_in_510(u0_col_in_510),
    .col_in_511(u0_col_in_511),
    .col_in_512(u0_col_in_512),
    .col_in_513(u0_col_in_513),
    .col_in_514(u0_col_in_514),
    .col_in_515(u0_col_in_515),
    .col_in_516(u0_col_in_516),
    .col_in_517(u0_col_in_517),
    .col_in_518(u0_col_in_518),
    .col_in_519(u0_col_in_519),
    .col_in_520(u0_col_in_520),
    .col_in_521(u0_col_in_521),
    .col_in_522(u0_col_in_522),
    .col_in_523(u0_col_in_523),
    .col_in_524(u0_col_in_524),
    .col_in_525(u0_col_in_525),
    .col_in_526(u0_col_in_526),
    .col_in_527(u0_col_in_527),
    .col_in_528(u0_col_in_528),
    .col_in_529(u0_col_in_529),
    .col_in_530(u0_col_in_530),
    .col_in_531(u0_col_in_531),
    .col_in_532(u0_col_in_532),
    .col_in_533(u0_col_in_533),
    .col_in_534(u0_col_in_534),
    .col_in_535(u0_col_in_535),
    .col_in_536(u0_col_in_536),
    .col_in_537(u0_col_in_537),
    .col_in_538(u0_col_in_538),
    .col_in_539(u0_col_in_539),
    .col_in_540(u0_col_in_540),
    .col_in_541(u0_col_in_541),
    .col_in_542(u0_col_in_542),
    .col_in_543(u0_col_in_543),
    .col_in_544(u0_col_in_544),
    .col_in_545(u0_col_in_545),
    .col_in_546(u0_col_in_546),
    .col_in_547(u0_col_in_547),
    .col_in_548(u0_col_in_548),
    .col_in_549(u0_col_in_549),
    .col_in_550(u0_col_in_550),
    .col_in_551(u0_col_in_551),
    .col_in_552(u0_col_in_552),
    .col_in_553(u0_col_in_553),
    .col_in_554(u0_col_in_554),
    .col_in_555(u0_col_in_555),
    .col_in_556(u0_col_in_556),
    .col_in_557(u0_col_in_557),
    .col_in_558(u0_col_in_558),
    .col_in_559(u0_col_in_559),
    .col_in_560(u0_col_in_560),
    .col_in_561(u0_col_in_561),
    .col_in_562(u0_col_in_562),
    .col_in_563(u0_col_in_563),
    .col_in_564(u0_col_in_564),
    .col_in_565(u0_col_in_565),
    .col_in_566(u0_col_in_566),
    .col_in_567(u0_col_in_567),
    .col_in_568(u0_col_in_568),
    .col_in_569(u0_col_in_569),
    .col_in_570(u0_col_in_570),
    .col_in_571(u0_col_in_571),
    .col_in_572(u0_col_in_572),
    .col_in_573(u0_col_in_573),
    .col_in_574(u0_col_in_574),
    .col_in_575(u0_col_in_575),
    .col_in_576(u0_col_in_576),
    .col_in_577(u0_col_in_577),
    .col_in_578(u0_col_in_578),
    .col_in_579(u0_col_in_579),
    .col_in_580(u0_col_in_580),
    .col_in_581(u0_col_in_581),
    .col_in_582(u0_col_in_582),
    .col_in_583(u0_col_in_583),
    .col_in_584(u0_col_in_584),
    .col_in_585(u0_col_in_585),
    .col_in_586(u0_col_in_586),
    .col_in_587(u0_col_in_587),
    .col_in_588(u0_col_in_588),
    .col_in_589(u0_col_in_589),
    .col_in_590(u0_col_in_590),
    .col_in_591(u0_col_in_591),
    .col_in_592(u0_col_in_592),
    .col_in_593(u0_col_in_593),
    .col_in_594(u0_col_in_594),
    .col_in_595(u0_col_in_595),
    .col_in_596(u0_col_in_596),
    .col_in_597(u0_col_in_597),
    .col_in_598(u0_col_in_598),
    .col_in_599(u0_col_in_599),
    .col_in_600(u0_col_in_600),
    .col_in_601(u0_col_in_601),
    .col_in_602(u0_col_in_602),
    .col_in_603(u0_col_in_603),
    .col_in_604(u0_col_in_604),
    .col_in_605(u0_col_in_605),
    .col_in_606(u0_col_in_606),
    .col_in_607(u0_col_in_607),
    .col_in_608(u0_col_in_608),
    .col_in_609(u0_col_in_609),
    .col_in_610(u0_col_in_610),
    .col_in_611(u0_col_in_611),
    .col_in_612(u0_col_in_612),
    .col_in_613(u0_col_in_613),
    .col_in_614(u0_col_in_614),
    .col_in_615(u0_col_in_615),
    .col_in_616(u0_col_in_616),
    .col_in_617(u0_col_in_617),
    .col_in_618(u0_col_in_618),
    .col_in_619(u0_col_in_619),
    .col_in_620(u0_col_in_620),
    .col_in_621(u0_col_in_621),
    .col_in_622(u0_col_in_622),
    .col_in_623(u0_col_in_623),
    .col_in_624(u0_col_in_624),
    .col_in_625(u0_col_in_625),
    .col_in_626(u0_col_in_626),
    .col_in_627(u0_col_in_627),
    .col_in_628(u0_col_in_628),
    .col_in_629(u0_col_in_629),
    .col_in_630(u0_col_in_630),
    .col_in_631(u0_col_in_631),
    .col_in_632(u0_col_in_632),
    .col_in_633(u0_col_in_633),
    .col_in_634(u0_col_in_634),
    .col_in_635(u0_col_in_635),
    .col_in_636(u0_col_in_636),
    .col_in_637(u0_col_in_637),
    .col_in_638(u0_col_in_638),
    .col_in_639(u0_col_in_639),
    .col_in_640(u0_col_in_640),
    .col_in_641(u0_col_in_641),
    .col_in_642(u0_col_in_642),
    .col_in_643(u0_col_in_643),
    .col_in_644(u0_col_in_644),
    .col_in_645(u0_col_in_645),
    .col_in_646(u0_col_in_646),
    .col_in_647(u0_col_in_647),
    .col_in_648(u0_col_in_648),
    .col_in_649(u0_col_in_649),
    .col_in_650(u0_col_in_650),
    .col_in_651(u0_col_in_651),
    .col_in_652(u0_col_in_652),
    .col_in_653(u0_col_in_653),
    .col_in_654(u0_col_in_654),
    .col_in_655(u0_col_in_655),
    .col_in_656(u0_col_in_656),
    .col_in_657(u0_col_in_657),
    .col_in_658(u0_col_in_658),
    .col_in_659(u0_col_in_659),
    .col_in_660(u0_col_in_660),
    .col_in_661(u0_col_in_661),
    .col_in_662(u0_col_in_662),
    .col_in_663(u0_col_in_663),
    .col_in_664(u0_col_in_664),
    .col_in_665(u0_col_in_665),
    .col_in_666(u0_col_in_666),
    .col_in_667(u0_col_in_667),
    .col_in_668(u0_col_in_668),
    .col_in_669(u0_col_in_669),
    .col_in_670(u0_col_in_670),
    .col_in_671(u0_col_in_671),
    .col_in_672(u0_col_in_672),
    .col_in_673(u0_col_in_673),
    .col_in_674(u0_col_in_674),
    .col_in_675(u0_col_in_675),
    .col_in_676(u0_col_in_676),
    .col_in_677(u0_col_in_677),
    .col_in_678(u0_col_in_678),
    .col_in_679(u0_col_in_679),
    .col_in_680(u0_col_in_680),
    .col_in_681(u0_col_in_681),
    .col_in_682(u0_col_in_682),
    .col_in_683(u0_col_in_683),
    .col_in_684(u0_col_in_684),
    .col_in_685(u0_col_in_685),
    .col_in_686(u0_col_in_686),
    .col_in_687(u0_col_in_687),
    .col_in_688(u0_col_in_688),
    .col_in_689(u0_col_in_689),
    .col_in_690(u0_col_in_690),
    .col_in_691(u0_col_in_691),
    .col_in_692(u0_col_in_692),
    .col_in_693(u0_col_in_693),
    .col_in_694(u0_col_in_694),
    .col_in_695(u0_col_in_695),
    .col_in_696(u0_col_in_696),
    .col_in_697(u0_col_in_697),
    .col_in_698(u0_col_in_698),
    .col_in_699(u0_col_in_699),
    .col_in_700(u0_col_in_700),
    .col_in_701(u0_col_in_701),
    .col_in_702(u0_col_in_702),
    .col_in_703(u0_col_in_703),
    .col_in_704(u0_col_in_704),
    .col_in_705(u0_col_in_705),
    .col_in_706(u0_col_in_706),
    .col_in_707(u0_col_in_707),
    .col_in_708(u0_col_in_708),
    .col_in_709(u0_col_in_709),
    .col_in_710(u0_col_in_710),
    .col_in_711(u0_col_in_711),
    .col_in_712(u0_col_in_712),
    .col_in_713(u0_col_in_713),
    .col_in_714(u0_col_in_714),
    .col_in_715(u0_col_in_715),
    .col_in_716(u0_col_in_716),
    .col_in_717(u0_col_in_717),
    .col_in_718(u0_col_in_718),
    .col_in_719(u0_col_in_719),
    .col_in_720(u0_col_in_720),
    .col_in_721(u0_col_in_721),
    .col_in_722(u0_col_in_722),
    .col_in_723(u0_col_in_723),
    .col_in_724(u0_col_in_724),
    .col_in_725(u0_col_in_725),
    .col_in_726(u0_col_in_726),
    .col_in_727(u0_col_in_727),
    .col_in_728(u0_col_in_728),
    .col_in_729(u0_col_in_729),
    .col_in_730(u0_col_in_730),
    .col_in_731(u0_col_in_731),
    .col_in_732(u0_col_in_732),
    .col_in_733(u0_col_in_733),
    .col_in_734(u0_col_in_734),
    .col_in_735(u0_col_in_735),
    .col_in_736(u0_col_in_736),
    .col_in_737(u0_col_in_737),
    .col_in_738(u0_col_in_738),
    .col_in_739(u0_col_in_739),
    .col_in_740(u0_col_in_740),
    .col_in_741(u0_col_in_741),
    .col_in_742(u0_col_in_742),
    .col_in_743(u0_col_in_743),
    .col_in_744(u0_col_in_744),
    .col_in_745(u0_col_in_745),
    .col_in_746(u0_col_in_746),
    .col_in_747(u0_col_in_747),
    .col_in_748(u0_col_in_748),
    .col_in_749(u0_col_in_749),
    .col_in_750(u0_col_in_750),
    .col_in_751(u0_col_in_751),
    .col_in_752(u0_col_in_752),
    .col_in_753(u0_col_in_753),
    .col_in_754(u0_col_in_754),
    .col_in_755(u0_col_in_755),
    .col_in_756(u0_col_in_756),
    .col_in_757(u0_col_in_757),
    .col_in_758(u0_col_in_758),
    .col_in_759(u0_col_in_759),
    .col_in_760(u0_col_in_760),
    .col_in_761(u0_col_in_761),
    .col_in_762(u0_col_in_762),
    .col_in_763(u0_col_in_763),
    .col_in_764(u0_col_in_764),
    .col_in_765(u0_col_in_765),
    .col_in_766(u0_col_in_766),
    .col_in_767(u0_col_in_767),
    .col_in_768(u0_col_in_768),
    .col_in_769(u0_col_in_769),
    .col_in_770(u0_col_in_770),
    .col_in_771(u0_col_in_771),
    .col_in_772(u0_col_in_772),
    .col_in_773(u0_col_in_773),
    .col_in_774(u0_col_in_774),
    .col_in_775(u0_col_in_775),
    .col_in_776(u0_col_in_776),
    .col_in_777(u0_col_in_777),
    .col_in_778(u0_col_in_778),
    .col_in_779(u0_col_in_779),
    .col_in_780(u0_col_in_780),
    .col_in_781(u0_col_in_781),
    .col_in_782(u0_col_in_782),
    .col_in_783(u0_col_in_783),
    .col_in_784(u0_col_in_784),
    .col_in_785(u0_col_in_785),
    .col_in_786(u0_col_in_786),
    .col_in_787(u0_col_in_787),
    .col_in_788(u0_col_in_788),
    .col_in_789(u0_col_in_789),
    .col_in_790(u0_col_in_790),
    .col_in_791(u0_col_in_791),
    .col_in_792(u0_col_in_792),
    .col_in_793(u0_col_in_793),
    .col_in_794(u0_col_in_794),
    .col_in_795(u0_col_in_795),
    .col_in_796(u0_col_in_796),
    .col_in_797(u0_col_in_797),
    .col_in_798(u0_col_in_798),
    .col_in_799(u0_col_in_799),
    .col_in_800(u0_col_in_800),
    .col_in_801(u0_col_in_801),
    .col_in_802(u0_col_in_802),
    .col_in_803(u0_col_in_803),
    .col_in_804(u0_col_in_804),
    .col_in_805(u0_col_in_805),
    .col_in_806(u0_col_in_806),
    .col_in_807(u0_col_in_807),
    .col_in_808(u0_col_in_808),
    .col_in_809(u0_col_in_809),
    .col_in_810(u0_col_in_810),
    .col_in_811(u0_col_in_811),
    .col_in_812(u0_col_in_812),
    .col_in_813(u0_col_in_813),
    .col_in_814(u0_col_in_814),
    .col_in_815(u0_col_in_815),
    .col_in_816(u0_col_in_816),
    .col_in_817(u0_col_in_817),
    .col_in_818(u0_col_in_818),
    .col_in_819(u0_col_in_819),
    .col_in_820(u0_col_in_820),
    .col_in_821(u0_col_in_821),
    .col_in_822(u0_col_in_822),
    .col_in_823(u0_col_in_823),
    .col_in_824(u0_col_in_824),
    .col_in_825(u0_col_in_825),
    .col_in_826(u0_col_in_826),
    .col_in_827(u0_col_in_827),
    .col_in_828(u0_col_in_828),
    .col_in_829(u0_col_in_829),
    .col_in_830(u0_col_in_830),
    .col_in_831(u0_col_in_831),
    .col_in_832(u0_col_in_832),
    .col_in_833(u0_col_in_833),
    .col_in_834(u0_col_in_834),
    .col_in_835(u0_col_in_835),
    .col_in_836(u0_col_in_836),
    .col_in_837(u0_col_in_837),
    .col_in_838(u0_col_in_838),
    .col_in_839(u0_col_in_839),
    .col_in_840(u0_col_in_840),
    .col_in_841(u0_col_in_841),
    .col_in_842(u0_col_in_842),
    .col_in_843(u0_col_in_843),
    .col_in_844(u0_col_in_844),
    .col_in_845(u0_col_in_845),
    .col_in_846(u0_col_in_846),
    .col_in_847(u0_col_in_847),
    .col_in_848(u0_col_in_848),
    .col_in_849(u0_col_in_849),
    .col_in_850(u0_col_in_850),
    .col_in_851(u0_col_in_851),
    .col_in_852(u0_col_in_852),
    .col_in_853(u0_col_in_853),
    .col_in_854(u0_col_in_854),
    .col_in_855(u0_col_in_855),
    .col_in_856(u0_col_in_856),
    .col_in_857(u0_col_in_857),
    .col_in_858(u0_col_in_858),
    .col_in_859(u0_col_in_859),
    .col_in_860(u0_col_in_860),
    .col_in_861(u0_col_in_861),
    .col_in_862(u0_col_in_862),
    .col_in_863(u0_col_in_863),
    .col_in_864(u0_col_in_864),
    .col_in_865(u0_col_in_865),
    .col_in_866(u0_col_in_866),
    .col_in_867(u0_col_in_867),
    .col_in_868(u0_col_in_868),
    .col_in_869(u0_col_in_869),
    .col_in_870(u0_col_in_870),
    .col_in_871(u0_col_in_871),
    .col_in_872(u0_col_in_872),
    .col_in_873(u0_col_in_873),
    .col_in_874(u0_col_in_874),
    .col_in_875(u0_col_in_875),
    .col_in_876(u0_col_in_876),
    .col_in_877(u0_col_in_877),
    .col_in_878(u0_col_in_878),
    .col_in_879(u0_col_in_879),
    .col_in_880(u0_col_in_880),
    .col_in_881(u0_col_in_881),
    .col_in_882(u0_col_in_882),
    .col_in_883(u0_col_in_883),
    .col_in_884(u0_col_in_884),
    .col_in_885(u0_col_in_885),
    .col_in_886(u0_col_in_886),
    .col_in_887(u0_col_in_887),
    .col_in_888(u0_col_in_888),
    .col_in_889(u0_col_in_889),
    .col_in_890(u0_col_in_890),
    .col_in_891(u0_col_in_891),
    .col_in_892(u0_col_in_892),
    .col_in_893(u0_col_in_893),
    .col_in_894(u0_col_in_894),
    .col_in_895(u0_col_in_895),
    .col_in_896(u0_col_in_896),
    .col_in_897(u0_col_in_897),
    .col_in_898(u0_col_in_898),
    .col_in_899(u0_col_in_899),
    .col_in_900(u0_col_in_900),
    .col_in_901(u0_col_in_901),
    .col_in_902(u0_col_in_902),
    .col_in_903(u0_col_in_903),
    .col_in_904(u0_col_in_904),
    .col_in_905(u0_col_in_905),
    .col_in_906(u0_col_in_906),
    .col_in_907(u0_col_in_907),
    .col_in_908(u0_col_in_908),
    .col_in_909(u0_col_in_909),
    .col_in_910(u0_col_in_910),
    .col_in_911(u0_col_in_911),
    .col_in_912(u0_col_in_912),
    .col_in_913(u0_col_in_913),
    .col_in_914(u0_col_in_914),
    .col_in_915(u0_col_in_915),
    .col_in_916(u0_col_in_916),
    .col_in_917(u0_col_in_917),
    .col_in_918(u0_col_in_918),
    .col_in_919(u0_col_in_919),
    .col_in_920(u0_col_in_920),
    .col_in_921(u0_col_in_921),
    .col_in_922(u0_col_in_922),
    .col_in_923(u0_col_in_923),
    .col_in_924(u0_col_in_924),
    .col_in_925(u0_col_in_925),
    .col_in_926(u0_col_in_926),
    .col_in_927(u0_col_in_927),
    .col_in_928(u0_col_in_928),
    .col_in_929(u0_col_in_929),
    .col_in_930(u0_col_in_930),
    .col_in_931(u0_col_in_931),
    .col_in_932(u0_col_in_932),
    .col_in_933(u0_col_in_933),
    .col_in_934(u0_col_in_934),
    .col_in_935(u0_col_in_935),
    .col_in_936(u0_col_in_936),
    .col_in_937(u0_col_in_937),
    .col_in_938(u0_col_in_938),
    .col_in_939(u0_col_in_939),
    .col_in_940(u0_col_in_940),
    .col_in_941(u0_col_in_941),
    .col_in_942(u0_col_in_942),
    .col_in_943(u0_col_in_943),
    .col_in_944(u0_col_in_944),
    .col_in_945(u0_col_in_945),
    .col_in_946(u0_col_in_946),
    .col_in_947(u0_col_in_947),
    .col_in_948(u0_col_in_948),
    .col_in_949(u0_col_in_949),
    .col_in_950(u0_col_in_950),
    .col_in_951(u0_col_in_951),
    .col_in_952(u0_col_in_952),
    .col_in_953(u0_col_in_953),
    .col_in_954(u0_col_in_954),
    .col_in_955(u0_col_in_955),
    .col_in_956(u0_col_in_956),
    .col_in_957(u0_col_in_957),
    .col_in_958(u0_col_in_958),
    .col_in_959(u0_col_in_959),
    .col_in_960(u0_col_in_960),
    .col_in_961(u0_col_in_961),
    .col_in_962(u0_col_in_962),
    .col_in_963(u0_col_in_963),
    .col_in_964(u0_col_in_964),
    .col_in_965(u0_col_in_965),
    .col_in_966(u0_col_in_966),
    .col_in_967(u0_col_in_967),
    .col_in_968(u0_col_in_968),
    .col_in_969(u0_col_in_969),
    .col_in_970(u0_col_in_970),
    .col_in_971(u0_col_in_971),
    .col_in_972(u0_col_in_972),
    .col_in_973(u0_col_in_973),
    .col_in_974(u0_col_in_974),
    .col_in_975(u0_col_in_975),
    .col_in_976(u0_col_in_976),
    .col_in_977(u0_col_in_977),
    .col_in_978(u0_col_in_978),
    .col_in_979(u0_col_in_979),
    .col_in_980(u0_col_in_980),
    .col_in_981(u0_col_in_981),
    .col_in_982(u0_col_in_982),
    .col_in_983(u0_col_in_983),
    .col_in_984(u0_col_in_984),
    .col_in_985(u0_col_in_985),
    .col_in_986(u0_col_in_986),
    .col_in_987(u0_col_in_987),
    .col_in_988(u0_col_in_988),
    .col_in_989(u0_col_in_989),
    .col_in_990(u0_col_in_990),
    .col_in_991(u0_col_in_991),
    .col_in_992(u0_col_in_992),
    .col_in_993(u0_col_in_993),
    .col_in_994(u0_col_in_994),
    .col_in_995(u0_col_in_995),
    .col_in_996(u0_col_in_996),
    .col_in_997(u0_col_in_997),
    .col_in_998(u0_col_in_998),
    .col_in_999(u0_col_in_999),
    .col_in_1000(u0_col_in_1000),
    .col_in_1001(u0_col_in_1001),
    .col_in_1002(u0_col_in_1002),
    .col_in_1003(u0_col_in_1003),
    .col_in_1004(u0_col_in_1004),
    .col_in_1005(u0_col_in_1005),
    .col_in_1006(u0_col_in_1006),
    .col_in_1007(u0_col_in_1007),
    .col_in_1008(u0_col_in_1008),
    .col_in_1009(u0_col_in_1009),
    .col_in_1010(u0_col_in_1010),
    .col_in_1011(u0_col_in_1011),
    .col_in_1012(u0_col_in_1012),
    .col_in_1013(u0_col_in_1013),
    .col_in_1014(u0_col_in_1014),
    .col_in_1015(u0_col_in_1015),
    .col_in_1016(u0_col_in_1016),
    .col_in_1017(u0_col_in_1017),
    .col_in_1018(u0_col_in_1018),
    .col_in_1019(u0_col_in_1019),
    .col_in_1020(u0_col_in_1020),
    .col_in_1021(u0_col_in_1021),
    .col_in_1022(u0_col_in_1022),
    .col_in_1023(u0_col_in_1023),

    .col_out_0(u0_col_out_0),
    .col_out_1(u0_col_out_1),
    .col_out_2(u0_col_out_2),
    .col_out_3(u0_col_out_3),
    .col_out_4(u0_col_out_4),
    .col_out_5(u0_col_out_5),
    .col_out_6(u0_col_out_6),
    .col_out_7(u0_col_out_7),
    .col_out_8(u0_col_out_8),
    .col_out_9(u0_col_out_9),
    .col_out_10(u0_col_out_10),
    .col_out_11(u0_col_out_11),
    .col_out_12(u0_col_out_12),
    .col_out_13(u0_col_out_13),
    .col_out_14(u0_col_out_14),
    .col_out_15(u0_col_out_15),
    .col_out_16(u0_col_out_16),
    .col_out_17(u0_col_out_17),
    .col_out_18(u0_col_out_18),
    .col_out_19(u0_col_out_19),
    .col_out_20(u0_col_out_20),
    .col_out_21(u0_col_out_21),
    .col_out_22(u0_col_out_22),
    .col_out_23(u0_col_out_23),
    .col_out_24(u0_col_out_24),
    .col_out_25(u0_col_out_25),
    .col_out_26(u0_col_out_26),
    .col_out_27(u0_col_out_27),
    .col_out_28(u0_col_out_28),
    .col_out_29(u0_col_out_29),
    .col_out_30(u0_col_out_30),
    .col_out_31(u0_col_out_31),
    .col_out_32(u0_col_out_32),
    .col_out_33(u0_col_out_33),
    .col_out_34(u0_col_out_34),
    .col_out_35(u0_col_out_35),
    .col_out_36(u0_col_out_36),
    .col_out_37(u0_col_out_37),
    .col_out_38(u0_col_out_38),
    .col_out_39(u0_col_out_39),
    .col_out_40(u0_col_out_40),
    .col_out_41(u0_col_out_41),
    .col_out_42(u0_col_out_42),
    .col_out_43(u0_col_out_43),
    .col_out_44(u0_col_out_44),
    .col_out_45(u0_col_out_45),
    .col_out_46(u0_col_out_46),
    .col_out_47(u0_col_out_47),
    .col_out_48(u0_col_out_48),
    .col_out_49(u0_col_out_49),
    .col_out_50(u0_col_out_50),
    .col_out_51(u0_col_out_51),
    .col_out_52(u0_col_out_52),
    .col_out_53(u0_col_out_53),
    .col_out_54(u0_col_out_54),
    .col_out_55(u0_col_out_55),
    .col_out_56(u0_col_out_56),
    .col_out_57(u0_col_out_57),
    .col_out_58(u0_col_out_58),
    .col_out_59(u0_col_out_59),
    .col_out_60(u0_col_out_60),
    .col_out_61(u0_col_out_61),
    .col_out_62(u0_col_out_62),
    .col_out_63(u0_col_out_63),
    .col_out_64(u0_col_out_64),
    .col_out_65(u0_col_out_65),
    .col_out_66(u0_col_out_66),
    .col_out_67(u0_col_out_67),
    .col_out_68(u0_col_out_68),
    .col_out_69(u0_col_out_69),
    .col_out_70(u0_col_out_70),
    .col_out_71(u0_col_out_71),
    .col_out_72(u0_col_out_72),
    .col_out_73(u0_col_out_73),
    .col_out_74(u0_col_out_74),
    .col_out_75(u0_col_out_75),
    .col_out_76(u0_col_out_76),
    .col_out_77(u0_col_out_77),
    .col_out_78(u0_col_out_78),
    .col_out_79(u0_col_out_79),
    .col_out_80(u0_col_out_80),
    .col_out_81(u0_col_out_81),
    .col_out_82(u0_col_out_82),
    .col_out_83(u0_col_out_83),
    .col_out_84(u0_col_out_84),
    .col_out_85(u0_col_out_85),
    .col_out_86(u0_col_out_86),
    .col_out_87(u0_col_out_87),
    .col_out_88(u0_col_out_88),
    .col_out_89(u0_col_out_89),
    .col_out_90(u0_col_out_90),
    .col_out_91(u0_col_out_91),
    .col_out_92(u0_col_out_92),
    .col_out_93(u0_col_out_93),
    .col_out_94(u0_col_out_94),
    .col_out_95(u0_col_out_95),
    .col_out_96(u0_col_out_96),
    .col_out_97(u0_col_out_97),
    .col_out_98(u0_col_out_98),
    .col_out_99(u0_col_out_99),
    .col_out_100(u0_col_out_100),
    .col_out_101(u0_col_out_101),
    .col_out_102(u0_col_out_102),
    .col_out_103(u0_col_out_103),
    .col_out_104(u0_col_out_104),
    .col_out_105(u0_col_out_105),
    .col_out_106(u0_col_out_106),
    .col_out_107(u0_col_out_107),
    .col_out_108(u0_col_out_108),
    .col_out_109(u0_col_out_109),
    .col_out_110(u0_col_out_110),
    .col_out_111(u0_col_out_111),
    .col_out_112(u0_col_out_112),
    .col_out_113(u0_col_out_113),
    .col_out_114(u0_col_out_114),
    .col_out_115(u0_col_out_115),
    .col_out_116(u0_col_out_116),
    .col_out_117(u0_col_out_117),
    .col_out_118(u0_col_out_118),
    .col_out_119(u0_col_out_119),
    .col_out_120(u0_col_out_120),
    .col_out_121(u0_col_out_121),
    .col_out_122(u0_col_out_122),
    .col_out_123(u0_col_out_123),
    .col_out_124(u0_col_out_124),
    .col_out_125(u0_col_out_125),
    .col_out_126(u0_col_out_126),
    .col_out_127(u0_col_out_127),
    .col_out_128(u0_col_out_128),
    .col_out_129(u0_col_out_129),
    .col_out_130(u0_col_out_130),
    .col_out_131(u0_col_out_131),
    .col_out_132(u0_col_out_132),
    .col_out_133(u0_col_out_133),
    .col_out_134(u0_col_out_134),
    .col_out_135(u0_col_out_135),
    .col_out_136(u0_col_out_136),
    .col_out_137(u0_col_out_137),
    .col_out_138(u0_col_out_138),
    .col_out_139(u0_col_out_139),
    .col_out_140(u0_col_out_140),
    .col_out_141(u0_col_out_141),
    .col_out_142(u0_col_out_142),
    .col_out_143(u0_col_out_143),
    .col_out_144(u0_col_out_144),
    .col_out_145(u0_col_out_145),
    .col_out_146(u0_col_out_146),
    .col_out_147(u0_col_out_147),
    .col_out_148(u0_col_out_148),
    .col_out_149(u0_col_out_149),
    .col_out_150(u0_col_out_150),
    .col_out_151(u0_col_out_151),
    .col_out_152(u0_col_out_152),
    .col_out_153(u0_col_out_153),
    .col_out_154(u0_col_out_154),
    .col_out_155(u0_col_out_155),
    .col_out_156(u0_col_out_156),
    .col_out_157(u0_col_out_157),
    .col_out_158(u0_col_out_158),
    .col_out_159(u0_col_out_159),
    .col_out_160(u0_col_out_160),
    .col_out_161(u0_col_out_161),
    .col_out_162(u0_col_out_162),
    .col_out_163(u0_col_out_163),
    .col_out_164(u0_col_out_164),
    .col_out_165(u0_col_out_165),
    .col_out_166(u0_col_out_166),
    .col_out_167(u0_col_out_167),
    .col_out_168(u0_col_out_168),
    .col_out_169(u0_col_out_169),
    .col_out_170(u0_col_out_170),
    .col_out_171(u0_col_out_171),
    .col_out_172(u0_col_out_172),
    .col_out_173(u0_col_out_173),
    .col_out_174(u0_col_out_174),
    .col_out_175(u0_col_out_175),
    .col_out_176(u0_col_out_176),
    .col_out_177(u0_col_out_177),
    .col_out_178(u0_col_out_178),
    .col_out_179(u0_col_out_179),
    .col_out_180(u0_col_out_180),
    .col_out_181(u0_col_out_181),
    .col_out_182(u0_col_out_182),
    .col_out_183(u0_col_out_183),
    .col_out_184(u0_col_out_184),
    .col_out_185(u0_col_out_185),
    .col_out_186(u0_col_out_186),
    .col_out_187(u0_col_out_187),
    .col_out_188(u0_col_out_188),
    .col_out_189(u0_col_out_189),
    .col_out_190(u0_col_out_190),
    .col_out_191(u0_col_out_191),
    .col_out_192(u0_col_out_192),
    .col_out_193(u0_col_out_193),
    .col_out_194(u0_col_out_194),
    .col_out_195(u0_col_out_195),
    .col_out_196(u0_col_out_196),
    .col_out_197(u0_col_out_197),
    .col_out_198(u0_col_out_198),
    .col_out_199(u0_col_out_199),
    .col_out_200(u0_col_out_200),
    .col_out_201(u0_col_out_201),
    .col_out_202(u0_col_out_202),
    .col_out_203(u0_col_out_203),
    .col_out_204(u0_col_out_204),
    .col_out_205(u0_col_out_205),
    .col_out_206(u0_col_out_206),
    .col_out_207(u0_col_out_207),
    .col_out_208(u0_col_out_208),
    .col_out_209(u0_col_out_209),
    .col_out_210(u0_col_out_210),
    .col_out_211(u0_col_out_211),
    .col_out_212(u0_col_out_212),
    .col_out_213(u0_col_out_213),
    .col_out_214(u0_col_out_214),
    .col_out_215(u0_col_out_215),
    .col_out_216(u0_col_out_216),
    .col_out_217(u0_col_out_217),
    .col_out_218(u0_col_out_218),
    .col_out_219(u0_col_out_219),
    .col_out_220(u0_col_out_220),
    .col_out_221(u0_col_out_221),
    .col_out_222(u0_col_out_222),
    .col_out_223(u0_col_out_223),
    .col_out_224(u0_col_out_224),
    .col_out_225(u0_col_out_225),
    .col_out_226(u0_col_out_226),
    .col_out_227(u0_col_out_227),
    .col_out_228(u0_col_out_228),
    .col_out_229(u0_col_out_229),
    .col_out_230(u0_col_out_230),
    .col_out_231(u0_col_out_231),
    .col_out_232(u0_col_out_232),
    .col_out_233(u0_col_out_233),
    .col_out_234(u0_col_out_234),
    .col_out_235(u0_col_out_235),
    .col_out_236(u0_col_out_236),
    .col_out_237(u0_col_out_237),
    .col_out_238(u0_col_out_238),
    .col_out_239(u0_col_out_239),
    .col_out_240(u0_col_out_240),
    .col_out_241(u0_col_out_241),
    .col_out_242(u0_col_out_242),
    .col_out_243(u0_col_out_243),
    .col_out_244(u0_col_out_244),
    .col_out_245(u0_col_out_245),
    .col_out_246(u0_col_out_246),
    .col_out_247(u0_col_out_247),
    .col_out_248(u0_col_out_248),
    .col_out_249(u0_col_out_249),
    .col_out_250(u0_col_out_250),
    .col_out_251(u0_col_out_251),
    .col_out_252(u0_col_out_252),
    .col_out_253(u0_col_out_253),
    .col_out_254(u0_col_out_254),
    .col_out_255(u0_col_out_255),
    .col_out_256(u0_col_out_256),
    .col_out_257(u0_col_out_257),
    .col_out_258(u0_col_out_258),
    .col_out_259(u0_col_out_259),
    .col_out_260(u0_col_out_260),
    .col_out_261(u0_col_out_261),
    .col_out_262(u0_col_out_262),
    .col_out_263(u0_col_out_263),
    .col_out_264(u0_col_out_264),
    .col_out_265(u0_col_out_265),
    .col_out_266(u0_col_out_266),
    .col_out_267(u0_col_out_267),
    .col_out_268(u0_col_out_268),
    .col_out_269(u0_col_out_269),
    .col_out_270(u0_col_out_270),
    .col_out_271(u0_col_out_271),
    .col_out_272(u0_col_out_272),
    .col_out_273(u0_col_out_273),
    .col_out_274(u0_col_out_274),
    .col_out_275(u0_col_out_275),
    .col_out_276(u0_col_out_276),
    .col_out_277(u0_col_out_277),
    .col_out_278(u0_col_out_278),
    .col_out_279(u0_col_out_279),
    .col_out_280(u0_col_out_280),
    .col_out_281(u0_col_out_281),
    .col_out_282(u0_col_out_282),
    .col_out_283(u0_col_out_283),
    .col_out_284(u0_col_out_284),
    .col_out_285(u0_col_out_285),
    .col_out_286(u0_col_out_286),
    .col_out_287(u0_col_out_287),
    .col_out_288(u0_col_out_288),
    .col_out_289(u0_col_out_289),
    .col_out_290(u0_col_out_290),
    .col_out_291(u0_col_out_291),
    .col_out_292(u0_col_out_292),
    .col_out_293(u0_col_out_293),
    .col_out_294(u0_col_out_294),
    .col_out_295(u0_col_out_295),
    .col_out_296(u0_col_out_296),
    .col_out_297(u0_col_out_297),
    .col_out_298(u0_col_out_298),
    .col_out_299(u0_col_out_299),
    .col_out_300(u0_col_out_300),
    .col_out_301(u0_col_out_301),
    .col_out_302(u0_col_out_302),
    .col_out_303(u0_col_out_303),
    .col_out_304(u0_col_out_304),
    .col_out_305(u0_col_out_305),
    .col_out_306(u0_col_out_306),
    .col_out_307(u0_col_out_307),
    .col_out_308(u0_col_out_308),
    .col_out_309(u0_col_out_309),
    .col_out_310(u0_col_out_310),
    .col_out_311(u0_col_out_311),
    .col_out_312(u0_col_out_312),
    .col_out_313(u0_col_out_313),
    .col_out_314(u0_col_out_314),
    .col_out_315(u0_col_out_315),
    .col_out_316(u0_col_out_316),
    .col_out_317(u0_col_out_317),
    .col_out_318(u0_col_out_318),
    .col_out_319(u0_col_out_319),
    .col_out_320(u0_col_out_320),
    .col_out_321(u0_col_out_321),
    .col_out_322(u0_col_out_322),
    .col_out_323(u0_col_out_323),
    .col_out_324(u0_col_out_324),
    .col_out_325(u0_col_out_325),
    .col_out_326(u0_col_out_326),
    .col_out_327(u0_col_out_327),
    .col_out_328(u0_col_out_328),
    .col_out_329(u0_col_out_329),
    .col_out_330(u0_col_out_330),
    .col_out_331(u0_col_out_331),
    .col_out_332(u0_col_out_332),
    .col_out_333(u0_col_out_333),
    .col_out_334(u0_col_out_334),
    .col_out_335(u0_col_out_335),
    .col_out_336(u0_col_out_336),
    .col_out_337(u0_col_out_337),
    .col_out_338(u0_col_out_338),
    .col_out_339(u0_col_out_339),
    .col_out_340(u0_col_out_340),
    .col_out_341(u0_col_out_341),
    .col_out_342(u0_col_out_342),
    .col_out_343(u0_col_out_343),
    .col_out_344(u0_col_out_344),
    .col_out_345(u0_col_out_345),
    .col_out_346(u0_col_out_346),
    .col_out_347(u0_col_out_347),
    .col_out_348(u0_col_out_348),
    .col_out_349(u0_col_out_349),
    .col_out_350(u0_col_out_350),
    .col_out_351(u0_col_out_351),
    .col_out_352(u0_col_out_352),
    .col_out_353(u0_col_out_353),
    .col_out_354(u0_col_out_354),
    .col_out_355(u0_col_out_355),
    .col_out_356(u0_col_out_356),
    .col_out_357(u0_col_out_357),
    .col_out_358(u0_col_out_358),
    .col_out_359(u0_col_out_359),
    .col_out_360(u0_col_out_360),
    .col_out_361(u0_col_out_361),
    .col_out_362(u0_col_out_362),
    .col_out_363(u0_col_out_363),
    .col_out_364(u0_col_out_364),
    .col_out_365(u0_col_out_365),
    .col_out_366(u0_col_out_366),
    .col_out_367(u0_col_out_367),
    .col_out_368(u0_col_out_368),
    .col_out_369(u0_col_out_369),
    .col_out_370(u0_col_out_370),
    .col_out_371(u0_col_out_371),
    .col_out_372(u0_col_out_372),
    .col_out_373(u0_col_out_373),
    .col_out_374(u0_col_out_374),
    .col_out_375(u0_col_out_375),
    .col_out_376(u0_col_out_376),
    .col_out_377(u0_col_out_377),
    .col_out_378(u0_col_out_378),
    .col_out_379(u0_col_out_379),
    .col_out_380(u0_col_out_380),
    .col_out_381(u0_col_out_381),
    .col_out_382(u0_col_out_382),
    .col_out_383(u0_col_out_383),
    .col_out_384(u0_col_out_384),
    .col_out_385(u0_col_out_385),
    .col_out_386(u0_col_out_386),
    .col_out_387(u0_col_out_387),
    .col_out_388(u0_col_out_388),
    .col_out_389(u0_col_out_389),
    .col_out_390(u0_col_out_390),
    .col_out_391(u0_col_out_391),
    .col_out_392(u0_col_out_392),
    .col_out_393(u0_col_out_393),
    .col_out_394(u0_col_out_394),
    .col_out_395(u0_col_out_395),
    .col_out_396(u0_col_out_396),
    .col_out_397(u0_col_out_397),
    .col_out_398(u0_col_out_398),
    .col_out_399(u0_col_out_399),
    .col_out_400(u0_col_out_400),
    .col_out_401(u0_col_out_401),
    .col_out_402(u0_col_out_402),
    .col_out_403(u0_col_out_403),
    .col_out_404(u0_col_out_404),
    .col_out_405(u0_col_out_405),
    .col_out_406(u0_col_out_406),
    .col_out_407(u0_col_out_407),
    .col_out_408(u0_col_out_408),
    .col_out_409(u0_col_out_409),
    .col_out_410(u0_col_out_410),
    .col_out_411(u0_col_out_411),
    .col_out_412(u0_col_out_412),
    .col_out_413(u0_col_out_413),
    .col_out_414(u0_col_out_414),
    .col_out_415(u0_col_out_415),
    .col_out_416(u0_col_out_416),
    .col_out_417(u0_col_out_417),
    .col_out_418(u0_col_out_418),
    .col_out_419(u0_col_out_419),
    .col_out_420(u0_col_out_420),
    .col_out_421(u0_col_out_421),
    .col_out_422(u0_col_out_422),
    .col_out_423(u0_col_out_423),
    .col_out_424(u0_col_out_424),
    .col_out_425(u0_col_out_425),
    .col_out_426(u0_col_out_426),
    .col_out_427(u0_col_out_427),
    .col_out_428(u0_col_out_428),
    .col_out_429(u0_col_out_429),
    .col_out_430(u0_col_out_430),
    .col_out_431(u0_col_out_431),
    .col_out_432(u0_col_out_432),
    .col_out_433(u0_col_out_433),
    .col_out_434(u0_col_out_434),
    .col_out_435(u0_col_out_435),
    .col_out_436(u0_col_out_436),
    .col_out_437(u0_col_out_437),
    .col_out_438(u0_col_out_438),
    .col_out_439(u0_col_out_439),
    .col_out_440(u0_col_out_440),
    .col_out_441(u0_col_out_441),
    .col_out_442(u0_col_out_442),
    .col_out_443(u0_col_out_443),
    .col_out_444(u0_col_out_444),
    .col_out_445(u0_col_out_445),
    .col_out_446(u0_col_out_446),
    .col_out_447(u0_col_out_447),
    .col_out_448(u0_col_out_448),
    .col_out_449(u0_col_out_449),
    .col_out_450(u0_col_out_450),
    .col_out_451(u0_col_out_451),
    .col_out_452(u0_col_out_452),
    .col_out_453(u0_col_out_453),
    .col_out_454(u0_col_out_454),
    .col_out_455(u0_col_out_455),
    .col_out_456(u0_col_out_456),
    .col_out_457(u0_col_out_457),
    .col_out_458(u0_col_out_458),
    .col_out_459(u0_col_out_459),
    .col_out_460(u0_col_out_460),
    .col_out_461(u0_col_out_461),
    .col_out_462(u0_col_out_462),
    .col_out_463(u0_col_out_463),
    .col_out_464(u0_col_out_464),
    .col_out_465(u0_col_out_465),
    .col_out_466(u0_col_out_466),
    .col_out_467(u0_col_out_467),
    .col_out_468(u0_col_out_468),
    .col_out_469(u0_col_out_469),
    .col_out_470(u0_col_out_470),
    .col_out_471(u0_col_out_471),
    .col_out_472(u0_col_out_472),
    .col_out_473(u0_col_out_473),
    .col_out_474(u0_col_out_474),
    .col_out_475(u0_col_out_475),
    .col_out_476(u0_col_out_476),
    .col_out_477(u0_col_out_477),
    .col_out_478(u0_col_out_478),
    .col_out_479(u0_col_out_479),
    .col_out_480(u0_col_out_480),
    .col_out_481(u0_col_out_481),
    .col_out_482(u0_col_out_482),
    .col_out_483(u0_col_out_483),
    .col_out_484(u0_col_out_484),
    .col_out_485(u0_col_out_485),
    .col_out_486(u0_col_out_486),
    .col_out_487(u0_col_out_487),
    .col_out_488(u0_col_out_488),
    .col_out_489(u0_col_out_489),
    .col_out_490(u0_col_out_490),
    .col_out_491(u0_col_out_491),
    .col_out_492(u0_col_out_492),
    .col_out_493(u0_col_out_493),
    .col_out_494(u0_col_out_494),
    .col_out_495(u0_col_out_495),
    .col_out_496(u0_col_out_496),
    .col_out_497(u0_col_out_497),
    .col_out_498(u0_col_out_498),
    .col_out_499(u0_col_out_499),
    .col_out_500(u0_col_out_500),
    .col_out_501(u0_col_out_501),
    .col_out_502(u0_col_out_502),
    .col_out_503(u0_col_out_503),
    .col_out_504(u0_col_out_504),
    .col_out_505(u0_col_out_505),
    .col_out_506(u0_col_out_506),
    .col_out_507(u0_col_out_507),
    .col_out_508(u0_col_out_508),
    .col_out_509(u0_col_out_509),
    .col_out_510(u0_col_out_510),
    .col_out_511(u0_col_out_511),
    .col_out_512(u0_col_out_512),
    .col_out_513(u0_col_out_513),
    .col_out_514(u0_col_out_514),
    .col_out_515(u0_col_out_515),
    .col_out_516(u0_col_out_516),
    .col_out_517(u0_col_out_517),
    .col_out_518(u0_col_out_518),
    .col_out_519(u0_col_out_519),
    .col_out_520(u0_col_out_520),
    .col_out_521(u0_col_out_521),
    .col_out_522(u0_col_out_522),
    .col_out_523(u0_col_out_523),
    .col_out_524(u0_col_out_524),
    .col_out_525(u0_col_out_525),
    .col_out_526(u0_col_out_526),
    .col_out_527(u0_col_out_527),
    .col_out_528(u0_col_out_528),
    .col_out_529(u0_col_out_529),
    .col_out_530(u0_col_out_530),
    .col_out_531(u0_col_out_531),
    .col_out_532(u0_col_out_532),
    .col_out_533(u0_col_out_533),
    .col_out_534(u0_col_out_534),
    .col_out_535(u0_col_out_535),
    .col_out_536(u0_col_out_536),
    .col_out_537(u0_col_out_537),
    .col_out_538(u0_col_out_538),
    .col_out_539(u0_col_out_539),
    .col_out_540(u0_col_out_540),
    .col_out_541(u0_col_out_541),
    .col_out_542(u0_col_out_542),
    .col_out_543(u0_col_out_543),
    .col_out_544(u0_col_out_544),
    .col_out_545(u0_col_out_545),
    .col_out_546(u0_col_out_546),
    .col_out_547(u0_col_out_547),
    .col_out_548(u0_col_out_548),
    .col_out_549(u0_col_out_549),
    .col_out_550(u0_col_out_550),
    .col_out_551(u0_col_out_551),
    .col_out_552(u0_col_out_552),
    .col_out_553(u0_col_out_553),
    .col_out_554(u0_col_out_554),
    .col_out_555(u0_col_out_555),
    .col_out_556(u0_col_out_556),
    .col_out_557(u0_col_out_557),
    .col_out_558(u0_col_out_558),
    .col_out_559(u0_col_out_559),
    .col_out_560(u0_col_out_560),
    .col_out_561(u0_col_out_561),
    .col_out_562(u0_col_out_562),
    .col_out_563(u0_col_out_563),
    .col_out_564(u0_col_out_564),
    .col_out_565(u0_col_out_565),
    .col_out_566(u0_col_out_566),
    .col_out_567(u0_col_out_567),
    .col_out_568(u0_col_out_568),
    .col_out_569(u0_col_out_569),
    .col_out_570(u0_col_out_570),
    .col_out_571(u0_col_out_571),
    .col_out_572(u0_col_out_572),
    .col_out_573(u0_col_out_573),
    .col_out_574(u0_col_out_574),
    .col_out_575(u0_col_out_575),
    .col_out_576(u0_col_out_576),
    .col_out_577(u0_col_out_577),
    .col_out_578(u0_col_out_578),
    .col_out_579(u0_col_out_579),
    .col_out_580(u0_col_out_580),
    .col_out_581(u0_col_out_581),
    .col_out_582(u0_col_out_582),
    .col_out_583(u0_col_out_583),
    .col_out_584(u0_col_out_584),
    .col_out_585(u0_col_out_585),
    .col_out_586(u0_col_out_586),
    .col_out_587(u0_col_out_587),
    .col_out_588(u0_col_out_588),
    .col_out_589(u0_col_out_589),
    .col_out_590(u0_col_out_590),
    .col_out_591(u0_col_out_591),
    .col_out_592(u0_col_out_592),
    .col_out_593(u0_col_out_593),
    .col_out_594(u0_col_out_594),
    .col_out_595(u0_col_out_595),
    .col_out_596(u0_col_out_596),
    .col_out_597(u0_col_out_597),
    .col_out_598(u0_col_out_598),
    .col_out_599(u0_col_out_599),
    .col_out_600(u0_col_out_600),
    .col_out_601(u0_col_out_601),
    .col_out_602(u0_col_out_602),
    .col_out_603(u0_col_out_603),
    .col_out_604(u0_col_out_604),
    .col_out_605(u0_col_out_605),
    .col_out_606(u0_col_out_606),
    .col_out_607(u0_col_out_607),
    .col_out_608(u0_col_out_608),
    .col_out_609(u0_col_out_609),
    .col_out_610(u0_col_out_610),
    .col_out_611(u0_col_out_611),
    .col_out_612(u0_col_out_612),
    .col_out_613(u0_col_out_613),
    .col_out_614(u0_col_out_614),
    .col_out_615(u0_col_out_615),
    .col_out_616(u0_col_out_616),
    .col_out_617(u0_col_out_617),
    .col_out_618(u0_col_out_618),
    .col_out_619(u0_col_out_619),
    .col_out_620(u0_col_out_620),
    .col_out_621(u0_col_out_621),
    .col_out_622(u0_col_out_622),
    .col_out_623(u0_col_out_623),
    .col_out_624(u0_col_out_624),
    .col_out_625(u0_col_out_625),
    .col_out_626(u0_col_out_626),
    .col_out_627(u0_col_out_627),
    .col_out_628(u0_col_out_628),
    .col_out_629(u0_col_out_629),
    .col_out_630(u0_col_out_630),
    .col_out_631(u0_col_out_631),
    .col_out_632(u0_col_out_632),
    .col_out_633(u0_col_out_633),
    .col_out_634(u0_col_out_634),
    .col_out_635(u0_col_out_635),
    .col_out_636(u0_col_out_636),
    .col_out_637(u0_col_out_637),
    .col_out_638(u0_col_out_638),
    .col_out_639(u0_col_out_639),
    .col_out_640(u0_col_out_640),
    .col_out_641(u0_col_out_641),
    .col_out_642(u0_col_out_642),
    .col_out_643(u0_col_out_643),
    .col_out_644(u0_col_out_644),
    .col_out_645(u0_col_out_645),
    .col_out_646(u0_col_out_646),
    .col_out_647(u0_col_out_647),
    .col_out_648(u0_col_out_648),
    .col_out_649(u0_col_out_649),
    .col_out_650(u0_col_out_650),
    .col_out_651(u0_col_out_651),
    .col_out_652(u0_col_out_652),
    .col_out_653(u0_col_out_653),
    .col_out_654(u0_col_out_654),
    .col_out_655(u0_col_out_655),
    .col_out_656(u0_col_out_656),
    .col_out_657(u0_col_out_657),
    .col_out_658(u0_col_out_658),
    .col_out_659(u0_col_out_659),
    .col_out_660(u0_col_out_660),
    .col_out_661(u0_col_out_661),
    .col_out_662(u0_col_out_662),
    .col_out_663(u0_col_out_663),
    .col_out_664(u0_col_out_664),
    .col_out_665(u0_col_out_665),
    .col_out_666(u0_col_out_666),
    .col_out_667(u0_col_out_667),
    .col_out_668(u0_col_out_668),
    .col_out_669(u0_col_out_669),
    .col_out_670(u0_col_out_670),
    .col_out_671(u0_col_out_671),
    .col_out_672(u0_col_out_672),
    .col_out_673(u0_col_out_673),
    .col_out_674(u0_col_out_674),
    .col_out_675(u0_col_out_675),
    .col_out_676(u0_col_out_676),
    .col_out_677(u0_col_out_677),
    .col_out_678(u0_col_out_678),
    .col_out_679(u0_col_out_679),
    .col_out_680(u0_col_out_680),
    .col_out_681(u0_col_out_681),
    .col_out_682(u0_col_out_682),
    .col_out_683(u0_col_out_683),
    .col_out_684(u0_col_out_684),
    .col_out_685(u0_col_out_685),
    .col_out_686(u0_col_out_686),
    .col_out_687(u0_col_out_687),
    .col_out_688(u0_col_out_688),
    .col_out_689(u0_col_out_689),
    .col_out_690(u0_col_out_690),
    .col_out_691(u0_col_out_691),
    .col_out_692(u0_col_out_692),
    .col_out_693(u0_col_out_693),
    .col_out_694(u0_col_out_694),
    .col_out_695(u0_col_out_695),
    .col_out_696(u0_col_out_696),
    .col_out_697(u0_col_out_697),
    .col_out_698(u0_col_out_698),
    .col_out_699(u0_col_out_699),
    .col_out_700(u0_col_out_700),
    .col_out_701(u0_col_out_701),
    .col_out_702(u0_col_out_702),
    .col_out_703(u0_col_out_703),
    .col_out_704(u0_col_out_704),
    .col_out_705(u0_col_out_705),
    .col_out_706(u0_col_out_706),
    .col_out_707(u0_col_out_707),
    .col_out_708(u0_col_out_708),
    .col_out_709(u0_col_out_709),
    .col_out_710(u0_col_out_710),
    .col_out_711(u0_col_out_711),
    .col_out_712(u0_col_out_712),
    .col_out_713(u0_col_out_713),
    .col_out_714(u0_col_out_714),
    .col_out_715(u0_col_out_715),
    .col_out_716(u0_col_out_716),
    .col_out_717(u0_col_out_717),
    .col_out_718(u0_col_out_718),
    .col_out_719(u0_col_out_719),
    .col_out_720(u0_col_out_720),
    .col_out_721(u0_col_out_721),
    .col_out_722(u0_col_out_722),
    .col_out_723(u0_col_out_723),
    .col_out_724(u0_col_out_724),
    .col_out_725(u0_col_out_725),
    .col_out_726(u0_col_out_726),
    .col_out_727(u0_col_out_727),
    .col_out_728(u0_col_out_728),
    .col_out_729(u0_col_out_729),
    .col_out_730(u0_col_out_730),
    .col_out_731(u0_col_out_731),
    .col_out_732(u0_col_out_732),
    .col_out_733(u0_col_out_733),
    .col_out_734(u0_col_out_734),
    .col_out_735(u0_col_out_735),
    .col_out_736(u0_col_out_736),
    .col_out_737(u0_col_out_737),
    .col_out_738(u0_col_out_738),
    .col_out_739(u0_col_out_739),
    .col_out_740(u0_col_out_740),
    .col_out_741(u0_col_out_741),
    .col_out_742(u0_col_out_742),
    .col_out_743(u0_col_out_743),
    .col_out_744(u0_col_out_744),
    .col_out_745(u0_col_out_745),
    .col_out_746(u0_col_out_746),
    .col_out_747(u0_col_out_747),
    .col_out_748(u0_col_out_748),
    .col_out_749(u0_col_out_749),
    .col_out_750(u0_col_out_750),
    .col_out_751(u0_col_out_751),
    .col_out_752(u0_col_out_752),
    .col_out_753(u0_col_out_753),
    .col_out_754(u0_col_out_754),
    .col_out_755(u0_col_out_755),
    .col_out_756(u0_col_out_756),
    .col_out_757(u0_col_out_757),
    .col_out_758(u0_col_out_758),
    .col_out_759(u0_col_out_759),
    .col_out_760(u0_col_out_760),
    .col_out_761(u0_col_out_761),
    .col_out_762(u0_col_out_762),
    .col_out_763(u0_col_out_763),
    .col_out_764(u0_col_out_764),
    .col_out_765(u0_col_out_765),
    .col_out_766(u0_col_out_766),
    .col_out_767(u0_col_out_767),
    .col_out_768(u0_col_out_768),
    .col_out_769(u0_col_out_769),
    .col_out_770(u0_col_out_770),
    .col_out_771(u0_col_out_771),
    .col_out_772(u0_col_out_772),
    .col_out_773(u0_col_out_773),
    .col_out_774(u0_col_out_774),
    .col_out_775(u0_col_out_775),
    .col_out_776(u0_col_out_776),
    .col_out_777(u0_col_out_777),
    .col_out_778(u0_col_out_778),
    .col_out_779(u0_col_out_779),
    .col_out_780(u0_col_out_780),
    .col_out_781(u0_col_out_781),
    .col_out_782(u0_col_out_782),
    .col_out_783(u0_col_out_783),
    .col_out_784(u0_col_out_784),
    .col_out_785(u0_col_out_785),
    .col_out_786(u0_col_out_786),
    .col_out_787(u0_col_out_787),
    .col_out_788(u0_col_out_788),
    .col_out_789(u0_col_out_789),
    .col_out_790(u0_col_out_790),
    .col_out_791(u0_col_out_791),
    .col_out_792(u0_col_out_792),
    .col_out_793(u0_col_out_793),
    .col_out_794(u0_col_out_794),
    .col_out_795(u0_col_out_795),
    .col_out_796(u0_col_out_796),
    .col_out_797(u0_col_out_797),
    .col_out_798(u0_col_out_798),
    .col_out_799(u0_col_out_799),
    .col_out_800(u0_col_out_800),
    .col_out_801(u0_col_out_801),
    .col_out_802(u0_col_out_802),
    .col_out_803(u0_col_out_803),
    .col_out_804(u0_col_out_804),
    .col_out_805(u0_col_out_805),
    .col_out_806(u0_col_out_806),
    .col_out_807(u0_col_out_807),
    .col_out_808(u0_col_out_808),
    .col_out_809(u0_col_out_809),
    .col_out_810(u0_col_out_810),
    .col_out_811(u0_col_out_811),
    .col_out_812(u0_col_out_812),
    .col_out_813(u0_col_out_813),
    .col_out_814(u0_col_out_814),
    .col_out_815(u0_col_out_815),
    .col_out_816(u0_col_out_816),
    .col_out_817(u0_col_out_817),
    .col_out_818(u0_col_out_818),
    .col_out_819(u0_col_out_819),
    .col_out_820(u0_col_out_820),
    .col_out_821(u0_col_out_821),
    .col_out_822(u0_col_out_822),
    .col_out_823(u0_col_out_823),
    .col_out_824(u0_col_out_824),
    .col_out_825(u0_col_out_825),
    .col_out_826(u0_col_out_826),
    .col_out_827(u0_col_out_827),
    .col_out_828(u0_col_out_828),
    .col_out_829(u0_col_out_829),
    .col_out_830(u0_col_out_830),
    .col_out_831(u0_col_out_831),
    .col_out_832(u0_col_out_832),
    .col_out_833(u0_col_out_833),
    .col_out_834(u0_col_out_834),
    .col_out_835(u0_col_out_835),
    .col_out_836(u0_col_out_836),
    .col_out_837(u0_col_out_837),
    .col_out_838(u0_col_out_838),
    .col_out_839(u0_col_out_839),
    .col_out_840(u0_col_out_840),
    .col_out_841(u0_col_out_841),
    .col_out_842(u0_col_out_842),
    .col_out_843(u0_col_out_843),
    .col_out_844(u0_col_out_844),
    .col_out_845(u0_col_out_845),
    .col_out_846(u0_col_out_846),
    .col_out_847(u0_col_out_847),
    .col_out_848(u0_col_out_848),
    .col_out_849(u0_col_out_849),
    .col_out_850(u0_col_out_850),
    .col_out_851(u0_col_out_851),
    .col_out_852(u0_col_out_852),
    .col_out_853(u0_col_out_853),
    .col_out_854(u0_col_out_854),
    .col_out_855(u0_col_out_855),
    .col_out_856(u0_col_out_856),
    .col_out_857(u0_col_out_857),
    .col_out_858(u0_col_out_858),
    .col_out_859(u0_col_out_859),
    .col_out_860(u0_col_out_860),
    .col_out_861(u0_col_out_861),
    .col_out_862(u0_col_out_862),
    .col_out_863(u0_col_out_863),
    .col_out_864(u0_col_out_864),
    .col_out_865(u0_col_out_865),
    .col_out_866(u0_col_out_866),
    .col_out_867(u0_col_out_867),
    .col_out_868(u0_col_out_868),
    .col_out_869(u0_col_out_869),
    .col_out_870(u0_col_out_870),
    .col_out_871(u0_col_out_871),
    .col_out_872(u0_col_out_872),
    .col_out_873(u0_col_out_873),
    .col_out_874(u0_col_out_874),
    .col_out_875(u0_col_out_875),
    .col_out_876(u0_col_out_876),
    .col_out_877(u0_col_out_877),
    .col_out_878(u0_col_out_878),
    .col_out_879(u0_col_out_879),
    .col_out_880(u0_col_out_880),
    .col_out_881(u0_col_out_881),
    .col_out_882(u0_col_out_882),
    .col_out_883(u0_col_out_883),
    .col_out_884(u0_col_out_884),
    .col_out_885(u0_col_out_885),
    .col_out_886(u0_col_out_886),
    .col_out_887(u0_col_out_887),
    .col_out_888(u0_col_out_888),
    .col_out_889(u0_col_out_889),
    .col_out_890(u0_col_out_890),
    .col_out_891(u0_col_out_891),
    .col_out_892(u0_col_out_892),
    .col_out_893(u0_col_out_893),
    .col_out_894(u0_col_out_894),
    .col_out_895(u0_col_out_895),
    .col_out_896(u0_col_out_896),
    .col_out_897(u0_col_out_897),
    .col_out_898(u0_col_out_898),
    .col_out_899(u0_col_out_899),
    .col_out_900(u0_col_out_900),
    .col_out_901(u0_col_out_901),
    .col_out_902(u0_col_out_902),
    .col_out_903(u0_col_out_903),
    .col_out_904(u0_col_out_904),
    .col_out_905(u0_col_out_905),
    .col_out_906(u0_col_out_906),
    .col_out_907(u0_col_out_907),
    .col_out_908(u0_col_out_908),
    .col_out_909(u0_col_out_909),
    .col_out_910(u0_col_out_910),
    .col_out_911(u0_col_out_911),
    .col_out_912(u0_col_out_912),
    .col_out_913(u0_col_out_913),
    .col_out_914(u0_col_out_914),
    .col_out_915(u0_col_out_915),
    .col_out_916(u0_col_out_916),
    .col_out_917(u0_col_out_917),
    .col_out_918(u0_col_out_918),
    .col_out_919(u0_col_out_919),
    .col_out_920(u0_col_out_920),
    .col_out_921(u0_col_out_921),
    .col_out_922(u0_col_out_922),
    .col_out_923(u0_col_out_923),
    .col_out_924(u0_col_out_924),
    .col_out_925(u0_col_out_925),
    .col_out_926(u0_col_out_926),
    .col_out_927(u0_col_out_927),
    .col_out_928(u0_col_out_928),
    .col_out_929(u0_col_out_929),
    .col_out_930(u0_col_out_930),
    .col_out_931(u0_col_out_931),
    .col_out_932(u0_col_out_932),
    .col_out_933(u0_col_out_933),
    .col_out_934(u0_col_out_934),
    .col_out_935(u0_col_out_935),
    .col_out_936(u0_col_out_936),
    .col_out_937(u0_col_out_937),
    .col_out_938(u0_col_out_938),
    .col_out_939(u0_col_out_939),
    .col_out_940(u0_col_out_940),
    .col_out_941(u0_col_out_941),
    .col_out_942(u0_col_out_942),
    .col_out_943(u0_col_out_943),
    .col_out_944(u0_col_out_944),
    .col_out_945(u0_col_out_945),
    .col_out_946(u0_col_out_946),
    .col_out_947(u0_col_out_947),
    .col_out_948(u0_col_out_948),
    .col_out_949(u0_col_out_949),
    .col_out_950(u0_col_out_950),
    .col_out_951(u0_col_out_951),
    .col_out_952(u0_col_out_952),
    .col_out_953(u0_col_out_953),
    .col_out_954(u0_col_out_954),
    .col_out_955(u0_col_out_955),
    .col_out_956(u0_col_out_956),
    .col_out_957(u0_col_out_957),
    .col_out_958(u0_col_out_958),
    .col_out_959(u0_col_out_959),
    .col_out_960(u0_col_out_960),
    .col_out_961(u0_col_out_961),
    .col_out_962(u0_col_out_962),
    .col_out_963(u0_col_out_963),
    .col_out_964(u0_col_out_964),
    .col_out_965(u0_col_out_965),
    .col_out_966(u0_col_out_966),
    .col_out_967(u0_col_out_967),
    .col_out_968(u0_col_out_968),
    .col_out_969(u0_col_out_969),
    .col_out_970(u0_col_out_970),
    .col_out_971(u0_col_out_971),
    .col_out_972(u0_col_out_972),
    .col_out_973(u0_col_out_973),
    .col_out_974(u0_col_out_974),
    .col_out_975(u0_col_out_975),
    .col_out_976(u0_col_out_976),
    .col_out_977(u0_col_out_977),
    .col_out_978(u0_col_out_978),
    .col_out_979(u0_col_out_979),
    .col_out_980(u0_col_out_980),
    .col_out_981(u0_col_out_981),
    .col_out_982(u0_col_out_982),
    .col_out_983(u0_col_out_983),
    .col_out_984(u0_col_out_984),
    .col_out_985(u0_col_out_985),
    .col_out_986(u0_col_out_986),
    .col_out_987(u0_col_out_987),
    .col_out_988(u0_col_out_988),
    .col_out_989(u0_col_out_989),
    .col_out_990(u0_col_out_990),
    .col_out_991(u0_col_out_991),
    .col_out_992(u0_col_out_992),
    .col_out_993(u0_col_out_993),
    .col_out_994(u0_col_out_994),
    .col_out_995(u0_col_out_995),
    .col_out_996(u0_col_out_996),
    .col_out_997(u0_col_out_997),
    .col_out_998(u0_col_out_998),
    .col_out_999(u0_col_out_999),
    .col_out_1000(u0_col_out_1000),
    .col_out_1001(u0_col_out_1001),
    .col_out_1002(u0_col_out_1002),
    .col_out_1003(u0_col_out_1003),
    .col_out_1004(u0_col_out_1004),
    .col_out_1005(u0_col_out_1005),
    .col_out_1006(u0_col_out_1006),
    .col_out_1007(u0_col_out_1007),
    .col_out_1008(u0_col_out_1008),
    .col_out_1009(u0_col_out_1009),
    .col_out_1010(u0_col_out_1010),
    .col_out_1011(u0_col_out_1011),
    .col_out_1012(u0_col_out_1012),
    .col_out_1013(u0_col_out_1013),
    .col_out_1014(u0_col_out_1014),
    .col_out_1015(u0_col_out_1015),
    .col_out_1016(u0_col_out_1016),
    .col_out_1017(u0_col_out_1017),
    .col_out_1018(u0_col_out_1018),
    .col_out_1019(u0_col_out_1019),
    .col_out_1020(u0_col_out_1020),
    .col_out_1021(u0_col_out_1021),
    .col_out_1022(u0_col_out_1022),
    .col_out_1023(u0_col_out_1023),
    .col_out_1024(u0_col_out_1024),
    .col_out_1025(u0_col_out_1025),
    .col_out_1026(u0_col_out_1026)
);
















//*****************************************************
//**************u1输入定义******************************
//*****************************************************
wire [151:0] u1_col_in_0;
wire [151:0] u1_col_in_1;
wire [151:0] u1_col_in_2;
wire [151:0] u1_col_in_3;
wire [151:0] u1_col_in_4;
wire [151:0] u1_col_in_5;
wire [151:0] u1_col_in_6;
wire [151:0] u1_col_in_7;
wire [151:0] u1_col_in_8;
wire [151:0] u1_col_in_9;
wire [151:0] u1_col_in_10;
wire [151:0] u1_col_in_11;
wire [151:0] u1_col_in_12;
wire [151:0] u1_col_in_13;
wire [151:0] u1_col_in_14;
wire [151:0] u1_col_in_15;
wire [151:0] u1_col_in_16;
wire [151:0] u1_col_in_17;
wire [151:0] u1_col_in_18;
wire [151:0] u1_col_in_19;
wire [151:0] u1_col_in_20;
wire [151:0] u1_col_in_21;
wire [151:0] u1_col_in_22;
wire [151:0] u1_col_in_23;
wire [151:0] u1_col_in_24;
wire [151:0] u1_col_in_25;
wire [151:0] u1_col_in_26;
wire [151:0] u1_col_in_27;
wire [151:0] u1_col_in_28;
wire [151:0] u1_col_in_29;
wire [151:0] u1_col_in_30;
wire [151:0] u1_col_in_31;
wire [151:0] u1_col_in_32;
wire [151:0] u1_col_in_33;
wire [151:0] u1_col_in_34;
wire [151:0] u1_col_in_35;
wire [151:0] u1_col_in_36;
wire [151:0] u1_col_in_37;
wire [151:0] u1_col_in_38;
wire [151:0] u1_col_in_39;
wire [151:0] u1_col_in_40;
wire [151:0] u1_col_in_41;
wire [151:0] u1_col_in_42;
wire [151:0] u1_col_in_43;
wire [151:0] u1_col_in_44;
wire [151:0] u1_col_in_45;
wire [151:0] u1_col_in_46;
wire [151:0] u1_col_in_47;
wire [151:0] u1_col_in_48;
wire [151:0] u1_col_in_49;
wire [151:0] u1_col_in_50;
wire [151:0] u1_col_in_51;
wire [151:0] u1_col_in_52;
wire [151:0] u1_col_in_53;
wire [151:0] u1_col_in_54;
wire [151:0] u1_col_in_55;
wire [151:0] u1_col_in_56;
wire [151:0] u1_col_in_57;
wire [151:0] u1_col_in_58;
wire [151:0] u1_col_in_59;
wire [151:0] u1_col_in_60;
wire [151:0] u1_col_in_61;
wire [151:0] u1_col_in_62;
wire [151:0] u1_col_in_63;
wire [151:0] u1_col_in_64;
wire [151:0] u1_col_in_65;
wire [151:0] u1_col_in_66;
wire [151:0] u1_col_in_67;
wire [151:0] u1_col_in_68;
wire [151:0] u1_col_in_69;
wire [151:0] u1_col_in_70;
wire [151:0] u1_col_in_71;
wire [151:0] u1_col_in_72;
wire [151:0] u1_col_in_73;
wire [151:0] u1_col_in_74;
wire [151:0] u1_col_in_75;
wire [151:0] u1_col_in_76;
wire [151:0] u1_col_in_77;
wire [151:0] u1_col_in_78;
wire [151:0] u1_col_in_79;
wire [151:0] u1_col_in_80;
wire [151:0] u1_col_in_81;
wire [151:0] u1_col_in_82;
wire [151:0] u1_col_in_83;
wire [151:0] u1_col_in_84;
wire [151:0] u1_col_in_85;
wire [151:0] u1_col_in_86;
wire [151:0] u1_col_in_87;
wire [151:0] u1_col_in_88;
wire [151:0] u1_col_in_89;
wire [151:0] u1_col_in_90;
wire [151:0] u1_col_in_91;
wire [151:0] u1_col_in_92;
wire [151:0] u1_col_in_93;
wire [151:0] u1_col_in_94;
wire [151:0] u1_col_in_95;
wire [151:0] u1_col_in_96;
wire [151:0] u1_col_in_97;
wire [151:0] u1_col_in_98;
wire [151:0] u1_col_in_99;
wire [151:0] u1_col_in_100;
wire [151:0] u1_col_in_101;
wire [151:0] u1_col_in_102;
wire [151:0] u1_col_in_103;
wire [151:0] u1_col_in_104;
wire [151:0] u1_col_in_105;
wire [151:0] u1_col_in_106;
wire [151:0] u1_col_in_107;
wire [151:0] u1_col_in_108;
wire [151:0] u1_col_in_109;
wire [151:0] u1_col_in_110;
wire [151:0] u1_col_in_111;
wire [151:0] u1_col_in_112;
wire [151:0] u1_col_in_113;
wire [151:0] u1_col_in_114;
wire [151:0] u1_col_in_115;
wire [151:0] u1_col_in_116;
wire [151:0] u1_col_in_117;
wire [151:0] u1_col_in_118;
wire [151:0] u1_col_in_119;
wire [151:0] u1_col_in_120;
wire [151:0] u1_col_in_121;
wire [151:0] u1_col_in_122;
wire [151:0] u1_col_in_123;
wire [151:0] u1_col_in_124;
wire [151:0] u1_col_in_125;
wire [151:0] u1_col_in_126;
wire [151:0] u1_col_in_127;
wire [151:0] u1_col_in_128;
wire [151:0] u1_col_in_129;
wire [151:0] u1_col_in_130;
wire [151:0] u1_col_in_131;
wire [151:0] u1_col_in_132;
wire [151:0] u1_col_in_133;
wire [151:0] u1_col_in_134;
wire [151:0] u1_col_in_135;
wire [151:0] u1_col_in_136;
wire [151:0] u1_col_in_137;
wire [151:0] u1_col_in_138;
wire [151:0] u1_col_in_139;
wire [151:0] u1_col_in_140;
wire [151:0] u1_col_in_141;
wire [151:0] u1_col_in_142;
wire [151:0] u1_col_in_143;
wire [151:0] u1_col_in_144;
wire [151:0] u1_col_in_145;
wire [151:0] u1_col_in_146;
wire [151:0] u1_col_in_147;
wire [151:0] u1_col_in_148;
wire [151:0] u1_col_in_149;
wire [151:0] u1_col_in_150;
wire [151:0] u1_col_in_151;
wire [151:0] u1_col_in_152;
wire [151:0] u1_col_in_153;
wire [151:0] u1_col_in_154;
wire [151:0] u1_col_in_155;
wire [151:0] u1_col_in_156;
wire [151:0] u1_col_in_157;
wire [151:0] u1_col_in_158;
wire [151:0] u1_col_in_159;
wire [151:0] u1_col_in_160;
wire [151:0] u1_col_in_161;
wire [151:0] u1_col_in_162;
wire [151:0] u1_col_in_163;
wire [151:0] u1_col_in_164;
wire [151:0] u1_col_in_165;
wire [151:0] u1_col_in_166;
wire [151:0] u1_col_in_167;
wire [151:0] u1_col_in_168;
wire [151:0] u1_col_in_169;
wire [151:0] u1_col_in_170;
wire [151:0] u1_col_in_171;
wire [151:0] u1_col_in_172;
wire [151:0] u1_col_in_173;
wire [151:0] u1_col_in_174;
wire [151:0] u1_col_in_175;
wire [151:0] u1_col_in_176;
wire [151:0] u1_col_in_177;
wire [151:0] u1_col_in_178;
wire [151:0] u1_col_in_179;
wire [151:0] u1_col_in_180;
wire [151:0] u1_col_in_181;
wire [151:0] u1_col_in_182;
wire [151:0] u1_col_in_183;
wire [151:0] u1_col_in_184;
wire [151:0] u1_col_in_185;
wire [151:0] u1_col_in_186;
wire [151:0] u1_col_in_187;
wire [151:0] u1_col_in_188;
wire [151:0] u1_col_in_189;
wire [151:0] u1_col_in_190;
wire [151:0] u1_col_in_191;
wire [151:0] u1_col_in_192;
wire [151:0] u1_col_in_193;
wire [151:0] u1_col_in_194;
wire [151:0] u1_col_in_195;
wire [151:0] u1_col_in_196;
wire [151:0] u1_col_in_197;
wire [151:0] u1_col_in_198;
wire [151:0] u1_col_in_199;
wire [151:0] u1_col_in_200;
wire [151:0] u1_col_in_201;
wire [151:0] u1_col_in_202;
wire [151:0] u1_col_in_203;
wire [151:0] u1_col_in_204;
wire [151:0] u1_col_in_205;
wire [151:0] u1_col_in_206;
wire [151:0] u1_col_in_207;
wire [151:0] u1_col_in_208;
wire [151:0] u1_col_in_209;
wire [151:0] u1_col_in_210;
wire [151:0] u1_col_in_211;
wire [151:0] u1_col_in_212;
wire [151:0] u1_col_in_213;
wire [151:0] u1_col_in_214;
wire [151:0] u1_col_in_215;
wire [151:0] u1_col_in_216;
wire [151:0] u1_col_in_217;
wire [151:0] u1_col_in_218;
wire [151:0] u1_col_in_219;
wire [151:0] u1_col_in_220;
wire [151:0] u1_col_in_221;
wire [151:0] u1_col_in_222;
wire [151:0] u1_col_in_223;
wire [151:0] u1_col_in_224;
wire [151:0] u1_col_in_225;
wire [151:0] u1_col_in_226;
wire [151:0] u1_col_in_227;
wire [151:0] u1_col_in_228;
wire [151:0] u1_col_in_229;
wire [151:0] u1_col_in_230;
wire [151:0] u1_col_in_231;
wire [151:0] u1_col_in_232;
wire [151:0] u1_col_in_233;
wire [151:0] u1_col_in_234;
wire [151:0] u1_col_in_235;
wire [151:0] u1_col_in_236;
wire [151:0] u1_col_in_237;
wire [151:0] u1_col_in_238;
wire [151:0] u1_col_in_239;
wire [151:0] u1_col_in_240;
wire [151:0] u1_col_in_241;
wire [151:0] u1_col_in_242;
wire [151:0] u1_col_in_243;
wire [151:0] u1_col_in_244;
wire [151:0] u1_col_in_245;
wire [151:0] u1_col_in_246;
wire [151:0] u1_col_in_247;
wire [151:0] u1_col_in_248;
wire [151:0] u1_col_in_249;
wire [151:0] u1_col_in_250;
wire [151:0] u1_col_in_251;
wire [151:0] u1_col_in_252;
wire [151:0] u1_col_in_253;
wire [151:0] u1_col_in_254;
wire [151:0] u1_col_in_255;
wire [151:0] u1_col_in_256;
wire [151:0] u1_col_in_257;
wire [151:0] u1_col_in_258;
wire [151:0] u1_col_in_259;
wire [151:0] u1_col_in_260;
wire [151:0] u1_col_in_261;
wire [151:0] u1_col_in_262;
wire [151:0] u1_col_in_263;
wire [151:0] u1_col_in_264;
wire [151:0] u1_col_in_265;
wire [151:0] u1_col_in_266;
wire [151:0] u1_col_in_267;
wire [151:0] u1_col_in_268;
wire [151:0] u1_col_in_269;
wire [151:0] u1_col_in_270;
wire [151:0] u1_col_in_271;
wire [151:0] u1_col_in_272;
wire [151:0] u1_col_in_273;
wire [151:0] u1_col_in_274;
wire [151:0] u1_col_in_275;
wire [151:0] u1_col_in_276;
wire [151:0] u1_col_in_277;
wire [151:0] u1_col_in_278;
wire [151:0] u1_col_in_279;
wire [151:0] u1_col_in_280;
wire [151:0] u1_col_in_281;
wire [151:0] u1_col_in_282;
wire [151:0] u1_col_in_283;
wire [151:0] u1_col_in_284;
wire [151:0] u1_col_in_285;
wire [151:0] u1_col_in_286;
wire [151:0] u1_col_in_287;
wire [151:0] u1_col_in_288;
wire [151:0] u1_col_in_289;
wire [151:0] u1_col_in_290;
wire [151:0] u1_col_in_291;
wire [151:0] u1_col_in_292;
wire [151:0] u1_col_in_293;
wire [151:0] u1_col_in_294;
wire [151:0] u1_col_in_295;
wire [151:0] u1_col_in_296;
wire [151:0] u1_col_in_297;
wire [151:0] u1_col_in_298;
wire [151:0] u1_col_in_299;
wire [151:0] u1_col_in_300;
wire [151:0] u1_col_in_301;
wire [151:0] u1_col_in_302;
wire [151:0] u1_col_in_303;
wire [151:0] u1_col_in_304;
wire [151:0] u1_col_in_305;
wire [151:0] u1_col_in_306;
wire [151:0] u1_col_in_307;
wire [151:0] u1_col_in_308;
wire [151:0] u1_col_in_309;
wire [151:0] u1_col_in_310;
wire [151:0] u1_col_in_311;
wire [151:0] u1_col_in_312;
wire [151:0] u1_col_in_313;
wire [151:0] u1_col_in_314;
wire [151:0] u1_col_in_315;
wire [151:0] u1_col_in_316;
wire [151:0] u1_col_in_317;
wire [151:0] u1_col_in_318;
wire [151:0] u1_col_in_319;
wire [151:0] u1_col_in_320;
wire [151:0] u1_col_in_321;
wire [151:0] u1_col_in_322;
wire [151:0] u1_col_in_323;
wire [151:0] u1_col_in_324;
wire [151:0] u1_col_in_325;
wire [151:0] u1_col_in_326;
wire [151:0] u1_col_in_327;
wire [151:0] u1_col_in_328;
wire [151:0] u1_col_in_329;
wire [151:0] u1_col_in_330;
wire [151:0] u1_col_in_331;
wire [151:0] u1_col_in_332;
wire [151:0] u1_col_in_333;
wire [151:0] u1_col_in_334;
wire [151:0] u1_col_in_335;
wire [151:0] u1_col_in_336;
wire [151:0] u1_col_in_337;
wire [151:0] u1_col_in_338;
wire [151:0] u1_col_in_339;
wire [151:0] u1_col_in_340;
wire [151:0] u1_col_in_341;
wire [151:0] u1_col_in_342;
wire [151:0] u1_col_in_343;
wire [151:0] u1_col_in_344;
wire [151:0] u1_col_in_345;
wire [151:0] u1_col_in_346;
wire [151:0] u1_col_in_347;
wire [151:0] u1_col_in_348;
wire [151:0] u1_col_in_349;
wire [151:0] u1_col_in_350;
wire [151:0] u1_col_in_351;
wire [151:0] u1_col_in_352;
wire [151:0] u1_col_in_353;
wire [151:0] u1_col_in_354;
wire [151:0] u1_col_in_355;
wire [151:0] u1_col_in_356;
wire [151:0] u1_col_in_357;
wire [151:0] u1_col_in_358;
wire [151:0] u1_col_in_359;
wire [151:0] u1_col_in_360;
wire [151:0] u1_col_in_361;
wire [151:0] u1_col_in_362;
wire [151:0] u1_col_in_363;
wire [151:0] u1_col_in_364;
wire [151:0] u1_col_in_365;
wire [151:0] u1_col_in_366;
wire [151:0] u1_col_in_367;
wire [151:0] u1_col_in_368;
wire [151:0] u1_col_in_369;
wire [151:0] u1_col_in_370;
wire [151:0] u1_col_in_371;
wire [151:0] u1_col_in_372;
wire [151:0] u1_col_in_373;
wire [151:0] u1_col_in_374;
wire [151:0] u1_col_in_375;
wire [151:0] u1_col_in_376;
wire [151:0] u1_col_in_377;
wire [151:0] u1_col_in_378;
wire [151:0] u1_col_in_379;
wire [151:0] u1_col_in_380;
wire [151:0] u1_col_in_381;
wire [151:0] u1_col_in_382;
wire [151:0] u1_col_in_383;
wire [151:0] u1_col_in_384;
wire [151:0] u1_col_in_385;
wire [151:0] u1_col_in_386;
wire [151:0] u1_col_in_387;
wire [151:0] u1_col_in_388;
wire [151:0] u1_col_in_389;
wire [151:0] u1_col_in_390;
wire [151:0] u1_col_in_391;
wire [151:0] u1_col_in_392;
wire [151:0] u1_col_in_393;
wire [151:0] u1_col_in_394;
wire [151:0] u1_col_in_395;
wire [151:0] u1_col_in_396;
wire [151:0] u1_col_in_397;
wire [151:0] u1_col_in_398;
wire [151:0] u1_col_in_399;
wire [151:0] u1_col_in_400;
wire [151:0] u1_col_in_401;
wire [151:0] u1_col_in_402;
wire [151:0] u1_col_in_403;
wire [151:0] u1_col_in_404;
wire [151:0] u1_col_in_405;
wire [151:0] u1_col_in_406;
wire [151:0] u1_col_in_407;
wire [151:0] u1_col_in_408;
wire [151:0] u1_col_in_409;
wire [151:0] u1_col_in_410;
wire [151:0] u1_col_in_411;
wire [151:0] u1_col_in_412;
wire [151:0] u1_col_in_413;
wire [151:0] u1_col_in_414;
wire [151:0] u1_col_in_415;
wire [151:0] u1_col_in_416;
wire [151:0] u1_col_in_417;
wire [151:0] u1_col_in_418;
wire [151:0] u1_col_in_419;
wire [151:0] u1_col_in_420;
wire [151:0] u1_col_in_421;
wire [151:0] u1_col_in_422;
wire [151:0] u1_col_in_423;
wire [151:0] u1_col_in_424;
wire [151:0] u1_col_in_425;
wire [151:0] u1_col_in_426;
wire [151:0] u1_col_in_427;
wire [151:0] u1_col_in_428;
wire [151:0] u1_col_in_429;
wire [151:0] u1_col_in_430;
wire [151:0] u1_col_in_431;
wire [151:0] u1_col_in_432;
wire [151:0] u1_col_in_433;
wire [151:0] u1_col_in_434;
wire [151:0] u1_col_in_435;
wire [151:0] u1_col_in_436;
wire [151:0] u1_col_in_437;
wire [151:0] u1_col_in_438;
wire [151:0] u1_col_in_439;
wire [151:0] u1_col_in_440;
wire [151:0] u1_col_in_441;
wire [151:0] u1_col_in_442;
wire [151:0] u1_col_in_443;
wire [151:0] u1_col_in_444;
wire [151:0] u1_col_in_445;
wire [151:0] u1_col_in_446;
wire [151:0] u1_col_in_447;
wire [151:0] u1_col_in_448;
wire [151:0] u1_col_in_449;
wire [151:0] u1_col_in_450;
wire [151:0] u1_col_in_451;
wire [151:0] u1_col_in_452;
wire [151:0] u1_col_in_453;
wire [151:0] u1_col_in_454;
wire [151:0] u1_col_in_455;
wire [151:0] u1_col_in_456;
wire [151:0] u1_col_in_457;
wire [151:0] u1_col_in_458;
wire [151:0] u1_col_in_459;
wire [151:0] u1_col_in_460;
wire [151:0] u1_col_in_461;
wire [151:0] u1_col_in_462;
wire [151:0] u1_col_in_463;
wire [151:0] u1_col_in_464;
wire [151:0] u1_col_in_465;
wire [151:0] u1_col_in_466;
wire [151:0] u1_col_in_467;
wire [151:0] u1_col_in_468;
wire [151:0] u1_col_in_469;
wire [151:0] u1_col_in_470;
wire [151:0] u1_col_in_471;
wire [151:0] u1_col_in_472;
wire [151:0] u1_col_in_473;
wire [151:0] u1_col_in_474;
wire [151:0] u1_col_in_475;
wire [151:0] u1_col_in_476;
wire [151:0] u1_col_in_477;
wire [151:0] u1_col_in_478;
wire [151:0] u1_col_in_479;
wire [151:0] u1_col_in_480;
wire [151:0] u1_col_in_481;
wire [151:0] u1_col_in_482;
wire [151:0] u1_col_in_483;
wire [151:0] u1_col_in_484;
wire [151:0] u1_col_in_485;
wire [151:0] u1_col_in_486;
wire [151:0] u1_col_in_487;
wire [151:0] u1_col_in_488;
wire [151:0] u1_col_in_489;
wire [151:0] u1_col_in_490;
wire [151:0] u1_col_in_491;
wire [151:0] u1_col_in_492;
wire [151:0] u1_col_in_493;
wire [151:0] u1_col_in_494;
wire [151:0] u1_col_in_495;
wire [151:0] u1_col_in_496;
wire [151:0] u1_col_in_497;
wire [151:0] u1_col_in_498;
wire [151:0] u1_col_in_499;
wire [151:0] u1_col_in_500;
wire [151:0] u1_col_in_501;
wire [151:0] u1_col_in_502;
wire [151:0] u1_col_in_503;
wire [151:0] u1_col_in_504;
wire [151:0] u1_col_in_505;
wire [151:0] u1_col_in_506;
wire [151:0] u1_col_in_507;
wire [151:0] u1_col_in_508;
wire [151:0] u1_col_in_509;
wire [151:0] u1_col_in_510;
wire [151:0] u1_col_in_511;
wire [151:0] u1_col_in_512;
wire [151:0] u1_col_in_513;
wire [151:0] u1_col_in_514;
wire [151:0] u1_col_in_515;
wire [151:0] u1_col_in_516;
wire [151:0] u1_col_in_517;
wire [151:0] u1_col_in_518;
wire [151:0] u1_col_in_519;
wire [151:0] u1_col_in_520;
wire [151:0] u1_col_in_521;
wire [151:0] u1_col_in_522;
wire [151:0] u1_col_in_523;
wire [151:0] u1_col_in_524;
wire [151:0] u1_col_in_525;
wire [151:0] u1_col_in_526;
wire [151:0] u1_col_in_527;
wire [151:0] u1_col_in_528;
wire [151:0] u1_col_in_529;
wire [151:0] u1_col_in_530;
wire [151:0] u1_col_in_531;
wire [151:0] u1_col_in_532;
wire [151:0] u1_col_in_533;
wire [151:0] u1_col_in_534;
wire [151:0] u1_col_in_535;
wire [151:0] u1_col_in_536;
wire [151:0] u1_col_in_537;
wire [151:0] u1_col_in_538;
wire [151:0] u1_col_in_539;
wire [151:0] u1_col_in_540;
wire [151:0] u1_col_in_541;
wire [151:0] u1_col_in_542;
wire [151:0] u1_col_in_543;
wire [151:0] u1_col_in_544;
wire [151:0] u1_col_in_545;
wire [151:0] u1_col_in_546;
wire [151:0] u1_col_in_547;
wire [151:0] u1_col_in_548;
wire [151:0] u1_col_in_549;
wire [151:0] u1_col_in_550;
wire [151:0] u1_col_in_551;
wire [151:0] u1_col_in_552;
wire [151:0] u1_col_in_553;
wire [151:0] u1_col_in_554;
wire [151:0] u1_col_in_555;
wire [151:0] u1_col_in_556;
wire [151:0] u1_col_in_557;
wire [151:0] u1_col_in_558;
wire [151:0] u1_col_in_559;
wire [151:0] u1_col_in_560;
wire [151:0] u1_col_in_561;
wire [151:0] u1_col_in_562;
wire [151:0] u1_col_in_563;
wire [151:0] u1_col_in_564;
wire [151:0] u1_col_in_565;
wire [151:0] u1_col_in_566;
wire [151:0] u1_col_in_567;
wire [151:0] u1_col_in_568;
wire [151:0] u1_col_in_569;
wire [151:0] u1_col_in_570;
wire [151:0] u1_col_in_571;
wire [151:0] u1_col_in_572;
wire [151:0] u1_col_in_573;
wire [151:0] u1_col_in_574;
wire [151:0] u1_col_in_575;
wire [151:0] u1_col_in_576;
wire [151:0] u1_col_in_577;
wire [151:0] u1_col_in_578;
wire [151:0] u1_col_in_579;
wire [151:0] u1_col_in_580;
wire [151:0] u1_col_in_581;
wire [151:0] u1_col_in_582;
wire [151:0] u1_col_in_583;
wire [151:0] u1_col_in_584;
wire [151:0] u1_col_in_585;
wire [151:0] u1_col_in_586;
wire [151:0] u1_col_in_587;
wire [151:0] u1_col_in_588;
wire [151:0] u1_col_in_589;
wire [151:0] u1_col_in_590;
wire [151:0] u1_col_in_591;
wire [151:0] u1_col_in_592;
wire [151:0] u1_col_in_593;
wire [151:0] u1_col_in_594;
wire [151:0] u1_col_in_595;
wire [151:0] u1_col_in_596;
wire [151:0] u1_col_in_597;
wire [151:0] u1_col_in_598;
wire [151:0] u1_col_in_599;
wire [151:0] u1_col_in_600;
wire [151:0] u1_col_in_601;
wire [151:0] u1_col_in_602;
wire [151:0] u1_col_in_603;
wire [151:0] u1_col_in_604;
wire [151:0] u1_col_in_605;
wire [151:0] u1_col_in_606;
wire [151:0] u1_col_in_607;
wire [151:0] u1_col_in_608;
wire [151:0] u1_col_in_609;
wire [151:0] u1_col_in_610;
wire [151:0] u1_col_in_611;
wire [151:0] u1_col_in_612;
wire [151:0] u1_col_in_613;
wire [151:0] u1_col_in_614;
wire [151:0] u1_col_in_615;
wire [151:0] u1_col_in_616;
wire [151:0] u1_col_in_617;
wire [151:0] u1_col_in_618;
wire [151:0] u1_col_in_619;
wire [151:0] u1_col_in_620;
wire [151:0] u1_col_in_621;
wire [151:0] u1_col_in_622;
wire [151:0] u1_col_in_623;
wire [151:0] u1_col_in_624;
wire [151:0] u1_col_in_625;
wire [151:0] u1_col_in_626;
wire [151:0] u1_col_in_627;
wire [151:0] u1_col_in_628;
wire [151:0] u1_col_in_629;
wire [151:0] u1_col_in_630;
wire [151:0] u1_col_in_631;
wire [151:0] u1_col_in_632;
wire [151:0] u1_col_in_633;
wire [151:0] u1_col_in_634;
wire [151:0] u1_col_in_635;
wire [151:0] u1_col_in_636;
wire [151:0] u1_col_in_637;
wire [151:0] u1_col_in_638;
wire [151:0] u1_col_in_639;
wire [151:0] u1_col_in_640;
wire [151:0] u1_col_in_641;
wire [151:0] u1_col_in_642;
wire [151:0] u1_col_in_643;
wire [151:0] u1_col_in_644;
wire [151:0] u1_col_in_645;
wire [151:0] u1_col_in_646;
wire [151:0] u1_col_in_647;
wire [151:0] u1_col_in_648;
wire [151:0] u1_col_in_649;
wire [151:0] u1_col_in_650;
wire [151:0] u1_col_in_651;
wire [151:0] u1_col_in_652;
wire [151:0] u1_col_in_653;
wire [151:0] u1_col_in_654;
wire [151:0] u1_col_in_655;
wire [151:0] u1_col_in_656;
wire [151:0] u1_col_in_657;
wire [151:0] u1_col_in_658;
wire [151:0] u1_col_in_659;
wire [151:0] u1_col_in_660;
wire [151:0] u1_col_in_661;
wire [151:0] u1_col_in_662;
wire [151:0] u1_col_in_663;
wire [151:0] u1_col_in_664;
wire [151:0] u1_col_in_665;
wire [151:0] u1_col_in_666;
wire [151:0] u1_col_in_667;
wire [151:0] u1_col_in_668;
wire [151:0] u1_col_in_669;
wire [151:0] u1_col_in_670;
wire [151:0] u1_col_in_671;
wire [151:0] u1_col_in_672;
wire [151:0] u1_col_in_673;
wire [151:0] u1_col_in_674;
wire [151:0] u1_col_in_675;
wire [151:0] u1_col_in_676;
wire [151:0] u1_col_in_677;
wire [151:0] u1_col_in_678;
wire [151:0] u1_col_in_679;
wire [151:0] u1_col_in_680;
wire [151:0] u1_col_in_681;
wire [151:0] u1_col_in_682;
wire [151:0] u1_col_in_683;
wire [151:0] u1_col_in_684;
wire [151:0] u1_col_in_685;
wire [151:0] u1_col_in_686;
wire [151:0] u1_col_in_687;
wire [151:0] u1_col_in_688;
wire [151:0] u1_col_in_689;
wire [151:0] u1_col_in_690;
wire [151:0] u1_col_in_691;
wire [151:0] u1_col_in_692;
wire [151:0] u1_col_in_693;
wire [151:0] u1_col_in_694;
wire [151:0] u1_col_in_695;
wire [151:0] u1_col_in_696;
wire [151:0] u1_col_in_697;
wire [151:0] u1_col_in_698;
wire [151:0] u1_col_in_699;
wire [151:0] u1_col_in_700;
wire [151:0] u1_col_in_701;
wire [151:0] u1_col_in_702;
wire [151:0] u1_col_in_703;
wire [151:0] u1_col_in_704;
wire [151:0] u1_col_in_705;
wire [151:0] u1_col_in_706;
wire [151:0] u1_col_in_707;
wire [151:0] u1_col_in_708;
wire [151:0] u1_col_in_709;
wire [151:0] u1_col_in_710;
wire [151:0] u1_col_in_711;
wire [151:0] u1_col_in_712;
wire [151:0] u1_col_in_713;
wire [151:0] u1_col_in_714;
wire [151:0] u1_col_in_715;
wire [151:0] u1_col_in_716;
wire [151:0] u1_col_in_717;
wire [151:0] u1_col_in_718;
wire [151:0] u1_col_in_719;
wire [151:0] u1_col_in_720;
wire [151:0] u1_col_in_721;
wire [151:0] u1_col_in_722;
wire [151:0] u1_col_in_723;
wire [151:0] u1_col_in_724;
wire [151:0] u1_col_in_725;
wire [151:0] u1_col_in_726;
wire [151:0] u1_col_in_727;
wire [151:0] u1_col_in_728;
wire [151:0] u1_col_in_729;
wire [151:0] u1_col_in_730;
wire [151:0] u1_col_in_731;
wire [151:0] u1_col_in_732;
wire [151:0] u1_col_in_733;
wire [151:0] u1_col_in_734;
wire [151:0] u1_col_in_735;
wire [151:0] u1_col_in_736;
wire [151:0] u1_col_in_737;
wire [151:0] u1_col_in_738;
wire [151:0] u1_col_in_739;
wire [151:0] u1_col_in_740;
wire [151:0] u1_col_in_741;
wire [151:0] u1_col_in_742;
wire [151:0] u1_col_in_743;
wire [151:0] u1_col_in_744;
wire [151:0] u1_col_in_745;
wire [151:0] u1_col_in_746;
wire [151:0] u1_col_in_747;
wire [151:0] u1_col_in_748;
wire [151:0] u1_col_in_749;
wire [151:0] u1_col_in_750;
wire [151:0] u1_col_in_751;
wire [151:0] u1_col_in_752;
wire [151:0] u1_col_in_753;
wire [151:0] u1_col_in_754;
wire [151:0] u1_col_in_755;
wire [151:0] u1_col_in_756;
wire [151:0] u1_col_in_757;
wire [151:0] u1_col_in_758;
wire [151:0] u1_col_in_759;
wire [151:0] u1_col_in_760;
wire [151:0] u1_col_in_761;
wire [151:0] u1_col_in_762;
wire [151:0] u1_col_in_763;
wire [151:0] u1_col_in_764;
wire [151:0] u1_col_in_765;
wire [151:0] u1_col_in_766;
wire [151:0] u1_col_in_767;
wire [151:0] u1_col_in_768;
wire [151:0] u1_col_in_769;
wire [151:0] u1_col_in_770;
wire [151:0] u1_col_in_771;
wire [151:0] u1_col_in_772;
wire [151:0] u1_col_in_773;
wire [151:0] u1_col_in_774;
wire [151:0] u1_col_in_775;
wire [151:0] u1_col_in_776;
wire [151:0] u1_col_in_777;
wire [151:0] u1_col_in_778;
wire [151:0] u1_col_in_779;
wire [151:0] u1_col_in_780;
wire [151:0] u1_col_in_781;
wire [151:0] u1_col_in_782;
wire [151:0] u1_col_in_783;
wire [151:0] u1_col_in_784;
wire [151:0] u1_col_in_785;
wire [151:0] u1_col_in_786;
wire [151:0] u1_col_in_787;
wire [151:0] u1_col_in_788;
wire [151:0] u1_col_in_789;
wire [151:0] u1_col_in_790;
wire [151:0] u1_col_in_791;
wire [151:0] u1_col_in_792;
wire [151:0] u1_col_in_793;
wire [151:0] u1_col_in_794;
wire [151:0] u1_col_in_795;
wire [151:0] u1_col_in_796;
wire [151:0] u1_col_in_797;
wire [151:0] u1_col_in_798;
wire [151:0] u1_col_in_799;
wire [151:0] u1_col_in_800;
wire [151:0] u1_col_in_801;
wire [151:0] u1_col_in_802;
wire [151:0] u1_col_in_803;
wire [151:0] u1_col_in_804;
wire [151:0] u1_col_in_805;
wire [151:0] u1_col_in_806;
wire [151:0] u1_col_in_807;
wire [151:0] u1_col_in_808;
wire [151:0] u1_col_in_809;
wire [151:0] u1_col_in_810;
wire [151:0] u1_col_in_811;
wire [151:0] u1_col_in_812;
wire [151:0] u1_col_in_813;
wire [151:0] u1_col_in_814;
wire [151:0] u1_col_in_815;
wire [151:0] u1_col_in_816;
wire [151:0] u1_col_in_817;
wire [151:0] u1_col_in_818;
wire [151:0] u1_col_in_819;
wire [151:0] u1_col_in_820;
wire [151:0] u1_col_in_821;
wire [151:0] u1_col_in_822;
wire [151:0] u1_col_in_823;
wire [151:0] u1_col_in_824;
wire [151:0] u1_col_in_825;
wire [151:0] u1_col_in_826;
wire [151:0] u1_col_in_827;
wire [151:0] u1_col_in_828;
wire [151:0] u1_col_in_829;
wire [151:0] u1_col_in_830;
wire [151:0] u1_col_in_831;
wire [151:0] u1_col_in_832;
wire [151:0] u1_col_in_833;
wire [151:0] u1_col_in_834;
wire [151:0] u1_col_in_835;
wire [151:0] u1_col_in_836;
wire [151:0] u1_col_in_837;
wire [151:0] u1_col_in_838;
wire [151:0] u1_col_in_839;
wire [151:0] u1_col_in_840;
wire [151:0] u1_col_in_841;
wire [151:0] u1_col_in_842;
wire [151:0] u1_col_in_843;
wire [151:0] u1_col_in_844;
wire [151:0] u1_col_in_845;
wire [151:0] u1_col_in_846;
wire [151:0] u1_col_in_847;
wire [151:0] u1_col_in_848;
wire [151:0] u1_col_in_849;
wire [151:0] u1_col_in_850;
wire [151:0] u1_col_in_851;
wire [151:0] u1_col_in_852;
wire [151:0] u1_col_in_853;
wire [151:0] u1_col_in_854;
wire [151:0] u1_col_in_855;
wire [151:0] u1_col_in_856;
wire [151:0] u1_col_in_857;
wire [151:0] u1_col_in_858;
wire [151:0] u1_col_in_859;
wire [151:0] u1_col_in_860;
wire [151:0] u1_col_in_861;
wire [151:0] u1_col_in_862;
wire [151:0] u1_col_in_863;
wire [151:0] u1_col_in_864;
wire [151:0] u1_col_in_865;
wire [151:0] u1_col_in_866;
wire [151:0] u1_col_in_867;
wire [151:0] u1_col_in_868;
wire [151:0] u1_col_in_869;
wire [151:0] u1_col_in_870;
wire [151:0] u1_col_in_871;
wire [151:0] u1_col_in_872;
wire [151:0] u1_col_in_873;
wire [151:0] u1_col_in_874;
wire [151:0] u1_col_in_875;
wire [151:0] u1_col_in_876;
wire [151:0] u1_col_in_877;
wire [151:0] u1_col_in_878;
wire [151:0] u1_col_in_879;
wire [151:0] u1_col_in_880;
wire [151:0] u1_col_in_881;
wire [151:0] u1_col_in_882;
wire [151:0] u1_col_in_883;
wire [151:0] u1_col_in_884;
wire [151:0] u1_col_in_885;
wire [151:0] u1_col_in_886;
wire [151:0] u1_col_in_887;
wire [151:0] u1_col_in_888;
wire [151:0] u1_col_in_889;
wire [151:0] u1_col_in_890;
wire [151:0] u1_col_in_891;
wire [151:0] u1_col_in_892;
wire [151:0] u1_col_in_893;
wire [151:0] u1_col_in_894;
wire [151:0] u1_col_in_895;
wire [151:0] u1_col_in_896;
wire [151:0] u1_col_in_897;
wire [151:0] u1_col_in_898;
wire [151:0] u1_col_in_899;
wire [151:0] u1_col_in_900;
wire [151:0] u1_col_in_901;
wire [151:0] u1_col_in_902;
wire [151:0] u1_col_in_903;
wire [151:0] u1_col_in_904;
wire [151:0] u1_col_in_905;
wire [151:0] u1_col_in_906;
wire [151:0] u1_col_in_907;
wire [151:0] u1_col_in_908;
wire [151:0] u1_col_in_909;
wire [151:0] u1_col_in_910;
wire [151:0] u1_col_in_911;
wire [151:0] u1_col_in_912;
wire [151:0] u1_col_in_913;
wire [151:0] u1_col_in_914;
wire [151:0] u1_col_in_915;
wire [151:0] u1_col_in_916;
wire [151:0] u1_col_in_917;
wire [151:0] u1_col_in_918;
wire [151:0] u1_col_in_919;
wire [151:0] u1_col_in_920;
wire [151:0] u1_col_in_921;
wire [151:0] u1_col_in_922;
wire [151:0] u1_col_in_923;
wire [151:0] u1_col_in_924;
wire [151:0] u1_col_in_925;
wire [151:0] u1_col_in_926;
wire [151:0] u1_col_in_927;
wire [151:0] u1_col_in_928;
wire [151:0] u1_col_in_929;
wire [151:0] u1_col_in_930;
wire [151:0] u1_col_in_931;
wire [151:0] u1_col_in_932;
wire [151:0] u1_col_in_933;
wire [151:0] u1_col_in_934;
wire [151:0] u1_col_in_935;
wire [151:0] u1_col_in_936;
wire [151:0] u1_col_in_937;
wire [151:0] u1_col_in_938;
wire [151:0] u1_col_in_939;
wire [151:0] u1_col_in_940;
wire [151:0] u1_col_in_941;
wire [151:0] u1_col_in_942;
wire [151:0] u1_col_in_943;
wire [151:0] u1_col_in_944;
wire [151:0] u1_col_in_945;
wire [151:0] u1_col_in_946;
wire [151:0] u1_col_in_947;
wire [151:0] u1_col_in_948;
wire [151:0] u1_col_in_949;
wire [151:0] u1_col_in_950;
wire [151:0] u1_col_in_951;
wire [151:0] u1_col_in_952;
wire [151:0] u1_col_in_953;
wire [151:0] u1_col_in_954;
wire [151:0] u1_col_in_955;
wire [151:0] u1_col_in_956;
wire [151:0] u1_col_in_957;
wire [151:0] u1_col_in_958;
wire [151:0] u1_col_in_959;
wire [151:0] u1_col_in_960;
wire [151:0] u1_col_in_961;
wire [151:0] u1_col_in_962;
wire [151:0] u1_col_in_963;
wire [151:0] u1_col_in_964;
wire [151:0] u1_col_in_965;
wire [151:0] u1_col_in_966;
wire [151:0] u1_col_in_967;
wire [151:0] u1_col_in_968;
wire [151:0] u1_col_in_969;
wire [151:0] u1_col_in_970;
wire [151:0] u1_col_in_971;
wire [151:0] u1_col_in_972;
wire [151:0] u1_col_in_973;
wire [151:0] u1_col_in_974;
wire [151:0] u1_col_in_975;
wire [151:0] u1_col_in_976;
wire [151:0] u1_col_in_977;
wire [151:0] u1_col_in_978;
wire [151:0] u1_col_in_979;
wire [151:0] u1_col_in_980;
wire [151:0] u1_col_in_981;
wire [151:0] u1_col_in_982;
wire [151:0] u1_col_in_983;
wire [151:0] u1_col_in_984;
wire [151:0] u1_col_in_985;
wire [151:0] u1_col_in_986;
wire [151:0] u1_col_in_987;
wire [151:0] u1_col_in_988;
wire [151:0] u1_col_in_989;
wire [151:0] u1_col_in_990;
wire [151:0] u1_col_in_991;
wire [151:0] u1_col_in_992;
wire [151:0] u1_col_in_993;
wire [151:0] u1_col_in_994;
wire [151:0] u1_col_in_995;
wire [151:0] u1_col_in_996;
wire [151:0] u1_col_in_997;
wire [151:0] u1_col_in_998;
wire [151:0] u1_col_in_999;
wire [151:0] u1_col_in_1000;
wire [151:0] u1_col_in_1001;
wire [151:0] u1_col_in_1002;
wire [151:0] u1_col_in_1003;
wire [151:0] u1_col_in_1004;
wire [151:0] u1_col_in_1005;
wire [151:0] u1_col_in_1006;
wire [151:0] u1_col_in_1007;
wire [151:0] u1_col_in_1008;
wire [151:0] u1_col_in_1009;
wire [151:0] u1_col_in_1010;
wire [151:0] u1_col_in_1011;
wire [151:0] u1_col_in_1012;
wire [151:0] u1_col_in_1013;
wire [151:0] u1_col_in_1014;
wire [151:0] u1_col_in_1015;
wire [151:0] u1_col_in_1016;
wire [151:0] u1_col_in_1017;
wire [151:0] u1_col_in_1018;
wire [151:0] u1_col_in_1019;
wire [151:0] u1_col_in_1020;
wire [151:0] u1_col_in_1021;
wire [151:0] u1_col_in_1022;
wire [151:0] u1_col_in_1023;
wire [151:0] u1_col_in_1024;
wire [151:0] u1_col_in_1025;
wire [151:0] u1_col_in_1026;




//*****************************************************
//**************u1输出定义******************************
//*****************************************************
wire [47:0] u1_col_out_0;
wire [47:0] u1_col_out_1;
wire [47:0] u1_col_out_2;
wire [47:0] u1_col_out_3;
wire [47:0] u1_col_out_4;
wire [47:0] u1_col_out_5;
wire [47:0] u1_col_out_6;
wire [47:0] u1_col_out_7;
wire [47:0] u1_col_out_8;
wire [47:0] u1_col_out_9;
wire [47:0] u1_col_out_10;
wire [47:0] u1_col_out_11;
wire [47:0] u1_col_out_12;
wire [47:0] u1_col_out_13;
wire [47:0] u1_col_out_14;
wire [47:0] u1_col_out_15;
wire [47:0] u1_col_out_16;
wire [47:0] u1_col_out_17;
wire [47:0] u1_col_out_18;
wire [47:0] u1_col_out_19;
wire [47:0] u1_col_out_20;
wire [47:0] u1_col_out_21;
wire [47:0] u1_col_out_22;
wire [47:0] u1_col_out_23;
wire [47:0] u1_col_out_24;
wire [47:0] u1_col_out_25;
wire [47:0] u1_col_out_26;
wire [47:0] u1_col_out_27;
wire [47:0] u1_col_out_28;
wire [47:0] u1_col_out_29;
wire [47:0] u1_col_out_30;
wire [47:0] u1_col_out_31;
wire [47:0] u1_col_out_32;
wire [47:0] u1_col_out_33;
wire [47:0] u1_col_out_34;
wire [47:0] u1_col_out_35;
wire [47:0] u1_col_out_36;
wire [47:0] u1_col_out_37;
wire [47:0] u1_col_out_38;
wire [47:0] u1_col_out_39;
wire [47:0] u1_col_out_40;
wire [47:0] u1_col_out_41;
wire [47:0] u1_col_out_42;
wire [47:0] u1_col_out_43;
wire [47:0] u1_col_out_44;
wire [47:0] u1_col_out_45;
wire [47:0] u1_col_out_46;
wire [47:0] u1_col_out_47;
wire [47:0] u1_col_out_48;
wire [47:0] u1_col_out_49;
wire [47:0] u1_col_out_50;
wire [47:0] u1_col_out_51;
wire [47:0] u1_col_out_52;
wire [47:0] u1_col_out_53;
wire [47:0] u1_col_out_54;
wire [47:0] u1_col_out_55;
wire [47:0] u1_col_out_56;
wire [47:0] u1_col_out_57;
wire [47:0] u1_col_out_58;
wire [47:0] u1_col_out_59;
wire [47:0] u1_col_out_60;
wire [47:0] u1_col_out_61;
wire [47:0] u1_col_out_62;
wire [47:0] u1_col_out_63;
wire [47:0] u1_col_out_64;
wire [47:0] u1_col_out_65;
wire [47:0] u1_col_out_66;
wire [47:0] u1_col_out_67;
wire [47:0] u1_col_out_68;
wire [47:0] u1_col_out_69;
wire [47:0] u1_col_out_70;
wire [47:0] u1_col_out_71;
wire [47:0] u1_col_out_72;
wire [47:0] u1_col_out_73;
wire [47:0] u1_col_out_74;
wire [47:0] u1_col_out_75;
wire [47:0] u1_col_out_76;
wire [47:0] u1_col_out_77;
wire [47:0] u1_col_out_78;
wire [47:0] u1_col_out_79;
wire [47:0] u1_col_out_80;
wire [47:0] u1_col_out_81;
wire [47:0] u1_col_out_82;
wire [47:0] u1_col_out_83;
wire [47:0] u1_col_out_84;
wire [47:0] u1_col_out_85;
wire [47:0] u1_col_out_86;
wire [47:0] u1_col_out_87;
wire [47:0] u1_col_out_88;
wire [47:0] u1_col_out_89;
wire [47:0] u1_col_out_90;
wire [47:0] u1_col_out_91;
wire [47:0] u1_col_out_92;
wire [47:0] u1_col_out_93;
wire [47:0] u1_col_out_94;
wire [47:0] u1_col_out_95;
wire [47:0] u1_col_out_96;
wire [47:0] u1_col_out_97;
wire [47:0] u1_col_out_98;
wire [47:0] u1_col_out_99;
wire [47:0] u1_col_out_100;
wire [47:0] u1_col_out_101;
wire [47:0] u1_col_out_102;
wire [47:0] u1_col_out_103;
wire [47:0] u1_col_out_104;
wire [47:0] u1_col_out_105;
wire [47:0] u1_col_out_106;
wire [47:0] u1_col_out_107;
wire [47:0] u1_col_out_108;
wire [47:0] u1_col_out_109;
wire [47:0] u1_col_out_110;
wire [47:0] u1_col_out_111;
wire [47:0] u1_col_out_112;
wire [47:0] u1_col_out_113;
wire [47:0] u1_col_out_114;
wire [47:0] u1_col_out_115;
wire [47:0] u1_col_out_116;
wire [47:0] u1_col_out_117;
wire [47:0] u1_col_out_118;
wire [47:0] u1_col_out_119;
wire [47:0] u1_col_out_120;
wire [47:0] u1_col_out_121;
wire [47:0] u1_col_out_122;
wire [47:0] u1_col_out_123;
wire [47:0] u1_col_out_124;
wire [47:0] u1_col_out_125;
wire [47:0] u1_col_out_126;
wire [47:0] u1_col_out_127;
wire [47:0] u1_col_out_128;
wire [47:0] u1_col_out_129;
wire [47:0] u1_col_out_130;
wire [47:0] u1_col_out_131;
wire [47:0] u1_col_out_132;
wire [47:0] u1_col_out_133;
wire [47:0] u1_col_out_134;
wire [47:0] u1_col_out_135;
wire [47:0] u1_col_out_136;
wire [47:0] u1_col_out_137;
wire [47:0] u1_col_out_138;
wire [47:0] u1_col_out_139;
wire [47:0] u1_col_out_140;
wire [47:0] u1_col_out_141;
wire [47:0] u1_col_out_142;
wire [47:0] u1_col_out_143;
wire [47:0] u1_col_out_144;
wire [47:0] u1_col_out_145;
wire [47:0] u1_col_out_146;
wire [47:0] u1_col_out_147;
wire [47:0] u1_col_out_148;
wire [47:0] u1_col_out_149;
wire [47:0] u1_col_out_150;
wire [47:0] u1_col_out_151;
wire [47:0] u1_col_out_152;
wire [47:0] u1_col_out_153;
wire [47:0] u1_col_out_154;
wire [47:0] u1_col_out_155;
wire [47:0] u1_col_out_156;
wire [47:0] u1_col_out_157;
wire [47:0] u1_col_out_158;
wire [47:0] u1_col_out_159;
wire [47:0] u1_col_out_160;
wire [47:0] u1_col_out_161;
wire [47:0] u1_col_out_162;
wire [47:0] u1_col_out_163;
wire [47:0] u1_col_out_164;
wire [47:0] u1_col_out_165;
wire [47:0] u1_col_out_166;
wire [47:0] u1_col_out_167;
wire [47:0] u1_col_out_168;
wire [47:0] u1_col_out_169;
wire [47:0] u1_col_out_170;
wire [47:0] u1_col_out_171;
wire [47:0] u1_col_out_172;
wire [47:0] u1_col_out_173;
wire [47:0] u1_col_out_174;
wire [47:0] u1_col_out_175;
wire [47:0] u1_col_out_176;
wire [47:0] u1_col_out_177;
wire [47:0] u1_col_out_178;
wire [47:0] u1_col_out_179;
wire [47:0] u1_col_out_180;
wire [47:0] u1_col_out_181;
wire [47:0] u1_col_out_182;
wire [47:0] u1_col_out_183;
wire [47:0] u1_col_out_184;
wire [47:0] u1_col_out_185;
wire [47:0] u1_col_out_186;
wire [47:0] u1_col_out_187;
wire [47:0] u1_col_out_188;
wire [47:0] u1_col_out_189;
wire [47:0] u1_col_out_190;
wire [47:0] u1_col_out_191;
wire [47:0] u1_col_out_192;
wire [47:0] u1_col_out_193;
wire [47:0] u1_col_out_194;
wire [47:0] u1_col_out_195;
wire [47:0] u1_col_out_196;
wire [47:0] u1_col_out_197;
wire [47:0] u1_col_out_198;
wire [47:0] u1_col_out_199;
wire [47:0] u1_col_out_200;
wire [47:0] u1_col_out_201;
wire [47:0] u1_col_out_202;
wire [47:0] u1_col_out_203;
wire [47:0] u1_col_out_204;
wire [47:0] u1_col_out_205;
wire [47:0] u1_col_out_206;
wire [47:0] u1_col_out_207;
wire [47:0] u1_col_out_208;
wire [47:0] u1_col_out_209;
wire [47:0] u1_col_out_210;
wire [47:0] u1_col_out_211;
wire [47:0] u1_col_out_212;
wire [47:0] u1_col_out_213;
wire [47:0] u1_col_out_214;
wire [47:0] u1_col_out_215;
wire [47:0] u1_col_out_216;
wire [47:0] u1_col_out_217;
wire [47:0] u1_col_out_218;
wire [47:0] u1_col_out_219;
wire [47:0] u1_col_out_220;
wire [47:0] u1_col_out_221;
wire [47:0] u1_col_out_222;
wire [47:0] u1_col_out_223;
wire [47:0] u1_col_out_224;
wire [47:0] u1_col_out_225;
wire [47:0] u1_col_out_226;
wire [47:0] u1_col_out_227;
wire [47:0] u1_col_out_228;
wire [47:0] u1_col_out_229;
wire [47:0] u1_col_out_230;
wire [47:0] u1_col_out_231;
wire [47:0] u1_col_out_232;
wire [47:0] u1_col_out_233;
wire [47:0] u1_col_out_234;
wire [47:0] u1_col_out_235;
wire [47:0] u1_col_out_236;
wire [47:0] u1_col_out_237;
wire [47:0] u1_col_out_238;
wire [47:0] u1_col_out_239;
wire [47:0] u1_col_out_240;
wire [47:0] u1_col_out_241;
wire [47:0] u1_col_out_242;
wire [47:0] u1_col_out_243;
wire [47:0] u1_col_out_244;
wire [47:0] u1_col_out_245;
wire [47:0] u1_col_out_246;
wire [47:0] u1_col_out_247;
wire [47:0] u1_col_out_248;
wire [47:0] u1_col_out_249;
wire [47:0] u1_col_out_250;
wire [47:0] u1_col_out_251;
wire [47:0] u1_col_out_252;
wire [47:0] u1_col_out_253;
wire [47:0] u1_col_out_254;
wire [47:0] u1_col_out_255;
wire [47:0] u1_col_out_256;
wire [47:0] u1_col_out_257;
wire [47:0] u1_col_out_258;
wire [47:0] u1_col_out_259;
wire [47:0] u1_col_out_260;
wire [47:0] u1_col_out_261;
wire [47:0] u1_col_out_262;
wire [47:0] u1_col_out_263;
wire [47:0] u1_col_out_264;
wire [47:0] u1_col_out_265;
wire [47:0] u1_col_out_266;
wire [47:0] u1_col_out_267;
wire [47:0] u1_col_out_268;
wire [47:0] u1_col_out_269;
wire [47:0] u1_col_out_270;
wire [47:0] u1_col_out_271;
wire [47:0] u1_col_out_272;
wire [47:0] u1_col_out_273;
wire [47:0] u1_col_out_274;
wire [47:0] u1_col_out_275;
wire [47:0] u1_col_out_276;
wire [47:0] u1_col_out_277;
wire [47:0] u1_col_out_278;
wire [47:0] u1_col_out_279;
wire [47:0] u1_col_out_280;
wire [47:0] u1_col_out_281;
wire [47:0] u1_col_out_282;
wire [47:0] u1_col_out_283;
wire [47:0] u1_col_out_284;
wire [47:0] u1_col_out_285;
wire [47:0] u1_col_out_286;
wire [47:0] u1_col_out_287;
wire [47:0] u1_col_out_288;
wire [47:0] u1_col_out_289;
wire [47:0] u1_col_out_290;
wire [47:0] u1_col_out_291;
wire [47:0] u1_col_out_292;
wire [47:0] u1_col_out_293;
wire [47:0] u1_col_out_294;
wire [47:0] u1_col_out_295;
wire [47:0] u1_col_out_296;
wire [47:0] u1_col_out_297;
wire [47:0] u1_col_out_298;
wire [47:0] u1_col_out_299;
wire [47:0] u1_col_out_300;
wire [47:0] u1_col_out_301;
wire [47:0] u1_col_out_302;
wire [47:0] u1_col_out_303;
wire [47:0] u1_col_out_304;
wire [47:0] u1_col_out_305;
wire [47:0] u1_col_out_306;
wire [47:0] u1_col_out_307;
wire [47:0] u1_col_out_308;
wire [47:0] u1_col_out_309;
wire [47:0] u1_col_out_310;
wire [47:0] u1_col_out_311;
wire [47:0] u1_col_out_312;
wire [47:0] u1_col_out_313;
wire [47:0] u1_col_out_314;
wire [47:0] u1_col_out_315;
wire [47:0] u1_col_out_316;
wire [47:0] u1_col_out_317;
wire [47:0] u1_col_out_318;
wire [47:0] u1_col_out_319;
wire [47:0] u1_col_out_320;
wire [47:0] u1_col_out_321;
wire [47:0] u1_col_out_322;
wire [47:0] u1_col_out_323;
wire [47:0] u1_col_out_324;
wire [47:0] u1_col_out_325;
wire [47:0] u1_col_out_326;
wire [47:0] u1_col_out_327;
wire [47:0] u1_col_out_328;
wire [47:0] u1_col_out_329;
wire [47:0] u1_col_out_330;
wire [47:0] u1_col_out_331;
wire [47:0] u1_col_out_332;
wire [47:0] u1_col_out_333;
wire [47:0] u1_col_out_334;
wire [47:0] u1_col_out_335;
wire [47:0] u1_col_out_336;
wire [47:0] u1_col_out_337;
wire [47:0] u1_col_out_338;
wire [47:0] u1_col_out_339;
wire [47:0] u1_col_out_340;
wire [47:0] u1_col_out_341;
wire [47:0] u1_col_out_342;
wire [47:0] u1_col_out_343;
wire [47:0] u1_col_out_344;
wire [47:0] u1_col_out_345;
wire [47:0] u1_col_out_346;
wire [47:0] u1_col_out_347;
wire [47:0] u1_col_out_348;
wire [47:0] u1_col_out_349;
wire [47:0] u1_col_out_350;
wire [47:0] u1_col_out_351;
wire [47:0] u1_col_out_352;
wire [47:0] u1_col_out_353;
wire [47:0] u1_col_out_354;
wire [47:0] u1_col_out_355;
wire [47:0] u1_col_out_356;
wire [47:0] u1_col_out_357;
wire [47:0] u1_col_out_358;
wire [47:0] u1_col_out_359;
wire [47:0] u1_col_out_360;
wire [47:0] u1_col_out_361;
wire [47:0] u1_col_out_362;
wire [47:0] u1_col_out_363;
wire [47:0] u1_col_out_364;
wire [47:0] u1_col_out_365;
wire [47:0] u1_col_out_366;
wire [47:0] u1_col_out_367;
wire [47:0] u1_col_out_368;
wire [47:0] u1_col_out_369;
wire [47:0] u1_col_out_370;
wire [47:0] u1_col_out_371;
wire [47:0] u1_col_out_372;
wire [47:0] u1_col_out_373;
wire [47:0] u1_col_out_374;
wire [47:0] u1_col_out_375;
wire [47:0] u1_col_out_376;
wire [47:0] u1_col_out_377;
wire [47:0] u1_col_out_378;
wire [47:0] u1_col_out_379;
wire [47:0] u1_col_out_380;
wire [47:0] u1_col_out_381;
wire [47:0] u1_col_out_382;
wire [47:0] u1_col_out_383;
wire [47:0] u1_col_out_384;
wire [47:0] u1_col_out_385;
wire [47:0] u1_col_out_386;
wire [47:0] u1_col_out_387;
wire [47:0] u1_col_out_388;
wire [47:0] u1_col_out_389;
wire [47:0] u1_col_out_390;
wire [47:0] u1_col_out_391;
wire [47:0] u1_col_out_392;
wire [47:0] u1_col_out_393;
wire [47:0] u1_col_out_394;
wire [47:0] u1_col_out_395;
wire [47:0] u1_col_out_396;
wire [47:0] u1_col_out_397;
wire [47:0] u1_col_out_398;
wire [47:0] u1_col_out_399;
wire [47:0] u1_col_out_400;
wire [47:0] u1_col_out_401;
wire [47:0] u1_col_out_402;
wire [47:0] u1_col_out_403;
wire [47:0] u1_col_out_404;
wire [47:0] u1_col_out_405;
wire [47:0] u1_col_out_406;
wire [47:0] u1_col_out_407;
wire [47:0] u1_col_out_408;
wire [47:0] u1_col_out_409;
wire [47:0] u1_col_out_410;
wire [47:0] u1_col_out_411;
wire [47:0] u1_col_out_412;
wire [47:0] u1_col_out_413;
wire [47:0] u1_col_out_414;
wire [47:0] u1_col_out_415;
wire [47:0] u1_col_out_416;
wire [47:0] u1_col_out_417;
wire [47:0] u1_col_out_418;
wire [47:0] u1_col_out_419;
wire [47:0] u1_col_out_420;
wire [47:0] u1_col_out_421;
wire [47:0] u1_col_out_422;
wire [47:0] u1_col_out_423;
wire [47:0] u1_col_out_424;
wire [47:0] u1_col_out_425;
wire [47:0] u1_col_out_426;
wire [47:0] u1_col_out_427;
wire [47:0] u1_col_out_428;
wire [47:0] u1_col_out_429;
wire [47:0] u1_col_out_430;
wire [47:0] u1_col_out_431;
wire [47:0] u1_col_out_432;
wire [47:0] u1_col_out_433;
wire [47:0] u1_col_out_434;
wire [47:0] u1_col_out_435;
wire [47:0] u1_col_out_436;
wire [47:0] u1_col_out_437;
wire [47:0] u1_col_out_438;
wire [47:0] u1_col_out_439;
wire [47:0] u1_col_out_440;
wire [47:0] u1_col_out_441;
wire [47:0] u1_col_out_442;
wire [47:0] u1_col_out_443;
wire [47:0] u1_col_out_444;
wire [47:0] u1_col_out_445;
wire [47:0] u1_col_out_446;
wire [47:0] u1_col_out_447;
wire [47:0] u1_col_out_448;
wire [47:0] u1_col_out_449;
wire [47:0] u1_col_out_450;
wire [47:0] u1_col_out_451;
wire [47:0] u1_col_out_452;
wire [47:0] u1_col_out_453;
wire [47:0] u1_col_out_454;
wire [47:0] u1_col_out_455;
wire [47:0] u1_col_out_456;
wire [47:0] u1_col_out_457;
wire [47:0] u1_col_out_458;
wire [47:0] u1_col_out_459;
wire [47:0] u1_col_out_460;
wire [47:0] u1_col_out_461;
wire [47:0] u1_col_out_462;
wire [47:0] u1_col_out_463;
wire [47:0] u1_col_out_464;
wire [47:0] u1_col_out_465;
wire [47:0] u1_col_out_466;
wire [47:0] u1_col_out_467;
wire [47:0] u1_col_out_468;
wire [47:0] u1_col_out_469;
wire [47:0] u1_col_out_470;
wire [47:0] u1_col_out_471;
wire [47:0] u1_col_out_472;
wire [47:0] u1_col_out_473;
wire [47:0] u1_col_out_474;
wire [47:0] u1_col_out_475;
wire [47:0] u1_col_out_476;
wire [47:0] u1_col_out_477;
wire [47:0] u1_col_out_478;
wire [47:0] u1_col_out_479;
wire [47:0] u1_col_out_480;
wire [47:0] u1_col_out_481;
wire [47:0] u1_col_out_482;
wire [47:0] u1_col_out_483;
wire [47:0] u1_col_out_484;
wire [47:0] u1_col_out_485;
wire [47:0] u1_col_out_486;
wire [47:0] u1_col_out_487;
wire [47:0] u1_col_out_488;
wire [47:0] u1_col_out_489;
wire [47:0] u1_col_out_490;
wire [47:0] u1_col_out_491;
wire [47:0] u1_col_out_492;
wire [47:0] u1_col_out_493;
wire [47:0] u1_col_out_494;
wire [47:0] u1_col_out_495;
wire [47:0] u1_col_out_496;
wire [47:0] u1_col_out_497;
wire [47:0] u1_col_out_498;
wire [47:0] u1_col_out_499;
wire [47:0] u1_col_out_500;
wire [47:0] u1_col_out_501;
wire [47:0] u1_col_out_502;
wire [47:0] u1_col_out_503;
wire [47:0] u1_col_out_504;
wire [47:0] u1_col_out_505;
wire [47:0] u1_col_out_506;
wire [47:0] u1_col_out_507;
wire [47:0] u1_col_out_508;
wire [47:0] u1_col_out_509;
wire [47:0] u1_col_out_510;
wire [47:0] u1_col_out_511;
wire [47:0] u1_col_out_512;
wire [47:0] u1_col_out_513;
wire [47:0] u1_col_out_514;
wire [47:0] u1_col_out_515;
wire [47:0] u1_col_out_516;
wire [47:0] u1_col_out_517;
wire [47:0] u1_col_out_518;
wire [47:0] u1_col_out_519;
wire [47:0] u1_col_out_520;
wire [47:0] u1_col_out_521;
wire [47:0] u1_col_out_522;
wire [47:0] u1_col_out_523;
wire [47:0] u1_col_out_524;
wire [47:0] u1_col_out_525;
wire [47:0] u1_col_out_526;
wire [47:0] u1_col_out_527;
wire [47:0] u1_col_out_528;
wire [47:0] u1_col_out_529;
wire [47:0] u1_col_out_530;
wire [47:0] u1_col_out_531;
wire [47:0] u1_col_out_532;
wire [47:0] u1_col_out_533;
wire [47:0] u1_col_out_534;
wire [47:0] u1_col_out_535;
wire [47:0] u1_col_out_536;
wire [47:0] u1_col_out_537;
wire [47:0] u1_col_out_538;
wire [47:0] u1_col_out_539;
wire [47:0] u1_col_out_540;
wire [47:0] u1_col_out_541;
wire [47:0] u1_col_out_542;
wire [47:0] u1_col_out_543;
wire [47:0] u1_col_out_544;
wire [47:0] u1_col_out_545;
wire [47:0] u1_col_out_546;
wire [47:0] u1_col_out_547;
wire [47:0] u1_col_out_548;
wire [47:0] u1_col_out_549;
wire [47:0] u1_col_out_550;
wire [47:0] u1_col_out_551;
wire [47:0] u1_col_out_552;
wire [47:0] u1_col_out_553;
wire [47:0] u1_col_out_554;
wire [47:0] u1_col_out_555;
wire [47:0] u1_col_out_556;
wire [47:0] u1_col_out_557;
wire [47:0] u1_col_out_558;
wire [47:0] u1_col_out_559;
wire [47:0] u1_col_out_560;
wire [47:0] u1_col_out_561;
wire [47:0] u1_col_out_562;
wire [47:0] u1_col_out_563;
wire [47:0] u1_col_out_564;
wire [47:0] u1_col_out_565;
wire [47:0] u1_col_out_566;
wire [47:0] u1_col_out_567;
wire [47:0] u1_col_out_568;
wire [47:0] u1_col_out_569;
wire [47:0] u1_col_out_570;
wire [47:0] u1_col_out_571;
wire [47:0] u1_col_out_572;
wire [47:0] u1_col_out_573;
wire [47:0] u1_col_out_574;
wire [47:0] u1_col_out_575;
wire [47:0] u1_col_out_576;
wire [47:0] u1_col_out_577;
wire [47:0] u1_col_out_578;
wire [47:0] u1_col_out_579;
wire [47:0] u1_col_out_580;
wire [47:0] u1_col_out_581;
wire [47:0] u1_col_out_582;
wire [47:0] u1_col_out_583;
wire [47:0] u1_col_out_584;
wire [47:0] u1_col_out_585;
wire [47:0] u1_col_out_586;
wire [47:0] u1_col_out_587;
wire [47:0] u1_col_out_588;
wire [47:0] u1_col_out_589;
wire [47:0] u1_col_out_590;
wire [47:0] u1_col_out_591;
wire [47:0] u1_col_out_592;
wire [47:0] u1_col_out_593;
wire [47:0] u1_col_out_594;
wire [47:0] u1_col_out_595;
wire [47:0] u1_col_out_596;
wire [47:0] u1_col_out_597;
wire [47:0] u1_col_out_598;
wire [47:0] u1_col_out_599;
wire [47:0] u1_col_out_600;
wire [47:0] u1_col_out_601;
wire [47:0] u1_col_out_602;
wire [47:0] u1_col_out_603;
wire [47:0] u1_col_out_604;
wire [47:0] u1_col_out_605;
wire [47:0] u1_col_out_606;
wire [47:0] u1_col_out_607;
wire [47:0] u1_col_out_608;
wire [47:0] u1_col_out_609;
wire [47:0] u1_col_out_610;
wire [47:0] u1_col_out_611;
wire [47:0] u1_col_out_612;
wire [47:0] u1_col_out_613;
wire [47:0] u1_col_out_614;
wire [47:0] u1_col_out_615;
wire [47:0] u1_col_out_616;
wire [47:0] u1_col_out_617;
wire [47:0] u1_col_out_618;
wire [47:0] u1_col_out_619;
wire [47:0] u1_col_out_620;
wire [47:0] u1_col_out_621;
wire [47:0] u1_col_out_622;
wire [47:0] u1_col_out_623;
wire [47:0] u1_col_out_624;
wire [47:0] u1_col_out_625;
wire [47:0] u1_col_out_626;
wire [47:0] u1_col_out_627;
wire [47:0] u1_col_out_628;
wire [47:0] u1_col_out_629;
wire [47:0] u1_col_out_630;
wire [47:0] u1_col_out_631;
wire [47:0] u1_col_out_632;
wire [47:0] u1_col_out_633;
wire [47:0] u1_col_out_634;
wire [47:0] u1_col_out_635;
wire [47:0] u1_col_out_636;
wire [47:0] u1_col_out_637;
wire [47:0] u1_col_out_638;
wire [47:0] u1_col_out_639;
wire [47:0] u1_col_out_640;
wire [47:0] u1_col_out_641;
wire [47:0] u1_col_out_642;
wire [47:0] u1_col_out_643;
wire [47:0] u1_col_out_644;
wire [47:0] u1_col_out_645;
wire [47:0] u1_col_out_646;
wire [47:0] u1_col_out_647;
wire [47:0] u1_col_out_648;
wire [47:0] u1_col_out_649;
wire [47:0] u1_col_out_650;
wire [47:0] u1_col_out_651;
wire [47:0] u1_col_out_652;
wire [47:0] u1_col_out_653;
wire [47:0] u1_col_out_654;
wire [47:0] u1_col_out_655;
wire [47:0] u1_col_out_656;
wire [47:0] u1_col_out_657;
wire [47:0] u1_col_out_658;
wire [47:0] u1_col_out_659;
wire [47:0] u1_col_out_660;
wire [47:0] u1_col_out_661;
wire [47:0] u1_col_out_662;
wire [47:0] u1_col_out_663;
wire [47:0] u1_col_out_664;
wire [47:0] u1_col_out_665;
wire [47:0] u1_col_out_666;
wire [47:0] u1_col_out_667;
wire [47:0] u1_col_out_668;
wire [47:0] u1_col_out_669;
wire [47:0] u1_col_out_670;
wire [47:0] u1_col_out_671;
wire [47:0] u1_col_out_672;
wire [47:0] u1_col_out_673;
wire [47:0] u1_col_out_674;
wire [47:0] u1_col_out_675;
wire [47:0] u1_col_out_676;
wire [47:0] u1_col_out_677;
wire [47:0] u1_col_out_678;
wire [47:0] u1_col_out_679;
wire [47:0] u1_col_out_680;
wire [47:0] u1_col_out_681;
wire [47:0] u1_col_out_682;
wire [47:0] u1_col_out_683;
wire [47:0] u1_col_out_684;
wire [47:0] u1_col_out_685;
wire [47:0] u1_col_out_686;
wire [47:0] u1_col_out_687;
wire [47:0] u1_col_out_688;
wire [47:0] u1_col_out_689;
wire [47:0] u1_col_out_690;
wire [47:0] u1_col_out_691;
wire [47:0] u1_col_out_692;
wire [47:0] u1_col_out_693;
wire [47:0] u1_col_out_694;
wire [47:0] u1_col_out_695;
wire [47:0] u1_col_out_696;
wire [47:0] u1_col_out_697;
wire [47:0] u1_col_out_698;
wire [47:0] u1_col_out_699;
wire [47:0] u1_col_out_700;
wire [47:0] u1_col_out_701;
wire [47:0] u1_col_out_702;
wire [47:0] u1_col_out_703;
wire [47:0] u1_col_out_704;
wire [47:0] u1_col_out_705;
wire [47:0] u1_col_out_706;
wire [47:0] u1_col_out_707;
wire [47:0] u1_col_out_708;
wire [47:0] u1_col_out_709;
wire [47:0] u1_col_out_710;
wire [47:0] u1_col_out_711;
wire [47:0] u1_col_out_712;
wire [47:0] u1_col_out_713;
wire [47:0] u1_col_out_714;
wire [47:0] u1_col_out_715;
wire [47:0] u1_col_out_716;
wire [47:0] u1_col_out_717;
wire [47:0] u1_col_out_718;
wire [47:0] u1_col_out_719;
wire [47:0] u1_col_out_720;
wire [47:0] u1_col_out_721;
wire [47:0] u1_col_out_722;
wire [47:0] u1_col_out_723;
wire [47:0] u1_col_out_724;
wire [47:0] u1_col_out_725;
wire [47:0] u1_col_out_726;
wire [47:0] u1_col_out_727;
wire [47:0] u1_col_out_728;
wire [47:0] u1_col_out_729;
wire [47:0] u1_col_out_730;
wire [47:0] u1_col_out_731;
wire [47:0] u1_col_out_732;
wire [47:0] u1_col_out_733;
wire [47:0] u1_col_out_734;
wire [47:0] u1_col_out_735;
wire [47:0] u1_col_out_736;
wire [47:0] u1_col_out_737;
wire [47:0] u1_col_out_738;
wire [47:0] u1_col_out_739;
wire [47:0] u1_col_out_740;
wire [47:0] u1_col_out_741;
wire [47:0] u1_col_out_742;
wire [47:0] u1_col_out_743;
wire [47:0] u1_col_out_744;
wire [47:0] u1_col_out_745;
wire [47:0] u1_col_out_746;
wire [47:0] u1_col_out_747;
wire [47:0] u1_col_out_748;
wire [47:0] u1_col_out_749;
wire [47:0] u1_col_out_750;
wire [47:0] u1_col_out_751;
wire [47:0] u1_col_out_752;
wire [47:0] u1_col_out_753;
wire [47:0] u1_col_out_754;
wire [47:0] u1_col_out_755;
wire [47:0] u1_col_out_756;
wire [47:0] u1_col_out_757;
wire [47:0] u1_col_out_758;
wire [47:0] u1_col_out_759;
wire [47:0] u1_col_out_760;
wire [47:0] u1_col_out_761;
wire [47:0] u1_col_out_762;
wire [47:0] u1_col_out_763;
wire [47:0] u1_col_out_764;
wire [47:0] u1_col_out_765;
wire [47:0] u1_col_out_766;
wire [47:0] u1_col_out_767;
wire [47:0] u1_col_out_768;
wire [47:0] u1_col_out_769;
wire [47:0] u1_col_out_770;
wire [47:0] u1_col_out_771;
wire [47:0] u1_col_out_772;
wire [47:0] u1_col_out_773;
wire [47:0] u1_col_out_774;
wire [47:0] u1_col_out_775;
wire [47:0] u1_col_out_776;
wire [47:0] u1_col_out_777;
wire [47:0] u1_col_out_778;
wire [47:0] u1_col_out_779;
wire [47:0] u1_col_out_780;
wire [47:0] u1_col_out_781;
wire [47:0] u1_col_out_782;
wire [47:0] u1_col_out_783;
wire [47:0] u1_col_out_784;
wire [47:0] u1_col_out_785;
wire [47:0] u1_col_out_786;
wire [47:0] u1_col_out_787;
wire [47:0] u1_col_out_788;
wire [47:0] u1_col_out_789;
wire [47:0] u1_col_out_790;
wire [47:0] u1_col_out_791;
wire [47:0] u1_col_out_792;
wire [47:0] u1_col_out_793;
wire [47:0] u1_col_out_794;
wire [47:0] u1_col_out_795;
wire [47:0] u1_col_out_796;
wire [47:0] u1_col_out_797;
wire [47:0] u1_col_out_798;
wire [47:0] u1_col_out_799;
wire [47:0] u1_col_out_800;
wire [47:0] u1_col_out_801;
wire [47:0] u1_col_out_802;
wire [47:0] u1_col_out_803;
wire [47:0] u1_col_out_804;
wire [47:0] u1_col_out_805;
wire [47:0] u1_col_out_806;
wire [47:0] u1_col_out_807;
wire [47:0] u1_col_out_808;
wire [47:0] u1_col_out_809;
wire [47:0] u1_col_out_810;
wire [47:0] u1_col_out_811;
wire [47:0] u1_col_out_812;
wire [47:0] u1_col_out_813;
wire [47:0] u1_col_out_814;
wire [47:0] u1_col_out_815;
wire [47:0] u1_col_out_816;
wire [47:0] u1_col_out_817;
wire [47:0] u1_col_out_818;
wire [47:0] u1_col_out_819;
wire [47:0] u1_col_out_820;
wire [47:0] u1_col_out_821;
wire [47:0] u1_col_out_822;
wire [47:0] u1_col_out_823;
wire [47:0] u1_col_out_824;
wire [47:0] u1_col_out_825;
wire [47:0] u1_col_out_826;
wire [47:0] u1_col_out_827;
wire [47:0] u1_col_out_828;
wire [47:0] u1_col_out_829;
wire [47:0] u1_col_out_830;
wire [47:0] u1_col_out_831;
wire [47:0] u1_col_out_832;
wire [47:0] u1_col_out_833;
wire [47:0] u1_col_out_834;
wire [47:0] u1_col_out_835;
wire [47:0] u1_col_out_836;
wire [47:0] u1_col_out_837;
wire [47:0] u1_col_out_838;
wire [47:0] u1_col_out_839;
wire [47:0] u1_col_out_840;
wire [47:0] u1_col_out_841;
wire [47:0] u1_col_out_842;
wire [47:0] u1_col_out_843;
wire [47:0] u1_col_out_844;
wire [47:0] u1_col_out_845;
wire [47:0] u1_col_out_846;
wire [47:0] u1_col_out_847;
wire [47:0] u1_col_out_848;
wire [47:0] u1_col_out_849;
wire [47:0] u1_col_out_850;
wire [47:0] u1_col_out_851;
wire [47:0] u1_col_out_852;
wire [47:0] u1_col_out_853;
wire [47:0] u1_col_out_854;
wire [47:0] u1_col_out_855;
wire [47:0] u1_col_out_856;
wire [47:0] u1_col_out_857;
wire [47:0] u1_col_out_858;
wire [47:0] u1_col_out_859;
wire [47:0] u1_col_out_860;
wire [47:0] u1_col_out_861;
wire [47:0] u1_col_out_862;
wire [47:0] u1_col_out_863;
wire [47:0] u1_col_out_864;
wire [47:0] u1_col_out_865;
wire [47:0] u1_col_out_866;
wire [47:0] u1_col_out_867;
wire [47:0] u1_col_out_868;
wire [47:0] u1_col_out_869;
wire [47:0] u1_col_out_870;
wire [47:0] u1_col_out_871;
wire [47:0] u1_col_out_872;
wire [47:0] u1_col_out_873;
wire [47:0] u1_col_out_874;
wire [47:0] u1_col_out_875;
wire [47:0] u1_col_out_876;
wire [47:0] u1_col_out_877;
wire [47:0] u1_col_out_878;
wire [47:0] u1_col_out_879;
wire [47:0] u1_col_out_880;
wire [47:0] u1_col_out_881;
wire [47:0] u1_col_out_882;
wire [47:0] u1_col_out_883;
wire [47:0] u1_col_out_884;
wire [47:0] u1_col_out_885;
wire [47:0] u1_col_out_886;
wire [47:0] u1_col_out_887;
wire [47:0] u1_col_out_888;
wire [47:0] u1_col_out_889;
wire [47:0] u1_col_out_890;
wire [47:0] u1_col_out_891;
wire [47:0] u1_col_out_892;
wire [47:0] u1_col_out_893;
wire [47:0] u1_col_out_894;
wire [47:0] u1_col_out_895;
wire [47:0] u1_col_out_896;
wire [47:0] u1_col_out_897;
wire [47:0] u1_col_out_898;
wire [47:0] u1_col_out_899;
wire [47:0] u1_col_out_900;
wire [47:0] u1_col_out_901;
wire [47:0] u1_col_out_902;
wire [47:0] u1_col_out_903;
wire [47:0] u1_col_out_904;
wire [47:0] u1_col_out_905;
wire [47:0] u1_col_out_906;
wire [47:0] u1_col_out_907;
wire [47:0] u1_col_out_908;
wire [47:0] u1_col_out_909;
wire [47:0] u1_col_out_910;
wire [47:0] u1_col_out_911;
wire [47:0] u1_col_out_912;
wire [47:0] u1_col_out_913;
wire [47:0] u1_col_out_914;
wire [47:0] u1_col_out_915;
wire [47:0] u1_col_out_916;
wire [47:0] u1_col_out_917;
wire [47:0] u1_col_out_918;
wire [47:0] u1_col_out_919;
wire [47:0] u1_col_out_920;
wire [47:0] u1_col_out_921;
wire [47:0] u1_col_out_922;
wire [47:0] u1_col_out_923;
wire [47:0] u1_col_out_924;
wire [47:0] u1_col_out_925;
wire [47:0] u1_col_out_926;
wire [47:0] u1_col_out_927;
wire [47:0] u1_col_out_928;
wire [47:0] u1_col_out_929;
wire [47:0] u1_col_out_930;
wire [47:0] u1_col_out_931;
wire [47:0] u1_col_out_932;
wire [47:0] u1_col_out_933;
wire [47:0] u1_col_out_934;
wire [47:0] u1_col_out_935;
wire [47:0] u1_col_out_936;
wire [47:0] u1_col_out_937;
wire [47:0] u1_col_out_938;
wire [47:0] u1_col_out_939;
wire [47:0] u1_col_out_940;
wire [47:0] u1_col_out_941;
wire [47:0] u1_col_out_942;
wire [47:0] u1_col_out_943;
wire [47:0] u1_col_out_944;
wire [47:0] u1_col_out_945;
wire [47:0] u1_col_out_946;
wire [47:0] u1_col_out_947;
wire [47:0] u1_col_out_948;
wire [47:0] u1_col_out_949;
wire [47:0] u1_col_out_950;
wire [47:0] u1_col_out_951;
wire [47:0] u1_col_out_952;
wire [47:0] u1_col_out_953;
wire [47:0] u1_col_out_954;
wire [47:0] u1_col_out_955;
wire [47:0] u1_col_out_956;
wire [47:0] u1_col_out_957;
wire [47:0] u1_col_out_958;
wire [47:0] u1_col_out_959;
wire [47:0] u1_col_out_960;
wire [47:0] u1_col_out_961;
wire [47:0] u1_col_out_962;
wire [47:0] u1_col_out_963;
wire [47:0] u1_col_out_964;
wire [47:0] u1_col_out_965;
wire [47:0] u1_col_out_966;
wire [47:0] u1_col_out_967;
wire [47:0] u1_col_out_968;
wire [47:0] u1_col_out_969;
wire [47:0] u1_col_out_970;
wire [47:0] u1_col_out_971;
wire [47:0] u1_col_out_972;
wire [47:0] u1_col_out_973;
wire [47:0] u1_col_out_974;
wire [47:0] u1_col_out_975;
wire [47:0] u1_col_out_976;
wire [47:0] u1_col_out_977;
wire [47:0] u1_col_out_978;
wire [47:0] u1_col_out_979;
wire [47:0] u1_col_out_980;
wire [47:0] u1_col_out_981;
wire [47:0] u1_col_out_982;
wire [47:0] u1_col_out_983;
wire [47:0] u1_col_out_984;
wire [47:0] u1_col_out_985;
wire [47:0] u1_col_out_986;
wire [47:0] u1_col_out_987;
wire [47:0] u1_col_out_988;
wire [47:0] u1_col_out_989;
wire [47:0] u1_col_out_990;
wire [47:0] u1_col_out_991;
wire [47:0] u1_col_out_992;
wire [47:0] u1_col_out_993;
wire [47:0] u1_col_out_994;
wire [47:0] u1_col_out_995;
wire [47:0] u1_col_out_996;
wire [47:0] u1_col_out_997;
wire [47:0] u1_col_out_998;
wire [47:0] u1_col_out_999;
wire [47:0] u1_col_out_1000;
wire [47:0] u1_col_out_1001;
wire [47:0] u1_col_out_1002;
wire [47:0] u1_col_out_1003;
wire [47:0] u1_col_out_1004;
wire [47:0] u1_col_out_1005;
wire [47:0] u1_col_out_1006;
wire [47:0] u1_col_out_1007;
wire [47:0] u1_col_out_1008;
wire [47:0] u1_col_out_1009;
wire [47:0] u1_col_out_1010;
wire [47:0] u1_col_out_1011;
wire [47:0] u1_col_out_1012;
wire [47:0] u1_col_out_1013;
wire [47:0] u1_col_out_1014;
wire [47:0] u1_col_out_1015;
wire [47:0] u1_col_out_1016;
wire [47:0] u1_col_out_1017;
wire [47:0] u1_col_out_1018;
wire [47:0] u1_col_out_1019;
wire [47:0] u1_col_out_1020;
wire [47:0] u1_col_out_1021;
wire [47:0] u1_col_out_1022;
wire [47:0] u1_col_out_1023;
wire [47:0] u1_col_out_1024;
wire [47:0] u1_col_out_1025;
wire [47:0] u1_col_out_1026;
wire [47:0] u1_col_out_1027;
wire [47:0] u1_col_out_1028;
wire [47:0] u1_col_out_1029;





//*****************************************************
//**************u1输入赋值******************************
//*****************************************************
assign u1_col_in_0 = u0_col_out_0;
assign u1_col_in_1 = u0_col_out_1;
assign u1_col_in_2 = u0_col_out_2;
assign u1_col_in_3 = u0_col_out_3;
assign u1_col_in_4 = u0_col_out_4;
assign u1_col_in_5 = u0_col_out_5;
assign u1_col_in_6 = u0_col_out_6;
assign u1_col_in_7 = u0_col_out_7;
assign u1_col_in_8 = u0_col_out_8;
assign u1_col_in_9 = u0_col_out_9;
assign u1_col_in_10 = u0_col_out_10;
assign u1_col_in_11 = u0_col_out_11;
assign u1_col_in_12 = u0_col_out_12;
assign u1_col_in_13 = u0_col_out_13;
assign u1_col_in_14 = u0_col_out_14;
assign u1_col_in_15 = u0_col_out_15;
assign u1_col_in_16 = u0_col_out_16;
assign u1_col_in_17 = u0_col_out_17;
assign u1_col_in_18 = u0_col_out_18;
assign u1_col_in_19 = u0_col_out_19;
assign u1_col_in_20 = u0_col_out_20;
assign u1_col_in_21 = u0_col_out_21;
assign u1_col_in_22 = u0_col_out_22;
assign u1_col_in_23 = u0_col_out_23;
assign u1_col_in_24 = u0_col_out_24;
assign u1_col_in_25 = u0_col_out_25;
assign u1_col_in_26 = u0_col_out_26;
assign u1_col_in_27 = u0_col_out_27;
assign u1_col_in_28 = u0_col_out_28;
assign u1_col_in_29 = u0_col_out_29;
assign u1_col_in_30 = u0_col_out_30;
assign u1_col_in_31 = u0_col_out_31;
assign u1_col_in_32 = u0_col_out_32;
assign u1_col_in_33 = u0_col_out_33;
assign u1_col_in_34 = u0_col_out_34;
assign u1_col_in_35 = u0_col_out_35;
assign u1_col_in_36 = u0_col_out_36;
assign u1_col_in_37 = u0_col_out_37;
assign u1_col_in_38 = u0_col_out_38;
assign u1_col_in_39 = u0_col_out_39;
assign u1_col_in_40 = u0_col_out_40;
assign u1_col_in_41 = u0_col_out_41;
assign u1_col_in_42 = u0_col_out_42;
assign u1_col_in_43 = u0_col_out_43;
assign u1_col_in_44 = u0_col_out_44;
assign u1_col_in_45 = u0_col_out_45;
assign u1_col_in_46 = u0_col_out_46;
assign u1_col_in_47 = u0_col_out_47;
assign u1_col_in_48 = u0_col_out_48;
assign u1_col_in_49 = u0_col_out_49;
assign u1_col_in_50 = u0_col_out_50;
assign u1_col_in_51 = u0_col_out_51;
assign u1_col_in_52 = u0_col_out_52;
assign u1_col_in_53 = u0_col_out_53;
assign u1_col_in_54 = u0_col_out_54;
assign u1_col_in_55 = u0_col_out_55;
assign u1_col_in_56 = u0_col_out_56;
assign u1_col_in_57 = u0_col_out_57;
assign u1_col_in_58 = u0_col_out_58;
assign u1_col_in_59 = u0_col_out_59;
assign u1_col_in_60 = u0_col_out_60;
assign u1_col_in_61 = u0_col_out_61;
assign u1_col_in_62 = u0_col_out_62;
assign u1_col_in_63 = u0_col_out_63;
assign u1_col_in_64 = u0_col_out_64;
assign u1_col_in_65 = u0_col_out_65;
assign u1_col_in_66 = u0_col_out_66;
assign u1_col_in_67 = u0_col_out_67;
assign u1_col_in_68 = u0_col_out_68;
assign u1_col_in_69 = u0_col_out_69;
assign u1_col_in_70 = u0_col_out_70;
assign u1_col_in_71 = u0_col_out_71;
assign u1_col_in_72 = u0_col_out_72;
assign u1_col_in_73 = u0_col_out_73;
assign u1_col_in_74 = u0_col_out_74;
assign u1_col_in_75 = u0_col_out_75;
assign u1_col_in_76 = u0_col_out_76;
assign u1_col_in_77 = u0_col_out_77;
assign u1_col_in_78 = u0_col_out_78;
assign u1_col_in_79 = u0_col_out_79;
assign u1_col_in_80 = u0_col_out_80;
assign u1_col_in_81 = u0_col_out_81;
assign u1_col_in_82 = u0_col_out_82;
assign u1_col_in_83 = u0_col_out_83;
assign u1_col_in_84 = u0_col_out_84;
assign u1_col_in_85 = u0_col_out_85;
assign u1_col_in_86 = u0_col_out_86;
assign u1_col_in_87 = u0_col_out_87;
assign u1_col_in_88 = u0_col_out_88;
assign u1_col_in_89 = u0_col_out_89;
assign u1_col_in_90 = u0_col_out_90;
assign u1_col_in_91 = u0_col_out_91;
assign u1_col_in_92 = u0_col_out_92;
assign u1_col_in_93 = u0_col_out_93;
assign u1_col_in_94 = u0_col_out_94;
assign u1_col_in_95 = u0_col_out_95;
assign u1_col_in_96 = u0_col_out_96;
assign u1_col_in_97 = u0_col_out_97;
assign u1_col_in_98 = u0_col_out_98;
assign u1_col_in_99 = u0_col_out_99;
assign u1_col_in_100 = u0_col_out_100;
assign u1_col_in_101 = u0_col_out_101;
assign u1_col_in_102 = u0_col_out_102;
assign u1_col_in_103 = u0_col_out_103;
assign u1_col_in_104 = u0_col_out_104;
assign u1_col_in_105 = u0_col_out_105;
assign u1_col_in_106 = u0_col_out_106;
assign u1_col_in_107 = u0_col_out_107;
assign u1_col_in_108 = u0_col_out_108;
assign u1_col_in_109 = u0_col_out_109;
assign u1_col_in_110 = u0_col_out_110;
assign u1_col_in_111 = u0_col_out_111;
assign u1_col_in_112 = u0_col_out_112;
assign u1_col_in_113 = u0_col_out_113;
assign u1_col_in_114 = u0_col_out_114;
assign u1_col_in_115 = u0_col_out_115;
assign u1_col_in_116 = u0_col_out_116;
assign u1_col_in_117 = u0_col_out_117;
assign u1_col_in_118 = u0_col_out_118;
assign u1_col_in_119 = u0_col_out_119;
assign u1_col_in_120 = u0_col_out_120;
assign u1_col_in_121 = u0_col_out_121;
assign u1_col_in_122 = u0_col_out_122;
assign u1_col_in_123 = u0_col_out_123;
assign u1_col_in_124 = u0_col_out_124;
assign u1_col_in_125 = u0_col_out_125;
assign u1_col_in_126 = u0_col_out_126;
assign u1_col_in_127 = u0_col_out_127;
assign u1_col_in_128 = u0_col_out_128;
assign u1_col_in_129 = u0_col_out_129;
assign u1_col_in_130 = u0_col_out_130;
assign u1_col_in_131 = u0_col_out_131;
assign u1_col_in_132 = u0_col_out_132;
assign u1_col_in_133 = u0_col_out_133;
assign u1_col_in_134 = u0_col_out_134;
assign u1_col_in_135 = u0_col_out_135;
assign u1_col_in_136 = u0_col_out_136;
assign u1_col_in_137 = u0_col_out_137;
assign u1_col_in_138 = u0_col_out_138;
assign u1_col_in_139 = u0_col_out_139;
assign u1_col_in_140 = u0_col_out_140;
assign u1_col_in_141 = u0_col_out_141;
assign u1_col_in_142 = u0_col_out_142;
assign u1_col_in_143 = u0_col_out_143;
assign u1_col_in_144 = u0_col_out_144;
assign u1_col_in_145 = u0_col_out_145;
assign u1_col_in_146 = u0_col_out_146;
assign u1_col_in_147 = u0_col_out_147;
assign u1_col_in_148 = u0_col_out_148;
assign u1_col_in_149 = u0_col_out_149;
assign u1_col_in_150 = u0_col_out_150;
assign u1_col_in_151 = u0_col_out_151;
assign u1_col_in_152 = u0_col_out_152;
assign u1_col_in_153 = u0_col_out_153;
assign u1_col_in_154 = u0_col_out_154;
assign u1_col_in_155 = u0_col_out_155;
assign u1_col_in_156 = u0_col_out_156;
assign u1_col_in_157 = u0_col_out_157;
assign u1_col_in_158 = u0_col_out_158;
assign u1_col_in_159 = u0_col_out_159;
assign u1_col_in_160 = u0_col_out_160;
assign u1_col_in_161 = u0_col_out_161;
assign u1_col_in_162 = u0_col_out_162;
assign u1_col_in_163 = u0_col_out_163;
assign u1_col_in_164 = u0_col_out_164;
assign u1_col_in_165 = u0_col_out_165;
assign u1_col_in_166 = u0_col_out_166;
assign u1_col_in_167 = u0_col_out_167;
assign u1_col_in_168 = u0_col_out_168;
assign u1_col_in_169 = u0_col_out_169;
assign u1_col_in_170 = u0_col_out_170;
assign u1_col_in_171 = u0_col_out_171;
assign u1_col_in_172 = u0_col_out_172;
assign u1_col_in_173 = u0_col_out_173;
assign u1_col_in_174 = u0_col_out_174;
assign u1_col_in_175 = u0_col_out_175;
assign u1_col_in_176 = u0_col_out_176;
assign u1_col_in_177 = u0_col_out_177;
assign u1_col_in_178 = u0_col_out_178;
assign u1_col_in_179 = u0_col_out_179;
assign u1_col_in_180 = u0_col_out_180;
assign u1_col_in_181 = u0_col_out_181;
assign u1_col_in_182 = u0_col_out_182;
assign u1_col_in_183 = u0_col_out_183;
assign u1_col_in_184 = u0_col_out_184;
assign u1_col_in_185 = u0_col_out_185;
assign u1_col_in_186 = u0_col_out_186;
assign u1_col_in_187 = u0_col_out_187;
assign u1_col_in_188 = u0_col_out_188;
assign u1_col_in_189 = u0_col_out_189;
assign u1_col_in_190 = u0_col_out_190;
assign u1_col_in_191 = u0_col_out_191;
assign u1_col_in_192 = u0_col_out_192;
assign u1_col_in_193 = u0_col_out_193;
assign u1_col_in_194 = u0_col_out_194;
assign u1_col_in_195 = u0_col_out_195;
assign u1_col_in_196 = u0_col_out_196;
assign u1_col_in_197 = u0_col_out_197;
assign u1_col_in_198 = u0_col_out_198;
assign u1_col_in_199 = u0_col_out_199;
assign u1_col_in_200 = u0_col_out_200;
assign u1_col_in_201 = u0_col_out_201;
assign u1_col_in_202 = u0_col_out_202;
assign u1_col_in_203 = u0_col_out_203;
assign u1_col_in_204 = u0_col_out_204;
assign u1_col_in_205 = u0_col_out_205;
assign u1_col_in_206 = u0_col_out_206;
assign u1_col_in_207 = u0_col_out_207;
assign u1_col_in_208 = u0_col_out_208;
assign u1_col_in_209 = u0_col_out_209;
assign u1_col_in_210 = u0_col_out_210;
assign u1_col_in_211 = u0_col_out_211;
assign u1_col_in_212 = u0_col_out_212;
assign u1_col_in_213 = u0_col_out_213;
assign u1_col_in_214 = u0_col_out_214;
assign u1_col_in_215 = u0_col_out_215;
assign u1_col_in_216 = u0_col_out_216;
assign u1_col_in_217 = u0_col_out_217;
assign u1_col_in_218 = u0_col_out_218;
assign u1_col_in_219 = u0_col_out_219;
assign u1_col_in_220 = u0_col_out_220;
assign u1_col_in_221 = u0_col_out_221;
assign u1_col_in_222 = u0_col_out_222;
assign u1_col_in_223 = u0_col_out_223;
assign u1_col_in_224 = u0_col_out_224;
assign u1_col_in_225 = u0_col_out_225;
assign u1_col_in_226 = u0_col_out_226;
assign u1_col_in_227 = u0_col_out_227;
assign u1_col_in_228 = u0_col_out_228;
assign u1_col_in_229 = u0_col_out_229;
assign u1_col_in_230 = u0_col_out_230;
assign u1_col_in_231 = u0_col_out_231;
assign u1_col_in_232 = u0_col_out_232;
assign u1_col_in_233 = u0_col_out_233;
assign u1_col_in_234 = u0_col_out_234;
assign u1_col_in_235 = u0_col_out_235;
assign u1_col_in_236 = u0_col_out_236;
assign u1_col_in_237 = u0_col_out_237;
assign u1_col_in_238 = u0_col_out_238;
assign u1_col_in_239 = u0_col_out_239;
assign u1_col_in_240 = u0_col_out_240;
assign u1_col_in_241 = u0_col_out_241;
assign u1_col_in_242 = u0_col_out_242;
assign u1_col_in_243 = u0_col_out_243;
assign u1_col_in_244 = u0_col_out_244;
assign u1_col_in_245 = u0_col_out_245;
assign u1_col_in_246 = u0_col_out_246;
assign u1_col_in_247 = u0_col_out_247;
assign u1_col_in_248 = u0_col_out_248;
assign u1_col_in_249 = u0_col_out_249;
assign u1_col_in_250 = u0_col_out_250;
assign u1_col_in_251 = u0_col_out_251;
assign u1_col_in_252 = u0_col_out_252;
assign u1_col_in_253 = u0_col_out_253;
assign u1_col_in_254 = u0_col_out_254;
assign u1_col_in_255 = u0_col_out_255;
assign u1_col_in_256 = u0_col_out_256;
assign u1_col_in_257 = u0_col_out_257;
assign u1_col_in_258 = u0_col_out_258;
assign u1_col_in_259 = u0_col_out_259;
assign u1_col_in_260 = u0_col_out_260;
assign u1_col_in_261 = u0_col_out_261;
assign u1_col_in_262 = u0_col_out_262;
assign u1_col_in_263 = u0_col_out_263;
assign u1_col_in_264 = u0_col_out_264;
assign u1_col_in_265 = u0_col_out_265;
assign u1_col_in_266 = u0_col_out_266;
assign u1_col_in_267 = u0_col_out_267;
assign u1_col_in_268 = u0_col_out_268;
assign u1_col_in_269 = u0_col_out_269;
assign u1_col_in_270 = u0_col_out_270;
assign u1_col_in_271 = u0_col_out_271;
assign u1_col_in_272 = u0_col_out_272;
assign u1_col_in_273 = u0_col_out_273;
assign u1_col_in_274 = u0_col_out_274;
assign u1_col_in_275 = u0_col_out_275;
assign u1_col_in_276 = u0_col_out_276;
assign u1_col_in_277 = u0_col_out_277;
assign u1_col_in_278 = u0_col_out_278;
assign u1_col_in_279 = u0_col_out_279;
assign u1_col_in_280 = u0_col_out_280;
assign u1_col_in_281 = u0_col_out_281;
assign u1_col_in_282 = u0_col_out_282;
assign u1_col_in_283 = u0_col_out_283;
assign u1_col_in_284 = u0_col_out_284;
assign u1_col_in_285 = u0_col_out_285;
assign u1_col_in_286 = u0_col_out_286;
assign u1_col_in_287 = u0_col_out_287;
assign u1_col_in_288 = u0_col_out_288;
assign u1_col_in_289 = u0_col_out_289;
assign u1_col_in_290 = u0_col_out_290;
assign u1_col_in_291 = u0_col_out_291;
assign u1_col_in_292 = u0_col_out_292;
assign u1_col_in_293 = u0_col_out_293;
assign u1_col_in_294 = u0_col_out_294;
assign u1_col_in_295 = u0_col_out_295;
assign u1_col_in_296 = u0_col_out_296;
assign u1_col_in_297 = u0_col_out_297;
assign u1_col_in_298 = u0_col_out_298;
assign u1_col_in_299 = u0_col_out_299;
assign u1_col_in_300 = u0_col_out_300;
assign u1_col_in_301 = u0_col_out_301;
assign u1_col_in_302 = u0_col_out_302;
assign u1_col_in_303 = u0_col_out_303;
assign u1_col_in_304 = u0_col_out_304;
assign u1_col_in_305 = u0_col_out_305;
assign u1_col_in_306 = u0_col_out_306;
assign u1_col_in_307 = u0_col_out_307;
assign u1_col_in_308 = u0_col_out_308;
assign u1_col_in_309 = u0_col_out_309;
assign u1_col_in_310 = u0_col_out_310;
assign u1_col_in_311 = u0_col_out_311;
assign u1_col_in_312 = u0_col_out_312;
assign u1_col_in_313 = u0_col_out_313;
assign u1_col_in_314 = u0_col_out_314;
assign u1_col_in_315 = u0_col_out_315;
assign u1_col_in_316 = u0_col_out_316;
assign u1_col_in_317 = u0_col_out_317;
assign u1_col_in_318 = u0_col_out_318;
assign u1_col_in_319 = u0_col_out_319;
assign u1_col_in_320 = u0_col_out_320;
assign u1_col_in_321 = u0_col_out_321;
assign u1_col_in_322 = u0_col_out_322;
assign u1_col_in_323 = u0_col_out_323;
assign u1_col_in_324 = u0_col_out_324;
assign u1_col_in_325 = u0_col_out_325;
assign u1_col_in_326 = u0_col_out_326;
assign u1_col_in_327 = u0_col_out_327;
assign u1_col_in_328 = u0_col_out_328;
assign u1_col_in_329 = u0_col_out_329;
assign u1_col_in_330 = u0_col_out_330;
assign u1_col_in_331 = u0_col_out_331;
assign u1_col_in_332 = u0_col_out_332;
assign u1_col_in_333 = u0_col_out_333;
assign u1_col_in_334 = u0_col_out_334;
assign u1_col_in_335 = u0_col_out_335;
assign u1_col_in_336 = u0_col_out_336;
assign u1_col_in_337 = u0_col_out_337;
assign u1_col_in_338 = u0_col_out_338;
assign u1_col_in_339 = u0_col_out_339;
assign u1_col_in_340 = u0_col_out_340;
assign u1_col_in_341 = u0_col_out_341;
assign u1_col_in_342 = u0_col_out_342;
assign u1_col_in_343 = u0_col_out_343;
assign u1_col_in_344 = u0_col_out_344;
assign u1_col_in_345 = u0_col_out_345;
assign u1_col_in_346 = u0_col_out_346;
assign u1_col_in_347 = u0_col_out_347;
assign u1_col_in_348 = u0_col_out_348;
assign u1_col_in_349 = u0_col_out_349;
assign u1_col_in_350 = u0_col_out_350;
assign u1_col_in_351 = u0_col_out_351;
assign u1_col_in_352 = u0_col_out_352;
assign u1_col_in_353 = u0_col_out_353;
assign u1_col_in_354 = u0_col_out_354;
assign u1_col_in_355 = u0_col_out_355;
assign u1_col_in_356 = u0_col_out_356;
assign u1_col_in_357 = u0_col_out_357;
assign u1_col_in_358 = u0_col_out_358;
assign u1_col_in_359 = u0_col_out_359;
assign u1_col_in_360 = u0_col_out_360;
assign u1_col_in_361 = u0_col_out_361;
assign u1_col_in_362 = u0_col_out_362;
assign u1_col_in_363 = u0_col_out_363;
assign u1_col_in_364 = u0_col_out_364;
assign u1_col_in_365 = u0_col_out_365;
assign u1_col_in_366 = u0_col_out_366;
assign u1_col_in_367 = u0_col_out_367;
assign u1_col_in_368 = u0_col_out_368;
assign u1_col_in_369 = u0_col_out_369;
assign u1_col_in_370 = u0_col_out_370;
assign u1_col_in_371 = u0_col_out_371;
assign u1_col_in_372 = u0_col_out_372;
assign u1_col_in_373 = u0_col_out_373;
assign u1_col_in_374 = u0_col_out_374;
assign u1_col_in_375 = u0_col_out_375;
assign u1_col_in_376 = u0_col_out_376;
assign u1_col_in_377 = u0_col_out_377;
assign u1_col_in_378 = u0_col_out_378;
assign u1_col_in_379 = u0_col_out_379;
assign u1_col_in_380 = u0_col_out_380;
assign u1_col_in_381 = u0_col_out_381;
assign u1_col_in_382 = u0_col_out_382;
assign u1_col_in_383 = u0_col_out_383;
assign u1_col_in_384 = u0_col_out_384;
assign u1_col_in_385 = u0_col_out_385;
assign u1_col_in_386 = u0_col_out_386;
assign u1_col_in_387 = u0_col_out_387;
assign u1_col_in_388 = u0_col_out_388;
assign u1_col_in_389 = u0_col_out_389;
assign u1_col_in_390 = u0_col_out_390;
assign u1_col_in_391 = u0_col_out_391;
assign u1_col_in_392 = u0_col_out_392;
assign u1_col_in_393 = u0_col_out_393;
assign u1_col_in_394 = u0_col_out_394;
assign u1_col_in_395 = u0_col_out_395;
assign u1_col_in_396 = u0_col_out_396;
assign u1_col_in_397 = u0_col_out_397;
assign u1_col_in_398 = u0_col_out_398;
assign u1_col_in_399 = u0_col_out_399;
assign u1_col_in_400 = u0_col_out_400;
assign u1_col_in_401 = u0_col_out_401;
assign u1_col_in_402 = u0_col_out_402;
assign u1_col_in_403 = u0_col_out_403;
assign u1_col_in_404 = u0_col_out_404;
assign u1_col_in_405 = u0_col_out_405;
assign u1_col_in_406 = u0_col_out_406;
assign u1_col_in_407 = u0_col_out_407;
assign u1_col_in_408 = u0_col_out_408;
assign u1_col_in_409 = u0_col_out_409;
assign u1_col_in_410 = u0_col_out_410;
assign u1_col_in_411 = u0_col_out_411;
assign u1_col_in_412 = u0_col_out_412;
assign u1_col_in_413 = u0_col_out_413;
assign u1_col_in_414 = u0_col_out_414;
assign u1_col_in_415 = u0_col_out_415;
assign u1_col_in_416 = u0_col_out_416;
assign u1_col_in_417 = u0_col_out_417;
assign u1_col_in_418 = u0_col_out_418;
assign u1_col_in_419 = u0_col_out_419;
assign u1_col_in_420 = u0_col_out_420;
assign u1_col_in_421 = u0_col_out_421;
assign u1_col_in_422 = u0_col_out_422;
assign u1_col_in_423 = u0_col_out_423;
assign u1_col_in_424 = u0_col_out_424;
assign u1_col_in_425 = u0_col_out_425;
assign u1_col_in_426 = u0_col_out_426;
assign u1_col_in_427 = u0_col_out_427;
assign u1_col_in_428 = u0_col_out_428;
assign u1_col_in_429 = u0_col_out_429;
assign u1_col_in_430 = u0_col_out_430;
assign u1_col_in_431 = u0_col_out_431;
assign u1_col_in_432 = u0_col_out_432;
assign u1_col_in_433 = u0_col_out_433;
assign u1_col_in_434 = u0_col_out_434;
assign u1_col_in_435 = u0_col_out_435;
assign u1_col_in_436 = u0_col_out_436;
assign u1_col_in_437 = u0_col_out_437;
assign u1_col_in_438 = u0_col_out_438;
assign u1_col_in_439 = u0_col_out_439;
assign u1_col_in_440 = u0_col_out_440;
assign u1_col_in_441 = u0_col_out_441;
assign u1_col_in_442 = u0_col_out_442;
assign u1_col_in_443 = u0_col_out_443;
assign u1_col_in_444 = u0_col_out_444;
assign u1_col_in_445 = u0_col_out_445;
assign u1_col_in_446 = u0_col_out_446;
assign u1_col_in_447 = u0_col_out_447;
assign u1_col_in_448 = u0_col_out_448;
assign u1_col_in_449 = u0_col_out_449;
assign u1_col_in_450 = u0_col_out_450;
assign u1_col_in_451 = u0_col_out_451;
assign u1_col_in_452 = u0_col_out_452;
assign u1_col_in_453 = u0_col_out_453;
assign u1_col_in_454 = u0_col_out_454;
assign u1_col_in_455 = u0_col_out_455;
assign u1_col_in_456 = u0_col_out_456;
assign u1_col_in_457 = u0_col_out_457;
assign u1_col_in_458 = u0_col_out_458;
assign u1_col_in_459 = u0_col_out_459;
assign u1_col_in_460 = u0_col_out_460;
assign u1_col_in_461 = u0_col_out_461;
assign u1_col_in_462 = u0_col_out_462;
assign u1_col_in_463 = u0_col_out_463;
assign u1_col_in_464 = u0_col_out_464;
assign u1_col_in_465 = u0_col_out_465;
assign u1_col_in_466 = u0_col_out_466;
assign u1_col_in_467 = u0_col_out_467;
assign u1_col_in_468 = u0_col_out_468;
assign u1_col_in_469 = u0_col_out_469;
assign u1_col_in_470 = u0_col_out_470;
assign u1_col_in_471 = u0_col_out_471;
assign u1_col_in_472 = u0_col_out_472;
assign u1_col_in_473 = u0_col_out_473;
assign u1_col_in_474 = u0_col_out_474;
assign u1_col_in_475 = u0_col_out_475;
assign u1_col_in_476 = u0_col_out_476;
assign u1_col_in_477 = u0_col_out_477;
assign u1_col_in_478 = u0_col_out_478;
assign u1_col_in_479 = u0_col_out_479;
assign u1_col_in_480 = u0_col_out_480;
assign u1_col_in_481 = u0_col_out_481;
assign u1_col_in_482 = u0_col_out_482;
assign u1_col_in_483 = u0_col_out_483;
assign u1_col_in_484 = u0_col_out_484;
assign u1_col_in_485 = u0_col_out_485;
assign u1_col_in_486 = u0_col_out_486;
assign u1_col_in_487 = u0_col_out_487;
assign u1_col_in_488 = u0_col_out_488;
assign u1_col_in_489 = u0_col_out_489;
assign u1_col_in_490 = u0_col_out_490;
assign u1_col_in_491 = u0_col_out_491;
assign u1_col_in_492 = u0_col_out_492;
assign u1_col_in_493 = u0_col_out_493;
assign u1_col_in_494 = u0_col_out_494;
assign u1_col_in_495 = u0_col_out_495;
assign u1_col_in_496 = u0_col_out_496;
assign u1_col_in_497 = u0_col_out_497;
assign u1_col_in_498 = u0_col_out_498;
assign u1_col_in_499 = u0_col_out_499;
assign u1_col_in_500 = u0_col_out_500;
assign u1_col_in_501 = u0_col_out_501;
assign u1_col_in_502 = u0_col_out_502;
assign u1_col_in_503 = u0_col_out_503;
assign u1_col_in_504 = u0_col_out_504;
assign u1_col_in_505 = u0_col_out_505;
assign u1_col_in_506 = u0_col_out_506;
assign u1_col_in_507 = u0_col_out_507;
assign u1_col_in_508 = u0_col_out_508;
assign u1_col_in_509 = u0_col_out_509;
assign u1_col_in_510 = u0_col_out_510;
assign u1_col_in_511 = u0_col_out_511;
assign u1_col_in_512 = u0_col_out_512;
assign u1_col_in_513 = u0_col_out_513;
assign u1_col_in_514 = u0_col_out_514;
assign u1_col_in_515 = u0_col_out_515;
assign u1_col_in_516 = u0_col_out_516;
assign u1_col_in_517 = u0_col_out_517;
assign u1_col_in_518 = u0_col_out_518;
assign u1_col_in_519 = u0_col_out_519;
assign u1_col_in_520 = u0_col_out_520;
assign u1_col_in_521 = u0_col_out_521;
assign u1_col_in_522 = u0_col_out_522;
assign u1_col_in_523 = u0_col_out_523;
assign u1_col_in_524 = u0_col_out_524;
assign u1_col_in_525 = u0_col_out_525;
assign u1_col_in_526 = u0_col_out_526;
assign u1_col_in_527 = u0_col_out_527;
assign u1_col_in_528 = u0_col_out_528;
assign u1_col_in_529 = u0_col_out_529;
assign u1_col_in_530 = u0_col_out_530;
assign u1_col_in_531 = u0_col_out_531;
assign u1_col_in_532 = u0_col_out_532;
assign u1_col_in_533 = u0_col_out_533;
assign u1_col_in_534 = u0_col_out_534;
assign u1_col_in_535 = u0_col_out_535;
assign u1_col_in_536 = u0_col_out_536;
assign u1_col_in_537 = u0_col_out_537;
assign u1_col_in_538 = u0_col_out_538;
assign u1_col_in_539 = u0_col_out_539;
assign u1_col_in_540 = u0_col_out_540;
assign u1_col_in_541 = u0_col_out_541;
assign u1_col_in_542 = u0_col_out_542;
assign u1_col_in_543 = u0_col_out_543;
assign u1_col_in_544 = u0_col_out_544;
assign u1_col_in_545 = u0_col_out_545;
assign u1_col_in_546 = u0_col_out_546;
assign u1_col_in_547 = u0_col_out_547;
assign u1_col_in_548 = u0_col_out_548;
assign u1_col_in_549 = u0_col_out_549;
assign u1_col_in_550 = u0_col_out_550;
assign u1_col_in_551 = u0_col_out_551;
assign u1_col_in_552 = u0_col_out_552;
assign u1_col_in_553 = u0_col_out_553;
assign u1_col_in_554 = u0_col_out_554;
assign u1_col_in_555 = u0_col_out_555;
assign u1_col_in_556 = u0_col_out_556;
assign u1_col_in_557 = u0_col_out_557;
assign u1_col_in_558 = u0_col_out_558;
assign u1_col_in_559 = u0_col_out_559;
assign u1_col_in_560 = u0_col_out_560;
assign u1_col_in_561 = u0_col_out_561;
assign u1_col_in_562 = u0_col_out_562;
assign u1_col_in_563 = u0_col_out_563;
assign u1_col_in_564 = u0_col_out_564;
assign u1_col_in_565 = u0_col_out_565;
assign u1_col_in_566 = u0_col_out_566;
assign u1_col_in_567 = u0_col_out_567;
assign u1_col_in_568 = u0_col_out_568;
assign u1_col_in_569 = u0_col_out_569;
assign u1_col_in_570 = u0_col_out_570;
assign u1_col_in_571 = u0_col_out_571;
assign u1_col_in_572 = u0_col_out_572;
assign u1_col_in_573 = u0_col_out_573;
assign u1_col_in_574 = u0_col_out_574;
assign u1_col_in_575 = u0_col_out_575;
assign u1_col_in_576 = u0_col_out_576;
assign u1_col_in_577 = u0_col_out_577;
assign u1_col_in_578 = u0_col_out_578;
assign u1_col_in_579 = u0_col_out_579;
assign u1_col_in_580 = u0_col_out_580;
assign u1_col_in_581 = u0_col_out_581;
assign u1_col_in_582 = u0_col_out_582;
assign u1_col_in_583 = u0_col_out_583;
assign u1_col_in_584 = u0_col_out_584;
assign u1_col_in_585 = u0_col_out_585;
assign u1_col_in_586 = u0_col_out_586;
assign u1_col_in_587 = u0_col_out_587;
assign u1_col_in_588 = u0_col_out_588;
assign u1_col_in_589 = u0_col_out_589;
assign u1_col_in_590 = u0_col_out_590;
assign u1_col_in_591 = u0_col_out_591;
assign u1_col_in_592 = u0_col_out_592;
assign u1_col_in_593 = u0_col_out_593;
assign u1_col_in_594 = u0_col_out_594;
assign u1_col_in_595 = u0_col_out_595;
assign u1_col_in_596 = u0_col_out_596;
assign u1_col_in_597 = u0_col_out_597;
assign u1_col_in_598 = u0_col_out_598;
assign u1_col_in_599 = u0_col_out_599;
assign u1_col_in_600 = u0_col_out_600;
assign u1_col_in_601 = u0_col_out_601;
assign u1_col_in_602 = u0_col_out_602;
assign u1_col_in_603 = u0_col_out_603;
assign u1_col_in_604 = u0_col_out_604;
assign u1_col_in_605 = u0_col_out_605;
assign u1_col_in_606 = u0_col_out_606;
assign u1_col_in_607 = u0_col_out_607;
assign u1_col_in_608 = u0_col_out_608;
assign u1_col_in_609 = u0_col_out_609;
assign u1_col_in_610 = u0_col_out_610;
assign u1_col_in_611 = u0_col_out_611;
assign u1_col_in_612 = u0_col_out_612;
assign u1_col_in_613 = u0_col_out_613;
assign u1_col_in_614 = u0_col_out_614;
assign u1_col_in_615 = u0_col_out_615;
assign u1_col_in_616 = u0_col_out_616;
assign u1_col_in_617 = u0_col_out_617;
assign u1_col_in_618 = u0_col_out_618;
assign u1_col_in_619 = u0_col_out_619;
assign u1_col_in_620 = u0_col_out_620;
assign u1_col_in_621 = u0_col_out_621;
assign u1_col_in_622 = u0_col_out_622;
assign u1_col_in_623 = u0_col_out_623;
assign u1_col_in_624 = u0_col_out_624;
assign u1_col_in_625 = u0_col_out_625;
assign u1_col_in_626 = u0_col_out_626;
assign u1_col_in_627 = u0_col_out_627;
assign u1_col_in_628 = u0_col_out_628;
assign u1_col_in_629 = u0_col_out_629;
assign u1_col_in_630 = u0_col_out_630;
assign u1_col_in_631 = u0_col_out_631;
assign u1_col_in_632 = u0_col_out_632;
assign u1_col_in_633 = u0_col_out_633;
assign u1_col_in_634 = u0_col_out_634;
assign u1_col_in_635 = u0_col_out_635;
assign u1_col_in_636 = u0_col_out_636;
assign u1_col_in_637 = u0_col_out_637;
assign u1_col_in_638 = u0_col_out_638;
assign u1_col_in_639 = u0_col_out_639;
assign u1_col_in_640 = u0_col_out_640;
assign u1_col_in_641 = u0_col_out_641;
assign u1_col_in_642 = u0_col_out_642;
assign u1_col_in_643 = u0_col_out_643;
assign u1_col_in_644 = u0_col_out_644;
assign u1_col_in_645 = u0_col_out_645;
assign u1_col_in_646 = u0_col_out_646;
assign u1_col_in_647 = u0_col_out_647;
assign u1_col_in_648 = u0_col_out_648;
assign u1_col_in_649 = u0_col_out_649;
assign u1_col_in_650 = u0_col_out_650;
assign u1_col_in_651 = u0_col_out_651;
assign u1_col_in_652 = u0_col_out_652;
assign u1_col_in_653 = u0_col_out_653;
assign u1_col_in_654 = u0_col_out_654;
assign u1_col_in_655 = u0_col_out_655;
assign u1_col_in_656 = u0_col_out_656;
assign u1_col_in_657 = u0_col_out_657;
assign u1_col_in_658 = u0_col_out_658;
assign u1_col_in_659 = u0_col_out_659;
assign u1_col_in_660 = u0_col_out_660;
assign u1_col_in_661 = u0_col_out_661;
assign u1_col_in_662 = u0_col_out_662;
assign u1_col_in_663 = u0_col_out_663;
assign u1_col_in_664 = u0_col_out_664;
assign u1_col_in_665 = u0_col_out_665;
assign u1_col_in_666 = u0_col_out_666;
assign u1_col_in_667 = u0_col_out_667;
assign u1_col_in_668 = u0_col_out_668;
assign u1_col_in_669 = u0_col_out_669;
assign u1_col_in_670 = u0_col_out_670;
assign u1_col_in_671 = u0_col_out_671;
assign u1_col_in_672 = u0_col_out_672;
assign u1_col_in_673 = u0_col_out_673;
assign u1_col_in_674 = u0_col_out_674;
assign u1_col_in_675 = u0_col_out_675;
assign u1_col_in_676 = u0_col_out_676;
assign u1_col_in_677 = u0_col_out_677;
assign u1_col_in_678 = u0_col_out_678;
assign u1_col_in_679 = u0_col_out_679;
assign u1_col_in_680 = u0_col_out_680;
assign u1_col_in_681 = u0_col_out_681;
assign u1_col_in_682 = u0_col_out_682;
assign u1_col_in_683 = u0_col_out_683;
assign u1_col_in_684 = u0_col_out_684;
assign u1_col_in_685 = u0_col_out_685;
assign u1_col_in_686 = u0_col_out_686;
assign u1_col_in_687 = u0_col_out_687;
assign u1_col_in_688 = u0_col_out_688;
assign u1_col_in_689 = u0_col_out_689;
assign u1_col_in_690 = u0_col_out_690;
assign u1_col_in_691 = u0_col_out_691;
assign u1_col_in_692 = u0_col_out_692;
assign u1_col_in_693 = u0_col_out_693;
assign u1_col_in_694 = u0_col_out_694;
assign u1_col_in_695 = u0_col_out_695;
assign u1_col_in_696 = u0_col_out_696;
assign u1_col_in_697 = u0_col_out_697;
assign u1_col_in_698 = u0_col_out_698;
assign u1_col_in_699 = u0_col_out_699;
assign u1_col_in_700 = u0_col_out_700;
assign u1_col_in_701 = u0_col_out_701;
assign u1_col_in_702 = u0_col_out_702;
assign u1_col_in_703 = u0_col_out_703;
assign u1_col_in_704 = u0_col_out_704;
assign u1_col_in_705 = u0_col_out_705;
assign u1_col_in_706 = u0_col_out_706;
assign u1_col_in_707 = u0_col_out_707;
assign u1_col_in_708 = u0_col_out_708;
assign u1_col_in_709 = u0_col_out_709;
assign u1_col_in_710 = u0_col_out_710;
assign u1_col_in_711 = u0_col_out_711;
assign u1_col_in_712 = u0_col_out_712;
assign u1_col_in_713 = u0_col_out_713;
assign u1_col_in_714 = u0_col_out_714;
assign u1_col_in_715 = u0_col_out_715;
assign u1_col_in_716 = u0_col_out_716;
assign u1_col_in_717 = u0_col_out_717;
assign u1_col_in_718 = u0_col_out_718;
assign u1_col_in_719 = u0_col_out_719;
assign u1_col_in_720 = u0_col_out_720;
assign u1_col_in_721 = u0_col_out_721;
assign u1_col_in_722 = u0_col_out_722;
assign u1_col_in_723 = u0_col_out_723;
assign u1_col_in_724 = u0_col_out_724;
assign u1_col_in_725 = u0_col_out_725;
assign u1_col_in_726 = u0_col_out_726;
assign u1_col_in_727 = u0_col_out_727;
assign u1_col_in_728 = u0_col_out_728;
assign u1_col_in_729 = u0_col_out_729;
assign u1_col_in_730 = u0_col_out_730;
assign u1_col_in_731 = u0_col_out_731;
assign u1_col_in_732 = u0_col_out_732;
assign u1_col_in_733 = u0_col_out_733;
assign u1_col_in_734 = u0_col_out_734;
assign u1_col_in_735 = u0_col_out_735;
assign u1_col_in_736 = u0_col_out_736;
assign u1_col_in_737 = u0_col_out_737;
assign u1_col_in_738 = u0_col_out_738;
assign u1_col_in_739 = u0_col_out_739;
assign u1_col_in_740 = u0_col_out_740;
assign u1_col_in_741 = u0_col_out_741;
assign u1_col_in_742 = u0_col_out_742;
assign u1_col_in_743 = u0_col_out_743;
assign u1_col_in_744 = u0_col_out_744;
assign u1_col_in_745 = u0_col_out_745;
assign u1_col_in_746 = u0_col_out_746;
assign u1_col_in_747 = u0_col_out_747;
assign u1_col_in_748 = u0_col_out_748;
assign u1_col_in_749 = u0_col_out_749;
assign u1_col_in_750 = u0_col_out_750;
assign u1_col_in_751 = u0_col_out_751;
assign u1_col_in_752 = u0_col_out_752;
assign u1_col_in_753 = u0_col_out_753;
assign u1_col_in_754 = u0_col_out_754;
assign u1_col_in_755 = u0_col_out_755;
assign u1_col_in_756 = u0_col_out_756;
assign u1_col_in_757 = u0_col_out_757;
assign u1_col_in_758 = u0_col_out_758;
assign u1_col_in_759 = u0_col_out_759;
assign u1_col_in_760 = u0_col_out_760;
assign u1_col_in_761 = u0_col_out_761;
assign u1_col_in_762 = u0_col_out_762;
assign u1_col_in_763 = u0_col_out_763;
assign u1_col_in_764 = u0_col_out_764;
assign u1_col_in_765 = u0_col_out_765;
assign u1_col_in_766 = u0_col_out_766;
assign u1_col_in_767 = u0_col_out_767;
assign u1_col_in_768 = u0_col_out_768;
assign u1_col_in_769 = u0_col_out_769;
assign u1_col_in_770 = u0_col_out_770;
assign u1_col_in_771 = u0_col_out_771;
assign u1_col_in_772 = u0_col_out_772;
assign u1_col_in_773 = u0_col_out_773;
assign u1_col_in_774 = u0_col_out_774;
assign u1_col_in_775 = u0_col_out_775;
assign u1_col_in_776 = u0_col_out_776;
assign u1_col_in_777 = u0_col_out_777;
assign u1_col_in_778 = u0_col_out_778;
assign u1_col_in_779 = u0_col_out_779;
assign u1_col_in_780 = u0_col_out_780;
assign u1_col_in_781 = u0_col_out_781;
assign u1_col_in_782 = u0_col_out_782;
assign u1_col_in_783 = u0_col_out_783;
assign u1_col_in_784 = u0_col_out_784;
assign u1_col_in_785 = u0_col_out_785;
assign u1_col_in_786 = u0_col_out_786;
assign u1_col_in_787 = u0_col_out_787;
assign u1_col_in_788 = u0_col_out_788;
assign u1_col_in_789 = u0_col_out_789;
assign u1_col_in_790 = u0_col_out_790;
assign u1_col_in_791 = u0_col_out_791;
assign u1_col_in_792 = u0_col_out_792;
assign u1_col_in_793 = u0_col_out_793;
assign u1_col_in_794 = u0_col_out_794;
assign u1_col_in_795 = u0_col_out_795;
assign u1_col_in_796 = u0_col_out_796;
assign u1_col_in_797 = u0_col_out_797;
assign u1_col_in_798 = u0_col_out_798;
assign u1_col_in_799 = u0_col_out_799;
assign u1_col_in_800 = u0_col_out_800;
assign u1_col_in_801 = u0_col_out_801;
assign u1_col_in_802 = u0_col_out_802;
assign u1_col_in_803 = u0_col_out_803;
assign u1_col_in_804 = u0_col_out_804;
assign u1_col_in_805 = u0_col_out_805;
assign u1_col_in_806 = u0_col_out_806;
assign u1_col_in_807 = u0_col_out_807;
assign u1_col_in_808 = u0_col_out_808;
assign u1_col_in_809 = u0_col_out_809;
assign u1_col_in_810 = u0_col_out_810;
assign u1_col_in_811 = u0_col_out_811;
assign u1_col_in_812 = u0_col_out_812;
assign u1_col_in_813 = u0_col_out_813;
assign u1_col_in_814 = u0_col_out_814;
assign u1_col_in_815 = u0_col_out_815;
assign u1_col_in_816 = u0_col_out_816;
assign u1_col_in_817 = u0_col_out_817;
assign u1_col_in_818 = u0_col_out_818;
assign u1_col_in_819 = u0_col_out_819;
assign u1_col_in_820 = u0_col_out_820;
assign u1_col_in_821 = u0_col_out_821;
assign u1_col_in_822 = u0_col_out_822;
assign u1_col_in_823 = u0_col_out_823;
assign u1_col_in_824 = u0_col_out_824;
assign u1_col_in_825 = u0_col_out_825;
assign u1_col_in_826 = u0_col_out_826;
assign u1_col_in_827 = u0_col_out_827;
assign u1_col_in_828 = u0_col_out_828;
assign u1_col_in_829 = u0_col_out_829;
assign u1_col_in_830 = u0_col_out_830;
assign u1_col_in_831 = u0_col_out_831;
assign u1_col_in_832 = u0_col_out_832;
assign u1_col_in_833 = u0_col_out_833;
assign u1_col_in_834 = u0_col_out_834;
assign u1_col_in_835 = u0_col_out_835;
assign u1_col_in_836 = u0_col_out_836;
assign u1_col_in_837 = u0_col_out_837;
assign u1_col_in_838 = u0_col_out_838;
assign u1_col_in_839 = u0_col_out_839;
assign u1_col_in_840 = u0_col_out_840;
assign u1_col_in_841 = u0_col_out_841;
assign u1_col_in_842 = u0_col_out_842;
assign u1_col_in_843 = u0_col_out_843;
assign u1_col_in_844 = u0_col_out_844;
assign u1_col_in_845 = u0_col_out_845;
assign u1_col_in_846 = u0_col_out_846;
assign u1_col_in_847 = u0_col_out_847;
assign u1_col_in_848 = u0_col_out_848;
assign u1_col_in_849 = u0_col_out_849;
assign u1_col_in_850 = u0_col_out_850;
assign u1_col_in_851 = u0_col_out_851;
assign u1_col_in_852 = u0_col_out_852;
assign u1_col_in_853 = u0_col_out_853;
assign u1_col_in_854 = u0_col_out_854;
assign u1_col_in_855 = u0_col_out_855;
assign u1_col_in_856 = u0_col_out_856;
assign u1_col_in_857 = u0_col_out_857;
assign u1_col_in_858 = u0_col_out_858;
assign u1_col_in_859 = u0_col_out_859;
assign u1_col_in_860 = u0_col_out_860;
assign u1_col_in_861 = u0_col_out_861;
assign u1_col_in_862 = u0_col_out_862;
assign u1_col_in_863 = u0_col_out_863;
assign u1_col_in_864 = u0_col_out_864;
assign u1_col_in_865 = u0_col_out_865;
assign u1_col_in_866 = u0_col_out_866;
assign u1_col_in_867 = u0_col_out_867;
assign u1_col_in_868 = u0_col_out_868;
assign u1_col_in_869 = u0_col_out_869;
assign u1_col_in_870 = u0_col_out_870;
assign u1_col_in_871 = u0_col_out_871;
assign u1_col_in_872 = u0_col_out_872;
assign u1_col_in_873 = u0_col_out_873;
assign u1_col_in_874 = u0_col_out_874;
assign u1_col_in_875 = u0_col_out_875;
assign u1_col_in_876 = u0_col_out_876;
assign u1_col_in_877 = u0_col_out_877;
assign u1_col_in_878 = u0_col_out_878;
assign u1_col_in_879 = u0_col_out_879;
assign u1_col_in_880 = u0_col_out_880;
assign u1_col_in_881 = u0_col_out_881;
assign u1_col_in_882 = u0_col_out_882;
assign u1_col_in_883 = u0_col_out_883;
assign u1_col_in_884 = u0_col_out_884;
assign u1_col_in_885 = u0_col_out_885;
assign u1_col_in_886 = u0_col_out_886;
assign u1_col_in_887 = u0_col_out_887;
assign u1_col_in_888 = u0_col_out_888;
assign u1_col_in_889 = u0_col_out_889;
assign u1_col_in_890 = u0_col_out_890;
assign u1_col_in_891 = u0_col_out_891;
assign u1_col_in_892 = u0_col_out_892;
assign u1_col_in_893 = u0_col_out_893;
assign u1_col_in_894 = u0_col_out_894;
assign u1_col_in_895 = u0_col_out_895;
assign u1_col_in_896 = u0_col_out_896;
assign u1_col_in_897 = u0_col_out_897;
assign u1_col_in_898 = u0_col_out_898;
assign u1_col_in_899 = u0_col_out_899;
assign u1_col_in_900 = u0_col_out_900;
assign u1_col_in_901 = u0_col_out_901;
assign u1_col_in_902 = u0_col_out_902;
assign u1_col_in_903 = u0_col_out_903;
assign u1_col_in_904 = u0_col_out_904;
assign u1_col_in_905 = u0_col_out_905;
assign u1_col_in_906 = u0_col_out_906;
assign u1_col_in_907 = u0_col_out_907;
assign u1_col_in_908 = u0_col_out_908;
assign u1_col_in_909 = u0_col_out_909;
assign u1_col_in_910 = u0_col_out_910;
assign u1_col_in_911 = u0_col_out_911;
assign u1_col_in_912 = u0_col_out_912;
assign u1_col_in_913 = u0_col_out_913;
assign u1_col_in_914 = u0_col_out_914;
assign u1_col_in_915 = u0_col_out_915;
assign u1_col_in_916 = u0_col_out_916;
assign u1_col_in_917 = u0_col_out_917;
assign u1_col_in_918 = u0_col_out_918;
assign u1_col_in_919 = u0_col_out_919;
assign u1_col_in_920 = u0_col_out_920;
assign u1_col_in_921 = u0_col_out_921;
assign u1_col_in_922 = u0_col_out_922;
assign u1_col_in_923 = u0_col_out_923;
assign u1_col_in_924 = u0_col_out_924;
assign u1_col_in_925 = u0_col_out_925;
assign u1_col_in_926 = u0_col_out_926;
assign u1_col_in_927 = u0_col_out_927;
assign u1_col_in_928 = u0_col_out_928;
assign u1_col_in_929 = u0_col_out_929;
assign u1_col_in_930 = u0_col_out_930;
assign u1_col_in_931 = u0_col_out_931;
assign u1_col_in_932 = u0_col_out_932;
assign u1_col_in_933 = u0_col_out_933;
assign u1_col_in_934 = u0_col_out_934;
assign u1_col_in_935 = u0_col_out_935;
assign u1_col_in_936 = u0_col_out_936;
assign u1_col_in_937 = u0_col_out_937;
assign u1_col_in_938 = u0_col_out_938;
assign u1_col_in_939 = u0_col_out_939;
assign u1_col_in_940 = u0_col_out_940;
assign u1_col_in_941 = u0_col_out_941;
assign u1_col_in_942 = u0_col_out_942;
assign u1_col_in_943 = u0_col_out_943;
assign u1_col_in_944 = u0_col_out_944;
assign u1_col_in_945 = u0_col_out_945;
assign u1_col_in_946 = u0_col_out_946;
assign u1_col_in_947 = u0_col_out_947;
assign u1_col_in_948 = u0_col_out_948;
assign u1_col_in_949 = u0_col_out_949;
assign u1_col_in_950 = u0_col_out_950;
assign u1_col_in_951 = u0_col_out_951;
assign u1_col_in_952 = u0_col_out_952;
assign u1_col_in_953 = u0_col_out_953;
assign u1_col_in_954 = u0_col_out_954;
assign u1_col_in_955 = u0_col_out_955;
assign u1_col_in_956 = u0_col_out_956;
assign u1_col_in_957 = u0_col_out_957;
assign u1_col_in_958 = u0_col_out_958;
assign u1_col_in_959 = u0_col_out_959;
assign u1_col_in_960 = u0_col_out_960;
assign u1_col_in_961 = u0_col_out_961;
assign u1_col_in_962 = u0_col_out_962;
assign u1_col_in_963 = u0_col_out_963;
assign u1_col_in_964 = u0_col_out_964;
assign u1_col_in_965 = u0_col_out_965;
assign u1_col_in_966 = u0_col_out_966;
assign u1_col_in_967 = u0_col_out_967;
assign u1_col_in_968 = u0_col_out_968;
assign u1_col_in_969 = u0_col_out_969;
assign u1_col_in_970 = u0_col_out_970;
assign u1_col_in_971 = u0_col_out_971;
assign u1_col_in_972 = u0_col_out_972;
assign u1_col_in_973 = u0_col_out_973;
assign u1_col_in_974 = u0_col_out_974;
assign u1_col_in_975 = u0_col_out_975;
assign u1_col_in_976 = u0_col_out_976;
assign u1_col_in_977 = u0_col_out_977;
assign u1_col_in_978 = u0_col_out_978;
assign u1_col_in_979 = u0_col_out_979;
assign u1_col_in_980 = u0_col_out_980;
assign u1_col_in_981 = u0_col_out_981;
assign u1_col_in_982 = u0_col_out_982;
assign u1_col_in_983 = u0_col_out_983;
assign u1_col_in_984 = u0_col_out_984;
assign u1_col_in_985 = u0_col_out_985;
assign u1_col_in_986 = u0_col_out_986;
assign u1_col_in_987 = u0_col_out_987;
assign u1_col_in_988 = u0_col_out_988;
assign u1_col_in_989 = u0_col_out_989;
assign u1_col_in_990 = u0_col_out_990;
assign u1_col_in_991 = u0_col_out_991;
assign u1_col_in_992 = u0_col_out_992;
assign u1_col_in_993 = u0_col_out_993;
assign u1_col_in_994 = u0_col_out_994;
assign u1_col_in_995 = u0_col_out_995;
assign u1_col_in_996 = u0_col_out_996;
assign u1_col_in_997 = u0_col_out_997;
assign u1_col_in_998 = u0_col_out_998;
assign u1_col_in_999 = u0_col_out_999;
assign u1_col_in_1000 = u0_col_out_1000;
assign u1_col_in_1001 = u0_col_out_1001;
assign u1_col_in_1002 = u0_col_out_1002;
assign u1_col_in_1003 = u0_col_out_1003;
assign u1_col_in_1004 = u0_col_out_1004;
assign u1_col_in_1005 = u0_col_out_1005;
assign u1_col_in_1006 = u0_col_out_1006;
assign u1_col_in_1007 = u0_col_out_1007;
assign u1_col_in_1008 = u0_col_out_1008;
assign u1_col_in_1009 = u0_col_out_1009;
assign u1_col_in_1010 = u0_col_out_1010;
assign u1_col_in_1011 = u0_col_out_1011;
assign u1_col_in_1012 = u0_col_out_1012;
assign u1_col_in_1013 = u0_col_out_1013;
assign u1_col_in_1014 = u0_col_out_1014;
assign u1_col_in_1015 = u0_col_out_1015;
assign u1_col_in_1016 = u0_col_out_1016;
assign u1_col_in_1017 = u0_col_out_1017;
assign u1_col_in_1018 = u0_col_out_1018;
assign u1_col_in_1019 = u0_col_out_1019;
assign u1_col_in_1020 = u0_col_out_1020;
assign u1_col_in_1021 = u0_col_out_1021;
assign u1_col_in_1022 = u0_col_out_1022;
assign u1_col_in_1023 = u0_col_out_1023;
assign u1_col_in_1024 = u0_col_out_1024;
assign u1_col_in_1025 = u0_col_out_1025;
assign u1_col_in_1026 = u0_col_out_1026;

//*****************************************************
//**************u1压缩阵列******************************
//*****************************************************
compressor_array_152_48_1027 u1_ca_152_48_1027
(
    .col_in_0(u1_col_in_0),
    .col_in_1(u1_col_in_1),
    .col_in_2(u1_col_in_2),
    .col_in_3(u1_col_in_3),
    .col_in_4(u1_col_in_4),
    .col_in_5(u1_col_in_5),
    .col_in_6(u1_col_in_6),
    .col_in_7(u1_col_in_7),
    .col_in_8(u1_col_in_8),
    .col_in_9(u1_col_in_9),
    .col_in_10(u1_col_in_10),
    .col_in_11(u1_col_in_11),
    .col_in_12(u1_col_in_12),
    .col_in_13(u1_col_in_13),
    .col_in_14(u1_col_in_14),
    .col_in_15(u1_col_in_15),
    .col_in_16(u1_col_in_16),
    .col_in_17(u1_col_in_17),
    .col_in_18(u1_col_in_18),
    .col_in_19(u1_col_in_19),
    .col_in_20(u1_col_in_20),
    .col_in_21(u1_col_in_21),
    .col_in_22(u1_col_in_22),
    .col_in_23(u1_col_in_23),
    .col_in_24(u1_col_in_24),
    .col_in_25(u1_col_in_25),
    .col_in_26(u1_col_in_26),
    .col_in_27(u1_col_in_27),
    .col_in_28(u1_col_in_28),
    .col_in_29(u1_col_in_29),
    .col_in_30(u1_col_in_30),
    .col_in_31(u1_col_in_31),
    .col_in_32(u1_col_in_32),
    .col_in_33(u1_col_in_33),
    .col_in_34(u1_col_in_34),
    .col_in_35(u1_col_in_35),
    .col_in_36(u1_col_in_36),
    .col_in_37(u1_col_in_37),
    .col_in_38(u1_col_in_38),
    .col_in_39(u1_col_in_39),
    .col_in_40(u1_col_in_40),
    .col_in_41(u1_col_in_41),
    .col_in_42(u1_col_in_42),
    .col_in_43(u1_col_in_43),
    .col_in_44(u1_col_in_44),
    .col_in_45(u1_col_in_45),
    .col_in_46(u1_col_in_46),
    .col_in_47(u1_col_in_47),
    .col_in_48(u1_col_in_48),
    .col_in_49(u1_col_in_49),
    .col_in_50(u1_col_in_50),
    .col_in_51(u1_col_in_51),
    .col_in_52(u1_col_in_52),
    .col_in_53(u1_col_in_53),
    .col_in_54(u1_col_in_54),
    .col_in_55(u1_col_in_55),
    .col_in_56(u1_col_in_56),
    .col_in_57(u1_col_in_57),
    .col_in_58(u1_col_in_58),
    .col_in_59(u1_col_in_59),
    .col_in_60(u1_col_in_60),
    .col_in_61(u1_col_in_61),
    .col_in_62(u1_col_in_62),
    .col_in_63(u1_col_in_63),
    .col_in_64(u1_col_in_64),
    .col_in_65(u1_col_in_65),
    .col_in_66(u1_col_in_66),
    .col_in_67(u1_col_in_67),
    .col_in_68(u1_col_in_68),
    .col_in_69(u1_col_in_69),
    .col_in_70(u1_col_in_70),
    .col_in_71(u1_col_in_71),
    .col_in_72(u1_col_in_72),
    .col_in_73(u1_col_in_73),
    .col_in_74(u1_col_in_74),
    .col_in_75(u1_col_in_75),
    .col_in_76(u1_col_in_76),
    .col_in_77(u1_col_in_77),
    .col_in_78(u1_col_in_78),
    .col_in_79(u1_col_in_79),
    .col_in_80(u1_col_in_80),
    .col_in_81(u1_col_in_81),
    .col_in_82(u1_col_in_82),
    .col_in_83(u1_col_in_83),
    .col_in_84(u1_col_in_84),
    .col_in_85(u1_col_in_85),
    .col_in_86(u1_col_in_86),
    .col_in_87(u1_col_in_87),
    .col_in_88(u1_col_in_88),
    .col_in_89(u1_col_in_89),
    .col_in_90(u1_col_in_90),
    .col_in_91(u1_col_in_91),
    .col_in_92(u1_col_in_92),
    .col_in_93(u1_col_in_93),
    .col_in_94(u1_col_in_94),
    .col_in_95(u1_col_in_95),
    .col_in_96(u1_col_in_96),
    .col_in_97(u1_col_in_97),
    .col_in_98(u1_col_in_98),
    .col_in_99(u1_col_in_99),
    .col_in_100(u1_col_in_100),
    .col_in_101(u1_col_in_101),
    .col_in_102(u1_col_in_102),
    .col_in_103(u1_col_in_103),
    .col_in_104(u1_col_in_104),
    .col_in_105(u1_col_in_105),
    .col_in_106(u1_col_in_106),
    .col_in_107(u1_col_in_107),
    .col_in_108(u1_col_in_108),
    .col_in_109(u1_col_in_109),
    .col_in_110(u1_col_in_110),
    .col_in_111(u1_col_in_111),
    .col_in_112(u1_col_in_112),
    .col_in_113(u1_col_in_113),
    .col_in_114(u1_col_in_114),
    .col_in_115(u1_col_in_115),
    .col_in_116(u1_col_in_116),
    .col_in_117(u1_col_in_117),
    .col_in_118(u1_col_in_118),
    .col_in_119(u1_col_in_119),
    .col_in_120(u1_col_in_120),
    .col_in_121(u1_col_in_121),
    .col_in_122(u1_col_in_122),
    .col_in_123(u1_col_in_123),
    .col_in_124(u1_col_in_124),
    .col_in_125(u1_col_in_125),
    .col_in_126(u1_col_in_126),
    .col_in_127(u1_col_in_127),
    .col_in_128(u1_col_in_128),
    .col_in_129(u1_col_in_129),
    .col_in_130(u1_col_in_130),
    .col_in_131(u1_col_in_131),
    .col_in_132(u1_col_in_132),
    .col_in_133(u1_col_in_133),
    .col_in_134(u1_col_in_134),
    .col_in_135(u1_col_in_135),
    .col_in_136(u1_col_in_136),
    .col_in_137(u1_col_in_137),
    .col_in_138(u1_col_in_138),
    .col_in_139(u1_col_in_139),
    .col_in_140(u1_col_in_140),
    .col_in_141(u1_col_in_141),
    .col_in_142(u1_col_in_142),
    .col_in_143(u1_col_in_143),
    .col_in_144(u1_col_in_144),
    .col_in_145(u1_col_in_145),
    .col_in_146(u1_col_in_146),
    .col_in_147(u1_col_in_147),
    .col_in_148(u1_col_in_148),
    .col_in_149(u1_col_in_149),
    .col_in_150(u1_col_in_150),
    .col_in_151(u1_col_in_151),
    .col_in_152(u1_col_in_152),
    .col_in_153(u1_col_in_153),
    .col_in_154(u1_col_in_154),
    .col_in_155(u1_col_in_155),
    .col_in_156(u1_col_in_156),
    .col_in_157(u1_col_in_157),
    .col_in_158(u1_col_in_158),
    .col_in_159(u1_col_in_159),
    .col_in_160(u1_col_in_160),
    .col_in_161(u1_col_in_161),
    .col_in_162(u1_col_in_162),
    .col_in_163(u1_col_in_163),
    .col_in_164(u1_col_in_164),
    .col_in_165(u1_col_in_165),
    .col_in_166(u1_col_in_166),
    .col_in_167(u1_col_in_167),
    .col_in_168(u1_col_in_168),
    .col_in_169(u1_col_in_169),
    .col_in_170(u1_col_in_170),
    .col_in_171(u1_col_in_171),
    .col_in_172(u1_col_in_172),
    .col_in_173(u1_col_in_173),
    .col_in_174(u1_col_in_174),
    .col_in_175(u1_col_in_175),
    .col_in_176(u1_col_in_176),
    .col_in_177(u1_col_in_177),
    .col_in_178(u1_col_in_178),
    .col_in_179(u1_col_in_179),
    .col_in_180(u1_col_in_180),
    .col_in_181(u1_col_in_181),
    .col_in_182(u1_col_in_182),
    .col_in_183(u1_col_in_183),
    .col_in_184(u1_col_in_184),
    .col_in_185(u1_col_in_185),
    .col_in_186(u1_col_in_186),
    .col_in_187(u1_col_in_187),
    .col_in_188(u1_col_in_188),
    .col_in_189(u1_col_in_189),
    .col_in_190(u1_col_in_190),
    .col_in_191(u1_col_in_191),
    .col_in_192(u1_col_in_192),
    .col_in_193(u1_col_in_193),
    .col_in_194(u1_col_in_194),
    .col_in_195(u1_col_in_195),
    .col_in_196(u1_col_in_196),
    .col_in_197(u1_col_in_197),
    .col_in_198(u1_col_in_198),
    .col_in_199(u1_col_in_199),
    .col_in_200(u1_col_in_200),
    .col_in_201(u1_col_in_201),
    .col_in_202(u1_col_in_202),
    .col_in_203(u1_col_in_203),
    .col_in_204(u1_col_in_204),
    .col_in_205(u1_col_in_205),
    .col_in_206(u1_col_in_206),
    .col_in_207(u1_col_in_207),
    .col_in_208(u1_col_in_208),
    .col_in_209(u1_col_in_209),
    .col_in_210(u1_col_in_210),
    .col_in_211(u1_col_in_211),
    .col_in_212(u1_col_in_212),
    .col_in_213(u1_col_in_213),
    .col_in_214(u1_col_in_214),
    .col_in_215(u1_col_in_215),
    .col_in_216(u1_col_in_216),
    .col_in_217(u1_col_in_217),
    .col_in_218(u1_col_in_218),
    .col_in_219(u1_col_in_219),
    .col_in_220(u1_col_in_220),
    .col_in_221(u1_col_in_221),
    .col_in_222(u1_col_in_222),
    .col_in_223(u1_col_in_223),
    .col_in_224(u1_col_in_224),
    .col_in_225(u1_col_in_225),
    .col_in_226(u1_col_in_226),
    .col_in_227(u1_col_in_227),
    .col_in_228(u1_col_in_228),
    .col_in_229(u1_col_in_229),
    .col_in_230(u1_col_in_230),
    .col_in_231(u1_col_in_231),
    .col_in_232(u1_col_in_232),
    .col_in_233(u1_col_in_233),
    .col_in_234(u1_col_in_234),
    .col_in_235(u1_col_in_235),
    .col_in_236(u1_col_in_236),
    .col_in_237(u1_col_in_237),
    .col_in_238(u1_col_in_238),
    .col_in_239(u1_col_in_239),
    .col_in_240(u1_col_in_240),
    .col_in_241(u1_col_in_241),
    .col_in_242(u1_col_in_242),
    .col_in_243(u1_col_in_243),
    .col_in_244(u1_col_in_244),
    .col_in_245(u1_col_in_245),
    .col_in_246(u1_col_in_246),
    .col_in_247(u1_col_in_247),
    .col_in_248(u1_col_in_248),
    .col_in_249(u1_col_in_249),
    .col_in_250(u1_col_in_250),
    .col_in_251(u1_col_in_251),
    .col_in_252(u1_col_in_252),
    .col_in_253(u1_col_in_253),
    .col_in_254(u1_col_in_254),
    .col_in_255(u1_col_in_255),
    .col_in_256(u1_col_in_256),
    .col_in_257(u1_col_in_257),
    .col_in_258(u1_col_in_258),
    .col_in_259(u1_col_in_259),
    .col_in_260(u1_col_in_260),
    .col_in_261(u1_col_in_261),
    .col_in_262(u1_col_in_262),
    .col_in_263(u1_col_in_263),
    .col_in_264(u1_col_in_264),
    .col_in_265(u1_col_in_265),
    .col_in_266(u1_col_in_266),
    .col_in_267(u1_col_in_267),
    .col_in_268(u1_col_in_268),
    .col_in_269(u1_col_in_269),
    .col_in_270(u1_col_in_270),
    .col_in_271(u1_col_in_271),
    .col_in_272(u1_col_in_272),
    .col_in_273(u1_col_in_273),
    .col_in_274(u1_col_in_274),
    .col_in_275(u1_col_in_275),
    .col_in_276(u1_col_in_276),
    .col_in_277(u1_col_in_277),
    .col_in_278(u1_col_in_278),
    .col_in_279(u1_col_in_279),
    .col_in_280(u1_col_in_280),
    .col_in_281(u1_col_in_281),
    .col_in_282(u1_col_in_282),
    .col_in_283(u1_col_in_283),
    .col_in_284(u1_col_in_284),
    .col_in_285(u1_col_in_285),
    .col_in_286(u1_col_in_286),
    .col_in_287(u1_col_in_287),
    .col_in_288(u1_col_in_288),
    .col_in_289(u1_col_in_289),
    .col_in_290(u1_col_in_290),
    .col_in_291(u1_col_in_291),
    .col_in_292(u1_col_in_292),
    .col_in_293(u1_col_in_293),
    .col_in_294(u1_col_in_294),
    .col_in_295(u1_col_in_295),
    .col_in_296(u1_col_in_296),
    .col_in_297(u1_col_in_297),
    .col_in_298(u1_col_in_298),
    .col_in_299(u1_col_in_299),
    .col_in_300(u1_col_in_300),
    .col_in_301(u1_col_in_301),
    .col_in_302(u1_col_in_302),
    .col_in_303(u1_col_in_303),
    .col_in_304(u1_col_in_304),
    .col_in_305(u1_col_in_305),
    .col_in_306(u1_col_in_306),
    .col_in_307(u1_col_in_307),
    .col_in_308(u1_col_in_308),
    .col_in_309(u1_col_in_309),
    .col_in_310(u1_col_in_310),
    .col_in_311(u1_col_in_311),
    .col_in_312(u1_col_in_312),
    .col_in_313(u1_col_in_313),
    .col_in_314(u1_col_in_314),
    .col_in_315(u1_col_in_315),
    .col_in_316(u1_col_in_316),
    .col_in_317(u1_col_in_317),
    .col_in_318(u1_col_in_318),
    .col_in_319(u1_col_in_319),
    .col_in_320(u1_col_in_320),
    .col_in_321(u1_col_in_321),
    .col_in_322(u1_col_in_322),
    .col_in_323(u1_col_in_323),
    .col_in_324(u1_col_in_324),
    .col_in_325(u1_col_in_325),
    .col_in_326(u1_col_in_326),
    .col_in_327(u1_col_in_327),
    .col_in_328(u1_col_in_328),
    .col_in_329(u1_col_in_329),
    .col_in_330(u1_col_in_330),
    .col_in_331(u1_col_in_331),
    .col_in_332(u1_col_in_332),
    .col_in_333(u1_col_in_333),
    .col_in_334(u1_col_in_334),
    .col_in_335(u1_col_in_335),
    .col_in_336(u1_col_in_336),
    .col_in_337(u1_col_in_337),
    .col_in_338(u1_col_in_338),
    .col_in_339(u1_col_in_339),
    .col_in_340(u1_col_in_340),
    .col_in_341(u1_col_in_341),
    .col_in_342(u1_col_in_342),
    .col_in_343(u1_col_in_343),
    .col_in_344(u1_col_in_344),
    .col_in_345(u1_col_in_345),
    .col_in_346(u1_col_in_346),
    .col_in_347(u1_col_in_347),
    .col_in_348(u1_col_in_348),
    .col_in_349(u1_col_in_349),
    .col_in_350(u1_col_in_350),
    .col_in_351(u1_col_in_351),
    .col_in_352(u1_col_in_352),
    .col_in_353(u1_col_in_353),
    .col_in_354(u1_col_in_354),
    .col_in_355(u1_col_in_355),
    .col_in_356(u1_col_in_356),
    .col_in_357(u1_col_in_357),
    .col_in_358(u1_col_in_358),
    .col_in_359(u1_col_in_359),
    .col_in_360(u1_col_in_360),
    .col_in_361(u1_col_in_361),
    .col_in_362(u1_col_in_362),
    .col_in_363(u1_col_in_363),
    .col_in_364(u1_col_in_364),
    .col_in_365(u1_col_in_365),
    .col_in_366(u1_col_in_366),
    .col_in_367(u1_col_in_367),
    .col_in_368(u1_col_in_368),
    .col_in_369(u1_col_in_369),
    .col_in_370(u1_col_in_370),
    .col_in_371(u1_col_in_371),
    .col_in_372(u1_col_in_372),
    .col_in_373(u1_col_in_373),
    .col_in_374(u1_col_in_374),
    .col_in_375(u1_col_in_375),
    .col_in_376(u1_col_in_376),
    .col_in_377(u1_col_in_377),
    .col_in_378(u1_col_in_378),
    .col_in_379(u1_col_in_379),
    .col_in_380(u1_col_in_380),
    .col_in_381(u1_col_in_381),
    .col_in_382(u1_col_in_382),
    .col_in_383(u1_col_in_383),
    .col_in_384(u1_col_in_384),
    .col_in_385(u1_col_in_385),
    .col_in_386(u1_col_in_386),
    .col_in_387(u1_col_in_387),
    .col_in_388(u1_col_in_388),
    .col_in_389(u1_col_in_389),
    .col_in_390(u1_col_in_390),
    .col_in_391(u1_col_in_391),
    .col_in_392(u1_col_in_392),
    .col_in_393(u1_col_in_393),
    .col_in_394(u1_col_in_394),
    .col_in_395(u1_col_in_395),
    .col_in_396(u1_col_in_396),
    .col_in_397(u1_col_in_397),
    .col_in_398(u1_col_in_398),
    .col_in_399(u1_col_in_399),
    .col_in_400(u1_col_in_400),
    .col_in_401(u1_col_in_401),
    .col_in_402(u1_col_in_402),
    .col_in_403(u1_col_in_403),
    .col_in_404(u1_col_in_404),
    .col_in_405(u1_col_in_405),
    .col_in_406(u1_col_in_406),
    .col_in_407(u1_col_in_407),
    .col_in_408(u1_col_in_408),
    .col_in_409(u1_col_in_409),
    .col_in_410(u1_col_in_410),
    .col_in_411(u1_col_in_411),
    .col_in_412(u1_col_in_412),
    .col_in_413(u1_col_in_413),
    .col_in_414(u1_col_in_414),
    .col_in_415(u1_col_in_415),
    .col_in_416(u1_col_in_416),
    .col_in_417(u1_col_in_417),
    .col_in_418(u1_col_in_418),
    .col_in_419(u1_col_in_419),
    .col_in_420(u1_col_in_420),
    .col_in_421(u1_col_in_421),
    .col_in_422(u1_col_in_422),
    .col_in_423(u1_col_in_423),
    .col_in_424(u1_col_in_424),
    .col_in_425(u1_col_in_425),
    .col_in_426(u1_col_in_426),
    .col_in_427(u1_col_in_427),
    .col_in_428(u1_col_in_428),
    .col_in_429(u1_col_in_429),
    .col_in_430(u1_col_in_430),
    .col_in_431(u1_col_in_431),
    .col_in_432(u1_col_in_432),
    .col_in_433(u1_col_in_433),
    .col_in_434(u1_col_in_434),
    .col_in_435(u1_col_in_435),
    .col_in_436(u1_col_in_436),
    .col_in_437(u1_col_in_437),
    .col_in_438(u1_col_in_438),
    .col_in_439(u1_col_in_439),
    .col_in_440(u1_col_in_440),
    .col_in_441(u1_col_in_441),
    .col_in_442(u1_col_in_442),
    .col_in_443(u1_col_in_443),
    .col_in_444(u1_col_in_444),
    .col_in_445(u1_col_in_445),
    .col_in_446(u1_col_in_446),
    .col_in_447(u1_col_in_447),
    .col_in_448(u1_col_in_448),
    .col_in_449(u1_col_in_449),
    .col_in_450(u1_col_in_450),
    .col_in_451(u1_col_in_451),
    .col_in_452(u1_col_in_452),
    .col_in_453(u1_col_in_453),
    .col_in_454(u1_col_in_454),
    .col_in_455(u1_col_in_455),
    .col_in_456(u1_col_in_456),
    .col_in_457(u1_col_in_457),
    .col_in_458(u1_col_in_458),
    .col_in_459(u1_col_in_459),
    .col_in_460(u1_col_in_460),
    .col_in_461(u1_col_in_461),
    .col_in_462(u1_col_in_462),
    .col_in_463(u1_col_in_463),
    .col_in_464(u1_col_in_464),
    .col_in_465(u1_col_in_465),
    .col_in_466(u1_col_in_466),
    .col_in_467(u1_col_in_467),
    .col_in_468(u1_col_in_468),
    .col_in_469(u1_col_in_469),
    .col_in_470(u1_col_in_470),
    .col_in_471(u1_col_in_471),
    .col_in_472(u1_col_in_472),
    .col_in_473(u1_col_in_473),
    .col_in_474(u1_col_in_474),
    .col_in_475(u1_col_in_475),
    .col_in_476(u1_col_in_476),
    .col_in_477(u1_col_in_477),
    .col_in_478(u1_col_in_478),
    .col_in_479(u1_col_in_479),
    .col_in_480(u1_col_in_480),
    .col_in_481(u1_col_in_481),
    .col_in_482(u1_col_in_482),
    .col_in_483(u1_col_in_483),
    .col_in_484(u1_col_in_484),
    .col_in_485(u1_col_in_485),
    .col_in_486(u1_col_in_486),
    .col_in_487(u1_col_in_487),
    .col_in_488(u1_col_in_488),
    .col_in_489(u1_col_in_489),
    .col_in_490(u1_col_in_490),
    .col_in_491(u1_col_in_491),
    .col_in_492(u1_col_in_492),
    .col_in_493(u1_col_in_493),
    .col_in_494(u1_col_in_494),
    .col_in_495(u1_col_in_495),
    .col_in_496(u1_col_in_496),
    .col_in_497(u1_col_in_497),
    .col_in_498(u1_col_in_498),
    .col_in_499(u1_col_in_499),
    .col_in_500(u1_col_in_500),
    .col_in_501(u1_col_in_501),
    .col_in_502(u1_col_in_502),
    .col_in_503(u1_col_in_503),
    .col_in_504(u1_col_in_504),
    .col_in_505(u1_col_in_505),
    .col_in_506(u1_col_in_506),
    .col_in_507(u1_col_in_507),
    .col_in_508(u1_col_in_508),
    .col_in_509(u1_col_in_509),
    .col_in_510(u1_col_in_510),
    .col_in_511(u1_col_in_511),
    .col_in_512(u1_col_in_512),
    .col_in_513(u1_col_in_513),
    .col_in_514(u1_col_in_514),
    .col_in_515(u1_col_in_515),
    .col_in_516(u1_col_in_516),
    .col_in_517(u1_col_in_517),
    .col_in_518(u1_col_in_518),
    .col_in_519(u1_col_in_519),
    .col_in_520(u1_col_in_520),
    .col_in_521(u1_col_in_521),
    .col_in_522(u1_col_in_522),
    .col_in_523(u1_col_in_523),
    .col_in_524(u1_col_in_524),
    .col_in_525(u1_col_in_525),
    .col_in_526(u1_col_in_526),
    .col_in_527(u1_col_in_527),
    .col_in_528(u1_col_in_528),
    .col_in_529(u1_col_in_529),
    .col_in_530(u1_col_in_530),
    .col_in_531(u1_col_in_531),
    .col_in_532(u1_col_in_532),
    .col_in_533(u1_col_in_533),
    .col_in_534(u1_col_in_534),
    .col_in_535(u1_col_in_535),
    .col_in_536(u1_col_in_536),
    .col_in_537(u1_col_in_537),
    .col_in_538(u1_col_in_538),
    .col_in_539(u1_col_in_539),
    .col_in_540(u1_col_in_540),
    .col_in_541(u1_col_in_541),
    .col_in_542(u1_col_in_542),
    .col_in_543(u1_col_in_543),
    .col_in_544(u1_col_in_544),
    .col_in_545(u1_col_in_545),
    .col_in_546(u1_col_in_546),
    .col_in_547(u1_col_in_547),
    .col_in_548(u1_col_in_548),
    .col_in_549(u1_col_in_549),
    .col_in_550(u1_col_in_550),
    .col_in_551(u1_col_in_551),
    .col_in_552(u1_col_in_552),
    .col_in_553(u1_col_in_553),
    .col_in_554(u1_col_in_554),
    .col_in_555(u1_col_in_555),
    .col_in_556(u1_col_in_556),
    .col_in_557(u1_col_in_557),
    .col_in_558(u1_col_in_558),
    .col_in_559(u1_col_in_559),
    .col_in_560(u1_col_in_560),
    .col_in_561(u1_col_in_561),
    .col_in_562(u1_col_in_562),
    .col_in_563(u1_col_in_563),
    .col_in_564(u1_col_in_564),
    .col_in_565(u1_col_in_565),
    .col_in_566(u1_col_in_566),
    .col_in_567(u1_col_in_567),
    .col_in_568(u1_col_in_568),
    .col_in_569(u1_col_in_569),
    .col_in_570(u1_col_in_570),
    .col_in_571(u1_col_in_571),
    .col_in_572(u1_col_in_572),
    .col_in_573(u1_col_in_573),
    .col_in_574(u1_col_in_574),
    .col_in_575(u1_col_in_575),
    .col_in_576(u1_col_in_576),
    .col_in_577(u1_col_in_577),
    .col_in_578(u1_col_in_578),
    .col_in_579(u1_col_in_579),
    .col_in_580(u1_col_in_580),
    .col_in_581(u1_col_in_581),
    .col_in_582(u1_col_in_582),
    .col_in_583(u1_col_in_583),
    .col_in_584(u1_col_in_584),
    .col_in_585(u1_col_in_585),
    .col_in_586(u1_col_in_586),
    .col_in_587(u1_col_in_587),
    .col_in_588(u1_col_in_588),
    .col_in_589(u1_col_in_589),
    .col_in_590(u1_col_in_590),
    .col_in_591(u1_col_in_591),
    .col_in_592(u1_col_in_592),
    .col_in_593(u1_col_in_593),
    .col_in_594(u1_col_in_594),
    .col_in_595(u1_col_in_595),
    .col_in_596(u1_col_in_596),
    .col_in_597(u1_col_in_597),
    .col_in_598(u1_col_in_598),
    .col_in_599(u1_col_in_599),
    .col_in_600(u1_col_in_600),
    .col_in_601(u1_col_in_601),
    .col_in_602(u1_col_in_602),
    .col_in_603(u1_col_in_603),
    .col_in_604(u1_col_in_604),
    .col_in_605(u1_col_in_605),
    .col_in_606(u1_col_in_606),
    .col_in_607(u1_col_in_607),
    .col_in_608(u1_col_in_608),
    .col_in_609(u1_col_in_609),
    .col_in_610(u1_col_in_610),
    .col_in_611(u1_col_in_611),
    .col_in_612(u1_col_in_612),
    .col_in_613(u1_col_in_613),
    .col_in_614(u1_col_in_614),
    .col_in_615(u1_col_in_615),
    .col_in_616(u1_col_in_616),
    .col_in_617(u1_col_in_617),
    .col_in_618(u1_col_in_618),
    .col_in_619(u1_col_in_619),
    .col_in_620(u1_col_in_620),
    .col_in_621(u1_col_in_621),
    .col_in_622(u1_col_in_622),
    .col_in_623(u1_col_in_623),
    .col_in_624(u1_col_in_624),
    .col_in_625(u1_col_in_625),
    .col_in_626(u1_col_in_626),
    .col_in_627(u1_col_in_627),
    .col_in_628(u1_col_in_628),
    .col_in_629(u1_col_in_629),
    .col_in_630(u1_col_in_630),
    .col_in_631(u1_col_in_631),
    .col_in_632(u1_col_in_632),
    .col_in_633(u1_col_in_633),
    .col_in_634(u1_col_in_634),
    .col_in_635(u1_col_in_635),
    .col_in_636(u1_col_in_636),
    .col_in_637(u1_col_in_637),
    .col_in_638(u1_col_in_638),
    .col_in_639(u1_col_in_639),
    .col_in_640(u1_col_in_640),
    .col_in_641(u1_col_in_641),
    .col_in_642(u1_col_in_642),
    .col_in_643(u1_col_in_643),
    .col_in_644(u1_col_in_644),
    .col_in_645(u1_col_in_645),
    .col_in_646(u1_col_in_646),
    .col_in_647(u1_col_in_647),
    .col_in_648(u1_col_in_648),
    .col_in_649(u1_col_in_649),
    .col_in_650(u1_col_in_650),
    .col_in_651(u1_col_in_651),
    .col_in_652(u1_col_in_652),
    .col_in_653(u1_col_in_653),
    .col_in_654(u1_col_in_654),
    .col_in_655(u1_col_in_655),
    .col_in_656(u1_col_in_656),
    .col_in_657(u1_col_in_657),
    .col_in_658(u1_col_in_658),
    .col_in_659(u1_col_in_659),
    .col_in_660(u1_col_in_660),
    .col_in_661(u1_col_in_661),
    .col_in_662(u1_col_in_662),
    .col_in_663(u1_col_in_663),
    .col_in_664(u1_col_in_664),
    .col_in_665(u1_col_in_665),
    .col_in_666(u1_col_in_666),
    .col_in_667(u1_col_in_667),
    .col_in_668(u1_col_in_668),
    .col_in_669(u1_col_in_669),
    .col_in_670(u1_col_in_670),
    .col_in_671(u1_col_in_671),
    .col_in_672(u1_col_in_672),
    .col_in_673(u1_col_in_673),
    .col_in_674(u1_col_in_674),
    .col_in_675(u1_col_in_675),
    .col_in_676(u1_col_in_676),
    .col_in_677(u1_col_in_677),
    .col_in_678(u1_col_in_678),
    .col_in_679(u1_col_in_679),
    .col_in_680(u1_col_in_680),
    .col_in_681(u1_col_in_681),
    .col_in_682(u1_col_in_682),
    .col_in_683(u1_col_in_683),
    .col_in_684(u1_col_in_684),
    .col_in_685(u1_col_in_685),
    .col_in_686(u1_col_in_686),
    .col_in_687(u1_col_in_687),
    .col_in_688(u1_col_in_688),
    .col_in_689(u1_col_in_689),
    .col_in_690(u1_col_in_690),
    .col_in_691(u1_col_in_691),
    .col_in_692(u1_col_in_692),
    .col_in_693(u1_col_in_693),
    .col_in_694(u1_col_in_694),
    .col_in_695(u1_col_in_695),
    .col_in_696(u1_col_in_696),
    .col_in_697(u1_col_in_697),
    .col_in_698(u1_col_in_698),
    .col_in_699(u1_col_in_699),
    .col_in_700(u1_col_in_700),
    .col_in_701(u1_col_in_701),
    .col_in_702(u1_col_in_702),
    .col_in_703(u1_col_in_703),
    .col_in_704(u1_col_in_704),
    .col_in_705(u1_col_in_705),
    .col_in_706(u1_col_in_706),
    .col_in_707(u1_col_in_707),
    .col_in_708(u1_col_in_708),
    .col_in_709(u1_col_in_709),
    .col_in_710(u1_col_in_710),
    .col_in_711(u1_col_in_711),
    .col_in_712(u1_col_in_712),
    .col_in_713(u1_col_in_713),
    .col_in_714(u1_col_in_714),
    .col_in_715(u1_col_in_715),
    .col_in_716(u1_col_in_716),
    .col_in_717(u1_col_in_717),
    .col_in_718(u1_col_in_718),
    .col_in_719(u1_col_in_719),
    .col_in_720(u1_col_in_720),
    .col_in_721(u1_col_in_721),
    .col_in_722(u1_col_in_722),
    .col_in_723(u1_col_in_723),
    .col_in_724(u1_col_in_724),
    .col_in_725(u1_col_in_725),
    .col_in_726(u1_col_in_726),
    .col_in_727(u1_col_in_727),
    .col_in_728(u1_col_in_728),
    .col_in_729(u1_col_in_729),
    .col_in_730(u1_col_in_730),
    .col_in_731(u1_col_in_731),
    .col_in_732(u1_col_in_732),
    .col_in_733(u1_col_in_733),
    .col_in_734(u1_col_in_734),
    .col_in_735(u1_col_in_735),
    .col_in_736(u1_col_in_736),
    .col_in_737(u1_col_in_737),
    .col_in_738(u1_col_in_738),
    .col_in_739(u1_col_in_739),
    .col_in_740(u1_col_in_740),
    .col_in_741(u1_col_in_741),
    .col_in_742(u1_col_in_742),
    .col_in_743(u1_col_in_743),
    .col_in_744(u1_col_in_744),
    .col_in_745(u1_col_in_745),
    .col_in_746(u1_col_in_746),
    .col_in_747(u1_col_in_747),
    .col_in_748(u1_col_in_748),
    .col_in_749(u1_col_in_749),
    .col_in_750(u1_col_in_750),
    .col_in_751(u1_col_in_751),
    .col_in_752(u1_col_in_752),
    .col_in_753(u1_col_in_753),
    .col_in_754(u1_col_in_754),
    .col_in_755(u1_col_in_755),
    .col_in_756(u1_col_in_756),
    .col_in_757(u1_col_in_757),
    .col_in_758(u1_col_in_758),
    .col_in_759(u1_col_in_759),
    .col_in_760(u1_col_in_760),
    .col_in_761(u1_col_in_761),
    .col_in_762(u1_col_in_762),
    .col_in_763(u1_col_in_763),
    .col_in_764(u1_col_in_764),
    .col_in_765(u1_col_in_765),
    .col_in_766(u1_col_in_766),
    .col_in_767(u1_col_in_767),
    .col_in_768(u1_col_in_768),
    .col_in_769(u1_col_in_769),
    .col_in_770(u1_col_in_770),
    .col_in_771(u1_col_in_771),
    .col_in_772(u1_col_in_772),
    .col_in_773(u1_col_in_773),
    .col_in_774(u1_col_in_774),
    .col_in_775(u1_col_in_775),
    .col_in_776(u1_col_in_776),
    .col_in_777(u1_col_in_777),
    .col_in_778(u1_col_in_778),
    .col_in_779(u1_col_in_779),
    .col_in_780(u1_col_in_780),
    .col_in_781(u1_col_in_781),
    .col_in_782(u1_col_in_782),
    .col_in_783(u1_col_in_783),
    .col_in_784(u1_col_in_784),
    .col_in_785(u1_col_in_785),
    .col_in_786(u1_col_in_786),
    .col_in_787(u1_col_in_787),
    .col_in_788(u1_col_in_788),
    .col_in_789(u1_col_in_789),
    .col_in_790(u1_col_in_790),
    .col_in_791(u1_col_in_791),
    .col_in_792(u1_col_in_792),
    .col_in_793(u1_col_in_793),
    .col_in_794(u1_col_in_794),
    .col_in_795(u1_col_in_795),
    .col_in_796(u1_col_in_796),
    .col_in_797(u1_col_in_797),
    .col_in_798(u1_col_in_798),
    .col_in_799(u1_col_in_799),
    .col_in_800(u1_col_in_800),
    .col_in_801(u1_col_in_801),
    .col_in_802(u1_col_in_802),
    .col_in_803(u1_col_in_803),
    .col_in_804(u1_col_in_804),
    .col_in_805(u1_col_in_805),
    .col_in_806(u1_col_in_806),
    .col_in_807(u1_col_in_807),
    .col_in_808(u1_col_in_808),
    .col_in_809(u1_col_in_809),
    .col_in_810(u1_col_in_810),
    .col_in_811(u1_col_in_811),
    .col_in_812(u1_col_in_812),
    .col_in_813(u1_col_in_813),
    .col_in_814(u1_col_in_814),
    .col_in_815(u1_col_in_815),
    .col_in_816(u1_col_in_816),
    .col_in_817(u1_col_in_817),
    .col_in_818(u1_col_in_818),
    .col_in_819(u1_col_in_819),
    .col_in_820(u1_col_in_820),
    .col_in_821(u1_col_in_821),
    .col_in_822(u1_col_in_822),
    .col_in_823(u1_col_in_823),
    .col_in_824(u1_col_in_824),
    .col_in_825(u1_col_in_825),
    .col_in_826(u1_col_in_826),
    .col_in_827(u1_col_in_827),
    .col_in_828(u1_col_in_828),
    .col_in_829(u1_col_in_829),
    .col_in_830(u1_col_in_830),
    .col_in_831(u1_col_in_831),
    .col_in_832(u1_col_in_832),
    .col_in_833(u1_col_in_833),
    .col_in_834(u1_col_in_834),
    .col_in_835(u1_col_in_835),
    .col_in_836(u1_col_in_836),
    .col_in_837(u1_col_in_837),
    .col_in_838(u1_col_in_838),
    .col_in_839(u1_col_in_839),
    .col_in_840(u1_col_in_840),
    .col_in_841(u1_col_in_841),
    .col_in_842(u1_col_in_842),
    .col_in_843(u1_col_in_843),
    .col_in_844(u1_col_in_844),
    .col_in_845(u1_col_in_845),
    .col_in_846(u1_col_in_846),
    .col_in_847(u1_col_in_847),
    .col_in_848(u1_col_in_848),
    .col_in_849(u1_col_in_849),
    .col_in_850(u1_col_in_850),
    .col_in_851(u1_col_in_851),
    .col_in_852(u1_col_in_852),
    .col_in_853(u1_col_in_853),
    .col_in_854(u1_col_in_854),
    .col_in_855(u1_col_in_855),
    .col_in_856(u1_col_in_856),
    .col_in_857(u1_col_in_857),
    .col_in_858(u1_col_in_858),
    .col_in_859(u1_col_in_859),
    .col_in_860(u1_col_in_860),
    .col_in_861(u1_col_in_861),
    .col_in_862(u1_col_in_862),
    .col_in_863(u1_col_in_863),
    .col_in_864(u1_col_in_864),
    .col_in_865(u1_col_in_865),
    .col_in_866(u1_col_in_866),
    .col_in_867(u1_col_in_867),
    .col_in_868(u1_col_in_868),
    .col_in_869(u1_col_in_869),
    .col_in_870(u1_col_in_870),
    .col_in_871(u1_col_in_871),
    .col_in_872(u1_col_in_872),
    .col_in_873(u1_col_in_873),
    .col_in_874(u1_col_in_874),
    .col_in_875(u1_col_in_875),
    .col_in_876(u1_col_in_876),
    .col_in_877(u1_col_in_877),
    .col_in_878(u1_col_in_878),
    .col_in_879(u1_col_in_879),
    .col_in_880(u1_col_in_880),
    .col_in_881(u1_col_in_881),
    .col_in_882(u1_col_in_882),
    .col_in_883(u1_col_in_883),
    .col_in_884(u1_col_in_884),
    .col_in_885(u1_col_in_885),
    .col_in_886(u1_col_in_886),
    .col_in_887(u1_col_in_887),
    .col_in_888(u1_col_in_888),
    .col_in_889(u1_col_in_889),
    .col_in_890(u1_col_in_890),
    .col_in_891(u1_col_in_891),
    .col_in_892(u1_col_in_892),
    .col_in_893(u1_col_in_893),
    .col_in_894(u1_col_in_894),
    .col_in_895(u1_col_in_895),
    .col_in_896(u1_col_in_896),
    .col_in_897(u1_col_in_897),
    .col_in_898(u1_col_in_898),
    .col_in_899(u1_col_in_899),
    .col_in_900(u1_col_in_900),
    .col_in_901(u1_col_in_901),
    .col_in_902(u1_col_in_902),
    .col_in_903(u1_col_in_903),
    .col_in_904(u1_col_in_904),
    .col_in_905(u1_col_in_905),
    .col_in_906(u1_col_in_906),
    .col_in_907(u1_col_in_907),
    .col_in_908(u1_col_in_908),
    .col_in_909(u1_col_in_909),
    .col_in_910(u1_col_in_910),
    .col_in_911(u1_col_in_911),
    .col_in_912(u1_col_in_912),
    .col_in_913(u1_col_in_913),
    .col_in_914(u1_col_in_914),
    .col_in_915(u1_col_in_915),
    .col_in_916(u1_col_in_916),
    .col_in_917(u1_col_in_917),
    .col_in_918(u1_col_in_918),
    .col_in_919(u1_col_in_919),
    .col_in_920(u1_col_in_920),
    .col_in_921(u1_col_in_921),
    .col_in_922(u1_col_in_922),
    .col_in_923(u1_col_in_923),
    .col_in_924(u1_col_in_924),
    .col_in_925(u1_col_in_925),
    .col_in_926(u1_col_in_926),
    .col_in_927(u1_col_in_927),
    .col_in_928(u1_col_in_928),
    .col_in_929(u1_col_in_929),
    .col_in_930(u1_col_in_930),
    .col_in_931(u1_col_in_931),
    .col_in_932(u1_col_in_932),
    .col_in_933(u1_col_in_933),
    .col_in_934(u1_col_in_934),
    .col_in_935(u1_col_in_935),
    .col_in_936(u1_col_in_936),
    .col_in_937(u1_col_in_937),
    .col_in_938(u1_col_in_938),
    .col_in_939(u1_col_in_939),
    .col_in_940(u1_col_in_940),
    .col_in_941(u1_col_in_941),
    .col_in_942(u1_col_in_942),
    .col_in_943(u1_col_in_943),
    .col_in_944(u1_col_in_944),
    .col_in_945(u1_col_in_945),
    .col_in_946(u1_col_in_946),
    .col_in_947(u1_col_in_947),
    .col_in_948(u1_col_in_948),
    .col_in_949(u1_col_in_949),
    .col_in_950(u1_col_in_950),
    .col_in_951(u1_col_in_951),
    .col_in_952(u1_col_in_952),
    .col_in_953(u1_col_in_953),
    .col_in_954(u1_col_in_954),
    .col_in_955(u1_col_in_955),
    .col_in_956(u1_col_in_956),
    .col_in_957(u1_col_in_957),
    .col_in_958(u1_col_in_958),
    .col_in_959(u1_col_in_959),
    .col_in_960(u1_col_in_960),
    .col_in_961(u1_col_in_961),
    .col_in_962(u1_col_in_962),
    .col_in_963(u1_col_in_963),
    .col_in_964(u1_col_in_964),
    .col_in_965(u1_col_in_965),
    .col_in_966(u1_col_in_966),
    .col_in_967(u1_col_in_967),
    .col_in_968(u1_col_in_968),
    .col_in_969(u1_col_in_969),
    .col_in_970(u1_col_in_970),
    .col_in_971(u1_col_in_971),
    .col_in_972(u1_col_in_972),
    .col_in_973(u1_col_in_973),
    .col_in_974(u1_col_in_974),
    .col_in_975(u1_col_in_975),
    .col_in_976(u1_col_in_976),
    .col_in_977(u1_col_in_977),
    .col_in_978(u1_col_in_978),
    .col_in_979(u1_col_in_979),
    .col_in_980(u1_col_in_980),
    .col_in_981(u1_col_in_981),
    .col_in_982(u1_col_in_982),
    .col_in_983(u1_col_in_983),
    .col_in_984(u1_col_in_984),
    .col_in_985(u1_col_in_985),
    .col_in_986(u1_col_in_986),
    .col_in_987(u1_col_in_987),
    .col_in_988(u1_col_in_988),
    .col_in_989(u1_col_in_989),
    .col_in_990(u1_col_in_990),
    .col_in_991(u1_col_in_991),
    .col_in_992(u1_col_in_992),
    .col_in_993(u1_col_in_993),
    .col_in_994(u1_col_in_994),
    .col_in_995(u1_col_in_995),
    .col_in_996(u1_col_in_996),
    .col_in_997(u1_col_in_997),
    .col_in_998(u1_col_in_998),
    .col_in_999(u1_col_in_999),
    .col_in_1000(u1_col_in_1000),
    .col_in_1001(u1_col_in_1001),
    .col_in_1002(u1_col_in_1002),
    .col_in_1003(u1_col_in_1003),
    .col_in_1004(u1_col_in_1004),
    .col_in_1005(u1_col_in_1005),
    .col_in_1006(u1_col_in_1006),
    .col_in_1007(u1_col_in_1007),
    .col_in_1008(u1_col_in_1008),
    .col_in_1009(u1_col_in_1009),
    .col_in_1010(u1_col_in_1010),
    .col_in_1011(u1_col_in_1011),
    .col_in_1012(u1_col_in_1012),
    .col_in_1013(u1_col_in_1013),
    .col_in_1014(u1_col_in_1014),
    .col_in_1015(u1_col_in_1015),
    .col_in_1016(u1_col_in_1016),
    .col_in_1017(u1_col_in_1017),
    .col_in_1018(u1_col_in_1018),
    .col_in_1019(u1_col_in_1019),
    .col_in_1020(u1_col_in_1020),
    .col_in_1021(u1_col_in_1021),
    .col_in_1022(u1_col_in_1022),
    .col_in_1023(u1_col_in_1023),
    .col_in_1024(u1_col_in_1024),
    .col_in_1025(u1_col_in_1025),
    .col_in_1026(u1_col_in_1026),

    .col_out_0(u1_col_out_0),
    .col_out_1(u1_col_out_1),
    .col_out_2(u1_col_out_2),
    .col_out_3(u1_col_out_3),
    .col_out_4(u1_col_out_4),
    .col_out_5(u1_col_out_5),
    .col_out_6(u1_col_out_6),
    .col_out_7(u1_col_out_7),
    .col_out_8(u1_col_out_8),
    .col_out_9(u1_col_out_9),
    .col_out_10(u1_col_out_10),
    .col_out_11(u1_col_out_11),
    .col_out_12(u1_col_out_12),
    .col_out_13(u1_col_out_13),
    .col_out_14(u1_col_out_14),
    .col_out_15(u1_col_out_15),
    .col_out_16(u1_col_out_16),
    .col_out_17(u1_col_out_17),
    .col_out_18(u1_col_out_18),
    .col_out_19(u1_col_out_19),
    .col_out_20(u1_col_out_20),
    .col_out_21(u1_col_out_21),
    .col_out_22(u1_col_out_22),
    .col_out_23(u1_col_out_23),
    .col_out_24(u1_col_out_24),
    .col_out_25(u1_col_out_25),
    .col_out_26(u1_col_out_26),
    .col_out_27(u1_col_out_27),
    .col_out_28(u1_col_out_28),
    .col_out_29(u1_col_out_29),
    .col_out_30(u1_col_out_30),
    .col_out_31(u1_col_out_31),
    .col_out_32(u1_col_out_32),
    .col_out_33(u1_col_out_33),
    .col_out_34(u1_col_out_34),
    .col_out_35(u1_col_out_35),
    .col_out_36(u1_col_out_36),
    .col_out_37(u1_col_out_37),
    .col_out_38(u1_col_out_38),
    .col_out_39(u1_col_out_39),
    .col_out_40(u1_col_out_40),
    .col_out_41(u1_col_out_41),
    .col_out_42(u1_col_out_42),
    .col_out_43(u1_col_out_43),
    .col_out_44(u1_col_out_44),
    .col_out_45(u1_col_out_45),
    .col_out_46(u1_col_out_46),
    .col_out_47(u1_col_out_47),
    .col_out_48(u1_col_out_48),
    .col_out_49(u1_col_out_49),
    .col_out_50(u1_col_out_50),
    .col_out_51(u1_col_out_51),
    .col_out_52(u1_col_out_52),
    .col_out_53(u1_col_out_53),
    .col_out_54(u1_col_out_54),
    .col_out_55(u1_col_out_55),
    .col_out_56(u1_col_out_56),
    .col_out_57(u1_col_out_57),
    .col_out_58(u1_col_out_58),
    .col_out_59(u1_col_out_59),
    .col_out_60(u1_col_out_60),
    .col_out_61(u1_col_out_61),
    .col_out_62(u1_col_out_62),
    .col_out_63(u1_col_out_63),
    .col_out_64(u1_col_out_64),
    .col_out_65(u1_col_out_65),
    .col_out_66(u1_col_out_66),
    .col_out_67(u1_col_out_67),
    .col_out_68(u1_col_out_68),
    .col_out_69(u1_col_out_69),
    .col_out_70(u1_col_out_70),
    .col_out_71(u1_col_out_71),
    .col_out_72(u1_col_out_72),
    .col_out_73(u1_col_out_73),
    .col_out_74(u1_col_out_74),
    .col_out_75(u1_col_out_75),
    .col_out_76(u1_col_out_76),
    .col_out_77(u1_col_out_77),
    .col_out_78(u1_col_out_78),
    .col_out_79(u1_col_out_79),
    .col_out_80(u1_col_out_80),
    .col_out_81(u1_col_out_81),
    .col_out_82(u1_col_out_82),
    .col_out_83(u1_col_out_83),
    .col_out_84(u1_col_out_84),
    .col_out_85(u1_col_out_85),
    .col_out_86(u1_col_out_86),
    .col_out_87(u1_col_out_87),
    .col_out_88(u1_col_out_88),
    .col_out_89(u1_col_out_89),
    .col_out_90(u1_col_out_90),
    .col_out_91(u1_col_out_91),
    .col_out_92(u1_col_out_92),
    .col_out_93(u1_col_out_93),
    .col_out_94(u1_col_out_94),
    .col_out_95(u1_col_out_95),
    .col_out_96(u1_col_out_96),
    .col_out_97(u1_col_out_97),
    .col_out_98(u1_col_out_98),
    .col_out_99(u1_col_out_99),
    .col_out_100(u1_col_out_100),
    .col_out_101(u1_col_out_101),
    .col_out_102(u1_col_out_102),
    .col_out_103(u1_col_out_103),
    .col_out_104(u1_col_out_104),
    .col_out_105(u1_col_out_105),
    .col_out_106(u1_col_out_106),
    .col_out_107(u1_col_out_107),
    .col_out_108(u1_col_out_108),
    .col_out_109(u1_col_out_109),
    .col_out_110(u1_col_out_110),
    .col_out_111(u1_col_out_111),
    .col_out_112(u1_col_out_112),
    .col_out_113(u1_col_out_113),
    .col_out_114(u1_col_out_114),
    .col_out_115(u1_col_out_115),
    .col_out_116(u1_col_out_116),
    .col_out_117(u1_col_out_117),
    .col_out_118(u1_col_out_118),
    .col_out_119(u1_col_out_119),
    .col_out_120(u1_col_out_120),
    .col_out_121(u1_col_out_121),
    .col_out_122(u1_col_out_122),
    .col_out_123(u1_col_out_123),
    .col_out_124(u1_col_out_124),
    .col_out_125(u1_col_out_125),
    .col_out_126(u1_col_out_126),
    .col_out_127(u1_col_out_127),
    .col_out_128(u1_col_out_128),
    .col_out_129(u1_col_out_129),
    .col_out_130(u1_col_out_130),
    .col_out_131(u1_col_out_131),
    .col_out_132(u1_col_out_132),
    .col_out_133(u1_col_out_133),
    .col_out_134(u1_col_out_134),
    .col_out_135(u1_col_out_135),
    .col_out_136(u1_col_out_136),
    .col_out_137(u1_col_out_137),
    .col_out_138(u1_col_out_138),
    .col_out_139(u1_col_out_139),
    .col_out_140(u1_col_out_140),
    .col_out_141(u1_col_out_141),
    .col_out_142(u1_col_out_142),
    .col_out_143(u1_col_out_143),
    .col_out_144(u1_col_out_144),
    .col_out_145(u1_col_out_145),
    .col_out_146(u1_col_out_146),
    .col_out_147(u1_col_out_147),
    .col_out_148(u1_col_out_148),
    .col_out_149(u1_col_out_149),
    .col_out_150(u1_col_out_150),
    .col_out_151(u1_col_out_151),
    .col_out_152(u1_col_out_152),
    .col_out_153(u1_col_out_153),
    .col_out_154(u1_col_out_154),
    .col_out_155(u1_col_out_155),
    .col_out_156(u1_col_out_156),
    .col_out_157(u1_col_out_157),
    .col_out_158(u1_col_out_158),
    .col_out_159(u1_col_out_159),
    .col_out_160(u1_col_out_160),
    .col_out_161(u1_col_out_161),
    .col_out_162(u1_col_out_162),
    .col_out_163(u1_col_out_163),
    .col_out_164(u1_col_out_164),
    .col_out_165(u1_col_out_165),
    .col_out_166(u1_col_out_166),
    .col_out_167(u1_col_out_167),
    .col_out_168(u1_col_out_168),
    .col_out_169(u1_col_out_169),
    .col_out_170(u1_col_out_170),
    .col_out_171(u1_col_out_171),
    .col_out_172(u1_col_out_172),
    .col_out_173(u1_col_out_173),
    .col_out_174(u1_col_out_174),
    .col_out_175(u1_col_out_175),
    .col_out_176(u1_col_out_176),
    .col_out_177(u1_col_out_177),
    .col_out_178(u1_col_out_178),
    .col_out_179(u1_col_out_179),
    .col_out_180(u1_col_out_180),
    .col_out_181(u1_col_out_181),
    .col_out_182(u1_col_out_182),
    .col_out_183(u1_col_out_183),
    .col_out_184(u1_col_out_184),
    .col_out_185(u1_col_out_185),
    .col_out_186(u1_col_out_186),
    .col_out_187(u1_col_out_187),
    .col_out_188(u1_col_out_188),
    .col_out_189(u1_col_out_189),
    .col_out_190(u1_col_out_190),
    .col_out_191(u1_col_out_191),
    .col_out_192(u1_col_out_192),
    .col_out_193(u1_col_out_193),
    .col_out_194(u1_col_out_194),
    .col_out_195(u1_col_out_195),
    .col_out_196(u1_col_out_196),
    .col_out_197(u1_col_out_197),
    .col_out_198(u1_col_out_198),
    .col_out_199(u1_col_out_199),
    .col_out_200(u1_col_out_200),
    .col_out_201(u1_col_out_201),
    .col_out_202(u1_col_out_202),
    .col_out_203(u1_col_out_203),
    .col_out_204(u1_col_out_204),
    .col_out_205(u1_col_out_205),
    .col_out_206(u1_col_out_206),
    .col_out_207(u1_col_out_207),
    .col_out_208(u1_col_out_208),
    .col_out_209(u1_col_out_209),
    .col_out_210(u1_col_out_210),
    .col_out_211(u1_col_out_211),
    .col_out_212(u1_col_out_212),
    .col_out_213(u1_col_out_213),
    .col_out_214(u1_col_out_214),
    .col_out_215(u1_col_out_215),
    .col_out_216(u1_col_out_216),
    .col_out_217(u1_col_out_217),
    .col_out_218(u1_col_out_218),
    .col_out_219(u1_col_out_219),
    .col_out_220(u1_col_out_220),
    .col_out_221(u1_col_out_221),
    .col_out_222(u1_col_out_222),
    .col_out_223(u1_col_out_223),
    .col_out_224(u1_col_out_224),
    .col_out_225(u1_col_out_225),
    .col_out_226(u1_col_out_226),
    .col_out_227(u1_col_out_227),
    .col_out_228(u1_col_out_228),
    .col_out_229(u1_col_out_229),
    .col_out_230(u1_col_out_230),
    .col_out_231(u1_col_out_231),
    .col_out_232(u1_col_out_232),
    .col_out_233(u1_col_out_233),
    .col_out_234(u1_col_out_234),
    .col_out_235(u1_col_out_235),
    .col_out_236(u1_col_out_236),
    .col_out_237(u1_col_out_237),
    .col_out_238(u1_col_out_238),
    .col_out_239(u1_col_out_239),
    .col_out_240(u1_col_out_240),
    .col_out_241(u1_col_out_241),
    .col_out_242(u1_col_out_242),
    .col_out_243(u1_col_out_243),
    .col_out_244(u1_col_out_244),
    .col_out_245(u1_col_out_245),
    .col_out_246(u1_col_out_246),
    .col_out_247(u1_col_out_247),
    .col_out_248(u1_col_out_248),
    .col_out_249(u1_col_out_249),
    .col_out_250(u1_col_out_250),
    .col_out_251(u1_col_out_251),
    .col_out_252(u1_col_out_252),
    .col_out_253(u1_col_out_253),
    .col_out_254(u1_col_out_254),
    .col_out_255(u1_col_out_255),
    .col_out_256(u1_col_out_256),
    .col_out_257(u1_col_out_257),
    .col_out_258(u1_col_out_258),
    .col_out_259(u1_col_out_259),
    .col_out_260(u1_col_out_260),
    .col_out_261(u1_col_out_261),
    .col_out_262(u1_col_out_262),
    .col_out_263(u1_col_out_263),
    .col_out_264(u1_col_out_264),
    .col_out_265(u1_col_out_265),
    .col_out_266(u1_col_out_266),
    .col_out_267(u1_col_out_267),
    .col_out_268(u1_col_out_268),
    .col_out_269(u1_col_out_269),
    .col_out_270(u1_col_out_270),
    .col_out_271(u1_col_out_271),
    .col_out_272(u1_col_out_272),
    .col_out_273(u1_col_out_273),
    .col_out_274(u1_col_out_274),
    .col_out_275(u1_col_out_275),
    .col_out_276(u1_col_out_276),
    .col_out_277(u1_col_out_277),
    .col_out_278(u1_col_out_278),
    .col_out_279(u1_col_out_279),
    .col_out_280(u1_col_out_280),
    .col_out_281(u1_col_out_281),
    .col_out_282(u1_col_out_282),
    .col_out_283(u1_col_out_283),
    .col_out_284(u1_col_out_284),
    .col_out_285(u1_col_out_285),
    .col_out_286(u1_col_out_286),
    .col_out_287(u1_col_out_287),
    .col_out_288(u1_col_out_288),
    .col_out_289(u1_col_out_289),
    .col_out_290(u1_col_out_290),
    .col_out_291(u1_col_out_291),
    .col_out_292(u1_col_out_292),
    .col_out_293(u1_col_out_293),
    .col_out_294(u1_col_out_294),
    .col_out_295(u1_col_out_295),
    .col_out_296(u1_col_out_296),
    .col_out_297(u1_col_out_297),
    .col_out_298(u1_col_out_298),
    .col_out_299(u1_col_out_299),
    .col_out_300(u1_col_out_300),
    .col_out_301(u1_col_out_301),
    .col_out_302(u1_col_out_302),
    .col_out_303(u1_col_out_303),
    .col_out_304(u1_col_out_304),
    .col_out_305(u1_col_out_305),
    .col_out_306(u1_col_out_306),
    .col_out_307(u1_col_out_307),
    .col_out_308(u1_col_out_308),
    .col_out_309(u1_col_out_309),
    .col_out_310(u1_col_out_310),
    .col_out_311(u1_col_out_311),
    .col_out_312(u1_col_out_312),
    .col_out_313(u1_col_out_313),
    .col_out_314(u1_col_out_314),
    .col_out_315(u1_col_out_315),
    .col_out_316(u1_col_out_316),
    .col_out_317(u1_col_out_317),
    .col_out_318(u1_col_out_318),
    .col_out_319(u1_col_out_319),
    .col_out_320(u1_col_out_320),
    .col_out_321(u1_col_out_321),
    .col_out_322(u1_col_out_322),
    .col_out_323(u1_col_out_323),
    .col_out_324(u1_col_out_324),
    .col_out_325(u1_col_out_325),
    .col_out_326(u1_col_out_326),
    .col_out_327(u1_col_out_327),
    .col_out_328(u1_col_out_328),
    .col_out_329(u1_col_out_329),
    .col_out_330(u1_col_out_330),
    .col_out_331(u1_col_out_331),
    .col_out_332(u1_col_out_332),
    .col_out_333(u1_col_out_333),
    .col_out_334(u1_col_out_334),
    .col_out_335(u1_col_out_335),
    .col_out_336(u1_col_out_336),
    .col_out_337(u1_col_out_337),
    .col_out_338(u1_col_out_338),
    .col_out_339(u1_col_out_339),
    .col_out_340(u1_col_out_340),
    .col_out_341(u1_col_out_341),
    .col_out_342(u1_col_out_342),
    .col_out_343(u1_col_out_343),
    .col_out_344(u1_col_out_344),
    .col_out_345(u1_col_out_345),
    .col_out_346(u1_col_out_346),
    .col_out_347(u1_col_out_347),
    .col_out_348(u1_col_out_348),
    .col_out_349(u1_col_out_349),
    .col_out_350(u1_col_out_350),
    .col_out_351(u1_col_out_351),
    .col_out_352(u1_col_out_352),
    .col_out_353(u1_col_out_353),
    .col_out_354(u1_col_out_354),
    .col_out_355(u1_col_out_355),
    .col_out_356(u1_col_out_356),
    .col_out_357(u1_col_out_357),
    .col_out_358(u1_col_out_358),
    .col_out_359(u1_col_out_359),
    .col_out_360(u1_col_out_360),
    .col_out_361(u1_col_out_361),
    .col_out_362(u1_col_out_362),
    .col_out_363(u1_col_out_363),
    .col_out_364(u1_col_out_364),
    .col_out_365(u1_col_out_365),
    .col_out_366(u1_col_out_366),
    .col_out_367(u1_col_out_367),
    .col_out_368(u1_col_out_368),
    .col_out_369(u1_col_out_369),
    .col_out_370(u1_col_out_370),
    .col_out_371(u1_col_out_371),
    .col_out_372(u1_col_out_372),
    .col_out_373(u1_col_out_373),
    .col_out_374(u1_col_out_374),
    .col_out_375(u1_col_out_375),
    .col_out_376(u1_col_out_376),
    .col_out_377(u1_col_out_377),
    .col_out_378(u1_col_out_378),
    .col_out_379(u1_col_out_379),
    .col_out_380(u1_col_out_380),
    .col_out_381(u1_col_out_381),
    .col_out_382(u1_col_out_382),
    .col_out_383(u1_col_out_383),
    .col_out_384(u1_col_out_384),
    .col_out_385(u1_col_out_385),
    .col_out_386(u1_col_out_386),
    .col_out_387(u1_col_out_387),
    .col_out_388(u1_col_out_388),
    .col_out_389(u1_col_out_389),
    .col_out_390(u1_col_out_390),
    .col_out_391(u1_col_out_391),
    .col_out_392(u1_col_out_392),
    .col_out_393(u1_col_out_393),
    .col_out_394(u1_col_out_394),
    .col_out_395(u1_col_out_395),
    .col_out_396(u1_col_out_396),
    .col_out_397(u1_col_out_397),
    .col_out_398(u1_col_out_398),
    .col_out_399(u1_col_out_399),
    .col_out_400(u1_col_out_400),
    .col_out_401(u1_col_out_401),
    .col_out_402(u1_col_out_402),
    .col_out_403(u1_col_out_403),
    .col_out_404(u1_col_out_404),
    .col_out_405(u1_col_out_405),
    .col_out_406(u1_col_out_406),
    .col_out_407(u1_col_out_407),
    .col_out_408(u1_col_out_408),
    .col_out_409(u1_col_out_409),
    .col_out_410(u1_col_out_410),
    .col_out_411(u1_col_out_411),
    .col_out_412(u1_col_out_412),
    .col_out_413(u1_col_out_413),
    .col_out_414(u1_col_out_414),
    .col_out_415(u1_col_out_415),
    .col_out_416(u1_col_out_416),
    .col_out_417(u1_col_out_417),
    .col_out_418(u1_col_out_418),
    .col_out_419(u1_col_out_419),
    .col_out_420(u1_col_out_420),
    .col_out_421(u1_col_out_421),
    .col_out_422(u1_col_out_422),
    .col_out_423(u1_col_out_423),
    .col_out_424(u1_col_out_424),
    .col_out_425(u1_col_out_425),
    .col_out_426(u1_col_out_426),
    .col_out_427(u1_col_out_427),
    .col_out_428(u1_col_out_428),
    .col_out_429(u1_col_out_429),
    .col_out_430(u1_col_out_430),
    .col_out_431(u1_col_out_431),
    .col_out_432(u1_col_out_432),
    .col_out_433(u1_col_out_433),
    .col_out_434(u1_col_out_434),
    .col_out_435(u1_col_out_435),
    .col_out_436(u1_col_out_436),
    .col_out_437(u1_col_out_437),
    .col_out_438(u1_col_out_438),
    .col_out_439(u1_col_out_439),
    .col_out_440(u1_col_out_440),
    .col_out_441(u1_col_out_441),
    .col_out_442(u1_col_out_442),
    .col_out_443(u1_col_out_443),
    .col_out_444(u1_col_out_444),
    .col_out_445(u1_col_out_445),
    .col_out_446(u1_col_out_446),
    .col_out_447(u1_col_out_447),
    .col_out_448(u1_col_out_448),
    .col_out_449(u1_col_out_449),
    .col_out_450(u1_col_out_450),
    .col_out_451(u1_col_out_451),
    .col_out_452(u1_col_out_452),
    .col_out_453(u1_col_out_453),
    .col_out_454(u1_col_out_454),
    .col_out_455(u1_col_out_455),
    .col_out_456(u1_col_out_456),
    .col_out_457(u1_col_out_457),
    .col_out_458(u1_col_out_458),
    .col_out_459(u1_col_out_459),
    .col_out_460(u1_col_out_460),
    .col_out_461(u1_col_out_461),
    .col_out_462(u1_col_out_462),
    .col_out_463(u1_col_out_463),
    .col_out_464(u1_col_out_464),
    .col_out_465(u1_col_out_465),
    .col_out_466(u1_col_out_466),
    .col_out_467(u1_col_out_467),
    .col_out_468(u1_col_out_468),
    .col_out_469(u1_col_out_469),
    .col_out_470(u1_col_out_470),
    .col_out_471(u1_col_out_471),
    .col_out_472(u1_col_out_472),
    .col_out_473(u1_col_out_473),
    .col_out_474(u1_col_out_474),
    .col_out_475(u1_col_out_475),
    .col_out_476(u1_col_out_476),
    .col_out_477(u1_col_out_477),
    .col_out_478(u1_col_out_478),
    .col_out_479(u1_col_out_479),
    .col_out_480(u1_col_out_480),
    .col_out_481(u1_col_out_481),
    .col_out_482(u1_col_out_482),
    .col_out_483(u1_col_out_483),
    .col_out_484(u1_col_out_484),
    .col_out_485(u1_col_out_485),
    .col_out_486(u1_col_out_486),
    .col_out_487(u1_col_out_487),
    .col_out_488(u1_col_out_488),
    .col_out_489(u1_col_out_489),
    .col_out_490(u1_col_out_490),
    .col_out_491(u1_col_out_491),
    .col_out_492(u1_col_out_492),
    .col_out_493(u1_col_out_493),
    .col_out_494(u1_col_out_494),
    .col_out_495(u1_col_out_495),
    .col_out_496(u1_col_out_496),
    .col_out_497(u1_col_out_497),
    .col_out_498(u1_col_out_498),
    .col_out_499(u1_col_out_499),
    .col_out_500(u1_col_out_500),
    .col_out_501(u1_col_out_501),
    .col_out_502(u1_col_out_502),
    .col_out_503(u1_col_out_503),
    .col_out_504(u1_col_out_504),
    .col_out_505(u1_col_out_505),
    .col_out_506(u1_col_out_506),
    .col_out_507(u1_col_out_507),
    .col_out_508(u1_col_out_508),
    .col_out_509(u1_col_out_509),
    .col_out_510(u1_col_out_510),
    .col_out_511(u1_col_out_511),
    .col_out_512(u1_col_out_512),
    .col_out_513(u1_col_out_513),
    .col_out_514(u1_col_out_514),
    .col_out_515(u1_col_out_515),
    .col_out_516(u1_col_out_516),
    .col_out_517(u1_col_out_517),
    .col_out_518(u1_col_out_518),
    .col_out_519(u1_col_out_519),
    .col_out_520(u1_col_out_520),
    .col_out_521(u1_col_out_521),
    .col_out_522(u1_col_out_522),
    .col_out_523(u1_col_out_523),
    .col_out_524(u1_col_out_524),
    .col_out_525(u1_col_out_525),
    .col_out_526(u1_col_out_526),
    .col_out_527(u1_col_out_527),
    .col_out_528(u1_col_out_528),
    .col_out_529(u1_col_out_529),
    .col_out_530(u1_col_out_530),
    .col_out_531(u1_col_out_531),
    .col_out_532(u1_col_out_532),
    .col_out_533(u1_col_out_533),
    .col_out_534(u1_col_out_534),
    .col_out_535(u1_col_out_535),
    .col_out_536(u1_col_out_536),
    .col_out_537(u1_col_out_537),
    .col_out_538(u1_col_out_538),
    .col_out_539(u1_col_out_539),
    .col_out_540(u1_col_out_540),
    .col_out_541(u1_col_out_541),
    .col_out_542(u1_col_out_542),
    .col_out_543(u1_col_out_543),
    .col_out_544(u1_col_out_544),
    .col_out_545(u1_col_out_545),
    .col_out_546(u1_col_out_546),
    .col_out_547(u1_col_out_547),
    .col_out_548(u1_col_out_548),
    .col_out_549(u1_col_out_549),
    .col_out_550(u1_col_out_550),
    .col_out_551(u1_col_out_551),
    .col_out_552(u1_col_out_552),
    .col_out_553(u1_col_out_553),
    .col_out_554(u1_col_out_554),
    .col_out_555(u1_col_out_555),
    .col_out_556(u1_col_out_556),
    .col_out_557(u1_col_out_557),
    .col_out_558(u1_col_out_558),
    .col_out_559(u1_col_out_559),
    .col_out_560(u1_col_out_560),
    .col_out_561(u1_col_out_561),
    .col_out_562(u1_col_out_562),
    .col_out_563(u1_col_out_563),
    .col_out_564(u1_col_out_564),
    .col_out_565(u1_col_out_565),
    .col_out_566(u1_col_out_566),
    .col_out_567(u1_col_out_567),
    .col_out_568(u1_col_out_568),
    .col_out_569(u1_col_out_569),
    .col_out_570(u1_col_out_570),
    .col_out_571(u1_col_out_571),
    .col_out_572(u1_col_out_572),
    .col_out_573(u1_col_out_573),
    .col_out_574(u1_col_out_574),
    .col_out_575(u1_col_out_575),
    .col_out_576(u1_col_out_576),
    .col_out_577(u1_col_out_577),
    .col_out_578(u1_col_out_578),
    .col_out_579(u1_col_out_579),
    .col_out_580(u1_col_out_580),
    .col_out_581(u1_col_out_581),
    .col_out_582(u1_col_out_582),
    .col_out_583(u1_col_out_583),
    .col_out_584(u1_col_out_584),
    .col_out_585(u1_col_out_585),
    .col_out_586(u1_col_out_586),
    .col_out_587(u1_col_out_587),
    .col_out_588(u1_col_out_588),
    .col_out_589(u1_col_out_589),
    .col_out_590(u1_col_out_590),
    .col_out_591(u1_col_out_591),
    .col_out_592(u1_col_out_592),
    .col_out_593(u1_col_out_593),
    .col_out_594(u1_col_out_594),
    .col_out_595(u1_col_out_595),
    .col_out_596(u1_col_out_596),
    .col_out_597(u1_col_out_597),
    .col_out_598(u1_col_out_598),
    .col_out_599(u1_col_out_599),
    .col_out_600(u1_col_out_600),
    .col_out_601(u1_col_out_601),
    .col_out_602(u1_col_out_602),
    .col_out_603(u1_col_out_603),
    .col_out_604(u1_col_out_604),
    .col_out_605(u1_col_out_605),
    .col_out_606(u1_col_out_606),
    .col_out_607(u1_col_out_607),
    .col_out_608(u1_col_out_608),
    .col_out_609(u1_col_out_609),
    .col_out_610(u1_col_out_610),
    .col_out_611(u1_col_out_611),
    .col_out_612(u1_col_out_612),
    .col_out_613(u1_col_out_613),
    .col_out_614(u1_col_out_614),
    .col_out_615(u1_col_out_615),
    .col_out_616(u1_col_out_616),
    .col_out_617(u1_col_out_617),
    .col_out_618(u1_col_out_618),
    .col_out_619(u1_col_out_619),
    .col_out_620(u1_col_out_620),
    .col_out_621(u1_col_out_621),
    .col_out_622(u1_col_out_622),
    .col_out_623(u1_col_out_623),
    .col_out_624(u1_col_out_624),
    .col_out_625(u1_col_out_625),
    .col_out_626(u1_col_out_626),
    .col_out_627(u1_col_out_627),
    .col_out_628(u1_col_out_628),
    .col_out_629(u1_col_out_629),
    .col_out_630(u1_col_out_630),
    .col_out_631(u1_col_out_631),
    .col_out_632(u1_col_out_632),
    .col_out_633(u1_col_out_633),
    .col_out_634(u1_col_out_634),
    .col_out_635(u1_col_out_635),
    .col_out_636(u1_col_out_636),
    .col_out_637(u1_col_out_637),
    .col_out_638(u1_col_out_638),
    .col_out_639(u1_col_out_639),
    .col_out_640(u1_col_out_640),
    .col_out_641(u1_col_out_641),
    .col_out_642(u1_col_out_642),
    .col_out_643(u1_col_out_643),
    .col_out_644(u1_col_out_644),
    .col_out_645(u1_col_out_645),
    .col_out_646(u1_col_out_646),
    .col_out_647(u1_col_out_647),
    .col_out_648(u1_col_out_648),
    .col_out_649(u1_col_out_649),
    .col_out_650(u1_col_out_650),
    .col_out_651(u1_col_out_651),
    .col_out_652(u1_col_out_652),
    .col_out_653(u1_col_out_653),
    .col_out_654(u1_col_out_654),
    .col_out_655(u1_col_out_655),
    .col_out_656(u1_col_out_656),
    .col_out_657(u1_col_out_657),
    .col_out_658(u1_col_out_658),
    .col_out_659(u1_col_out_659),
    .col_out_660(u1_col_out_660),
    .col_out_661(u1_col_out_661),
    .col_out_662(u1_col_out_662),
    .col_out_663(u1_col_out_663),
    .col_out_664(u1_col_out_664),
    .col_out_665(u1_col_out_665),
    .col_out_666(u1_col_out_666),
    .col_out_667(u1_col_out_667),
    .col_out_668(u1_col_out_668),
    .col_out_669(u1_col_out_669),
    .col_out_670(u1_col_out_670),
    .col_out_671(u1_col_out_671),
    .col_out_672(u1_col_out_672),
    .col_out_673(u1_col_out_673),
    .col_out_674(u1_col_out_674),
    .col_out_675(u1_col_out_675),
    .col_out_676(u1_col_out_676),
    .col_out_677(u1_col_out_677),
    .col_out_678(u1_col_out_678),
    .col_out_679(u1_col_out_679),
    .col_out_680(u1_col_out_680),
    .col_out_681(u1_col_out_681),
    .col_out_682(u1_col_out_682),
    .col_out_683(u1_col_out_683),
    .col_out_684(u1_col_out_684),
    .col_out_685(u1_col_out_685),
    .col_out_686(u1_col_out_686),
    .col_out_687(u1_col_out_687),
    .col_out_688(u1_col_out_688),
    .col_out_689(u1_col_out_689),
    .col_out_690(u1_col_out_690),
    .col_out_691(u1_col_out_691),
    .col_out_692(u1_col_out_692),
    .col_out_693(u1_col_out_693),
    .col_out_694(u1_col_out_694),
    .col_out_695(u1_col_out_695),
    .col_out_696(u1_col_out_696),
    .col_out_697(u1_col_out_697),
    .col_out_698(u1_col_out_698),
    .col_out_699(u1_col_out_699),
    .col_out_700(u1_col_out_700),
    .col_out_701(u1_col_out_701),
    .col_out_702(u1_col_out_702),
    .col_out_703(u1_col_out_703),
    .col_out_704(u1_col_out_704),
    .col_out_705(u1_col_out_705),
    .col_out_706(u1_col_out_706),
    .col_out_707(u1_col_out_707),
    .col_out_708(u1_col_out_708),
    .col_out_709(u1_col_out_709),
    .col_out_710(u1_col_out_710),
    .col_out_711(u1_col_out_711),
    .col_out_712(u1_col_out_712),
    .col_out_713(u1_col_out_713),
    .col_out_714(u1_col_out_714),
    .col_out_715(u1_col_out_715),
    .col_out_716(u1_col_out_716),
    .col_out_717(u1_col_out_717),
    .col_out_718(u1_col_out_718),
    .col_out_719(u1_col_out_719),
    .col_out_720(u1_col_out_720),
    .col_out_721(u1_col_out_721),
    .col_out_722(u1_col_out_722),
    .col_out_723(u1_col_out_723),
    .col_out_724(u1_col_out_724),
    .col_out_725(u1_col_out_725),
    .col_out_726(u1_col_out_726),
    .col_out_727(u1_col_out_727),
    .col_out_728(u1_col_out_728),
    .col_out_729(u1_col_out_729),
    .col_out_730(u1_col_out_730),
    .col_out_731(u1_col_out_731),
    .col_out_732(u1_col_out_732),
    .col_out_733(u1_col_out_733),
    .col_out_734(u1_col_out_734),
    .col_out_735(u1_col_out_735),
    .col_out_736(u1_col_out_736),
    .col_out_737(u1_col_out_737),
    .col_out_738(u1_col_out_738),
    .col_out_739(u1_col_out_739),
    .col_out_740(u1_col_out_740),
    .col_out_741(u1_col_out_741),
    .col_out_742(u1_col_out_742),
    .col_out_743(u1_col_out_743),
    .col_out_744(u1_col_out_744),
    .col_out_745(u1_col_out_745),
    .col_out_746(u1_col_out_746),
    .col_out_747(u1_col_out_747),
    .col_out_748(u1_col_out_748),
    .col_out_749(u1_col_out_749),
    .col_out_750(u1_col_out_750),
    .col_out_751(u1_col_out_751),
    .col_out_752(u1_col_out_752),
    .col_out_753(u1_col_out_753),
    .col_out_754(u1_col_out_754),
    .col_out_755(u1_col_out_755),
    .col_out_756(u1_col_out_756),
    .col_out_757(u1_col_out_757),
    .col_out_758(u1_col_out_758),
    .col_out_759(u1_col_out_759),
    .col_out_760(u1_col_out_760),
    .col_out_761(u1_col_out_761),
    .col_out_762(u1_col_out_762),
    .col_out_763(u1_col_out_763),
    .col_out_764(u1_col_out_764),
    .col_out_765(u1_col_out_765),
    .col_out_766(u1_col_out_766),
    .col_out_767(u1_col_out_767),
    .col_out_768(u1_col_out_768),
    .col_out_769(u1_col_out_769),
    .col_out_770(u1_col_out_770),
    .col_out_771(u1_col_out_771),
    .col_out_772(u1_col_out_772),
    .col_out_773(u1_col_out_773),
    .col_out_774(u1_col_out_774),
    .col_out_775(u1_col_out_775),
    .col_out_776(u1_col_out_776),
    .col_out_777(u1_col_out_777),
    .col_out_778(u1_col_out_778),
    .col_out_779(u1_col_out_779),
    .col_out_780(u1_col_out_780),
    .col_out_781(u1_col_out_781),
    .col_out_782(u1_col_out_782),
    .col_out_783(u1_col_out_783),
    .col_out_784(u1_col_out_784),
    .col_out_785(u1_col_out_785),
    .col_out_786(u1_col_out_786),
    .col_out_787(u1_col_out_787),
    .col_out_788(u1_col_out_788),
    .col_out_789(u1_col_out_789),
    .col_out_790(u1_col_out_790),
    .col_out_791(u1_col_out_791),
    .col_out_792(u1_col_out_792),
    .col_out_793(u1_col_out_793),
    .col_out_794(u1_col_out_794),
    .col_out_795(u1_col_out_795),
    .col_out_796(u1_col_out_796),
    .col_out_797(u1_col_out_797),
    .col_out_798(u1_col_out_798),
    .col_out_799(u1_col_out_799),
    .col_out_800(u1_col_out_800),
    .col_out_801(u1_col_out_801),
    .col_out_802(u1_col_out_802),
    .col_out_803(u1_col_out_803),
    .col_out_804(u1_col_out_804),
    .col_out_805(u1_col_out_805),
    .col_out_806(u1_col_out_806),
    .col_out_807(u1_col_out_807),
    .col_out_808(u1_col_out_808),
    .col_out_809(u1_col_out_809),
    .col_out_810(u1_col_out_810),
    .col_out_811(u1_col_out_811),
    .col_out_812(u1_col_out_812),
    .col_out_813(u1_col_out_813),
    .col_out_814(u1_col_out_814),
    .col_out_815(u1_col_out_815),
    .col_out_816(u1_col_out_816),
    .col_out_817(u1_col_out_817),
    .col_out_818(u1_col_out_818),
    .col_out_819(u1_col_out_819),
    .col_out_820(u1_col_out_820),
    .col_out_821(u1_col_out_821),
    .col_out_822(u1_col_out_822),
    .col_out_823(u1_col_out_823),
    .col_out_824(u1_col_out_824),
    .col_out_825(u1_col_out_825),
    .col_out_826(u1_col_out_826),
    .col_out_827(u1_col_out_827),
    .col_out_828(u1_col_out_828),
    .col_out_829(u1_col_out_829),
    .col_out_830(u1_col_out_830),
    .col_out_831(u1_col_out_831),
    .col_out_832(u1_col_out_832),
    .col_out_833(u1_col_out_833),
    .col_out_834(u1_col_out_834),
    .col_out_835(u1_col_out_835),
    .col_out_836(u1_col_out_836),
    .col_out_837(u1_col_out_837),
    .col_out_838(u1_col_out_838),
    .col_out_839(u1_col_out_839),
    .col_out_840(u1_col_out_840),
    .col_out_841(u1_col_out_841),
    .col_out_842(u1_col_out_842),
    .col_out_843(u1_col_out_843),
    .col_out_844(u1_col_out_844),
    .col_out_845(u1_col_out_845),
    .col_out_846(u1_col_out_846),
    .col_out_847(u1_col_out_847),
    .col_out_848(u1_col_out_848),
    .col_out_849(u1_col_out_849),
    .col_out_850(u1_col_out_850),
    .col_out_851(u1_col_out_851),
    .col_out_852(u1_col_out_852),
    .col_out_853(u1_col_out_853),
    .col_out_854(u1_col_out_854),
    .col_out_855(u1_col_out_855),
    .col_out_856(u1_col_out_856),
    .col_out_857(u1_col_out_857),
    .col_out_858(u1_col_out_858),
    .col_out_859(u1_col_out_859),
    .col_out_860(u1_col_out_860),
    .col_out_861(u1_col_out_861),
    .col_out_862(u1_col_out_862),
    .col_out_863(u1_col_out_863),
    .col_out_864(u1_col_out_864),
    .col_out_865(u1_col_out_865),
    .col_out_866(u1_col_out_866),
    .col_out_867(u1_col_out_867),
    .col_out_868(u1_col_out_868),
    .col_out_869(u1_col_out_869),
    .col_out_870(u1_col_out_870),
    .col_out_871(u1_col_out_871),
    .col_out_872(u1_col_out_872),
    .col_out_873(u1_col_out_873),
    .col_out_874(u1_col_out_874),
    .col_out_875(u1_col_out_875),
    .col_out_876(u1_col_out_876),
    .col_out_877(u1_col_out_877),
    .col_out_878(u1_col_out_878),
    .col_out_879(u1_col_out_879),
    .col_out_880(u1_col_out_880),
    .col_out_881(u1_col_out_881),
    .col_out_882(u1_col_out_882),
    .col_out_883(u1_col_out_883),
    .col_out_884(u1_col_out_884),
    .col_out_885(u1_col_out_885),
    .col_out_886(u1_col_out_886),
    .col_out_887(u1_col_out_887),
    .col_out_888(u1_col_out_888),
    .col_out_889(u1_col_out_889),
    .col_out_890(u1_col_out_890),
    .col_out_891(u1_col_out_891),
    .col_out_892(u1_col_out_892),
    .col_out_893(u1_col_out_893),
    .col_out_894(u1_col_out_894),
    .col_out_895(u1_col_out_895),
    .col_out_896(u1_col_out_896),
    .col_out_897(u1_col_out_897),
    .col_out_898(u1_col_out_898),
    .col_out_899(u1_col_out_899),
    .col_out_900(u1_col_out_900),
    .col_out_901(u1_col_out_901),
    .col_out_902(u1_col_out_902),
    .col_out_903(u1_col_out_903),
    .col_out_904(u1_col_out_904),
    .col_out_905(u1_col_out_905),
    .col_out_906(u1_col_out_906),
    .col_out_907(u1_col_out_907),
    .col_out_908(u1_col_out_908),
    .col_out_909(u1_col_out_909),
    .col_out_910(u1_col_out_910),
    .col_out_911(u1_col_out_911),
    .col_out_912(u1_col_out_912),
    .col_out_913(u1_col_out_913),
    .col_out_914(u1_col_out_914),
    .col_out_915(u1_col_out_915),
    .col_out_916(u1_col_out_916),
    .col_out_917(u1_col_out_917),
    .col_out_918(u1_col_out_918),
    .col_out_919(u1_col_out_919),
    .col_out_920(u1_col_out_920),
    .col_out_921(u1_col_out_921),
    .col_out_922(u1_col_out_922),
    .col_out_923(u1_col_out_923),
    .col_out_924(u1_col_out_924),
    .col_out_925(u1_col_out_925),
    .col_out_926(u1_col_out_926),
    .col_out_927(u1_col_out_927),
    .col_out_928(u1_col_out_928),
    .col_out_929(u1_col_out_929),
    .col_out_930(u1_col_out_930),
    .col_out_931(u1_col_out_931),
    .col_out_932(u1_col_out_932),
    .col_out_933(u1_col_out_933),
    .col_out_934(u1_col_out_934),
    .col_out_935(u1_col_out_935),
    .col_out_936(u1_col_out_936),
    .col_out_937(u1_col_out_937),
    .col_out_938(u1_col_out_938),
    .col_out_939(u1_col_out_939),
    .col_out_940(u1_col_out_940),
    .col_out_941(u1_col_out_941),
    .col_out_942(u1_col_out_942),
    .col_out_943(u1_col_out_943),
    .col_out_944(u1_col_out_944),
    .col_out_945(u1_col_out_945),
    .col_out_946(u1_col_out_946),
    .col_out_947(u1_col_out_947),
    .col_out_948(u1_col_out_948),
    .col_out_949(u1_col_out_949),
    .col_out_950(u1_col_out_950),
    .col_out_951(u1_col_out_951),
    .col_out_952(u1_col_out_952),
    .col_out_953(u1_col_out_953),
    .col_out_954(u1_col_out_954),
    .col_out_955(u1_col_out_955),
    .col_out_956(u1_col_out_956),
    .col_out_957(u1_col_out_957),
    .col_out_958(u1_col_out_958),
    .col_out_959(u1_col_out_959),
    .col_out_960(u1_col_out_960),
    .col_out_961(u1_col_out_961),
    .col_out_962(u1_col_out_962),
    .col_out_963(u1_col_out_963),
    .col_out_964(u1_col_out_964),
    .col_out_965(u1_col_out_965),
    .col_out_966(u1_col_out_966),
    .col_out_967(u1_col_out_967),
    .col_out_968(u1_col_out_968),
    .col_out_969(u1_col_out_969),
    .col_out_970(u1_col_out_970),
    .col_out_971(u1_col_out_971),
    .col_out_972(u1_col_out_972),
    .col_out_973(u1_col_out_973),
    .col_out_974(u1_col_out_974),
    .col_out_975(u1_col_out_975),
    .col_out_976(u1_col_out_976),
    .col_out_977(u1_col_out_977),
    .col_out_978(u1_col_out_978),
    .col_out_979(u1_col_out_979),
    .col_out_980(u1_col_out_980),
    .col_out_981(u1_col_out_981),
    .col_out_982(u1_col_out_982),
    .col_out_983(u1_col_out_983),
    .col_out_984(u1_col_out_984),
    .col_out_985(u1_col_out_985),
    .col_out_986(u1_col_out_986),
    .col_out_987(u1_col_out_987),
    .col_out_988(u1_col_out_988),
    .col_out_989(u1_col_out_989),
    .col_out_990(u1_col_out_990),
    .col_out_991(u1_col_out_991),
    .col_out_992(u1_col_out_992),
    .col_out_993(u1_col_out_993),
    .col_out_994(u1_col_out_994),
    .col_out_995(u1_col_out_995),
    .col_out_996(u1_col_out_996),
    .col_out_997(u1_col_out_997),
    .col_out_998(u1_col_out_998),
    .col_out_999(u1_col_out_999),
    .col_out_1000(u1_col_out_1000),
    .col_out_1001(u1_col_out_1001),
    .col_out_1002(u1_col_out_1002),
    .col_out_1003(u1_col_out_1003),
    .col_out_1004(u1_col_out_1004),
    .col_out_1005(u1_col_out_1005),
    .col_out_1006(u1_col_out_1006),
    .col_out_1007(u1_col_out_1007),
    .col_out_1008(u1_col_out_1008),
    .col_out_1009(u1_col_out_1009),
    .col_out_1010(u1_col_out_1010),
    .col_out_1011(u1_col_out_1011),
    .col_out_1012(u1_col_out_1012),
    .col_out_1013(u1_col_out_1013),
    .col_out_1014(u1_col_out_1014),
    .col_out_1015(u1_col_out_1015),
    .col_out_1016(u1_col_out_1016),
    .col_out_1017(u1_col_out_1017),
    .col_out_1018(u1_col_out_1018),
    .col_out_1019(u1_col_out_1019),
    .col_out_1020(u1_col_out_1020),
    .col_out_1021(u1_col_out_1021),
    .col_out_1022(u1_col_out_1022),
    .col_out_1023(u1_col_out_1023),
    .col_out_1024(u1_col_out_1024),
    .col_out_1025(u1_col_out_1025),
    .col_out_1026(u1_col_out_1026),
    .col_out_1027(u1_col_out_1027),
    .col_out_1028(u1_col_out_1028),
    .col_out_1029(u1_col_out_1029)
);




















//*****************************************************
//**************u2输入定义******************************
//*****************************************************
wire [47:0] u2_col_in_0;
wire [47:0] u2_col_in_1;
wire [47:0] u2_col_in_2;
wire [47:0] u2_col_in_3;
wire [47:0] u2_col_in_4;
wire [47:0] u2_col_in_5;
wire [47:0] u2_col_in_6;
wire [47:0] u2_col_in_7;
wire [47:0] u2_col_in_8;
wire [47:0] u2_col_in_9;
wire [47:0] u2_col_in_10;
wire [47:0] u2_col_in_11;
wire [47:0] u2_col_in_12;
wire [47:0] u2_col_in_13;
wire [47:0] u2_col_in_14;
wire [47:0] u2_col_in_15;
wire [47:0] u2_col_in_16;
wire [47:0] u2_col_in_17;
wire [47:0] u2_col_in_18;
wire [47:0] u2_col_in_19;
wire [47:0] u2_col_in_20;
wire [47:0] u2_col_in_21;
wire [47:0] u2_col_in_22;
wire [47:0] u2_col_in_23;
wire [47:0] u2_col_in_24;
wire [47:0] u2_col_in_25;
wire [47:0] u2_col_in_26;
wire [47:0] u2_col_in_27;
wire [47:0] u2_col_in_28;
wire [47:0] u2_col_in_29;
wire [47:0] u2_col_in_30;
wire [47:0] u2_col_in_31;
wire [47:0] u2_col_in_32;
wire [47:0] u2_col_in_33;
wire [47:0] u2_col_in_34;
wire [47:0] u2_col_in_35;
wire [47:0] u2_col_in_36;
wire [47:0] u2_col_in_37;
wire [47:0] u2_col_in_38;
wire [47:0] u2_col_in_39;
wire [47:0] u2_col_in_40;
wire [47:0] u2_col_in_41;
wire [47:0] u2_col_in_42;
wire [47:0] u2_col_in_43;
wire [47:0] u2_col_in_44;
wire [47:0] u2_col_in_45;
wire [47:0] u2_col_in_46;
wire [47:0] u2_col_in_47;
wire [47:0] u2_col_in_48;
wire [47:0] u2_col_in_49;
wire [47:0] u2_col_in_50;
wire [47:0] u2_col_in_51;
wire [47:0] u2_col_in_52;
wire [47:0] u2_col_in_53;
wire [47:0] u2_col_in_54;
wire [47:0] u2_col_in_55;
wire [47:0] u2_col_in_56;
wire [47:0] u2_col_in_57;
wire [47:0] u2_col_in_58;
wire [47:0] u2_col_in_59;
wire [47:0] u2_col_in_60;
wire [47:0] u2_col_in_61;
wire [47:0] u2_col_in_62;
wire [47:0] u2_col_in_63;
wire [47:0] u2_col_in_64;
wire [47:0] u2_col_in_65;
wire [47:0] u2_col_in_66;
wire [47:0] u2_col_in_67;
wire [47:0] u2_col_in_68;
wire [47:0] u2_col_in_69;
wire [47:0] u2_col_in_70;
wire [47:0] u2_col_in_71;
wire [47:0] u2_col_in_72;
wire [47:0] u2_col_in_73;
wire [47:0] u2_col_in_74;
wire [47:0] u2_col_in_75;
wire [47:0] u2_col_in_76;
wire [47:0] u2_col_in_77;
wire [47:0] u2_col_in_78;
wire [47:0] u2_col_in_79;
wire [47:0] u2_col_in_80;
wire [47:0] u2_col_in_81;
wire [47:0] u2_col_in_82;
wire [47:0] u2_col_in_83;
wire [47:0] u2_col_in_84;
wire [47:0] u2_col_in_85;
wire [47:0] u2_col_in_86;
wire [47:0] u2_col_in_87;
wire [47:0] u2_col_in_88;
wire [47:0] u2_col_in_89;
wire [47:0] u2_col_in_90;
wire [47:0] u2_col_in_91;
wire [47:0] u2_col_in_92;
wire [47:0] u2_col_in_93;
wire [47:0] u2_col_in_94;
wire [47:0] u2_col_in_95;
wire [47:0] u2_col_in_96;
wire [47:0] u2_col_in_97;
wire [47:0] u2_col_in_98;
wire [47:0] u2_col_in_99;
wire [47:0] u2_col_in_100;
wire [47:0] u2_col_in_101;
wire [47:0] u2_col_in_102;
wire [47:0] u2_col_in_103;
wire [47:0] u2_col_in_104;
wire [47:0] u2_col_in_105;
wire [47:0] u2_col_in_106;
wire [47:0] u2_col_in_107;
wire [47:0] u2_col_in_108;
wire [47:0] u2_col_in_109;
wire [47:0] u2_col_in_110;
wire [47:0] u2_col_in_111;
wire [47:0] u2_col_in_112;
wire [47:0] u2_col_in_113;
wire [47:0] u2_col_in_114;
wire [47:0] u2_col_in_115;
wire [47:0] u2_col_in_116;
wire [47:0] u2_col_in_117;
wire [47:0] u2_col_in_118;
wire [47:0] u2_col_in_119;
wire [47:0] u2_col_in_120;
wire [47:0] u2_col_in_121;
wire [47:0] u2_col_in_122;
wire [47:0] u2_col_in_123;
wire [47:0] u2_col_in_124;
wire [47:0] u2_col_in_125;
wire [47:0] u2_col_in_126;
wire [47:0] u2_col_in_127;
wire [47:0] u2_col_in_128;
wire [47:0] u2_col_in_129;
wire [47:0] u2_col_in_130;
wire [47:0] u2_col_in_131;
wire [47:0] u2_col_in_132;
wire [47:0] u2_col_in_133;
wire [47:0] u2_col_in_134;
wire [47:0] u2_col_in_135;
wire [47:0] u2_col_in_136;
wire [47:0] u2_col_in_137;
wire [47:0] u2_col_in_138;
wire [47:0] u2_col_in_139;
wire [47:0] u2_col_in_140;
wire [47:0] u2_col_in_141;
wire [47:0] u2_col_in_142;
wire [47:0] u2_col_in_143;
wire [47:0] u2_col_in_144;
wire [47:0] u2_col_in_145;
wire [47:0] u2_col_in_146;
wire [47:0] u2_col_in_147;
wire [47:0] u2_col_in_148;
wire [47:0] u2_col_in_149;
wire [47:0] u2_col_in_150;
wire [47:0] u2_col_in_151;
wire [47:0] u2_col_in_152;
wire [47:0] u2_col_in_153;
wire [47:0] u2_col_in_154;
wire [47:0] u2_col_in_155;
wire [47:0] u2_col_in_156;
wire [47:0] u2_col_in_157;
wire [47:0] u2_col_in_158;
wire [47:0] u2_col_in_159;
wire [47:0] u2_col_in_160;
wire [47:0] u2_col_in_161;
wire [47:0] u2_col_in_162;
wire [47:0] u2_col_in_163;
wire [47:0] u2_col_in_164;
wire [47:0] u2_col_in_165;
wire [47:0] u2_col_in_166;
wire [47:0] u2_col_in_167;
wire [47:0] u2_col_in_168;
wire [47:0] u2_col_in_169;
wire [47:0] u2_col_in_170;
wire [47:0] u2_col_in_171;
wire [47:0] u2_col_in_172;
wire [47:0] u2_col_in_173;
wire [47:0] u2_col_in_174;
wire [47:0] u2_col_in_175;
wire [47:0] u2_col_in_176;
wire [47:0] u2_col_in_177;
wire [47:0] u2_col_in_178;
wire [47:0] u2_col_in_179;
wire [47:0] u2_col_in_180;
wire [47:0] u2_col_in_181;
wire [47:0] u2_col_in_182;
wire [47:0] u2_col_in_183;
wire [47:0] u2_col_in_184;
wire [47:0] u2_col_in_185;
wire [47:0] u2_col_in_186;
wire [47:0] u2_col_in_187;
wire [47:0] u2_col_in_188;
wire [47:0] u2_col_in_189;
wire [47:0] u2_col_in_190;
wire [47:0] u2_col_in_191;
wire [47:0] u2_col_in_192;
wire [47:0] u2_col_in_193;
wire [47:0] u2_col_in_194;
wire [47:0] u2_col_in_195;
wire [47:0] u2_col_in_196;
wire [47:0] u2_col_in_197;
wire [47:0] u2_col_in_198;
wire [47:0] u2_col_in_199;
wire [47:0] u2_col_in_200;
wire [47:0] u2_col_in_201;
wire [47:0] u2_col_in_202;
wire [47:0] u2_col_in_203;
wire [47:0] u2_col_in_204;
wire [47:0] u2_col_in_205;
wire [47:0] u2_col_in_206;
wire [47:0] u2_col_in_207;
wire [47:0] u2_col_in_208;
wire [47:0] u2_col_in_209;
wire [47:0] u2_col_in_210;
wire [47:0] u2_col_in_211;
wire [47:0] u2_col_in_212;
wire [47:0] u2_col_in_213;
wire [47:0] u2_col_in_214;
wire [47:0] u2_col_in_215;
wire [47:0] u2_col_in_216;
wire [47:0] u2_col_in_217;
wire [47:0] u2_col_in_218;
wire [47:0] u2_col_in_219;
wire [47:0] u2_col_in_220;
wire [47:0] u2_col_in_221;
wire [47:0] u2_col_in_222;
wire [47:0] u2_col_in_223;
wire [47:0] u2_col_in_224;
wire [47:0] u2_col_in_225;
wire [47:0] u2_col_in_226;
wire [47:0] u2_col_in_227;
wire [47:0] u2_col_in_228;
wire [47:0] u2_col_in_229;
wire [47:0] u2_col_in_230;
wire [47:0] u2_col_in_231;
wire [47:0] u2_col_in_232;
wire [47:0] u2_col_in_233;
wire [47:0] u2_col_in_234;
wire [47:0] u2_col_in_235;
wire [47:0] u2_col_in_236;
wire [47:0] u2_col_in_237;
wire [47:0] u2_col_in_238;
wire [47:0] u2_col_in_239;
wire [47:0] u2_col_in_240;
wire [47:0] u2_col_in_241;
wire [47:0] u2_col_in_242;
wire [47:0] u2_col_in_243;
wire [47:0] u2_col_in_244;
wire [47:0] u2_col_in_245;
wire [47:0] u2_col_in_246;
wire [47:0] u2_col_in_247;
wire [47:0] u2_col_in_248;
wire [47:0] u2_col_in_249;
wire [47:0] u2_col_in_250;
wire [47:0] u2_col_in_251;
wire [47:0] u2_col_in_252;
wire [47:0] u2_col_in_253;
wire [47:0] u2_col_in_254;
wire [47:0] u2_col_in_255;
wire [47:0] u2_col_in_256;
wire [47:0] u2_col_in_257;
wire [47:0] u2_col_in_258;
wire [47:0] u2_col_in_259;
wire [47:0] u2_col_in_260;
wire [47:0] u2_col_in_261;
wire [47:0] u2_col_in_262;
wire [47:0] u2_col_in_263;
wire [47:0] u2_col_in_264;
wire [47:0] u2_col_in_265;
wire [47:0] u2_col_in_266;
wire [47:0] u2_col_in_267;
wire [47:0] u2_col_in_268;
wire [47:0] u2_col_in_269;
wire [47:0] u2_col_in_270;
wire [47:0] u2_col_in_271;
wire [47:0] u2_col_in_272;
wire [47:0] u2_col_in_273;
wire [47:0] u2_col_in_274;
wire [47:0] u2_col_in_275;
wire [47:0] u2_col_in_276;
wire [47:0] u2_col_in_277;
wire [47:0] u2_col_in_278;
wire [47:0] u2_col_in_279;
wire [47:0] u2_col_in_280;
wire [47:0] u2_col_in_281;
wire [47:0] u2_col_in_282;
wire [47:0] u2_col_in_283;
wire [47:0] u2_col_in_284;
wire [47:0] u2_col_in_285;
wire [47:0] u2_col_in_286;
wire [47:0] u2_col_in_287;
wire [47:0] u2_col_in_288;
wire [47:0] u2_col_in_289;
wire [47:0] u2_col_in_290;
wire [47:0] u2_col_in_291;
wire [47:0] u2_col_in_292;
wire [47:0] u2_col_in_293;
wire [47:0] u2_col_in_294;
wire [47:0] u2_col_in_295;
wire [47:0] u2_col_in_296;
wire [47:0] u2_col_in_297;
wire [47:0] u2_col_in_298;
wire [47:0] u2_col_in_299;
wire [47:0] u2_col_in_300;
wire [47:0] u2_col_in_301;
wire [47:0] u2_col_in_302;
wire [47:0] u2_col_in_303;
wire [47:0] u2_col_in_304;
wire [47:0] u2_col_in_305;
wire [47:0] u2_col_in_306;
wire [47:0] u2_col_in_307;
wire [47:0] u2_col_in_308;
wire [47:0] u2_col_in_309;
wire [47:0] u2_col_in_310;
wire [47:0] u2_col_in_311;
wire [47:0] u2_col_in_312;
wire [47:0] u2_col_in_313;
wire [47:0] u2_col_in_314;
wire [47:0] u2_col_in_315;
wire [47:0] u2_col_in_316;
wire [47:0] u2_col_in_317;
wire [47:0] u2_col_in_318;
wire [47:0] u2_col_in_319;
wire [47:0] u2_col_in_320;
wire [47:0] u2_col_in_321;
wire [47:0] u2_col_in_322;
wire [47:0] u2_col_in_323;
wire [47:0] u2_col_in_324;
wire [47:0] u2_col_in_325;
wire [47:0] u2_col_in_326;
wire [47:0] u2_col_in_327;
wire [47:0] u2_col_in_328;
wire [47:0] u2_col_in_329;
wire [47:0] u2_col_in_330;
wire [47:0] u2_col_in_331;
wire [47:0] u2_col_in_332;
wire [47:0] u2_col_in_333;
wire [47:0] u2_col_in_334;
wire [47:0] u2_col_in_335;
wire [47:0] u2_col_in_336;
wire [47:0] u2_col_in_337;
wire [47:0] u2_col_in_338;
wire [47:0] u2_col_in_339;
wire [47:0] u2_col_in_340;
wire [47:0] u2_col_in_341;
wire [47:0] u2_col_in_342;
wire [47:0] u2_col_in_343;
wire [47:0] u2_col_in_344;
wire [47:0] u2_col_in_345;
wire [47:0] u2_col_in_346;
wire [47:0] u2_col_in_347;
wire [47:0] u2_col_in_348;
wire [47:0] u2_col_in_349;
wire [47:0] u2_col_in_350;
wire [47:0] u2_col_in_351;
wire [47:0] u2_col_in_352;
wire [47:0] u2_col_in_353;
wire [47:0] u2_col_in_354;
wire [47:0] u2_col_in_355;
wire [47:0] u2_col_in_356;
wire [47:0] u2_col_in_357;
wire [47:0] u2_col_in_358;
wire [47:0] u2_col_in_359;
wire [47:0] u2_col_in_360;
wire [47:0] u2_col_in_361;
wire [47:0] u2_col_in_362;
wire [47:0] u2_col_in_363;
wire [47:0] u2_col_in_364;
wire [47:0] u2_col_in_365;
wire [47:0] u2_col_in_366;
wire [47:0] u2_col_in_367;
wire [47:0] u2_col_in_368;
wire [47:0] u2_col_in_369;
wire [47:0] u2_col_in_370;
wire [47:0] u2_col_in_371;
wire [47:0] u2_col_in_372;
wire [47:0] u2_col_in_373;
wire [47:0] u2_col_in_374;
wire [47:0] u2_col_in_375;
wire [47:0] u2_col_in_376;
wire [47:0] u2_col_in_377;
wire [47:0] u2_col_in_378;
wire [47:0] u2_col_in_379;
wire [47:0] u2_col_in_380;
wire [47:0] u2_col_in_381;
wire [47:0] u2_col_in_382;
wire [47:0] u2_col_in_383;
wire [47:0] u2_col_in_384;
wire [47:0] u2_col_in_385;
wire [47:0] u2_col_in_386;
wire [47:0] u2_col_in_387;
wire [47:0] u2_col_in_388;
wire [47:0] u2_col_in_389;
wire [47:0] u2_col_in_390;
wire [47:0] u2_col_in_391;
wire [47:0] u2_col_in_392;
wire [47:0] u2_col_in_393;
wire [47:0] u2_col_in_394;
wire [47:0] u2_col_in_395;
wire [47:0] u2_col_in_396;
wire [47:0] u2_col_in_397;
wire [47:0] u2_col_in_398;
wire [47:0] u2_col_in_399;
wire [47:0] u2_col_in_400;
wire [47:0] u2_col_in_401;
wire [47:0] u2_col_in_402;
wire [47:0] u2_col_in_403;
wire [47:0] u2_col_in_404;
wire [47:0] u2_col_in_405;
wire [47:0] u2_col_in_406;
wire [47:0] u2_col_in_407;
wire [47:0] u2_col_in_408;
wire [47:0] u2_col_in_409;
wire [47:0] u2_col_in_410;
wire [47:0] u2_col_in_411;
wire [47:0] u2_col_in_412;
wire [47:0] u2_col_in_413;
wire [47:0] u2_col_in_414;
wire [47:0] u2_col_in_415;
wire [47:0] u2_col_in_416;
wire [47:0] u2_col_in_417;
wire [47:0] u2_col_in_418;
wire [47:0] u2_col_in_419;
wire [47:0] u2_col_in_420;
wire [47:0] u2_col_in_421;
wire [47:0] u2_col_in_422;
wire [47:0] u2_col_in_423;
wire [47:0] u2_col_in_424;
wire [47:0] u2_col_in_425;
wire [47:0] u2_col_in_426;
wire [47:0] u2_col_in_427;
wire [47:0] u2_col_in_428;
wire [47:0] u2_col_in_429;
wire [47:0] u2_col_in_430;
wire [47:0] u2_col_in_431;
wire [47:0] u2_col_in_432;
wire [47:0] u2_col_in_433;
wire [47:0] u2_col_in_434;
wire [47:0] u2_col_in_435;
wire [47:0] u2_col_in_436;
wire [47:0] u2_col_in_437;
wire [47:0] u2_col_in_438;
wire [47:0] u2_col_in_439;
wire [47:0] u2_col_in_440;
wire [47:0] u2_col_in_441;
wire [47:0] u2_col_in_442;
wire [47:0] u2_col_in_443;
wire [47:0] u2_col_in_444;
wire [47:0] u2_col_in_445;
wire [47:0] u2_col_in_446;
wire [47:0] u2_col_in_447;
wire [47:0] u2_col_in_448;
wire [47:0] u2_col_in_449;
wire [47:0] u2_col_in_450;
wire [47:0] u2_col_in_451;
wire [47:0] u2_col_in_452;
wire [47:0] u2_col_in_453;
wire [47:0] u2_col_in_454;
wire [47:0] u2_col_in_455;
wire [47:0] u2_col_in_456;
wire [47:0] u2_col_in_457;
wire [47:0] u2_col_in_458;
wire [47:0] u2_col_in_459;
wire [47:0] u2_col_in_460;
wire [47:0] u2_col_in_461;
wire [47:0] u2_col_in_462;
wire [47:0] u2_col_in_463;
wire [47:0] u2_col_in_464;
wire [47:0] u2_col_in_465;
wire [47:0] u2_col_in_466;
wire [47:0] u2_col_in_467;
wire [47:0] u2_col_in_468;
wire [47:0] u2_col_in_469;
wire [47:0] u2_col_in_470;
wire [47:0] u2_col_in_471;
wire [47:0] u2_col_in_472;
wire [47:0] u2_col_in_473;
wire [47:0] u2_col_in_474;
wire [47:0] u2_col_in_475;
wire [47:0] u2_col_in_476;
wire [47:0] u2_col_in_477;
wire [47:0] u2_col_in_478;
wire [47:0] u2_col_in_479;
wire [47:0] u2_col_in_480;
wire [47:0] u2_col_in_481;
wire [47:0] u2_col_in_482;
wire [47:0] u2_col_in_483;
wire [47:0] u2_col_in_484;
wire [47:0] u2_col_in_485;
wire [47:0] u2_col_in_486;
wire [47:0] u2_col_in_487;
wire [47:0] u2_col_in_488;
wire [47:0] u2_col_in_489;
wire [47:0] u2_col_in_490;
wire [47:0] u2_col_in_491;
wire [47:0] u2_col_in_492;
wire [47:0] u2_col_in_493;
wire [47:0] u2_col_in_494;
wire [47:0] u2_col_in_495;
wire [47:0] u2_col_in_496;
wire [47:0] u2_col_in_497;
wire [47:0] u2_col_in_498;
wire [47:0] u2_col_in_499;
wire [47:0] u2_col_in_500;
wire [47:0] u2_col_in_501;
wire [47:0] u2_col_in_502;
wire [47:0] u2_col_in_503;
wire [47:0] u2_col_in_504;
wire [47:0] u2_col_in_505;
wire [47:0] u2_col_in_506;
wire [47:0] u2_col_in_507;
wire [47:0] u2_col_in_508;
wire [47:0] u2_col_in_509;
wire [47:0] u2_col_in_510;
wire [47:0] u2_col_in_511;
wire [47:0] u2_col_in_512;
wire [47:0] u2_col_in_513;
wire [47:0] u2_col_in_514;
wire [47:0] u2_col_in_515;
wire [47:0] u2_col_in_516;
wire [47:0] u2_col_in_517;
wire [47:0] u2_col_in_518;
wire [47:0] u2_col_in_519;
wire [47:0] u2_col_in_520;
wire [47:0] u2_col_in_521;
wire [47:0] u2_col_in_522;
wire [47:0] u2_col_in_523;
wire [47:0] u2_col_in_524;
wire [47:0] u2_col_in_525;
wire [47:0] u2_col_in_526;
wire [47:0] u2_col_in_527;
wire [47:0] u2_col_in_528;
wire [47:0] u2_col_in_529;
wire [47:0] u2_col_in_530;
wire [47:0] u2_col_in_531;
wire [47:0] u2_col_in_532;
wire [47:0] u2_col_in_533;
wire [47:0] u2_col_in_534;
wire [47:0] u2_col_in_535;
wire [47:0] u2_col_in_536;
wire [47:0] u2_col_in_537;
wire [47:0] u2_col_in_538;
wire [47:0] u2_col_in_539;
wire [47:0] u2_col_in_540;
wire [47:0] u2_col_in_541;
wire [47:0] u2_col_in_542;
wire [47:0] u2_col_in_543;
wire [47:0] u2_col_in_544;
wire [47:0] u2_col_in_545;
wire [47:0] u2_col_in_546;
wire [47:0] u2_col_in_547;
wire [47:0] u2_col_in_548;
wire [47:0] u2_col_in_549;
wire [47:0] u2_col_in_550;
wire [47:0] u2_col_in_551;
wire [47:0] u2_col_in_552;
wire [47:0] u2_col_in_553;
wire [47:0] u2_col_in_554;
wire [47:0] u2_col_in_555;
wire [47:0] u2_col_in_556;
wire [47:0] u2_col_in_557;
wire [47:0] u2_col_in_558;
wire [47:0] u2_col_in_559;
wire [47:0] u2_col_in_560;
wire [47:0] u2_col_in_561;
wire [47:0] u2_col_in_562;
wire [47:0] u2_col_in_563;
wire [47:0] u2_col_in_564;
wire [47:0] u2_col_in_565;
wire [47:0] u2_col_in_566;
wire [47:0] u2_col_in_567;
wire [47:0] u2_col_in_568;
wire [47:0] u2_col_in_569;
wire [47:0] u2_col_in_570;
wire [47:0] u2_col_in_571;
wire [47:0] u2_col_in_572;
wire [47:0] u2_col_in_573;
wire [47:0] u2_col_in_574;
wire [47:0] u2_col_in_575;
wire [47:0] u2_col_in_576;
wire [47:0] u2_col_in_577;
wire [47:0] u2_col_in_578;
wire [47:0] u2_col_in_579;
wire [47:0] u2_col_in_580;
wire [47:0] u2_col_in_581;
wire [47:0] u2_col_in_582;
wire [47:0] u2_col_in_583;
wire [47:0] u2_col_in_584;
wire [47:0] u2_col_in_585;
wire [47:0] u2_col_in_586;
wire [47:0] u2_col_in_587;
wire [47:0] u2_col_in_588;
wire [47:0] u2_col_in_589;
wire [47:0] u2_col_in_590;
wire [47:0] u2_col_in_591;
wire [47:0] u2_col_in_592;
wire [47:0] u2_col_in_593;
wire [47:0] u2_col_in_594;
wire [47:0] u2_col_in_595;
wire [47:0] u2_col_in_596;
wire [47:0] u2_col_in_597;
wire [47:0] u2_col_in_598;
wire [47:0] u2_col_in_599;
wire [47:0] u2_col_in_600;
wire [47:0] u2_col_in_601;
wire [47:0] u2_col_in_602;
wire [47:0] u2_col_in_603;
wire [47:0] u2_col_in_604;
wire [47:0] u2_col_in_605;
wire [47:0] u2_col_in_606;
wire [47:0] u2_col_in_607;
wire [47:0] u2_col_in_608;
wire [47:0] u2_col_in_609;
wire [47:0] u2_col_in_610;
wire [47:0] u2_col_in_611;
wire [47:0] u2_col_in_612;
wire [47:0] u2_col_in_613;
wire [47:0] u2_col_in_614;
wire [47:0] u2_col_in_615;
wire [47:0] u2_col_in_616;
wire [47:0] u2_col_in_617;
wire [47:0] u2_col_in_618;
wire [47:0] u2_col_in_619;
wire [47:0] u2_col_in_620;
wire [47:0] u2_col_in_621;
wire [47:0] u2_col_in_622;
wire [47:0] u2_col_in_623;
wire [47:0] u2_col_in_624;
wire [47:0] u2_col_in_625;
wire [47:0] u2_col_in_626;
wire [47:0] u2_col_in_627;
wire [47:0] u2_col_in_628;
wire [47:0] u2_col_in_629;
wire [47:0] u2_col_in_630;
wire [47:0] u2_col_in_631;
wire [47:0] u2_col_in_632;
wire [47:0] u2_col_in_633;
wire [47:0] u2_col_in_634;
wire [47:0] u2_col_in_635;
wire [47:0] u2_col_in_636;
wire [47:0] u2_col_in_637;
wire [47:0] u2_col_in_638;
wire [47:0] u2_col_in_639;
wire [47:0] u2_col_in_640;
wire [47:0] u2_col_in_641;
wire [47:0] u2_col_in_642;
wire [47:0] u2_col_in_643;
wire [47:0] u2_col_in_644;
wire [47:0] u2_col_in_645;
wire [47:0] u2_col_in_646;
wire [47:0] u2_col_in_647;
wire [47:0] u2_col_in_648;
wire [47:0] u2_col_in_649;
wire [47:0] u2_col_in_650;
wire [47:0] u2_col_in_651;
wire [47:0] u2_col_in_652;
wire [47:0] u2_col_in_653;
wire [47:0] u2_col_in_654;
wire [47:0] u2_col_in_655;
wire [47:0] u2_col_in_656;
wire [47:0] u2_col_in_657;
wire [47:0] u2_col_in_658;
wire [47:0] u2_col_in_659;
wire [47:0] u2_col_in_660;
wire [47:0] u2_col_in_661;
wire [47:0] u2_col_in_662;
wire [47:0] u2_col_in_663;
wire [47:0] u2_col_in_664;
wire [47:0] u2_col_in_665;
wire [47:0] u2_col_in_666;
wire [47:0] u2_col_in_667;
wire [47:0] u2_col_in_668;
wire [47:0] u2_col_in_669;
wire [47:0] u2_col_in_670;
wire [47:0] u2_col_in_671;
wire [47:0] u2_col_in_672;
wire [47:0] u2_col_in_673;
wire [47:0] u2_col_in_674;
wire [47:0] u2_col_in_675;
wire [47:0] u2_col_in_676;
wire [47:0] u2_col_in_677;
wire [47:0] u2_col_in_678;
wire [47:0] u2_col_in_679;
wire [47:0] u2_col_in_680;
wire [47:0] u2_col_in_681;
wire [47:0] u2_col_in_682;
wire [47:0] u2_col_in_683;
wire [47:0] u2_col_in_684;
wire [47:0] u2_col_in_685;
wire [47:0] u2_col_in_686;
wire [47:0] u2_col_in_687;
wire [47:0] u2_col_in_688;
wire [47:0] u2_col_in_689;
wire [47:0] u2_col_in_690;
wire [47:0] u2_col_in_691;
wire [47:0] u2_col_in_692;
wire [47:0] u2_col_in_693;
wire [47:0] u2_col_in_694;
wire [47:0] u2_col_in_695;
wire [47:0] u2_col_in_696;
wire [47:0] u2_col_in_697;
wire [47:0] u2_col_in_698;
wire [47:0] u2_col_in_699;
wire [47:0] u2_col_in_700;
wire [47:0] u2_col_in_701;
wire [47:0] u2_col_in_702;
wire [47:0] u2_col_in_703;
wire [47:0] u2_col_in_704;
wire [47:0] u2_col_in_705;
wire [47:0] u2_col_in_706;
wire [47:0] u2_col_in_707;
wire [47:0] u2_col_in_708;
wire [47:0] u2_col_in_709;
wire [47:0] u2_col_in_710;
wire [47:0] u2_col_in_711;
wire [47:0] u2_col_in_712;
wire [47:0] u2_col_in_713;
wire [47:0] u2_col_in_714;
wire [47:0] u2_col_in_715;
wire [47:0] u2_col_in_716;
wire [47:0] u2_col_in_717;
wire [47:0] u2_col_in_718;
wire [47:0] u2_col_in_719;
wire [47:0] u2_col_in_720;
wire [47:0] u2_col_in_721;
wire [47:0] u2_col_in_722;
wire [47:0] u2_col_in_723;
wire [47:0] u2_col_in_724;
wire [47:0] u2_col_in_725;
wire [47:0] u2_col_in_726;
wire [47:0] u2_col_in_727;
wire [47:0] u2_col_in_728;
wire [47:0] u2_col_in_729;
wire [47:0] u2_col_in_730;
wire [47:0] u2_col_in_731;
wire [47:0] u2_col_in_732;
wire [47:0] u2_col_in_733;
wire [47:0] u2_col_in_734;
wire [47:0] u2_col_in_735;
wire [47:0] u2_col_in_736;
wire [47:0] u2_col_in_737;
wire [47:0] u2_col_in_738;
wire [47:0] u2_col_in_739;
wire [47:0] u2_col_in_740;
wire [47:0] u2_col_in_741;
wire [47:0] u2_col_in_742;
wire [47:0] u2_col_in_743;
wire [47:0] u2_col_in_744;
wire [47:0] u2_col_in_745;
wire [47:0] u2_col_in_746;
wire [47:0] u2_col_in_747;
wire [47:0] u2_col_in_748;
wire [47:0] u2_col_in_749;
wire [47:0] u2_col_in_750;
wire [47:0] u2_col_in_751;
wire [47:0] u2_col_in_752;
wire [47:0] u2_col_in_753;
wire [47:0] u2_col_in_754;
wire [47:0] u2_col_in_755;
wire [47:0] u2_col_in_756;
wire [47:0] u2_col_in_757;
wire [47:0] u2_col_in_758;
wire [47:0] u2_col_in_759;
wire [47:0] u2_col_in_760;
wire [47:0] u2_col_in_761;
wire [47:0] u2_col_in_762;
wire [47:0] u2_col_in_763;
wire [47:0] u2_col_in_764;
wire [47:0] u2_col_in_765;
wire [47:0] u2_col_in_766;
wire [47:0] u2_col_in_767;
wire [47:0] u2_col_in_768;
wire [47:0] u2_col_in_769;
wire [47:0] u2_col_in_770;
wire [47:0] u2_col_in_771;
wire [47:0] u2_col_in_772;
wire [47:0] u2_col_in_773;
wire [47:0] u2_col_in_774;
wire [47:0] u2_col_in_775;
wire [47:0] u2_col_in_776;
wire [47:0] u2_col_in_777;
wire [47:0] u2_col_in_778;
wire [47:0] u2_col_in_779;
wire [47:0] u2_col_in_780;
wire [47:0] u2_col_in_781;
wire [47:0] u2_col_in_782;
wire [47:0] u2_col_in_783;
wire [47:0] u2_col_in_784;
wire [47:0] u2_col_in_785;
wire [47:0] u2_col_in_786;
wire [47:0] u2_col_in_787;
wire [47:0] u2_col_in_788;
wire [47:0] u2_col_in_789;
wire [47:0] u2_col_in_790;
wire [47:0] u2_col_in_791;
wire [47:0] u2_col_in_792;
wire [47:0] u2_col_in_793;
wire [47:0] u2_col_in_794;
wire [47:0] u2_col_in_795;
wire [47:0] u2_col_in_796;
wire [47:0] u2_col_in_797;
wire [47:0] u2_col_in_798;
wire [47:0] u2_col_in_799;
wire [47:0] u2_col_in_800;
wire [47:0] u2_col_in_801;
wire [47:0] u2_col_in_802;
wire [47:0] u2_col_in_803;
wire [47:0] u2_col_in_804;
wire [47:0] u2_col_in_805;
wire [47:0] u2_col_in_806;
wire [47:0] u2_col_in_807;
wire [47:0] u2_col_in_808;
wire [47:0] u2_col_in_809;
wire [47:0] u2_col_in_810;
wire [47:0] u2_col_in_811;
wire [47:0] u2_col_in_812;
wire [47:0] u2_col_in_813;
wire [47:0] u2_col_in_814;
wire [47:0] u2_col_in_815;
wire [47:0] u2_col_in_816;
wire [47:0] u2_col_in_817;
wire [47:0] u2_col_in_818;
wire [47:0] u2_col_in_819;
wire [47:0] u2_col_in_820;
wire [47:0] u2_col_in_821;
wire [47:0] u2_col_in_822;
wire [47:0] u2_col_in_823;
wire [47:0] u2_col_in_824;
wire [47:0] u2_col_in_825;
wire [47:0] u2_col_in_826;
wire [47:0] u2_col_in_827;
wire [47:0] u2_col_in_828;
wire [47:0] u2_col_in_829;
wire [47:0] u2_col_in_830;
wire [47:0] u2_col_in_831;
wire [47:0] u2_col_in_832;
wire [47:0] u2_col_in_833;
wire [47:0] u2_col_in_834;
wire [47:0] u2_col_in_835;
wire [47:0] u2_col_in_836;
wire [47:0] u2_col_in_837;
wire [47:0] u2_col_in_838;
wire [47:0] u2_col_in_839;
wire [47:0] u2_col_in_840;
wire [47:0] u2_col_in_841;
wire [47:0] u2_col_in_842;
wire [47:0] u2_col_in_843;
wire [47:0] u2_col_in_844;
wire [47:0] u2_col_in_845;
wire [47:0] u2_col_in_846;
wire [47:0] u2_col_in_847;
wire [47:0] u2_col_in_848;
wire [47:0] u2_col_in_849;
wire [47:0] u2_col_in_850;
wire [47:0] u2_col_in_851;
wire [47:0] u2_col_in_852;
wire [47:0] u2_col_in_853;
wire [47:0] u2_col_in_854;
wire [47:0] u2_col_in_855;
wire [47:0] u2_col_in_856;
wire [47:0] u2_col_in_857;
wire [47:0] u2_col_in_858;
wire [47:0] u2_col_in_859;
wire [47:0] u2_col_in_860;
wire [47:0] u2_col_in_861;
wire [47:0] u2_col_in_862;
wire [47:0] u2_col_in_863;
wire [47:0] u2_col_in_864;
wire [47:0] u2_col_in_865;
wire [47:0] u2_col_in_866;
wire [47:0] u2_col_in_867;
wire [47:0] u2_col_in_868;
wire [47:0] u2_col_in_869;
wire [47:0] u2_col_in_870;
wire [47:0] u2_col_in_871;
wire [47:0] u2_col_in_872;
wire [47:0] u2_col_in_873;
wire [47:0] u2_col_in_874;
wire [47:0] u2_col_in_875;
wire [47:0] u2_col_in_876;
wire [47:0] u2_col_in_877;
wire [47:0] u2_col_in_878;
wire [47:0] u2_col_in_879;
wire [47:0] u2_col_in_880;
wire [47:0] u2_col_in_881;
wire [47:0] u2_col_in_882;
wire [47:0] u2_col_in_883;
wire [47:0] u2_col_in_884;
wire [47:0] u2_col_in_885;
wire [47:0] u2_col_in_886;
wire [47:0] u2_col_in_887;
wire [47:0] u2_col_in_888;
wire [47:0] u2_col_in_889;
wire [47:0] u2_col_in_890;
wire [47:0] u2_col_in_891;
wire [47:0] u2_col_in_892;
wire [47:0] u2_col_in_893;
wire [47:0] u2_col_in_894;
wire [47:0] u2_col_in_895;
wire [47:0] u2_col_in_896;
wire [47:0] u2_col_in_897;
wire [47:0] u2_col_in_898;
wire [47:0] u2_col_in_899;
wire [47:0] u2_col_in_900;
wire [47:0] u2_col_in_901;
wire [47:0] u2_col_in_902;
wire [47:0] u2_col_in_903;
wire [47:0] u2_col_in_904;
wire [47:0] u2_col_in_905;
wire [47:0] u2_col_in_906;
wire [47:0] u2_col_in_907;
wire [47:0] u2_col_in_908;
wire [47:0] u2_col_in_909;
wire [47:0] u2_col_in_910;
wire [47:0] u2_col_in_911;
wire [47:0] u2_col_in_912;
wire [47:0] u2_col_in_913;
wire [47:0] u2_col_in_914;
wire [47:0] u2_col_in_915;
wire [47:0] u2_col_in_916;
wire [47:0] u2_col_in_917;
wire [47:0] u2_col_in_918;
wire [47:0] u2_col_in_919;
wire [47:0] u2_col_in_920;
wire [47:0] u2_col_in_921;
wire [47:0] u2_col_in_922;
wire [47:0] u2_col_in_923;
wire [47:0] u2_col_in_924;
wire [47:0] u2_col_in_925;
wire [47:0] u2_col_in_926;
wire [47:0] u2_col_in_927;
wire [47:0] u2_col_in_928;
wire [47:0] u2_col_in_929;
wire [47:0] u2_col_in_930;
wire [47:0] u2_col_in_931;
wire [47:0] u2_col_in_932;
wire [47:0] u2_col_in_933;
wire [47:0] u2_col_in_934;
wire [47:0] u2_col_in_935;
wire [47:0] u2_col_in_936;
wire [47:0] u2_col_in_937;
wire [47:0] u2_col_in_938;
wire [47:0] u2_col_in_939;
wire [47:0] u2_col_in_940;
wire [47:0] u2_col_in_941;
wire [47:0] u2_col_in_942;
wire [47:0] u2_col_in_943;
wire [47:0] u2_col_in_944;
wire [47:0] u2_col_in_945;
wire [47:0] u2_col_in_946;
wire [47:0] u2_col_in_947;
wire [47:0] u2_col_in_948;
wire [47:0] u2_col_in_949;
wire [47:0] u2_col_in_950;
wire [47:0] u2_col_in_951;
wire [47:0] u2_col_in_952;
wire [47:0] u2_col_in_953;
wire [47:0] u2_col_in_954;
wire [47:0] u2_col_in_955;
wire [47:0] u2_col_in_956;
wire [47:0] u2_col_in_957;
wire [47:0] u2_col_in_958;
wire [47:0] u2_col_in_959;
wire [47:0] u2_col_in_960;
wire [47:0] u2_col_in_961;
wire [47:0] u2_col_in_962;
wire [47:0] u2_col_in_963;
wire [47:0] u2_col_in_964;
wire [47:0] u2_col_in_965;
wire [47:0] u2_col_in_966;
wire [47:0] u2_col_in_967;
wire [47:0] u2_col_in_968;
wire [47:0] u2_col_in_969;
wire [47:0] u2_col_in_970;
wire [47:0] u2_col_in_971;
wire [47:0] u2_col_in_972;
wire [47:0] u2_col_in_973;
wire [47:0] u2_col_in_974;
wire [47:0] u2_col_in_975;
wire [47:0] u2_col_in_976;
wire [47:0] u2_col_in_977;
wire [47:0] u2_col_in_978;
wire [47:0] u2_col_in_979;
wire [47:0] u2_col_in_980;
wire [47:0] u2_col_in_981;
wire [47:0] u2_col_in_982;
wire [47:0] u2_col_in_983;
wire [47:0] u2_col_in_984;
wire [47:0] u2_col_in_985;
wire [47:0] u2_col_in_986;
wire [47:0] u2_col_in_987;
wire [47:0] u2_col_in_988;
wire [47:0] u2_col_in_989;
wire [47:0] u2_col_in_990;
wire [47:0] u2_col_in_991;
wire [47:0] u2_col_in_992;
wire [47:0] u2_col_in_993;
wire [47:0] u2_col_in_994;
wire [47:0] u2_col_in_995;
wire [47:0] u2_col_in_996;
wire [47:0] u2_col_in_997;
wire [47:0] u2_col_in_998;
wire [47:0] u2_col_in_999;
wire [47:0] u2_col_in_1000;
wire [47:0] u2_col_in_1001;
wire [47:0] u2_col_in_1002;
wire [47:0] u2_col_in_1003;
wire [47:0] u2_col_in_1004;
wire [47:0] u2_col_in_1005;
wire [47:0] u2_col_in_1006;
wire [47:0] u2_col_in_1007;
wire [47:0] u2_col_in_1008;
wire [47:0] u2_col_in_1009;
wire [47:0] u2_col_in_1010;
wire [47:0] u2_col_in_1011;
wire [47:0] u2_col_in_1012;
wire [47:0] u2_col_in_1013;
wire [47:0] u2_col_in_1014;
wire [47:0] u2_col_in_1015;
wire [47:0] u2_col_in_1016;
wire [47:0] u2_col_in_1017;
wire [47:0] u2_col_in_1018;
wire [47:0] u2_col_in_1019;
wire [47:0] u2_col_in_1020;
wire [47:0] u2_col_in_1021;
wire [47:0] u2_col_in_1022;
wire [47:0] u2_col_in_1023;
wire [47:0] u2_col_in_1024;
wire [47:0] u2_col_in_1025;
wire [47:0] u2_col_in_1026;
wire [47:0] u2_col_in_1027;
wire [47:0] u2_col_in_1028;
wire [47:0] u2_col_in_1029;



//*****************************************************
//**************u2输出定义******************************
//*****************************************************
wire [15:0] u2_col_out_0;
wire [15:0] u2_col_out_1;
wire [15:0] u2_col_out_2;
wire [15:0] u2_col_out_3;
wire [15:0] u2_col_out_4;
wire [15:0] u2_col_out_5;
wire [15:0] u2_col_out_6;
wire [15:0] u2_col_out_7;
wire [15:0] u2_col_out_8;
wire [15:0] u2_col_out_9;
wire [15:0] u2_col_out_10;
wire [15:0] u2_col_out_11;
wire [15:0] u2_col_out_12;
wire [15:0] u2_col_out_13;
wire [15:0] u2_col_out_14;
wire [15:0] u2_col_out_15;
wire [15:0] u2_col_out_16;
wire [15:0] u2_col_out_17;
wire [15:0] u2_col_out_18;
wire [15:0] u2_col_out_19;
wire [15:0] u2_col_out_20;
wire [15:0] u2_col_out_21;
wire [15:0] u2_col_out_22;
wire [15:0] u2_col_out_23;
wire [15:0] u2_col_out_24;
wire [15:0] u2_col_out_25;
wire [15:0] u2_col_out_26;
wire [15:0] u2_col_out_27;
wire [15:0] u2_col_out_28;
wire [15:0] u2_col_out_29;
wire [15:0] u2_col_out_30;
wire [15:0] u2_col_out_31;
wire [15:0] u2_col_out_32;
wire [15:0] u2_col_out_33;
wire [15:0] u2_col_out_34;
wire [15:0] u2_col_out_35;
wire [15:0] u2_col_out_36;
wire [15:0] u2_col_out_37;
wire [15:0] u2_col_out_38;
wire [15:0] u2_col_out_39;
wire [15:0] u2_col_out_40;
wire [15:0] u2_col_out_41;
wire [15:0] u2_col_out_42;
wire [15:0] u2_col_out_43;
wire [15:0] u2_col_out_44;
wire [15:0] u2_col_out_45;
wire [15:0] u2_col_out_46;
wire [15:0] u2_col_out_47;
wire [15:0] u2_col_out_48;
wire [15:0] u2_col_out_49;
wire [15:0] u2_col_out_50;
wire [15:0] u2_col_out_51;
wire [15:0] u2_col_out_52;
wire [15:0] u2_col_out_53;
wire [15:0] u2_col_out_54;
wire [15:0] u2_col_out_55;
wire [15:0] u2_col_out_56;
wire [15:0] u2_col_out_57;
wire [15:0] u2_col_out_58;
wire [15:0] u2_col_out_59;
wire [15:0] u2_col_out_60;
wire [15:0] u2_col_out_61;
wire [15:0] u2_col_out_62;
wire [15:0] u2_col_out_63;
wire [15:0] u2_col_out_64;
wire [15:0] u2_col_out_65;
wire [15:0] u2_col_out_66;
wire [15:0] u2_col_out_67;
wire [15:0] u2_col_out_68;
wire [15:0] u2_col_out_69;
wire [15:0] u2_col_out_70;
wire [15:0] u2_col_out_71;
wire [15:0] u2_col_out_72;
wire [15:0] u2_col_out_73;
wire [15:0] u2_col_out_74;
wire [15:0] u2_col_out_75;
wire [15:0] u2_col_out_76;
wire [15:0] u2_col_out_77;
wire [15:0] u2_col_out_78;
wire [15:0] u2_col_out_79;
wire [15:0] u2_col_out_80;
wire [15:0] u2_col_out_81;
wire [15:0] u2_col_out_82;
wire [15:0] u2_col_out_83;
wire [15:0] u2_col_out_84;
wire [15:0] u2_col_out_85;
wire [15:0] u2_col_out_86;
wire [15:0] u2_col_out_87;
wire [15:0] u2_col_out_88;
wire [15:0] u2_col_out_89;
wire [15:0] u2_col_out_90;
wire [15:0] u2_col_out_91;
wire [15:0] u2_col_out_92;
wire [15:0] u2_col_out_93;
wire [15:0] u2_col_out_94;
wire [15:0] u2_col_out_95;
wire [15:0] u2_col_out_96;
wire [15:0] u2_col_out_97;
wire [15:0] u2_col_out_98;
wire [15:0] u2_col_out_99;
wire [15:0] u2_col_out_100;
wire [15:0] u2_col_out_101;
wire [15:0] u2_col_out_102;
wire [15:0] u2_col_out_103;
wire [15:0] u2_col_out_104;
wire [15:0] u2_col_out_105;
wire [15:0] u2_col_out_106;
wire [15:0] u2_col_out_107;
wire [15:0] u2_col_out_108;
wire [15:0] u2_col_out_109;
wire [15:0] u2_col_out_110;
wire [15:0] u2_col_out_111;
wire [15:0] u2_col_out_112;
wire [15:0] u2_col_out_113;
wire [15:0] u2_col_out_114;
wire [15:0] u2_col_out_115;
wire [15:0] u2_col_out_116;
wire [15:0] u2_col_out_117;
wire [15:0] u2_col_out_118;
wire [15:0] u2_col_out_119;
wire [15:0] u2_col_out_120;
wire [15:0] u2_col_out_121;
wire [15:0] u2_col_out_122;
wire [15:0] u2_col_out_123;
wire [15:0] u2_col_out_124;
wire [15:0] u2_col_out_125;
wire [15:0] u2_col_out_126;
wire [15:0] u2_col_out_127;
wire [15:0] u2_col_out_128;
wire [15:0] u2_col_out_129;
wire [15:0] u2_col_out_130;
wire [15:0] u2_col_out_131;
wire [15:0] u2_col_out_132;
wire [15:0] u2_col_out_133;
wire [15:0] u2_col_out_134;
wire [15:0] u2_col_out_135;
wire [15:0] u2_col_out_136;
wire [15:0] u2_col_out_137;
wire [15:0] u2_col_out_138;
wire [15:0] u2_col_out_139;
wire [15:0] u2_col_out_140;
wire [15:0] u2_col_out_141;
wire [15:0] u2_col_out_142;
wire [15:0] u2_col_out_143;
wire [15:0] u2_col_out_144;
wire [15:0] u2_col_out_145;
wire [15:0] u2_col_out_146;
wire [15:0] u2_col_out_147;
wire [15:0] u2_col_out_148;
wire [15:0] u2_col_out_149;
wire [15:0] u2_col_out_150;
wire [15:0] u2_col_out_151;
wire [15:0] u2_col_out_152;
wire [15:0] u2_col_out_153;
wire [15:0] u2_col_out_154;
wire [15:0] u2_col_out_155;
wire [15:0] u2_col_out_156;
wire [15:0] u2_col_out_157;
wire [15:0] u2_col_out_158;
wire [15:0] u2_col_out_159;
wire [15:0] u2_col_out_160;
wire [15:0] u2_col_out_161;
wire [15:0] u2_col_out_162;
wire [15:0] u2_col_out_163;
wire [15:0] u2_col_out_164;
wire [15:0] u2_col_out_165;
wire [15:0] u2_col_out_166;
wire [15:0] u2_col_out_167;
wire [15:0] u2_col_out_168;
wire [15:0] u2_col_out_169;
wire [15:0] u2_col_out_170;
wire [15:0] u2_col_out_171;
wire [15:0] u2_col_out_172;
wire [15:0] u2_col_out_173;
wire [15:0] u2_col_out_174;
wire [15:0] u2_col_out_175;
wire [15:0] u2_col_out_176;
wire [15:0] u2_col_out_177;
wire [15:0] u2_col_out_178;
wire [15:0] u2_col_out_179;
wire [15:0] u2_col_out_180;
wire [15:0] u2_col_out_181;
wire [15:0] u2_col_out_182;
wire [15:0] u2_col_out_183;
wire [15:0] u2_col_out_184;
wire [15:0] u2_col_out_185;
wire [15:0] u2_col_out_186;
wire [15:0] u2_col_out_187;
wire [15:0] u2_col_out_188;
wire [15:0] u2_col_out_189;
wire [15:0] u2_col_out_190;
wire [15:0] u2_col_out_191;
wire [15:0] u2_col_out_192;
wire [15:0] u2_col_out_193;
wire [15:0] u2_col_out_194;
wire [15:0] u2_col_out_195;
wire [15:0] u2_col_out_196;
wire [15:0] u2_col_out_197;
wire [15:0] u2_col_out_198;
wire [15:0] u2_col_out_199;
wire [15:0] u2_col_out_200;
wire [15:0] u2_col_out_201;
wire [15:0] u2_col_out_202;
wire [15:0] u2_col_out_203;
wire [15:0] u2_col_out_204;
wire [15:0] u2_col_out_205;
wire [15:0] u2_col_out_206;
wire [15:0] u2_col_out_207;
wire [15:0] u2_col_out_208;
wire [15:0] u2_col_out_209;
wire [15:0] u2_col_out_210;
wire [15:0] u2_col_out_211;
wire [15:0] u2_col_out_212;
wire [15:0] u2_col_out_213;
wire [15:0] u2_col_out_214;
wire [15:0] u2_col_out_215;
wire [15:0] u2_col_out_216;
wire [15:0] u2_col_out_217;
wire [15:0] u2_col_out_218;
wire [15:0] u2_col_out_219;
wire [15:0] u2_col_out_220;
wire [15:0] u2_col_out_221;
wire [15:0] u2_col_out_222;
wire [15:0] u2_col_out_223;
wire [15:0] u2_col_out_224;
wire [15:0] u2_col_out_225;
wire [15:0] u2_col_out_226;
wire [15:0] u2_col_out_227;
wire [15:0] u2_col_out_228;
wire [15:0] u2_col_out_229;
wire [15:0] u2_col_out_230;
wire [15:0] u2_col_out_231;
wire [15:0] u2_col_out_232;
wire [15:0] u2_col_out_233;
wire [15:0] u2_col_out_234;
wire [15:0] u2_col_out_235;
wire [15:0] u2_col_out_236;
wire [15:0] u2_col_out_237;
wire [15:0] u2_col_out_238;
wire [15:0] u2_col_out_239;
wire [15:0] u2_col_out_240;
wire [15:0] u2_col_out_241;
wire [15:0] u2_col_out_242;
wire [15:0] u2_col_out_243;
wire [15:0] u2_col_out_244;
wire [15:0] u2_col_out_245;
wire [15:0] u2_col_out_246;
wire [15:0] u2_col_out_247;
wire [15:0] u2_col_out_248;
wire [15:0] u2_col_out_249;
wire [15:0] u2_col_out_250;
wire [15:0] u2_col_out_251;
wire [15:0] u2_col_out_252;
wire [15:0] u2_col_out_253;
wire [15:0] u2_col_out_254;
wire [15:0] u2_col_out_255;
wire [15:0] u2_col_out_256;
wire [15:0] u2_col_out_257;
wire [15:0] u2_col_out_258;
wire [15:0] u2_col_out_259;
wire [15:0] u2_col_out_260;
wire [15:0] u2_col_out_261;
wire [15:0] u2_col_out_262;
wire [15:0] u2_col_out_263;
wire [15:0] u2_col_out_264;
wire [15:0] u2_col_out_265;
wire [15:0] u2_col_out_266;
wire [15:0] u2_col_out_267;
wire [15:0] u2_col_out_268;
wire [15:0] u2_col_out_269;
wire [15:0] u2_col_out_270;
wire [15:0] u2_col_out_271;
wire [15:0] u2_col_out_272;
wire [15:0] u2_col_out_273;
wire [15:0] u2_col_out_274;
wire [15:0] u2_col_out_275;
wire [15:0] u2_col_out_276;
wire [15:0] u2_col_out_277;
wire [15:0] u2_col_out_278;
wire [15:0] u2_col_out_279;
wire [15:0] u2_col_out_280;
wire [15:0] u2_col_out_281;
wire [15:0] u2_col_out_282;
wire [15:0] u2_col_out_283;
wire [15:0] u2_col_out_284;
wire [15:0] u2_col_out_285;
wire [15:0] u2_col_out_286;
wire [15:0] u2_col_out_287;
wire [15:0] u2_col_out_288;
wire [15:0] u2_col_out_289;
wire [15:0] u2_col_out_290;
wire [15:0] u2_col_out_291;
wire [15:0] u2_col_out_292;
wire [15:0] u2_col_out_293;
wire [15:0] u2_col_out_294;
wire [15:0] u2_col_out_295;
wire [15:0] u2_col_out_296;
wire [15:0] u2_col_out_297;
wire [15:0] u2_col_out_298;
wire [15:0] u2_col_out_299;
wire [15:0] u2_col_out_300;
wire [15:0] u2_col_out_301;
wire [15:0] u2_col_out_302;
wire [15:0] u2_col_out_303;
wire [15:0] u2_col_out_304;
wire [15:0] u2_col_out_305;
wire [15:0] u2_col_out_306;
wire [15:0] u2_col_out_307;
wire [15:0] u2_col_out_308;
wire [15:0] u2_col_out_309;
wire [15:0] u2_col_out_310;
wire [15:0] u2_col_out_311;
wire [15:0] u2_col_out_312;
wire [15:0] u2_col_out_313;
wire [15:0] u2_col_out_314;
wire [15:0] u2_col_out_315;
wire [15:0] u2_col_out_316;
wire [15:0] u2_col_out_317;
wire [15:0] u2_col_out_318;
wire [15:0] u2_col_out_319;
wire [15:0] u2_col_out_320;
wire [15:0] u2_col_out_321;
wire [15:0] u2_col_out_322;
wire [15:0] u2_col_out_323;
wire [15:0] u2_col_out_324;
wire [15:0] u2_col_out_325;
wire [15:0] u2_col_out_326;
wire [15:0] u2_col_out_327;
wire [15:0] u2_col_out_328;
wire [15:0] u2_col_out_329;
wire [15:0] u2_col_out_330;
wire [15:0] u2_col_out_331;
wire [15:0] u2_col_out_332;
wire [15:0] u2_col_out_333;
wire [15:0] u2_col_out_334;
wire [15:0] u2_col_out_335;
wire [15:0] u2_col_out_336;
wire [15:0] u2_col_out_337;
wire [15:0] u2_col_out_338;
wire [15:0] u2_col_out_339;
wire [15:0] u2_col_out_340;
wire [15:0] u2_col_out_341;
wire [15:0] u2_col_out_342;
wire [15:0] u2_col_out_343;
wire [15:0] u2_col_out_344;
wire [15:0] u2_col_out_345;
wire [15:0] u2_col_out_346;
wire [15:0] u2_col_out_347;
wire [15:0] u2_col_out_348;
wire [15:0] u2_col_out_349;
wire [15:0] u2_col_out_350;
wire [15:0] u2_col_out_351;
wire [15:0] u2_col_out_352;
wire [15:0] u2_col_out_353;
wire [15:0] u2_col_out_354;
wire [15:0] u2_col_out_355;
wire [15:0] u2_col_out_356;
wire [15:0] u2_col_out_357;
wire [15:0] u2_col_out_358;
wire [15:0] u2_col_out_359;
wire [15:0] u2_col_out_360;
wire [15:0] u2_col_out_361;
wire [15:0] u2_col_out_362;
wire [15:0] u2_col_out_363;
wire [15:0] u2_col_out_364;
wire [15:0] u2_col_out_365;
wire [15:0] u2_col_out_366;
wire [15:0] u2_col_out_367;
wire [15:0] u2_col_out_368;
wire [15:0] u2_col_out_369;
wire [15:0] u2_col_out_370;
wire [15:0] u2_col_out_371;
wire [15:0] u2_col_out_372;
wire [15:0] u2_col_out_373;
wire [15:0] u2_col_out_374;
wire [15:0] u2_col_out_375;
wire [15:0] u2_col_out_376;
wire [15:0] u2_col_out_377;
wire [15:0] u2_col_out_378;
wire [15:0] u2_col_out_379;
wire [15:0] u2_col_out_380;
wire [15:0] u2_col_out_381;
wire [15:0] u2_col_out_382;
wire [15:0] u2_col_out_383;
wire [15:0] u2_col_out_384;
wire [15:0] u2_col_out_385;
wire [15:0] u2_col_out_386;
wire [15:0] u2_col_out_387;
wire [15:0] u2_col_out_388;
wire [15:0] u2_col_out_389;
wire [15:0] u2_col_out_390;
wire [15:0] u2_col_out_391;
wire [15:0] u2_col_out_392;
wire [15:0] u2_col_out_393;
wire [15:0] u2_col_out_394;
wire [15:0] u2_col_out_395;
wire [15:0] u2_col_out_396;
wire [15:0] u2_col_out_397;
wire [15:0] u2_col_out_398;
wire [15:0] u2_col_out_399;
wire [15:0] u2_col_out_400;
wire [15:0] u2_col_out_401;
wire [15:0] u2_col_out_402;
wire [15:0] u2_col_out_403;
wire [15:0] u2_col_out_404;
wire [15:0] u2_col_out_405;
wire [15:0] u2_col_out_406;
wire [15:0] u2_col_out_407;
wire [15:0] u2_col_out_408;
wire [15:0] u2_col_out_409;
wire [15:0] u2_col_out_410;
wire [15:0] u2_col_out_411;
wire [15:0] u2_col_out_412;
wire [15:0] u2_col_out_413;
wire [15:0] u2_col_out_414;
wire [15:0] u2_col_out_415;
wire [15:0] u2_col_out_416;
wire [15:0] u2_col_out_417;
wire [15:0] u2_col_out_418;
wire [15:0] u2_col_out_419;
wire [15:0] u2_col_out_420;
wire [15:0] u2_col_out_421;
wire [15:0] u2_col_out_422;
wire [15:0] u2_col_out_423;
wire [15:0] u2_col_out_424;
wire [15:0] u2_col_out_425;
wire [15:0] u2_col_out_426;
wire [15:0] u2_col_out_427;
wire [15:0] u2_col_out_428;
wire [15:0] u2_col_out_429;
wire [15:0] u2_col_out_430;
wire [15:0] u2_col_out_431;
wire [15:0] u2_col_out_432;
wire [15:0] u2_col_out_433;
wire [15:0] u2_col_out_434;
wire [15:0] u2_col_out_435;
wire [15:0] u2_col_out_436;
wire [15:0] u2_col_out_437;
wire [15:0] u2_col_out_438;
wire [15:0] u2_col_out_439;
wire [15:0] u2_col_out_440;
wire [15:0] u2_col_out_441;
wire [15:0] u2_col_out_442;
wire [15:0] u2_col_out_443;
wire [15:0] u2_col_out_444;
wire [15:0] u2_col_out_445;
wire [15:0] u2_col_out_446;
wire [15:0] u2_col_out_447;
wire [15:0] u2_col_out_448;
wire [15:0] u2_col_out_449;
wire [15:0] u2_col_out_450;
wire [15:0] u2_col_out_451;
wire [15:0] u2_col_out_452;
wire [15:0] u2_col_out_453;
wire [15:0] u2_col_out_454;
wire [15:0] u2_col_out_455;
wire [15:0] u2_col_out_456;
wire [15:0] u2_col_out_457;
wire [15:0] u2_col_out_458;
wire [15:0] u2_col_out_459;
wire [15:0] u2_col_out_460;
wire [15:0] u2_col_out_461;
wire [15:0] u2_col_out_462;
wire [15:0] u2_col_out_463;
wire [15:0] u2_col_out_464;
wire [15:0] u2_col_out_465;
wire [15:0] u2_col_out_466;
wire [15:0] u2_col_out_467;
wire [15:0] u2_col_out_468;
wire [15:0] u2_col_out_469;
wire [15:0] u2_col_out_470;
wire [15:0] u2_col_out_471;
wire [15:0] u2_col_out_472;
wire [15:0] u2_col_out_473;
wire [15:0] u2_col_out_474;
wire [15:0] u2_col_out_475;
wire [15:0] u2_col_out_476;
wire [15:0] u2_col_out_477;
wire [15:0] u2_col_out_478;
wire [15:0] u2_col_out_479;
wire [15:0] u2_col_out_480;
wire [15:0] u2_col_out_481;
wire [15:0] u2_col_out_482;
wire [15:0] u2_col_out_483;
wire [15:0] u2_col_out_484;
wire [15:0] u2_col_out_485;
wire [15:0] u2_col_out_486;
wire [15:0] u2_col_out_487;
wire [15:0] u2_col_out_488;
wire [15:0] u2_col_out_489;
wire [15:0] u2_col_out_490;
wire [15:0] u2_col_out_491;
wire [15:0] u2_col_out_492;
wire [15:0] u2_col_out_493;
wire [15:0] u2_col_out_494;
wire [15:0] u2_col_out_495;
wire [15:0] u2_col_out_496;
wire [15:0] u2_col_out_497;
wire [15:0] u2_col_out_498;
wire [15:0] u2_col_out_499;
wire [15:0] u2_col_out_500;
wire [15:0] u2_col_out_501;
wire [15:0] u2_col_out_502;
wire [15:0] u2_col_out_503;
wire [15:0] u2_col_out_504;
wire [15:0] u2_col_out_505;
wire [15:0] u2_col_out_506;
wire [15:0] u2_col_out_507;
wire [15:0] u2_col_out_508;
wire [15:0] u2_col_out_509;
wire [15:0] u2_col_out_510;
wire [15:0] u2_col_out_511;
wire [15:0] u2_col_out_512;
wire [15:0] u2_col_out_513;
wire [15:0] u2_col_out_514;
wire [15:0] u2_col_out_515;
wire [15:0] u2_col_out_516;
wire [15:0] u2_col_out_517;
wire [15:0] u2_col_out_518;
wire [15:0] u2_col_out_519;
wire [15:0] u2_col_out_520;
wire [15:0] u2_col_out_521;
wire [15:0] u2_col_out_522;
wire [15:0] u2_col_out_523;
wire [15:0] u2_col_out_524;
wire [15:0] u2_col_out_525;
wire [15:0] u2_col_out_526;
wire [15:0] u2_col_out_527;
wire [15:0] u2_col_out_528;
wire [15:0] u2_col_out_529;
wire [15:0] u2_col_out_530;
wire [15:0] u2_col_out_531;
wire [15:0] u2_col_out_532;
wire [15:0] u2_col_out_533;
wire [15:0] u2_col_out_534;
wire [15:0] u2_col_out_535;
wire [15:0] u2_col_out_536;
wire [15:0] u2_col_out_537;
wire [15:0] u2_col_out_538;
wire [15:0] u2_col_out_539;
wire [15:0] u2_col_out_540;
wire [15:0] u2_col_out_541;
wire [15:0] u2_col_out_542;
wire [15:0] u2_col_out_543;
wire [15:0] u2_col_out_544;
wire [15:0] u2_col_out_545;
wire [15:0] u2_col_out_546;
wire [15:0] u2_col_out_547;
wire [15:0] u2_col_out_548;
wire [15:0] u2_col_out_549;
wire [15:0] u2_col_out_550;
wire [15:0] u2_col_out_551;
wire [15:0] u2_col_out_552;
wire [15:0] u2_col_out_553;
wire [15:0] u2_col_out_554;
wire [15:0] u2_col_out_555;
wire [15:0] u2_col_out_556;
wire [15:0] u2_col_out_557;
wire [15:0] u2_col_out_558;
wire [15:0] u2_col_out_559;
wire [15:0] u2_col_out_560;
wire [15:0] u2_col_out_561;
wire [15:0] u2_col_out_562;
wire [15:0] u2_col_out_563;
wire [15:0] u2_col_out_564;
wire [15:0] u2_col_out_565;
wire [15:0] u2_col_out_566;
wire [15:0] u2_col_out_567;
wire [15:0] u2_col_out_568;
wire [15:0] u2_col_out_569;
wire [15:0] u2_col_out_570;
wire [15:0] u2_col_out_571;
wire [15:0] u2_col_out_572;
wire [15:0] u2_col_out_573;
wire [15:0] u2_col_out_574;
wire [15:0] u2_col_out_575;
wire [15:0] u2_col_out_576;
wire [15:0] u2_col_out_577;
wire [15:0] u2_col_out_578;
wire [15:0] u2_col_out_579;
wire [15:0] u2_col_out_580;
wire [15:0] u2_col_out_581;
wire [15:0] u2_col_out_582;
wire [15:0] u2_col_out_583;
wire [15:0] u2_col_out_584;
wire [15:0] u2_col_out_585;
wire [15:0] u2_col_out_586;
wire [15:0] u2_col_out_587;
wire [15:0] u2_col_out_588;
wire [15:0] u2_col_out_589;
wire [15:0] u2_col_out_590;
wire [15:0] u2_col_out_591;
wire [15:0] u2_col_out_592;
wire [15:0] u2_col_out_593;
wire [15:0] u2_col_out_594;
wire [15:0] u2_col_out_595;
wire [15:0] u2_col_out_596;
wire [15:0] u2_col_out_597;
wire [15:0] u2_col_out_598;
wire [15:0] u2_col_out_599;
wire [15:0] u2_col_out_600;
wire [15:0] u2_col_out_601;
wire [15:0] u2_col_out_602;
wire [15:0] u2_col_out_603;
wire [15:0] u2_col_out_604;
wire [15:0] u2_col_out_605;
wire [15:0] u2_col_out_606;
wire [15:0] u2_col_out_607;
wire [15:0] u2_col_out_608;
wire [15:0] u2_col_out_609;
wire [15:0] u2_col_out_610;
wire [15:0] u2_col_out_611;
wire [15:0] u2_col_out_612;
wire [15:0] u2_col_out_613;
wire [15:0] u2_col_out_614;
wire [15:0] u2_col_out_615;
wire [15:0] u2_col_out_616;
wire [15:0] u2_col_out_617;
wire [15:0] u2_col_out_618;
wire [15:0] u2_col_out_619;
wire [15:0] u2_col_out_620;
wire [15:0] u2_col_out_621;
wire [15:0] u2_col_out_622;
wire [15:0] u2_col_out_623;
wire [15:0] u2_col_out_624;
wire [15:0] u2_col_out_625;
wire [15:0] u2_col_out_626;
wire [15:0] u2_col_out_627;
wire [15:0] u2_col_out_628;
wire [15:0] u2_col_out_629;
wire [15:0] u2_col_out_630;
wire [15:0] u2_col_out_631;
wire [15:0] u2_col_out_632;
wire [15:0] u2_col_out_633;
wire [15:0] u2_col_out_634;
wire [15:0] u2_col_out_635;
wire [15:0] u2_col_out_636;
wire [15:0] u2_col_out_637;
wire [15:0] u2_col_out_638;
wire [15:0] u2_col_out_639;
wire [15:0] u2_col_out_640;
wire [15:0] u2_col_out_641;
wire [15:0] u2_col_out_642;
wire [15:0] u2_col_out_643;
wire [15:0] u2_col_out_644;
wire [15:0] u2_col_out_645;
wire [15:0] u2_col_out_646;
wire [15:0] u2_col_out_647;
wire [15:0] u2_col_out_648;
wire [15:0] u2_col_out_649;
wire [15:0] u2_col_out_650;
wire [15:0] u2_col_out_651;
wire [15:0] u2_col_out_652;
wire [15:0] u2_col_out_653;
wire [15:0] u2_col_out_654;
wire [15:0] u2_col_out_655;
wire [15:0] u2_col_out_656;
wire [15:0] u2_col_out_657;
wire [15:0] u2_col_out_658;
wire [15:0] u2_col_out_659;
wire [15:0] u2_col_out_660;
wire [15:0] u2_col_out_661;
wire [15:0] u2_col_out_662;
wire [15:0] u2_col_out_663;
wire [15:0] u2_col_out_664;
wire [15:0] u2_col_out_665;
wire [15:0] u2_col_out_666;
wire [15:0] u2_col_out_667;
wire [15:0] u2_col_out_668;
wire [15:0] u2_col_out_669;
wire [15:0] u2_col_out_670;
wire [15:0] u2_col_out_671;
wire [15:0] u2_col_out_672;
wire [15:0] u2_col_out_673;
wire [15:0] u2_col_out_674;
wire [15:0] u2_col_out_675;
wire [15:0] u2_col_out_676;
wire [15:0] u2_col_out_677;
wire [15:0] u2_col_out_678;
wire [15:0] u2_col_out_679;
wire [15:0] u2_col_out_680;
wire [15:0] u2_col_out_681;
wire [15:0] u2_col_out_682;
wire [15:0] u2_col_out_683;
wire [15:0] u2_col_out_684;
wire [15:0] u2_col_out_685;
wire [15:0] u2_col_out_686;
wire [15:0] u2_col_out_687;
wire [15:0] u2_col_out_688;
wire [15:0] u2_col_out_689;
wire [15:0] u2_col_out_690;
wire [15:0] u2_col_out_691;
wire [15:0] u2_col_out_692;
wire [15:0] u2_col_out_693;
wire [15:0] u2_col_out_694;
wire [15:0] u2_col_out_695;
wire [15:0] u2_col_out_696;
wire [15:0] u2_col_out_697;
wire [15:0] u2_col_out_698;
wire [15:0] u2_col_out_699;
wire [15:0] u2_col_out_700;
wire [15:0] u2_col_out_701;
wire [15:0] u2_col_out_702;
wire [15:0] u2_col_out_703;
wire [15:0] u2_col_out_704;
wire [15:0] u2_col_out_705;
wire [15:0] u2_col_out_706;
wire [15:0] u2_col_out_707;
wire [15:0] u2_col_out_708;
wire [15:0] u2_col_out_709;
wire [15:0] u2_col_out_710;
wire [15:0] u2_col_out_711;
wire [15:0] u2_col_out_712;
wire [15:0] u2_col_out_713;
wire [15:0] u2_col_out_714;
wire [15:0] u2_col_out_715;
wire [15:0] u2_col_out_716;
wire [15:0] u2_col_out_717;
wire [15:0] u2_col_out_718;
wire [15:0] u2_col_out_719;
wire [15:0] u2_col_out_720;
wire [15:0] u2_col_out_721;
wire [15:0] u2_col_out_722;
wire [15:0] u2_col_out_723;
wire [15:0] u2_col_out_724;
wire [15:0] u2_col_out_725;
wire [15:0] u2_col_out_726;
wire [15:0] u2_col_out_727;
wire [15:0] u2_col_out_728;
wire [15:0] u2_col_out_729;
wire [15:0] u2_col_out_730;
wire [15:0] u2_col_out_731;
wire [15:0] u2_col_out_732;
wire [15:0] u2_col_out_733;
wire [15:0] u2_col_out_734;
wire [15:0] u2_col_out_735;
wire [15:0] u2_col_out_736;
wire [15:0] u2_col_out_737;
wire [15:0] u2_col_out_738;
wire [15:0] u2_col_out_739;
wire [15:0] u2_col_out_740;
wire [15:0] u2_col_out_741;
wire [15:0] u2_col_out_742;
wire [15:0] u2_col_out_743;
wire [15:0] u2_col_out_744;
wire [15:0] u2_col_out_745;
wire [15:0] u2_col_out_746;
wire [15:0] u2_col_out_747;
wire [15:0] u2_col_out_748;
wire [15:0] u2_col_out_749;
wire [15:0] u2_col_out_750;
wire [15:0] u2_col_out_751;
wire [15:0] u2_col_out_752;
wire [15:0] u2_col_out_753;
wire [15:0] u2_col_out_754;
wire [15:0] u2_col_out_755;
wire [15:0] u2_col_out_756;
wire [15:0] u2_col_out_757;
wire [15:0] u2_col_out_758;
wire [15:0] u2_col_out_759;
wire [15:0] u2_col_out_760;
wire [15:0] u2_col_out_761;
wire [15:0] u2_col_out_762;
wire [15:0] u2_col_out_763;
wire [15:0] u2_col_out_764;
wire [15:0] u2_col_out_765;
wire [15:0] u2_col_out_766;
wire [15:0] u2_col_out_767;
wire [15:0] u2_col_out_768;
wire [15:0] u2_col_out_769;
wire [15:0] u2_col_out_770;
wire [15:0] u2_col_out_771;
wire [15:0] u2_col_out_772;
wire [15:0] u2_col_out_773;
wire [15:0] u2_col_out_774;
wire [15:0] u2_col_out_775;
wire [15:0] u2_col_out_776;
wire [15:0] u2_col_out_777;
wire [15:0] u2_col_out_778;
wire [15:0] u2_col_out_779;
wire [15:0] u2_col_out_780;
wire [15:0] u2_col_out_781;
wire [15:0] u2_col_out_782;
wire [15:0] u2_col_out_783;
wire [15:0] u2_col_out_784;
wire [15:0] u2_col_out_785;
wire [15:0] u2_col_out_786;
wire [15:0] u2_col_out_787;
wire [15:0] u2_col_out_788;
wire [15:0] u2_col_out_789;
wire [15:0] u2_col_out_790;
wire [15:0] u2_col_out_791;
wire [15:0] u2_col_out_792;
wire [15:0] u2_col_out_793;
wire [15:0] u2_col_out_794;
wire [15:0] u2_col_out_795;
wire [15:0] u2_col_out_796;
wire [15:0] u2_col_out_797;
wire [15:0] u2_col_out_798;
wire [15:0] u2_col_out_799;
wire [15:0] u2_col_out_800;
wire [15:0] u2_col_out_801;
wire [15:0] u2_col_out_802;
wire [15:0] u2_col_out_803;
wire [15:0] u2_col_out_804;
wire [15:0] u2_col_out_805;
wire [15:0] u2_col_out_806;
wire [15:0] u2_col_out_807;
wire [15:0] u2_col_out_808;
wire [15:0] u2_col_out_809;
wire [15:0] u2_col_out_810;
wire [15:0] u2_col_out_811;
wire [15:0] u2_col_out_812;
wire [15:0] u2_col_out_813;
wire [15:0] u2_col_out_814;
wire [15:0] u2_col_out_815;
wire [15:0] u2_col_out_816;
wire [15:0] u2_col_out_817;
wire [15:0] u2_col_out_818;
wire [15:0] u2_col_out_819;
wire [15:0] u2_col_out_820;
wire [15:0] u2_col_out_821;
wire [15:0] u2_col_out_822;
wire [15:0] u2_col_out_823;
wire [15:0] u2_col_out_824;
wire [15:0] u2_col_out_825;
wire [15:0] u2_col_out_826;
wire [15:0] u2_col_out_827;
wire [15:0] u2_col_out_828;
wire [15:0] u2_col_out_829;
wire [15:0] u2_col_out_830;
wire [15:0] u2_col_out_831;
wire [15:0] u2_col_out_832;
wire [15:0] u2_col_out_833;
wire [15:0] u2_col_out_834;
wire [15:0] u2_col_out_835;
wire [15:0] u2_col_out_836;
wire [15:0] u2_col_out_837;
wire [15:0] u2_col_out_838;
wire [15:0] u2_col_out_839;
wire [15:0] u2_col_out_840;
wire [15:0] u2_col_out_841;
wire [15:0] u2_col_out_842;
wire [15:0] u2_col_out_843;
wire [15:0] u2_col_out_844;
wire [15:0] u2_col_out_845;
wire [15:0] u2_col_out_846;
wire [15:0] u2_col_out_847;
wire [15:0] u2_col_out_848;
wire [15:0] u2_col_out_849;
wire [15:0] u2_col_out_850;
wire [15:0] u2_col_out_851;
wire [15:0] u2_col_out_852;
wire [15:0] u2_col_out_853;
wire [15:0] u2_col_out_854;
wire [15:0] u2_col_out_855;
wire [15:0] u2_col_out_856;
wire [15:0] u2_col_out_857;
wire [15:0] u2_col_out_858;
wire [15:0] u2_col_out_859;
wire [15:0] u2_col_out_860;
wire [15:0] u2_col_out_861;
wire [15:0] u2_col_out_862;
wire [15:0] u2_col_out_863;
wire [15:0] u2_col_out_864;
wire [15:0] u2_col_out_865;
wire [15:0] u2_col_out_866;
wire [15:0] u2_col_out_867;
wire [15:0] u2_col_out_868;
wire [15:0] u2_col_out_869;
wire [15:0] u2_col_out_870;
wire [15:0] u2_col_out_871;
wire [15:0] u2_col_out_872;
wire [15:0] u2_col_out_873;
wire [15:0] u2_col_out_874;
wire [15:0] u2_col_out_875;
wire [15:0] u2_col_out_876;
wire [15:0] u2_col_out_877;
wire [15:0] u2_col_out_878;
wire [15:0] u2_col_out_879;
wire [15:0] u2_col_out_880;
wire [15:0] u2_col_out_881;
wire [15:0] u2_col_out_882;
wire [15:0] u2_col_out_883;
wire [15:0] u2_col_out_884;
wire [15:0] u2_col_out_885;
wire [15:0] u2_col_out_886;
wire [15:0] u2_col_out_887;
wire [15:0] u2_col_out_888;
wire [15:0] u2_col_out_889;
wire [15:0] u2_col_out_890;
wire [15:0] u2_col_out_891;
wire [15:0] u2_col_out_892;
wire [15:0] u2_col_out_893;
wire [15:0] u2_col_out_894;
wire [15:0] u2_col_out_895;
wire [15:0] u2_col_out_896;
wire [15:0] u2_col_out_897;
wire [15:0] u2_col_out_898;
wire [15:0] u2_col_out_899;
wire [15:0] u2_col_out_900;
wire [15:0] u2_col_out_901;
wire [15:0] u2_col_out_902;
wire [15:0] u2_col_out_903;
wire [15:0] u2_col_out_904;
wire [15:0] u2_col_out_905;
wire [15:0] u2_col_out_906;
wire [15:0] u2_col_out_907;
wire [15:0] u2_col_out_908;
wire [15:0] u2_col_out_909;
wire [15:0] u2_col_out_910;
wire [15:0] u2_col_out_911;
wire [15:0] u2_col_out_912;
wire [15:0] u2_col_out_913;
wire [15:0] u2_col_out_914;
wire [15:0] u2_col_out_915;
wire [15:0] u2_col_out_916;
wire [15:0] u2_col_out_917;
wire [15:0] u2_col_out_918;
wire [15:0] u2_col_out_919;
wire [15:0] u2_col_out_920;
wire [15:0] u2_col_out_921;
wire [15:0] u2_col_out_922;
wire [15:0] u2_col_out_923;
wire [15:0] u2_col_out_924;
wire [15:0] u2_col_out_925;
wire [15:0] u2_col_out_926;
wire [15:0] u2_col_out_927;
wire [15:0] u2_col_out_928;
wire [15:0] u2_col_out_929;
wire [15:0] u2_col_out_930;
wire [15:0] u2_col_out_931;
wire [15:0] u2_col_out_932;
wire [15:0] u2_col_out_933;
wire [15:0] u2_col_out_934;
wire [15:0] u2_col_out_935;
wire [15:0] u2_col_out_936;
wire [15:0] u2_col_out_937;
wire [15:0] u2_col_out_938;
wire [15:0] u2_col_out_939;
wire [15:0] u2_col_out_940;
wire [15:0] u2_col_out_941;
wire [15:0] u2_col_out_942;
wire [15:0] u2_col_out_943;
wire [15:0] u2_col_out_944;
wire [15:0] u2_col_out_945;
wire [15:0] u2_col_out_946;
wire [15:0] u2_col_out_947;
wire [15:0] u2_col_out_948;
wire [15:0] u2_col_out_949;
wire [15:0] u2_col_out_950;
wire [15:0] u2_col_out_951;
wire [15:0] u2_col_out_952;
wire [15:0] u2_col_out_953;
wire [15:0] u2_col_out_954;
wire [15:0] u2_col_out_955;
wire [15:0] u2_col_out_956;
wire [15:0] u2_col_out_957;
wire [15:0] u2_col_out_958;
wire [15:0] u2_col_out_959;
wire [15:0] u2_col_out_960;
wire [15:0] u2_col_out_961;
wire [15:0] u2_col_out_962;
wire [15:0] u2_col_out_963;
wire [15:0] u2_col_out_964;
wire [15:0] u2_col_out_965;
wire [15:0] u2_col_out_966;
wire [15:0] u2_col_out_967;
wire [15:0] u2_col_out_968;
wire [15:0] u2_col_out_969;
wire [15:0] u2_col_out_970;
wire [15:0] u2_col_out_971;
wire [15:0] u2_col_out_972;
wire [15:0] u2_col_out_973;
wire [15:0] u2_col_out_974;
wire [15:0] u2_col_out_975;
wire [15:0] u2_col_out_976;
wire [15:0] u2_col_out_977;
wire [15:0] u2_col_out_978;
wire [15:0] u2_col_out_979;
wire [15:0] u2_col_out_980;
wire [15:0] u2_col_out_981;
wire [15:0] u2_col_out_982;
wire [15:0] u2_col_out_983;
wire [15:0] u2_col_out_984;
wire [15:0] u2_col_out_985;
wire [15:0] u2_col_out_986;
wire [15:0] u2_col_out_987;
wire [15:0] u2_col_out_988;
wire [15:0] u2_col_out_989;
wire [15:0] u2_col_out_990;
wire [15:0] u2_col_out_991;
wire [15:0] u2_col_out_992;
wire [15:0] u2_col_out_993;
wire [15:0] u2_col_out_994;
wire [15:0] u2_col_out_995;
wire [15:0] u2_col_out_996;
wire [15:0] u2_col_out_997;
wire [15:0] u2_col_out_998;
wire [15:0] u2_col_out_999;
wire [15:0] u2_col_out_1000;
wire [15:0] u2_col_out_1001;
wire [15:0] u2_col_out_1002;
wire [15:0] u2_col_out_1003;
wire [15:0] u2_col_out_1004;
wire [15:0] u2_col_out_1005;
wire [15:0] u2_col_out_1006;
wire [15:0] u2_col_out_1007;
wire [15:0] u2_col_out_1008;
wire [15:0] u2_col_out_1009;
wire [15:0] u2_col_out_1010;
wire [15:0] u2_col_out_1011;
wire [15:0] u2_col_out_1012;
wire [15:0] u2_col_out_1013;
wire [15:0] u2_col_out_1014;
wire [15:0] u2_col_out_1015;
wire [15:0] u2_col_out_1016;
wire [15:0] u2_col_out_1017;
wire [15:0] u2_col_out_1018;
wire [15:0] u2_col_out_1019;
wire [15:0] u2_col_out_1020;
wire [15:0] u2_col_out_1021;
wire [15:0] u2_col_out_1022;
wire [15:0] u2_col_out_1023;
wire [15:0] u2_col_out_1024;
wire [15:0] u2_col_out_1025;
wire [15:0] u2_col_out_1026;
wire [15:0] u2_col_out_1027;
wire [15:0] u2_col_out_1028;
wire [15:0] u2_col_out_1029;
wire [15:0] u2_col_out_1030;
wire [15:0] u2_col_out_1031;
wire [15:0] u2_col_out_1032;




//*****************************************************
//**************u2输入赋值******************************
//*****************************************************
assign u2_col_in_0 = u1_col_out_0;
assign u2_col_in_1 = u1_col_out_1;
assign u2_col_in_2 = u1_col_out_2;
assign u2_col_in_3 = u1_col_out_3;
assign u2_col_in_4 = u1_col_out_4;
assign u2_col_in_5 = u1_col_out_5;
assign u2_col_in_6 = u1_col_out_6;
assign u2_col_in_7 = u1_col_out_7;
assign u2_col_in_8 = u1_col_out_8;
assign u2_col_in_9 = u1_col_out_9;
assign u2_col_in_10 = u1_col_out_10;
assign u2_col_in_11 = u1_col_out_11;
assign u2_col_in_12 = u1_col_out_12;
assign u2_col_in_13 = u1_col_out_13;
assign u2_col_in_14 = u1_col_out_14;
assign u2_col_in_15 = u1_col_out_15;
assign u2_col_in_16 = u1_col_out_16;
assign u2_col_in_17 = u1_col_out_17;
assign u2_col_in_18 = u1_col_out_18;
assign u2_col_in_19 = u1_col_out_19;
assign u2_col_in_20 = u1_col_out_20;
assign u2_col_in_21 = u1_col_out_21;
assign u2_col_in_22 = u1_col_out_22;
assign u2_col_in_23 = u1_col_out_23;
assign u2_col_in_24 = u1_col_out_24;
assign u2_col_in_25 = u1_col_out_25;
assign u2_col_in_26 = u1_col_out_26;
assign u2_col_in_27 = u1_col_out_27;
assign u2_col_in_28 = u1_col_out_28;
assign u2_col_in_29 = u1_col_out_29;
assign u2_col_in_30 = u1_col_out_30;
assign u2_col_in_31 = u1_col_out_31;
assign u2_col_in_32 = u1_col_out_32;
assign u2_col_in_33 = u1_col_out_33;
assign u2_col_in_34 = u1_col_out_34;
assign u2_col_in_35 = u1_col_out_35;
assign u2_col_in_36 = u1_col_out_36;
assign u2_col_in_37 = u1_col_out_37;
assign u2_col_in_38 = u1_col_out_38;
assign u2_col_in_39 = u1_col_out_39;
assign u2_col_in_40 = u1_col_out_40;
assign u2_col_in_41 = u1_col_out_41;
assign u2_col_in_42 = u1_col_out_42;
assign u2_col_in_43 = u1_col_out_43;
assign u2_col_in_44 = u1_col_out_44;
assign u2_col_in_45 = u1_col_out_45;
assign u2_col_in_46 = u1_col_out_46;
assign u2_col_in_47 = u1_col_out_47;
assign u2_col_in_48 = u1_col_out_48;
assign u2_col_in_49 = u1_col_out_49;
assign u2_col_in_50 = u1_col_out_50;
assign u2_col_in_51 = u1_col_out_51;
assign u2_col_in_52 = u1_col_out_52;
assign u2_col_in_53 = u1_col_out_53;
assign u2_col_in_54 = u1_col_out_54;
assign u2_col_in_55 = u1_col_out_55;
assign u2_col_in_56 = u1_col_out_56;
assign u2_col_in_57 = u1_col_out_57;
assign u2_col_in_58 = u1_col_out_58;
assign u2_col_in_59 = u1_col_out_59;
assign u2_col_in_60 = u1_col_out_60;
assign u2_col_in_61 = u1_col_out_61;
assign u2_col_in_62 = u1_col_out_62;
assign u2_col_in_63 = u1_col_out_63;
assign u2_col_in_64 = u1_col_out_64;
assign u2_col_in_65 = u1_col_out_65;
assign u2_col_in_66 = u1_col_out_66;
assign u2_col_in_67 = u1_col_out_67;
assign u2_col_in_68 = u1_col_out_68;
assign u2_col_in_69 = u1_col_out_69;
assign u2_col_in_70 = u1_col_out_70;
assign u2_col_in_71 = u1_col_out_71;
assign u2_col_in_72 = u1_col_out_72;
assign u2_col_in_73 = u1_col_out_73;
assign u2_col_in_74 = u1_col_out_74;
assign u2_col_in_75 = u1_col_out_75;
assign u2_col_in_76 = u1_col_out_76;
assign u2_col_in_77 = u1_col_out_77;
assign u2_col_in_78 = u1_col_out_78;
assign u2_col_in_79 = u1_col_out_79;
assign u2_col_in_80 = u1_col_out_80;
assign u2_col_in_81 = u1_col_out_81;
assign u2_col_in_82 = u1_col_out_82;
assign u2_col_in_83 = u1_col_out_83;
assign u2_col_in_84 = u1_col_out_84;
assign u2_col_in_85 = u1_col_out_85;
assign u2_col_in_86 = u1_col_out_86;
assign u2_col_in_87 = u1_col_out_87;
assign u2_col_in_88 = u1_col_out_88;
assign u2_col_in_89 = u1_col_out_89;
assign u2_col_in_90 = u1_col_out_90;
assign u2_col_in_91 = u1_col_out_91;
assign u2_col_in_92 = u1_col_out_92;
assign u2_col_in_93 = u1_col_out_93;
assign u2_col_in_94 = u1_col_out_94;
assign u2_col_in_95 = u1_col_out_95;
assign u2_col_in_96 = u1_col_out_96;
assign u2_col_in_97 = u1_col_out_97;
assign u2_col_in_98 = u1_col_out_98;
assign u2_col_in_99 = u1_col_out_99;
assign u2_col_in_100 = u1_col_out_100;
assign u2_col_in_101 = u1_col_out_101;
assign u2_col_in_102 = u1_col_out_102;
assign u2_col_in_103 = u1_col_out_103;
assign u2_col_in_104 = u1_col_out_104;
assign u2_col_in_105 = u1_col_out_105;
assign u2_col_in_106 = u1_col_out_106;
assign u2_col_in_107 = u1_col_out_107;
assign u2_col_in_108 = u1_col_out_108;
assign u2_col_in_109 = u1_col_out_109;
assign u2_col_in_110 = u1_col_out_110;
assign u2_col_in_111 = u1_col_out_111;
assign u2_col_in_112 = u1_col_out_112;
assign u2_col_in_113 = u1_col_out_113;
assign u2_col_in_114 = u1_col_out_114;
assign u2_col_in_115 = u1_col_out_115;
assign u2_col_in_116 = u1_col_out_116;
assign u2_col_in_117 = u1_col_out_117;
assign u2_col_in_118 = u1_col_out_118;
assign u2_col_in_119 = u1_col_out_119;
assign u2_col_in_120 = u1_col_out_120;
assign u2_col_in_121 = u1_col_out_121;
assign u2_col_in_122 = u1_col_out_122;
assign u2_col_in_123 = u1_col_out_123;
assign u2_col_in_124 = u1_col_out_124;
assign u2_col_in_125 = u1_col_out_125;
assign u2_col_in_126 = u1_col_out_126;
assign u2_col_in_127 = u1_col_out_127;
assign u2_col_in_128 = u1_col_out_128;
assign u2_col_in_129 = u1_col_out_129;
assign u2_col_in_130 = u1_col_out_130;
assign u2_col_in_131 = u1_col_out_131;
assign u2_col_in_132 = u1_col_out_132;
assign u2_col_in_133 = u1_col_out_133;
assign u2_col_in_134 = u1_col_out_134;
assign u2_col_in_135 = u1_col_out_135;
assign u2_col_in_136 = u1_col_out_136;
assign u2_col_in_137 = u1_col_out_137;
assign u2_col_in_138 = u1_col_out_138;
assign u2_col_in_139 = u1_col_out_139;
assign u2_col_in_140 = u1_col_out_140;
assign u2_col_in_141 = u1_col_out_141;
assign u2_col_in_142 = u1_col_out_142;
assign u2_col_in_143 = u1_col_out_143;
assign u2_col_in_144 = u1_col_out_144;
assign u2_col_in_145 = u1_col_out_145;
assign u2_col_in_146 = u1_col_out_146;
assign u2_col_in_147 = u1_col_out_147;
assign u2_col_in_148 = u1_col_out_148;
assign u2_col_in_149 = u1_col_out_149;
assign u2_col_in_150 = u1_col_out_150;
assign u2_col_in_151 = u1_col_out_151;
assign u2_col_in_152 = u1_col_out_152;
assign u2_col_in_153 = u1_col_out_153;
assign u2_col_in_154 = u1_col_out_154;
assign u2_col_in_155 = u1_col_out_155;
assign u2_col_in_156 = u1_col_out_156;
assign u2_col_in_157 = u1_col_out_157;
assign u2_col_in_158 = u1_col_out_158;
assign u2_col_in_159 = u1_col_out_159;
assign u2_col_in_160 = u1_col_out_160;
assign u2_col_in_161 = u1_col_out_161;
assign u2_col_in_162 = u1_col_out_162;
assign u2_col_in_163 = u1_col_out_163;
assign u2_col_in_164 = u1_col_out_164;
assign u2_col_in_165 = u1_col_out_165;
assign u2_col_in_166 = u1_col_out_166;
assign u2_col_in_167 = u1_col_out_167;
assign u2_col_in_168 = u1_col_out_168;
assign u2_col_in_169 = u1_col_out_169;
assign u2_col_in_170 = u1_col_out_170;
assign u2_col_in_171 = u1_col_out_171;
assign u2_col_in_172 = u1_col_out_172;
assign u2_col_in_173 = u1_col_out_173;
assign u2_col_in_174 = u1_col_out_174;
assign u2_col_in_175 = u1_col_out_175;
assign u2_col_in_176 = u1_col_out_176;
assign u2_col_in_177 = u1_col_out_177;
assign u2_col_in_178 = u1_col_out_178;
assign u2_col_in_179 = u1_col_out_179;
assign u2_col_in_180 = u1_col_out_180;
assign u2_col_in_181 = u1_col_out_181;
assign u2_col_in_182 = u1_col_out_182;
assign u2_col_in_183 = u1_col_out_183;
assign u2_col_in_184 = u1_col_out_184;
assign u2_col_in_185 = u1_col_out_185;
assign u2_col_in_186 = u1_col_out_186;
assign u2_col_in_187 = u1_col_out_187;
assign u2_col_in_188 = u1_col_out_188;
assign u2_col_in_189 = u1_col_out_189;
assign u2_col_in_190 = u1_col_out_190;
assign u2_col_in_191 = u1_col_out_191;
assign u2_col_in_192 = u1_col_out_192;
assign u2_col_in_193 = u1_col_out_193;
assign u2_col_in_194 = u1_col_out_194;
assign u2_col_in_195 = u1_col_out_195;
assign u2_col_in_196 = u1_col_out_196;
assign u2_col_in_197 = u1_col_out_197;
assign u2_col_in_198 = u1_col_out_198;
assign u2_col_in_199 = u1_col_out_199;
assign u2_col_in_200 = u1_col_out_200;
assign u2_col_in_201 = u1_col_out_201;
assign u2_col_in_202 = u1_col_out_202;
assign u2_col_in_203 = u1_col_out_203;
assign u2_col_in_204 = u1_col_out_204;
assign u2_col_in_205 = u1_col_out_205;
assign u2_col_in_206 = u1_col_out_206;
assign u2_col_in_207 = u1_col_out_207;
assign u2_col_in_208 = u1_col_out_208;
assign u2_col_in_209 = u1_col_out_209;
assign u2_col_in_210 = u1_col_out_210;
assign u2_col_in_211 = u1_col_out_211;
assign u2_col_in_212 = u1_col_out_212;
assign u2_col_in_213 = u1_col_out_213;
assign u2_col_in_214 = u1_col_out_214;
assign u2_col_in_215 = u1_col_out_215;
assign u2_col_in_216 = u1_col_out_216;
assign u2_col_in_217 = u1_col_out_217;
assign u2_col_in_218 = u1_col_out_218;
assign u2_col_in_219 = u1_col_out_219;
assign u2_col_in_220 = u1_col_out_220;
assign u2_col_in_221 = u1_col_out_221;
assign u2_col_in_222 = u1_col_out_222;
assign u2_col_in_223 = u1_col_out_223;
assign u2_col_in_224 = u1_col_out_224;
assign u2_col_in_225 = u1_col_out_225;
assign u2_col_in_226 = u1_col_out_226;
assign u2_col_in_227 = u1_col_out_227;
assign u2_col_in_228 = u1_col_out_228;
assign u2_col_in_229 = u1_col_out_229;
assign u2_col_in_230 = u1_col_out_230;
assign u2_col_in_231 = u1_col_out_231;
assign u2_col_in_232 = u1_col_out_232;
assign u2_col_in_233 = u1_col_out_233;
assign u2_col_in_234 = u1_col_out_234;
assign u2_col_in_235 = u1_col_out_235;
assign u2_col_in_236 = u1_col_out_236;
assign u2_col_in_237 = u1_col_out_237;
assign u2_col_in_238 = u1_col_out_238;
assign u2_col_in_239 = u1_col_out_239;
assign u2_col_in_240 = u1_col_out_240;
assign u2_col_in_241 = u1_col_out_241;
assign u2_col_in_242 = u1_col_out_242;
assign u2_col_in_243 = u1_col_out_243;
assign u2_col_in_244 = u1_col_out_244;
assign u2_col_in_245 = u1_col_out_245;
assign u2_col_in_246 = u1_col_out_246;
assign u2_col_in_247 = u1_col_out_247;
assign u2_col_in_248 = u1_col_out_248;
assign u2_col_in_249 = u1_col_out_249;
assign u2_col_in_250 = u1_col_out_250;
assign u2_col_in_251 = u1_col_out_251;
assign u2_col_in_252 = u1_col_out_252;
assign u2_col_in_253 = u1_col_out_253;
assign u2_col_in_254 = u1_col_out_254;
assign u2_col_in_255 = u1_col_out_255;
assign u2_col_in_256 = u1_col_out_256;
assign u2_col_in_257 = u1_col_out_257;
assign u2_col_in_258 = u1_col_out_258;
assign u2_col_in_259 = u1_col_out_259;
assign u2_col_in_260 = u1_col_out_260;
assign u2_col_in_261 = u1_col_out_261;
assign u2_col_in_262 = u1_col_out_262;
assign u2_col_in_263 = u1_col_out_263;
assign u2_col_in_264 = u1_col_out_264;
assign u2_col_in_265 = u1_col_out_265;
assign u2_col_in_266 = u1_col_out_266;
assign u2_col_in_267 = u1_col_out_267;
assign u2_col_in_268 = u1_col_out_268;
assign u2_col_in_269 = u1_col_out_269;
assign u2_col_in_270 = u1_col_out_270;
assign u2_col_in_271 = u1_col_out_271;
assign u2_col_in_272 = u1_col_out_272;
assign u2_col_in_273 = u1_col_out_273;
assign u2_col_in_274 = u1_col_out_274;
assign u2_col_in_275 = u1_col_out_275;
assign u2_col_in_276 = u1_col_out_276;
assign u2_col_in_277 = u1_col_out_277;
assign u2_col_in_278 = u1_col_out_278;
assign u2_col_in_279 = u1_col_out_279;
assign u2_col_in_280 = u1_col_out_280;
assign u2_col_in_281 = u1_col_out_281;
assign u2_col_in_282 = u1_col_out_282;
assign u2_col_in_283 = u1_col_out_283;
assign u2_col_in_284 = u1_col_out_284;
assign u2_col_in_285 = u1_col_out_285;
assign u2_col_in_286 = u1_col_out_286;
assign u2_col_in_287 = u1_col_out_287;
assign u2_col_in_288 = u1_col_out_288;
assign u2_col_in_289 = u1_col_out_289;
assign u2_col_in_290 = u1_col_out_290;
assign u2_col_in_291 = u1_col_out_291;
assign u2_col_in_292 = u1_col_out_292;
assign u2_col_in_293 = u1_col_out_293;
assign u2_col_in_294 = u1_col_out_294;
assign u2_col_in_295 = u1_col_out_295;
assign u2_col_in_296 = u1_col_out_296;
assign u2_col_in_297 = u1_col_out_297;
assign u2_col_in_298 = u1_col_out_298;
assign u2_col_in_299 = u1_col_out_299;
assign u2_col_in_300 = u1_col_out_300;
assign u2_col_in_301 = u1_col_out_301;
assign u2_col_in_302 = u1_col_out_302;
assign u2_col_in_303 = u1_col_out_303;
assign u2_col_in_304 = u1_col_out_304;
assign u2_col_in_305 = u1_col_out_305;
assign u2_col_in_306 = u1_col_out_306;
assign u2_col_in_307 = u1_col_out_307;
assign u2_col_in_308 = u1_col_out_308;
assign u2_col_in_309 = u1_col_out_309;
assign u2_col_in_310 = u1_col_out_310;
assign u2_col_in_311 = u1_col_out_311;
assign u2_col_in_312 = u1_col_out_312;
assign u2_col_in_313 = u1_col_out_313;
assign u2_col_in_314 = u1_col_out_314;
assign u2_col_in_315 = u1_col_out_315;
assign u2_col_in_316 = u1_col_out_316;
assign u2_col_in_317 = u1_col_out_317;
assign u2_col_in_318 = u1_col_out_318;
assign u2_col_in_319 = u1_col_out_319;
assign u2_col_in_320 = u1_col_out_320;
assign u2_col_in_321 = u1_col_out_321;
assign u2_col_in_322 = u1_col_out_322;
assign u2_col_in_323 = u1_col_out_323;
assign u2_col_in_324 = u1_col_out_324;
assign u2_col_in_325 = u1_col_out_325;
assign u2_col_in_326 = u1_col_out_326;
assign u2_col_in_327 = u1_col_out_327;
assign u2_col_in_328 = u1_col_out_328;
assign u2_col_in_329 = u1_col_out_329;
assign u2_col_in_330 = u1_col_out_330;
assign u2_col_in_331 = u1_col_out_331;
assign u2_col_in_332 = u1_col_out_332;
assign u2_col_in_333 = u1_col_out_333;
assign u2_col_in_334 = u1_col_out_334;
assign u2_col_in_335 = u1_col_out_335;
assign u2_col_in_336 = u1_col_out_336;
assign u2_col_in_337 = u1_col_out_337;
assign u2_col_in_338 = u1_col_out_338;
assign u2_col_in_339 = u1_col_out_339;
assign u2_col_in_340 = u1_col_out_340;
assign u2_col_in_341 = u1_col_out_341;
assign u2_col_in_342 = u1_col_out_342;
assign u2_col_in_343 = u1_col_out_343;
assign u2_col_in_344 = u1_col_out_344;
assign u2_col_in_345 = u1_col_out_345;
assign u2_col_in_346 = u1_col_out_346;
assign u2_col_in_347 = u1_col_out_347;
assign u2_col_in_348 = u1_col_out_348;
assign u2_col_in_349 = u1_col_out_349;
assign u2_col_in_350 = u1_col_out_350;
assign u2_col_in_351 = u1_col_out_351;
assign u2_col_in_352 = u1_col_out_352;
assign u2_col_in_353 = u1_col_out_353;
assign u2_col_in_354 = u1_col_out_354;
assign u2_col_in_355 = u1_col_out_355;
assign u2_col_in_356 = u1_col_out_356;
assign u2_col_in_357 = u1_col_out_357;
assign u2_col_in_358 = u1_col_out_358;
assign u2_col_in_359 = u1_col_out_359;
assign u2_col_in_360 = u1_col_out_360;
assign u2_col_in_361 = u1_col_out_361;
assign u2_col_in_362 = u1_col_out_362;
assign u2_col_in_363 = u1_col_out_363;
assign u2_col_in_364 = u1_col_out_364;
assign u2_col_in_365 = u1_col_out_365;
assign u2_col_in_366 = u1_col_out_366;
assign u2_col_in_367 = u1_col_out_367;
assign u2_col_in_368 = u1_col_out_368;
assign u2_col_in_369 = u1_col_out_369;
assign u2_col_in_370 = u1_col_out_370;
assign u2_col_in_371 = u1_col_out_371;
assign u2_col_in_372 = u1_col_out_372;
assign u2_col_in_373 = u1_col_out_373;
assign u2_col_in_374 = u1_col_out_374;
assign u2_col_in_375 = u1_col_out_375;
assign u2_col_in_376 = u1_col_out_376;
assign u2_col_in_377 = u1_col_out_377;
assign u2_col_in_378 = u1_col_out_378;
assign u2_col_in_379 = u1_col_out_379;
assign u2_col_in_380 = u1_col_out_380;
assign u2_col_in_381 = u1_col_out_381;
assign u2_col_in_382 = u1_col_out_382;
assign u2_col_in_383 = u1_col_out_383;
assign u2_col_in_384 = u1_col_out_384;
assign u2_col_in_385 = u1_col_out_385;
assign u2_col_in_386 = u1_col_out_386;
assign u2_col_in_387 = u1_col_out_387;
assign u2_col_in_388 = u1_col_out_388;
assign u2_col_in_389 = u1_col_out_389;
assign u2_col_in_390 = u1_col_out_390;
assign u2_col_in_391 = u1_col_out_391;
assign u2_col_in_392 = u1_col_out_392;
assign u2_col_in_393 = u1_col_out_393;
assign u2_col_in_394 = u1_col_out_394;
assign u2_col_in_395 = u1_col_out_395;
assign u2_col_in_396 = u1_col_out_396;
assign u2_col_in_397 = u1_col_out_397;
assign u2_col_in_398 = u1_col_out_398;
assign u2_col_in_399 = u1_col_out_399;
assign u2_col_in_400 = u1_col_out_400;
assign u2_col_in_401 = u1_col_out_401;
assign u2_col_in_402 = u1_col_out_402;
assign u2_col_in_403 = u1_col_out_403;
assign u2_col_in_404 = u1_col_out_404;
assign u2_col_in_405 = u1_col_out_405;
assign u2_col_in_406 = u1_col_out_406;
assign u2_col_in_407 = u1_col_out_407;
assign u2_col_in_408 = u1_col_out_408;
assign u2_col_in_409 = u1_col_out_409;
assign u2_col_in_410 = u1_col_out_410;
assign u2_col_in_411 = u1_col_out_411;
assign u2_col_in_412 = u1_col_out_412;
assign u2_col_in_413 = u1_col_out_413;
assign u2_col_in_414 = u1_col_out_414;
assign u2_col_in_415 = u1_col_out_415;
assign u2_col_in_416 = u1_col_out_416;
assign u2_col_in_417 = u1_col_out_417;
assign u2_col_in_418 = u1_col_out_418;
assign u2_col_in_419 = u1_col_out_419;
assign u2_col_in_420 = u1_col_out_420;
assign u2_col_in_421 = u1_col_out_421;
assign u2_col_in_422 = u1_col_out_422;
assign u2_col_in_423 = u1_col_out_423;
assign u2_col_in_424 = u1_col_out_424;
assign u2_col_in_425 = u1_col_out_425;
assign u2_col_in_426 = u1_col_out_426;
assign u2_col_in_427 = u1_col_out_427;
assign u2_col_in_428 = u1_col_out_428;
assign u2_col_in_429 = u1_col_out_429;
assign u2_col_in_430 = u1_col_out_430;
assign u2_col_in_431 = u1_col_out_431;
assign u2_col_in_432 = u1_col_out_432;
assign u2_col_in_433 = u1_col_out_433;
assign u2_col_in_434 = u1_col_out_434;
assign u2_col_in_435 = u1_col_out_435;
assign u2_col_in_436 = u1_col_out_436;
assign u2_col_in_437 = u1_col_out_437;
assign u2_col_in_438 = u1_col_out_438;
assign u2_col_in_439 = u1_col_out_439;
assign u2_col_in_440 = u1_col_out_440;
assign u2_col_in_441 = u1_col_out_441;
assign u2_col_in_442 = u1_col_out_442;
assign u2_col_in_443 = u1_col_out_443;
assign u2_col_in_444 = u1_col_out_444;
assign u2_col_in_445 = u1_col_out_445;
assign u2_col_in_446 = u1_col_out_446;
assign u2_col_in_447 = u1_col_out_447;
assign u2_col_in_448 = u1_col_out_448;
assign u2_col_in_449 = u1_col_out_449;
assign u2_col_in_450 = u1_col_out_450;
assign u2_col_in_451 = u1_col_out_451;
assign u2_col_in_452 = u1_col_out_452;
assign u2_col_in_453 = u1_col_out_453;
assign u2_col_in_454 = u1_col_out_454;
assign u2_col_in_455 = u1_col_out_455;
assign u2_col_in_456 = u1_col_out_456;
assign u2_col_in_457 = u1_col_out_457;
assign u2_col_in_458 = u1_col_out_458;
assign u2_col_in_459 = u1_col_out_459;
assign u2_col_in_460 = u1_col_out_460;
assign u2_col_in_461 = u1_col_out_461;
assign u2_col_in_462 = u1_col_out_462;
assign u2_col_in_463 = u1_col_out_463;
assign u2_col_in_464 = u1_col_out_464;
assign u2_col_in_465 = u1_col_out_465;
assign u2_col_in_466 = u1_col_out_466;
assign u2_col_in_467 = u1_col_out_467;
assign u2_col_in_468 = u1_col_out_468;
assign u2_col_in_469 = u1_col_out_469;
assign u2_col_in_470 = u1_col_out_470;
assign u2_col_in_471 = u1_col_out_471;
assign u2_col_in_472 = u1_col_out_472;
assign u2_col_in_473 = u1_col_out_473;
assign u2_col_in_474 = u1_col_out_474;
assign u2_col_in_475 = u1_col_out_475;
assign u2_col_in_476 = u1_col_out_476;
assign u2_col_in_477 = u1_col_out_477;
assign u2_col_in_478 = u1_col_out_478;
assign u2_col_in_479 = u1_col_out_479;
assign u2_col_in_480 = u1_col_out_480;
assign u2_col_in_481 = u1_col_out_481;
assign u2_col_in_482 = u1_col_out_482;
assign u2_col_in_483 = u1_col_out_483;
assign u2_col_in_484 = u1_col_out_484;
assign u2_col_in_485 = u1_col_out_485;
assign u2_col_in_486 = u1_col_out_486;
assign u2_col_in_487 = u1_col_out_487;
assign u2_col_in_488 = u1_col_out_488;
assign u2_col_in_489 = u1_col_out_489;
assign u2_col_in_490 = u1_col_out_490;
assign u2_col_in_491 = u1_col_out_491;
assign u2_col_in_492 = u1_col_out_492;
assign u2_col_in_493 = u1_col_out_493;
assign u2_col_in_494 = u1_col_out_494;
assign u2_col_in_495 = u1_col_out_495;
assign u2_col_in_496 = u1_col_out_496;
assign u2_col_in_497 = u1_col_out_497;
assign u2_col_in_498 = u1_col_out_498;
assign u2_col_in_499 = u1_col_out_499;
assign u2_col_in_500 = u1_col_out_500;
assign u2_col_in_501 = u1_col_out_501;
assign u2_col_in_502 = u1_col_out_502;
assign u2_col_in_503 = u1_col_out_503;
assign u2_col_in_504 = u1_col_out_504;
assign u2_col_in_505 = u1_col_out_505;
assign u2_col_in_506 = u1_col_out_506;
assign u2_col_in_507 = u1_col_out_507;
assign u2_col_in_508 = u1_col_out_508;
assign u2_col_in_509 = u1_col_out_509;
assign u2_col_in_510 = u1_col_out_510;
assign u2_col_in_511 = u1_col_out_511;
assign u2_col_in_512 = u1_col_out_512;
assign u2_col_in_513 = u1_col_out_513;
assign u2_col_in_514 = u1_col_out_514;
assign u2_col_in_515 = u1_col_out_515;
assign u2_col_in_516 = u1_col_out_516;
assign u2_col_in_517 = u1_col_out_517;
assign u2_col_in_518 = u1_col_out_518;
assign u2_col_in_519 = u1_col_out_519;
assign u2_col_in_520 = u1_col_out_520;
assign u2_col_in_521 = u1_col_out_521;
assign u2_col_in_522 = u1_col_out_522;
assign u2_col_in_523 = u1_col_out_523;
assign u2_col_in_524 = u1_col_out_524;
assign u2_col_in_525 = u1_col_out_525;
assign u2_col_in_526 = u1_col_out_526;
assign u2_col_in_527 = u1_col_out_527;
assign u2_col_in_528 = u1_col_out_528;
assign u2_col_in_529 = u1_col_out_529;
assign u2_col_in_530 = u1_col_out_530;
assign u2_col_in_531 = u1_col_out_531;
assign u2_col_in_532 = u1_col_out_532;
assign u2_col_in_533 = u1_col_out_533;
assign u2_col_in_534 = u1_col_out_534;
assign u2_col_in_535 = u1_col_out_535;
assign u2_col_in_536 = u1_col_out_536;
assign u2_col_in_537 = u1_col_out_537;
assign u2_col_in_538 = u1_col_out_538;
assign u2_col_in_539 = u1_col_out_539;
assign u2_col_in_540 = u1_col_out_540;
assign u2_col_in_541 = u1_col_out_541;
assign u2_col_in_542 = u1_col_out_542;
assign u2_col_in_543 = u1_col_out_543;
assign u2_col_in_544 = u1_col_out_544;
assign u2_col_in_545 = u1_col_out_545;
assign u2_col_in_546 = u1_col_out_546;
assign u2_col_in_547 = u1_col_out_547;
assign u2_col_in_548 = u1_col_out_548;
assign u2_col_in_549 = u1_col_out_549;
assign u2_col_in_550 = u1_col_out_550;
assign u2_col_in_551 = u1_col_out_551;
assign u2_col_in_552 = u1_col_out_552;
assign u2_col_in_553 = u1_col_out_553;
assign u2_col_in_554 = u1_col_out_554;
assign u2_col_in_555 = u1_col_out_555;
assign u2_col_in_556 = u1_col_out_556;
assign u2_col_in_557 = u1_col_out_557;
assign u2_col_in_558 = u1_col_out_558;
assign u2_col_in_559 = u1_col_out_559;
assign u2_col_in_560 = u1_col_out_560;
assign u2_col_in_561 = u1_col_out_561;
assign u2_col_in_562 = u1_col_out_562;
assign u2_col_in_563 = u1_col_out_563;
assign u2_col_in_564 = u1_col_out_564;
assign u2_col_in_565 = u1_col_out_565;
assign u2_col_in_566 = u1_col_out_566;
assign u2_col_in_567 = u1_col_out_567;
assign u2_col_in_568 = u1_col_out_568;
assign u2_col_in_569 = u1_col_out_569;
assign u2_col_in_570 = u1_col_out_570;
assign u2_col_in_571 = u1_col_out_571;
assign u2_col_in_572 = u1_col_out_572;
assign u2_col_in_573 = u1_col_out_573;
assign u2_col_in_574 = u1_col_out_574;
assign u2_col_in_575 = u1_col_out_575;
assign u2_col_in_576 = u1_col_out_576;
assign u2_col_in_577 = u1_col_out_577;
assign u2_col_in_578 = u1_col_out_578;
assign u2_col_in_579 = u1_col_out_579;
assign u2_col_in_580 = u1_col_out_580;
assign u2_col_in_581 = u1_col_out_581;
assign u2_col_in_582 = u1_col_out_582;
assign u2_col_in_583 = u1_col_out_583;
assign u2_col_in_584 = u1_col_out_584;
assign u2_col_in_585 = u1_col_out_585;
assign u2_col_in_586 = u1_col_out_586;
assign u2_col_in_587 = u1_col_out_587;
assign u2_col_in_588 = u1_col_out_588;
assign u2_col_in_589 = u1_col_out_589;
assign u2_col_in_590 = u1_col_out_590;
assign u2_col_in_591 = u1_col_out_591;
assign u2_col_in_592 = u1_col_out_592;
assign u2_col_in_593 = u1_col_out_593;
assign u2_col_in_594 = u1_col_out_594;
assign u2_col_in_595 = u1_col_out_595;
assign u2_col_in_596 = u1_col_out_596;
assign u2_col_in_597 = u1_col_out_597;
assign u2_col_in_598 = u1_col_out_598;
assign u2_col_in_599 = u1_col_out_599;
assign u2_col_in_600 = u1_col_out_600;
assign u2_col_in_601 = u1_col_out_601;
assign u2_col_in_602 = u1_col_out_602;
assign u2_col_in_603 = u1_col_out_603;
assign u2_col_in_604 = u1_col_out_604;
assign u2_col_in_605 = u1_col_out_605;
assign u2_col_in_606 = u1_col_out_606;
assign u2_col_in_607 = u1_col_out_607;
assign u2_col_in_608 = u1_col_out_608;
assign u2_col_in_609 = u1_col_out_609;
assign u2_col_in_610 = u1_col_out_610;
assign u2_col_in_611 = u1_col_out_611;
assign u2_col_in_612 = u1_col_out_612;
assign u2_col_in_613 = u1_col_out_613;
assign u2_col_in_614 = u1_col_out_614;
assign u2_col_in_615 = u1_col_out_615;
assign u2_col_in_616 = u1_col_out_616;
assign u2_col_in_617 = u1_col_out_617;
assign u2_col_in_618 = u1_col_out_618;
assign u2_col_in_619 = u1_col_out_619;
assign u2_col_in_620 = u1_col_out_620;
assign u2_col_in_621 = u1_col_out_621;
assign u2_col_in_622 = u1_col_out_622;
assign u2_col_in_623 = u1_col_out_623;
assign u2_col_in_624 = u1_col_out_624;
assign u2_col_in_625 = u1_col_out_625;
assign u2_col_in_626 = u1_col_out_626;
assign u2_col_in_627 = u1_col_out_627;
assign u2_col_in_628 = u1_col_out_628;
assign u2_col_in_629 = u1_col_out_629;
assign u2_col_in_630 = u1_col_out_630;
assign u2_col_in_631 = u1_col_out_631;
assign u2_col_in_632 = u1_col_out_632;
assign u2_col_in_633 = u1_col_out_633;
assign u2_col_in_634 = u1_col_out_634;
assign u2_col_in_635 = u1_col_out_635;
assign u2_col_in_636 = u1_col_out_636;
assign u2_col_in_637 = u1_col_out_637;
assign u2_col_in_638 = u1_col_out_638;
assign u2_col_in_639 = u1_col_out_639;
assign u2_col_in_640 = u1_col_out_640;
assign u2_col_in_641 = u1_col_out_641;
assign u2_col_in_642 = u1_col_out_642;
assign u2_col_in_643 = u1_col_out_643;
assign u2_col_in_644 = u1_col_out_644;
assign u2_col_in_645 = u1_col_out_645;
assign u2_col_in_646 = u1_col_out_646;
assign u2_col_in_647 = u1_col_out_647;
assign u2_col_in_648 = u1_col_out_648;
assign u2_col_in_649 = u1_col_out_649;
assign u2_col_in_650 = u1_col_out_650;
assign u2_col_in_651 = u1_col_out_651;
assign u2_col_in_652 = u1_col_out_652;
assign u2_col_in_653 = u1_col_out_653;
assign u2_col_in_654 = u1_col_out_654;
assign u2_col_in_655 = u1_col_out_655;
assign u2_col_in_656 = u1_col_out_656;
assign u2_col_in_657 = u1_col_out_657;
assign u2_col_in_658 = u1_col_out_658;
assign u2_col_in_659 = u1_col_out_659;
assign u2_col_in_660 = u1_col_out_660;
assign u2_col_in_661 = u1_col_out_661;
assign u2_col_in_662 = u1_col_out_662;
assign u2_col_in_663 = u1_col_out_663;
assign u2_col_in_664 = u1_col_out_664;
assign u2_col_in_665 = u1_col_out_665;
assign u2_col_in_666 = u1_col_out_666;
assign u2_col_in_667 = u1_col_out_667;
assign u2_col_in_668 = u1_col_out_668;
assign u2_col_in_669 = u1_col_out_669;
assign u2_col_in_670 = u1_col_out_670;
assign u2_col_in_671 = u1_col_out_671;
assign u2_col_in_672 = u1_col_out_672;
assign u2_col_in_673 = u1_col_out_673;
assign u2_col_in_674 = u1_col_out_674;
assign u2_col_in_675 = u1_col_out_675;
assign u2_col_in_676 = u1_col_out_676;
assign u2_col_in_677 = u1_col_out_677;
assign u2_col_in_678 = u1_col_out_678;
assign u2_col_in_679 = u1_col_out_679;
assign u2_col_in_680 = u1_col_out_680;
assign u2_col_in_681 = u1_col_out_681;
assign u2_col_in_682 = u1_col_out_682;
assign u2_col_in_683 = u1_col_out_683;
assign u2_col_in_684 = u1_col_out_684;
assign u2_col_in_685 = u1_col_out_685;
assign u2_col_in_686 = u1_col_out_686;
assign u2_col_in_687 = u1_col_out_687;
assign u2_col_in_688 = u1_col_out_688;
assign u2_col_in_689 = u1_col_out_689;
assign u2_col_in_690 = u1_col_out_690;
assign u2_col_in_691 = u1_col_out_691;
assign u2_col_in_692 = u1_col_out_692;
assign u2_col_in_693 = u1_col_out_693;
assign u2_col_in_694 = u1_col_out_694;
assign u2_col_in_695 = u1_col_out_695;
assign u2_col_in_696 = u1_col_out_696;
assign u2_col_in_697 = u1_col_out_697;
assign u2_col_in_698 = u1_col_out_698;
assign u2_col_in_699 = u1_col_out_699;
assign u2_col_in_700 = u1_col_out_700;
assign u2_col_in_701 = u1_col_out_701;
assign u2_col_in_702 = u1_col_out_702;
assign u2_col_in_703 = u1_col_out_703;
assign u2_col_in_704 = u1_col_out_704;
assign u2_col_in_705 = u1_col_out_705;
assign u2_col_in_706 = u1_col_out_706;
assign u2_col_in_707 = u1_col_out_707;
assign u2_col_in_708 = u1_col_out_708;
assign u2_col_in_709 = u1_col_out_709;
assign u2_col_in_710 = u1_col_out_710;
assign u2_col_in_711 = u1_col_out_711;
assign u2_col_in_712 = u1_col_out_712;
assign u2_col_in_713 = u1_col_out_713;
assign u2_col_in_714 = u1_col_out_714;
assign u2_col_in_715 = u1_col_out_715;
assign u2_col_in_716 = u1_col_out_716;
assign u2_col_in_717 = u1_col_out_717;
assign u2_col_in_718 = u1_col_out_718;
assign u2_col_in_719 = u1_col_out_719;
assign u2_col_in_720 = u1_col_out_720;
assign u2_col_in_721 = u1_col_out_721;
assign u2_col_in_722 = u1_col_out_722;
assign u2_col_in_723 = u1_col_out_723;
assign u2_col_in_724 = u1_col_out_724;
assign u2_col_in_725 = u1_col_out_725;
assign u2_col_in_726 = u1_col_out_726;
assign u2_col_in_727 = u1_col_out_727;
assign u2_col_in_728 = u1_col_out_728;
assign u2_col_in_729 = u1_col_out_729;
assign u2_col_in_730 = u1_col_out_730;
assign u2_col_in_731 = u1_col_out_731;
assign u2_col_in_732 = u1_col_out_732;
assign u2_col_in_733 = u1_col_out_733;
assign u2_col_in_734 = u1_col_out_734;
assign u2_col_in_735 = u1_col_out_735;
assign u2_col_in_736 = u1_col_out_736;
assign u2_col_in_737 = u1_col_out_737;
assign u2_col_in_738 = u1_col_out_738;
assign u2_col_in_739 = u1_col_out_739;
assign u2_col_in_740 = u1_col_out_740;
assign u2_col_in_741 = u1_col_out_741;
assign u2_col_in_742 = u1_col_out_742;
assign u2_col_in_743 = u1_col_out_743;
assign u2_col_in_744 = u1_col_out_744;
assign u2_col_in_745 = u1_col_out_745;
assign u2_col_in_746 = u1_col_out_746;
assign u2_col_in_747 = u1_col_out_747;
assign u2_col_in_748 = u1_col_out_748;
assign u2_col_in_749 = u1_col_out_749;
assign u2_col_in_750 = u1_col_out_750;
assign u2_col_in_751 = u1_col_out_751;
assign u2_col_in_752 = u1_col_out_752;
assign u2_col_in_753 = u1_col_out_753;
assign u2_col_in_754 = u1_col_out_754;
assign u2_col_in_755 = u1_col_out_755;
assign u2_col_in_756 = u1_col_out_756;
assign u2_col_in_757 = u1_col_out_757;
assign u2_col_in_758 = u1_col_out_758;
assign u2_col_in_759 = u1_col_out_759;
assign u2_col_in_760 = u1_col_out_760;
assign u2_col_in_761 = u1_col_out_761;
assign u2_col_in_762 = u1_col_out_762;
assign u2_col_in_763 = u1_col_out_763;
assign u2_col_in_764 = u1_col_out_764;
assign u2_col_in_765 = u1_col_out_765;
assign u2_col_in_766 = u1_col_out_766;
assign u2_col_in_767 = u1_col_out_767;
assign u2_col_in_768 = u1_col_out_768;
assign u2_col_in_769 = u1_col_out_769;
assign u2_col_in_770 = u1_col_out_770;
assign u2_col_in_771 = u1_col_out_771;
assign u2_col_in_772 = u1_col_out_772;
assign u2_col_in_773 = u1_col_out_773;
assign u2_col_in_774 = u1_col_out_774;
assign u2_col_in_775 = u1_col_out_775;
assign u2_col_in_776 = u1_col_out_776;
assign u2_col_in_777 = u1_col_out_777;
assign u2_col_in_778 = u1_col_out_778;
assign u2_col_in_779 = u1_col_out_779;
assign u2_col_in_780 = u1_col_out_780;
assign u2_col_in_781 = u1_col_out_781;
assign u2_col_in_782 = u1_col_out_782;
assign u2_col_in_783 = u1_col_out_783;
assign u2_col_in_784 = u1_col_out_784;
assign u2_col_in_785 = u1_col_out_785;
assign u2_col_in_786 = u1_col_out_786;
assign u2_col_in_787 = u1_col_out_787;
assign u2_col_in_788 = u1_col_out_788;
assign u2_col_in_789 = u1_col_out_789;
assign u2_col_in_790 = u1_col_out_790;
assign u2_col_in_791 = u1_col_out_791;
assign u2_col_in_792 = u1_col_out_792;
assign u2_col_in_793 = u1_col_out_793;
assign u2_col_in_794 = u1_col_out_794;
assign u2_col_in_795 = u1_col_out_795;
assign u2_col_in_796 = u1_col_out_796;
assign u2_col_in_797 = u1_col_out_797;
assign u2_col_in_798 = u1_col_out_798;
assign u2_col_in_799 = u1_col_out_799;
assign u2_col_in_800 = u1_col_out_800;
assign u2_col_in_801 = u1_col_out_801;
assign u2_col_in_802 = u1_col_out_802;
assign u2_col_in_803 = u1_col_out_803;
assign u2_col_in_804 = u1_col_out_804;
assign u2_col_in_805 = u1_col_out_805;
assign u2_col_in_806 = u1_col_out_806;
assign u2_col_in_807 = u1_col_out_807;
assign u2_col_in_808 = u1_col_out_808;
assign u2_col_in_809 = u1_col_out_809;
assign u2_col_in_810 = u1_col_out_810;
assign u2_col_in_811 = u1_col_out_811;
assign u2_col_in_812 = u1_col_out_812;
assign u2_col_in_813 = u1_col_out_813;
assign u2_col_in_814 = u1_col_out_814;
assign u2_col_in_815 = u1_col_out_815;
assign u2_col_in_816 = u1_col_out_816;
assign u2_col_in_817 = u1_col_out_817;
assign u2_col_in_818 = u1_col_out_818;
assign u2_col_in_819 = u1_col_out_819;
assign u2_col_in_820 = u1_col_out_820;
assign u2_col_in_821 = u1_col_out_821;
assign u2_col_in_822 = u1_col_out_822;
assign u2_col_in_823 = u1_col_out_823;
assign u2_col_in_824 = u1_col_out_824;
assign u2_col_in_825 = u1_col_out_825;
assign u2_col_in_826 = u1_col_out_826;
assign u2_col_in_827 = u1_col_out_827;
assign u2_col_in_828 = u1_col_out_828;
assign u2_col_in_829 = u1_col_out_829;
assign u2_col_in_830 = u1_col_out_830;
assign u2_col_in_831 = u1_col_out_831;
assign u2_col_in_832 = u1_col_out_832;
assign u2_col_in_833 = u1_col_out_833;
assign u2_col_in_834 = u1_col_out_834;
assign u2_col_in_835 = u1_col_out_835;
assign u2_col_in_836 = u1_col_out_836;
assign u2_col_in_837 = u1_col_out_837;
assign u2_col_in_838 = u1_col_out_838;
assign u2_col_in_839 = u1_col_out_839;
assign u2_col_in_840 = u1_col_out_840;
assign u2_col_in_841 = u1_col_out_841;
assign u2_col_in_842 = u1_col_out_842;
assign u2_col_in_843 = u1_col_out_843;
assign u2_col_in_844 = u1_col_out_844;
assign u2_col_in_845 = u1_col_out_845;
assign u2_col_in_846 = u1_col_out_846;
assign u2_col_in_847 = u1_col_out_847;
assign u2_col_in_848 = u1_col_out_848;
assign u2_col_in_849 = u1_col_out_849;
assign u2_col_in_850 = u1_col_out_850;
assign u2_col_in_851 = u1_col_out_851;
assign u2_col_in_852 = u1_col_out_852;
assign u2_col_in_853 = u1_col_out_853;
assign u2_col_in_854 = u1_col_out_854;
assign u2_col_in_855 = u1_col_out_855;
assign u2_col_in_856 = u1_col_out_856;
assign u2_col_in_857 = u1_col_out_857;
assign u2_col_in_858 = u1_col_out_858;
assign u2_col_in_859 = u1_col_out_859;
assign u2_col_in_860 = u1_col_out_860;
assign u2_col_in_861 = u1_col_out_861;
assign u2_col_in_862 = u1_col_out_862;
assign u2_col_in_863 = u1_col_out_863;
assign u2_col_in_864 = u1_col_out_864;
assign u2_col_in_865 = u1_col_out_865;
assign u2_col_in_866 = u1_col_out_866;
assign u2_col_in_867 = u1_col_out_867;
assign u2_col_in_868 = u1_col_out_868;
assign u2_col_in_869 = u1_col_out_869;
assign u2_col_in_870 = u1_col_out_870;
assign u2_col_in_871 = u1_col_out_871;
assign u2_col_in_872 = u1_col_out_872;
assign u2_col_in_873 = u1_col_out_873;
assign u2_col_in_874 = u1_col_out_874;
assign u2_col_in_875 = u1_col_out_875;
assign u2_col_in_876 = u1_col_out_876;
assign u2_col_in_877 = u1_col_out_877;
assign u2_col_in_878 = u1_col_out_878;
assign u2_col_in_879 = u1_col_out_879;
assign u2_col_in_880 = u1_col_out_880;
assign u2_col_in_881 = u1_col_out_881;
assign u2_col_in_882 = u1_col_out_882;
assign u2_col_in_883 = u1_col_out_883;
assign u2_col_in_884 = u1_col_out_884;
assign u2_col_in_885 = u1_col_out_885;
assign u2_col_in_886 = u1_col_out_886;
assign u2_col_in_887 = u1_col_out_887;
assign u2_col_in_888 = u1_col_out_888;
assign u2_col_in_889 = u1_col_out_889;
assign u2_col_in_890 = u1_col_out_890;
assign u2_col_in_891 = u1_col_out_891;
assign u2_col_in_892 = u1_col_out_892;
assign u2_col_in_893 = u1_col_out_893;
assign u2_col_in_894 = u1_col_out_894;
assign u2_col_in_895 = u1_col_out_895;
assign u2_col_in_896 = u1_col_out_896;
assign u2_col_in_897 = u1_col_out_897;
assign u2_col_in_898 = u1_col_out_898;
assign u2_col_in_899 = u1_col_out_899;
assign u2_col_in_900 = u1_col_out_900;
assign u2_col_in_901 = u1_col_out_901;
assign u2_col_in_902 = u1_col_out_902;
assign u2_col_in_903 = u1_col_out_903;
assign u2_col_in_904 = u1_col_out_904;
assign u2_col_in_905 = u1_col_out_905;
assign u2_col_in_906 = u1_col_out_906;
assign u2_col_in_907 = u1_col_out_907;
assign u2_col_in_908 = u1_col_out_908;
assign u2_col_in_909 = u1_col_out_909;
assign u2_col_in_910 = u1_col_out_910;
assign u2_col_in_911 = u1_col_out_911;
assign u2_col_in_912 = u1_col_out_912;
assign u2_col_in_913 = u1_col_out_913;
assign u2_col_in_914 = u1_col_out_914;
assign u2_col_in_915 = u1_col_out_915;
assign u2_col_in_916 = u1_col_out_916;
assign u2_col_in_917 = u1_col_out_917;
assign u2_col_in_918 = u1_col_out_918;
assign u2_col_in_919 = u1_col_out_919;
assign u2_col_in_920 = u1_col_out_920;
assign u2_col_in_921 = u1_col_out_921;
assign u2_col_in_922 = u1_col_out_922;
assign u2_col_in_923 = u1_col_out_923;
assign u2_col_in_924 = u1_col_out_924;
assign u2_col_in_925 = u1_col_out_925;
assign u2_col_in_926 = u1_col_out_926;
assign u2_col_in_927 = u1_col_out_927;
assign u2_col_in_928 = u1_col_out_928;
assign u2_col_in_929 = u1_col_out_929;
assign u2_col_in_930 = u1_col_out_930;
assign u2_col_in_931 = u1_col_out_931;
assign u2_col_in_932 = u1_col_out_932;
assign u2_col_in_933 = u1_col_out_933;
assign u2_col_in_934 = u1_col_out_934;
assign u2_col_in_935 = u1_col_out_935;
assign u2_col_in_936 = u1_col_out_936;
assign u2_col_in_937 = u1_col_out_937;
assign u2_col_in_938 = u1_col_out_938;
assign u2_col_in_939 = u1_col_out_939;
assign u2_col_in_940 = u1_col_out_940;
assign u2_col_in_941 = u1_col_out_941;
assign u2_col_in_942 = u1_col_out_942;
assign u2_col_in_943 = u1_col_out_943;
assign u2_col_in_944 = u1_col_out_944;
assign u2_col_in_945 = u1_col_out_945;
assign u2_col_in_946 = u1_col_out_946;
assign u2_col_in_947 = u1_col_out_947;
assign u2_col_in_948 = u1_col_out_948;
assign u2_col_in_949 = u1_col_out_949;
assign u2_col_in_950 = u1_col_out_950;
assign u2_col_in_951 = u1_col_out_951;
assign u2_col_in_952 = u1_col_out_952;
assign u2_col_in_953 = u1_col_out_953;
assign u2_col_in_954 = u1_col_out_954;
assign u2_col_in_955 = u1_col_out_955;
assign u2_col_in_956 = u1_col_out_956;
assign u2_col_in_957 = u1_col_out_957;
assign u2_col_in_958 = u1_col_out_958;
assign u2_col_in_959 = u1_col_out_959;
assign u2_col_in_960 = u1_col_out_960;
assign u2_col_in_961 = u1_col_out_961;
assign u2_col_in_962 = u1_col_out_962;
assign u2_col_in_963 = u1_col_out_963;
assign u2_col_in_964 = u1_col_out_964;
assign u2_col_in_965 = u1_col_out_965;
assign u2_col_in_966 = u1_col_out_966;
assign u2_col_in_967 = u1_col_out_967;
assign u2_col_in_968 = u1_col_out_968;
assign u2_col_in_969 = u1_col_out_969;
assign u2_col_in_970 = u1_col_out_970;
assign u2_col_in_971 = u1_col_out_971;
assign u2_col_in_972 = u1_col_out_972;
assign u2_col_in_973 = u1_col_out_973;
assign u2_col_in_974 = u1_col_out_974;
assign u2_col_in_975 = u1_col_out_975;
assign u2_col_in_976 = u1_col_out_976;
assign u2_col_in_977 = u1_col_out_977;
assign u2_col_in_978 = u1_col_out_978;
assign u2_col_in_979 = u1_col_out_979;
assign u2_col_in_980 = u1_col_out_980;
assign u2_col_in_981 = u1_col_out_981;
assign u2_col_in_982 = u1_col_out_982;
assign u2_col_in_983 = u1_col_out_983;
assign u2_col_in_984 = u1_col_out_984;
assign u2_col_in_985 = u1_col_out_985;
assign u2_col_in_986 = u1_col_out_986;
assign u2_col_in_987 = u1_col_out_987;
assign u2_col_in_988 = u1_col_out_988;
assign u2_col_in_989 = u1_col_out_989;
assign u2_col_in_990 = u1_col_out_990;
assign u2_col_in_991 = u1_col_out_991;
assign u2_col_in_992 = u1_col_out_992;
assign u2_col_in_993 = u1_col_out_993;
assign u2_col_in_994 = u1_col_out_994;
assign u2_col_in_995 = u1_col_out_995;
assign u2_col_in_996 = u1_col_out_996;
assign u2_col_in_997 = u1_col_out_997;
assign u2_col_in_998 = u1_col_out_998;
assign u2_col_in_999 = u1_col_out_999;
assign u2_col_in_1000 = u1_col_out_1000;
assign u2_col_in_1001 = u1_col_out_1001;
assign u2_col_in_1002 = u1_col_out_1002;
assign u2_col_in_1003 = u1_col_out_1003;
assign u2_col_in_1004 = u1_col_out_1004;
assign u2_col_in_1005 = u1_col_out_1005;
assign u2_col_in_1006 = u1_col_out_1006;
assign u2_col_in_1007 = u1_col_out_1007;
assign u2_col_in_1008 = u1_col_out_1008;
assign u2_col_in_1009 = u1_col_out_1009;
assign u2_col_in_1010 = u1_col_out_1010;
assign u2_col_in_1011 = u1_col_out_1011;
assign u2_col_in_1012 = u1_col_out_1012;
assign u2_col_in_1013 = u1_col_out_1013;
assign u2_col_in_1014 = u1_col_out_1014;
assign u2_col_in_1015 = u1_col_out_1015;
assign u2_col_in_1016 = u1_col_out_1016;
assign u2_col_in_1017 = u1_col_out_1017;
assign u2_col_in_1018 = u1_col_out_1018;
assign u2_col_in_1019 = u1_col_out_1019;
assign u2_col_in_1020 = u1_col_out_1020;
assign u2_col_in_1021 = u1_col_out_1021;
assign u2_col_in_1022 = u1_col_out_1022;
assign u2_col_in_1023 = u1_col_out_1023;
assign u2_col_in_1024 = u1_col_out_1024;
assign u2_col_in_1025 = u1_col_out_1025;
assign u2_col_in_1026 = u1_col_out_1026;
assign u2_col_in_1027 = u1_col_out_1027;
assign u2_col_in_1028 = u1_col_out_1028;
assign u2_col_in_1029 = u1_col_out_1029;

//*****************************************************
//**************u2压缩阵列******************************
//*****************************************************
compressor_array_48_16_1030 u2_ca_48_17_1030
(
    .col_in_0(u2_col_in_0),
    .col_in_1(u2_col_in_1),
    .col_in_2(u2_col_in_2),
    .col_in_3(u2_col_in_3),
    .col_in_4(u2_col_in_4),
    .col_in_5(u2_col_in_5),
    .col_in_6(u2_col_in_6),
    .col_in_7(u2_col_in_7),
    .col_in_8(u2_col_in_8),
    .col_in_9(u2_col_in_9),
    .col_in_10(u2_col_in_10),
    .col_in_11(u2_col_in_11),
    .col_in_12(u2_col_in_12),
    .col_in_13(u2_col_in_13),
    .col_in_14(u2_col_in_14),
    .col_in_15(u2_col_in_15),
    .col_in_16(u2_col_in_16),
    .col_in_17(u2_col_in_17),
    .col_in_18(u2_col_in_18),
    .col_in_19(u2_col_in_19),
    .col_in_20(u2_col_in_20),
    .col_in_21(u2_col_in_21),
    .col_in_22(u2_col_in_22),
    .col_in_23(u2_col_in_23),
    .col_in_24(u2_col_in_24),
    .col_in_25(u2_col_in_25),
    .col_in_26(u2_col_in_26),
    .col_in_27(u2_col_in_27),
    .col_in_28(u2_col_in_28),
    .col_in_29(u2_col_in_29),
    .col_in_30(u2_col_in_30),
    .col_in_31(u2_col_in_31),
    .col_in_32(u2_col_in_32),
    .col_in_33(u2_col_in_33),
    .col_in_34(u2_col_in_34),
    .col_in_35(u2_col_in_35),
    .col_in_36(u2_col_in_36),
    .col_in_37(u2_col_in_37),
    .col_in_38(u2_col_in_38),
    .col_in_39(u2_col_in_39),
    .col_in_40(u2_col_in_40),
    .col_in_41(u2_col_in_41),
    .col_in_42(u2_col_in_42),
    .col_in_43(u2_col_in_43),
    .col_in_44(u2_col_in_44),
    .col_in_45(u2_col_in_45),
    .col_in_46(u2_col_in_46),
    .col_in_47(u2_col_in_47),
    .col_in_48(u2_col_in_48),
    .col_in_49(u2_col_in_49),
    .col_in_50(u2_col_in_50),
    .col_in_51(u2_col_in_51),
    .col_in_52(u2_col_in_52),
    .col_in_53(u2_col_in_53),
    .col_in_54(u2_col_in_54),
    .col_in_55(u2_col_in_55),
    .col_in_56(u2_col_in_56),
    .col_in_57(u2_col_in_57),
    .col_in_58(u2_col_in_58),
    .col_in_59(u2_col_in_59),
    .col_in_60(u2_col_in_60),
    .col_in_61(u2_col_in_61),
    .col_in_62(u2_col_in_62),
    .col_in_63(u2_col_in_63),
    .col_in_64(u2_col_in_64),
    .col_in_65(u2_col_in_65),
    .col_in_66(u2_col_in_66),
    .col_in_67(u2_col_in_67),
    .col_in_68(u2_col_in_68),
    .col_in_69(u2_col_in_69),
    .col_in_70(u2_col_in_70),
    .col_in_71(u2_col_in_71),
    .col_in_72(u2_col_in_72),
    .col_in_73(u2_col_in_73),
    .col_in_74(u2_col_in_74),
    .col_in_75(u2_col_in_75),
    .col_in_76(u2_col_in_76),
    .col_in_77(u2_col_in_77),
    .col_in_78(u2_col_in_78),
    .col_in_79(u2_col_in_79),
    .col_in_80(u2_col_in_80),
    .col_in_81(u2_col_in_81),
    .col_in_82(u2_col_in_82),
    .col_in_83(u2_col_in_83),
    .col_in_84(u2_col_in_84),
    .col_in_85(u2_col_in_85),
    .col_in_86(u2_col_in_86),
    .col_in_87(u2_col_in_87),
    .col_in_88(u2_col_in_88),
    .col_in_89(u2_col_in_89),
    .col_in_90(u2_col_in_90),
    .col_in_91(u2_col_in_91),
    .col_in_92(u2_col_in_92),
    .col_in_93(u2_col_in_93),
    .col_in_94(u2_col_in_94),
    .col_in_95(u2_col_in_95),
    .col_in_96(u2_col_in_96),
    .col_in_97(u2_col_in_97),
    .col_in_98(u2_col_in_98),
    .col_in_99(u2_col_in_99),
    .col_in_100(u2_col_in_100),
    .col_in_101(u2_col_in_101),
    .col_in_102(u2_col_in_102),
    .col_in_103(u2_col_in_103),
    .col_in_104(u2_col_in_104),
    .col_in_105(u2_col_in_105),
    .col_in_106(u2_col_in_106),
    .col_in_107(u2_col_in_107),
    .col_in_108(u2_col_in_108),
    .col_in_109(u2_col_in_109),
    .col_in_110(u2_col_in_110),
    .col_in_111(u2_col_in_111),
    .col_in_112(u2_col_in_112),
    .col_in_113(u2_col_in_113),
    .col_in_114(u2_col_in_114),
    .col_in_115(u2_col_in_115),
    .col_in_116(u2_col_in_116),
    .col_in_117(u2_col_in_117),
    .col_in_118(u2_col_in_118),
    .col_in_119(u2_col_in_119),
    .col_in_120(u2_col_in_120),
    .col_in_121(u2_col_in_121),
    .col_in_122(u2_col_in_122),
    .col_in_123(u2_col_in_123),
    .col_in_124(u2_col_in_124),
    .col_in_125(u2_col_in_125),
    .col_in_126(u2_col_in_126),
    .col_in_127(u2_col_in_127),
    .col_in_128(u2_col_in_128),
    .col_in_129(u2_col_in_129),
    .col_in_130(u2_col_in_130),
    .col_in_131(u2_col_in_131),
    .col_in_132(u2_col_in_132),
    .col_in_133(u2_col_in_133),
    .col_in_134(u2_col_in_134),
    .col_in_135(u2_col_in_135),
    .col_in_136(u2_col_in_136),
    .col_in_137(u2_col_in_137),
    .col_in_138(u2_col_in_138),
    .col_in_139(u2_col_in_139),
    .col_in_140(u2_col_in_140),
    .col_in_141(u2_col_in_141),
    .col_in_142(u2_col_in_142),
    .col_in_143(u2_col_in_143),
    .col_in_144(u2_col_in_144),
    .col_in_145(u2_col_in_145),
    .col_in_146(u2_col_in_146),
    .col_in_147(u2_col_in_147),
    .col_in_148(u2_col_in_148),
    .col_in_149(u2_col_in_149),
    .col_in_150(u2_col_in_150),
    .col_in_151(u2_col_in_151),
    .col_in_152(u2_col_in_152),
    .col_in_153(u2_col_in_153),
    .col_in_154(u2_col_in_154),
    .col_in_155(u2_col_in_155),
    .col_in_156(u2_col_in_156),
    .col_in_157(u2_col_in_157),
    .col_in_158(u2_col_in_158),
    .col_in_159(u2_col_in_159),
    .col_in_160(u2_col_in_160),
    .col_in_161(u2_col_in_161),
    .col_in_162(u2_col_in_162),
    .col_in_163(u2_col_in_163),
    .col_in_164(u2_col_in_164),
    .col_in_165(u2_col_in_165),
    .col_in_166(u2_col_in_166),
    .col_in_167(u2_col_in_167),
    .col_in_168(u2_col_in_168),
    .col_in_169(u2_col_in_169),
    .col_in_170(u2_col_in_170),
    .col_in_171(u2_col_in_171),
    .col_in_172(u2_col_in_172),
    .col_in_173(u2_col_in_173),
    .col_in_174(u2_col_in_174),
    .col_in_175(u2_col_in_175),
    .col_in_176(u2_col_in_176),
    .col_in_177(u2_col_in_177),
    .col_in_178(u2_col_in_178),
    .col_in_179(u2_col_in_179),
    .col_in_180(u2_col_in_180),
    .col_in_181(u2_col_in_181),
    .col_in_182(u2_col_in_182),
    .col_in_183(u2_col_in_183),
    .col_in_184(u2_col_in_184),
    .col_in_185(u2_col_in_185),
    .col_in_186(u2_col_in_186),
    .col_in_187(u2_col_in_187),
    .col_in_188(u2_col_in_188),
    .col_in_189(u2_col_in_189),
    .col_in_190(u2_col_in_190),
    .col_in_191(u2_col_in_191),
    .col_in_192(u2_col_in_192),
    .col_in_193(u2_col_in_193),
    .col_in_194(u2_col_in_194),
    .col_in_195(u2_col_in_195),
    .col_in_196(u2_col_in_196),
    .col_in_197(u2_col_in_197),
    .col_in_198(u2_col_in_198),
    .col_in_199(u2_col_in_199),
    .col_in_200(u2_col_in_200),
    .col_in_201(u2_col_in_201),
    .col_in_202(u2_col_in_202),
    .col_in_203(u2_col_in_203),
    .col_in_204(u2_col_in_204),
    .col_in_205(u2_col_in_205),
    .col_in_206(u2_col_in_206),
    .col_in_207(u2_col_in_207),
    .col_in_208(u2_col_in_208),
    .col_in_209(u2_col_in_209),
    .col_in_210(u2_col_in_210),
    .col_in_211(u2_col_in_211),
    .col_in_212(u2_col_in_212),
    .col_in_213(u2_col_in_213),
    .col_in_214(u2_col_in_214),
    .col_in_215(u2_col_in_215),
    .col_in_216(u2_col_in_216),
    .col_in_217(u2_col_in_217),
    .col_in_218(u2_col_in_218),
    .col_in_219(u2_col_in_219),
    .col_in_220(u2_col_in_220),
    .col_in_221(u2_col_in_221),
    .col_in_222(u2_col_in_222),
    .col_in_223(u2_col_in_223),
    .col_in_224(u2_col_in_224),
    .col_in_225(u2_col_in_225),
    .col_in_226(u2_col_in_226),
    .col_in_227(u2_col_in_227),
    .col_in_228(u2_col_in_228),
    .col_in_229(u2_col_in_229),
    .col_in_230(u2_col_in_230),
    .col_in_231(u2_col_in_231),
    .col_in_232(u2_col_in_232),
    .col_in_233(u2_col_in_233),
    .col_in_234(u2_col_in_234),
    .col_in_235(u2_col_in_235),
    .col_in_236(u2_col_in_236),
    .col_in_237(u2_col_in_237),
    .col_in_238(u2_col_in_238),
    .col_in_239(u2_col_in_239),
    .col_in_240(u2_col_in_240),
    .col_in_241(u2_col_in_241),
    .col_in_242(u2_col_in_242),
    .col_in_243(u2_col_in_243),
    .col_in_244(u2_col_in_244),
    .col_in_245(u2_col_in_245),
    .col_in_246(u2_col_in_246),
    .col_in_247(u2_col_in_247),
    .col_in_248(u2_col_in_248),
    .col_in_249(u2_col_in_249),
    .col_in_250(u2_col_in_250),
    .col_in_251(u2_col_in_251),
    .col_in_252(u2_col_in_252),
    .col_in_253(u2_col_in_253),
    .col_in_254(u2_col_in_254),
    .col_in_255(u2_col_in_255),
    .col_in_256(u2_col_in_256),
    .col_in_257(u2_col_in_257),
    .col_in_258(u2_col_in_258),
    .col_in_259(u2_col_in_259),
    .col_in_260(u2_col_in_260),
    .col_in_261(u2_col_in_261),
    .col_in_262(u2_col_in_262),
    .col_in_263(u2_col_in_263),
    .col_in_264(u2_col_in_264),
    .col_in_265(u2_col_in_265),
    .col_in_266(u2_col_in_266),
    .col_in_267(u2_col_in_267),
    .col_in_268(u2_col_in_268),
    .col_in_269(u2_col_in_269),
    .col_in_270(u2_col_in_270),
    .col_in_271(u2_col_in_271),
    .col_in_272(u2_col_in_272),
    .col_in_273(u2_col_in_273),
    .col_in_274(u2_col_in_274),
    .col_in_275(u2_col_in_275),
    .col_in_276(u2_col_in_276),
    .col_in_277(u2_col_in_277),
    .col_in_278(u2_col_in_278),
    .col_in_279(u2_col_in_279),
    .col_in_280(u2_col_in_280),
    .col_in_281(u2_col_in_281),
    .col_in_282(u2_col_in_282),
    .col_in_283(u2_col_in_283),
    .col_in_284(u2_col_in_284),
    .col_in_285(u2_col_in_285),
    .col_in_286(u2_col_in_286),
    .col_in_287(u2_col_in_287),
    .col_in_288(u2_col_in_288),
    .col_in_289(u2_col_in_289),
    .col_in_290(u2_col_in_290),
    .col_in_291(u2_col_in_291),
    .col_in_292(u2_col_in_292),
    .col_in_293(u2_col_in_293),
    .col_in_294(u2_col_in_294),
    .col_in_295(u2_col_in_295),
    .col_in_296(u2_col_in_296),
    .col_in_297(u2_col_in_297),
    .col_in_298(u2_col_in_298),
    .col_in_299(u2_col_in_299),
    .col_in_300(u2_col_in_300),
    .col_in_301(u2_col_in_301),
    .col_in_302(u2_col_in_302),
    .col_in_303(u2_col_in_303),
    .col_in_304(u2_col_in_304),
    .col_in_305(u2_col_in_305),
    .col_in_306(u2_col_in_306),
    .col_in_307(u2_col_in_307),
    .col_in_308(u2_col_in_308),
    .col_in_309(u2_col_in_309),
    .col_in_310(u2_col_in_310),
    .col_in_311(u2_col_in_311),
    .col_in_312(u2_col_in_312),
    .col_in_313(u2_col_in_313),
    .col_in_314(u2_col_in_314),
    .col_in_315(u2_col_in_315),
    .col_in_316(u2_col_in_316),
    .col_in_317(u2_col_in_317),
    .col_in_318(u2_col_in_318),
    .col_in_319(u2_col_in_319),
    .col_in_320(u2_col_in_320),
    .col_in_321(u2_col_in_321),
    .col_in_322(u2_col_in_322),
    .col_in_323(u2_col_in_323),
    .col_in_324(u2_col_in_324),
    .col_in_325(u2_col_in_325),
    .col_in_326(u2_col_in_326),
    .col_in_327(u2_col_in_327),
    .col_in_328(u2_col_in_328),
    .col_in_329(u2_col_in_329),
    .col_in_330(u2_col_in_330),
    .col_in_331(u2_col_in_331),
    .col_in_332(u2_col_in_332),
    .col_in_333(u2_col_in_333),
    .col_in_334(u2_col_in_334),
    .col_in_335(u2_col_in_335),
    .col_in_336(u2_col_in_336),
    .col_in_337(u2_col_in_337),
    .col_in_338(u2_col_in_338),
    .col_in_339(u2_col_in_339),
    .col_in_340(u2_col_in_340),
    .col_in_341(u2_col_in_341),
    .col_in_342(u2_col_in_342),
    .col_in_343(u2_col_in_343),
    .col_in_344(u2_col_in_344),
    .col_in_345(u2_col_in_345),
    .col_in_346(u2_col_in_346),
    .col_in_347(u2_col_in_347),
    .col_in_348(u2_col_in_348),
    .col_in_349(u2_col_in_349),
    .col_in_350(u2_col_in_350),
    .col_in_351(u2_col_in_351),
    .col_in_352(u2_col_in_352),
    .col_in_353(u2_col_in_353),
    .col_in_354(u2_col_in_354),
    .col_in_355(u2_col_in_355),
    .col_in_356(u2_col_in_356),
    .col_in_357(u2_col_in_357),
    .col_in_358(u2_col_in_358),
    .col_in_359(u2_col_in_359),
    .col_in_360(u2_col_in_360),
    .col_in_361(u2_col_in_361),
    .col_in_362(u2_col_in_362),
    .col_in_363(u2_col_in_363),
    .col_in_364(u2_col_in_364),
    .col_in_365(u2_col_in_365),
    .col_in_366(u2_col_in_366),
    .col_in_367(u2_col_in_367),
    .col_in_368(u2_col_in_368),
    .col_in_369(u2_col_in_369),
    .col_in_370(u2_col_in_370),
    .col_in_371(u2_col_in_371),
    .col_in_372(u2_col_in_372),
    .col_in_373(u2_col_in_373),
    .col_in_374(u2_col_in_374),
    .col_in_375(u2_col_in_375),
    .col_in_376(u2_col_in_376),
    .col_in_377(u2_col_in_377),
    .col_in_378(u2_col_in_378),
    .col_in_379(u2_col_in_379),
    .col_in_380(u2_col_in_380),
    .col_in_381(u2_col_in_381),
    .col_in_382(u2_col_in_382),
    .col_in_383(u2_col_in_383),
    .col_in_384(u2_col_in_384),
    .col_in_385(u2_col_in_385),
    .col_in_386(u2_col_in_386),
    .col_in_387(u2_col_in_387),
    .col_in_388(u2_col_in_388),
    .col_in_389(u2_col_in_389),
    .col_in_390(u2_col_in_390),
    .col_in_391(u2_col_in_391),
    .col_in_392(u2_col_in_392),
    .col_in_393(u2_col_in_393),
    .col_in_394(u2_col_in_394),
    .col_in_395(u2_col_in_395),
    .col_in_396(u2_col_in_396),
    .col_in_397(u2_col_in_397),
    .col_in_398(u2_col_in_398),
    .col_in_399(u2_col_in_399),
    .col_in_400(u2_col_in_400),
    .col_in_401(u2_col_in_401),
    .col_in_402(u2_col_in_402),
    .col_in_403(u2_col_in_403),
    .col_in_404(u2_col_in_404),
    .col_in_405(u2_col_in_405),
    .col_in_406(u2_col_in_406),
    .col_in_407(u2_col_in_407),
    .col_in_408(u2_col_in_408),
    .col_in_409(u2_col_in_409),
    .col_in_410(u2_col_in_410),
    .col_in_411(u2_col_in_411),
    .col_in_412(u2_col_in_412),
    .col_in_413(u2_col_in_413),
    .col_in_414(u2_col_in_414),
    .col_in_415(u2_col_in_415),
    .col_in_416(u2_col_in_416),
    .col_in_417(u2_col_in_417),
    .col_in_418(u2_col_in_418),
    .col_in_419(u2_col_in_419),
    .col_in_420(u2_col_in_420),
    .col_in_421(u2_col_in_421),
    .col_in_422(u2_col_in_422),
    .col_in_423(u2_col_in_423),
    .col_in_424(u2_col_in_424),
    .col_in_425(u2_col_in_425),
    .col_in_426(u2_col_in_426),
    .col_in_427(u2_col_in_427),
    .col_in_428(u2_col_in_428),
    .col_in_429(u2_col_in_429),
    .col_in_430(u2_col_in_430),
    .col_in_431(u2_col_in_431),
    .col_in_432(u2_col_in_432),
    .col_in_433(u2_col_in_433),
    .col_in_434(u2_col_in_434),
    .col_in_435(u2_col_in_435),
    .col_in_436(u2_col_in_436),
    .col_in_437(u2_col_in_437),
    .col_in_438(u2_col_in_438),
    .col_in_439(u2_col_in_439),
    .col_in_440(u2_col_in_440),
    .col_in_441(u2_col_in_441),
    .col_in_442(u2_col_in_442),
    .col_in_443(u2_col_in_443),
    .col_in_444(u2_col_in_444),
    .col_in_445(u2_col_in_445),
    .col_in_446(u2_col_in_446),
    .col_in_447(u2_col_in_447),
    .col_in_448(u2_col_in_448),
    .col_in_449(u2_col_in_449),
    .col_in_450(u2_col_in_450),
    .col_in_451(u2_col_in_451),
    .col_in_452(u2_col_in_452),
    .col_in_453(u2_col_in_453),
    .col_in_454(u2_col_in_454),
    .col_in_455(u2_col_in_455),
    .col_in_456(u2_col_in_456),
    .col_in_457(u2_col_in_457),
    .col_in_458(u2_col_in_458),
    .col_in_459(u2_col_in_459),
    .col_in_460(u2_col_in_460),
    .col_in_461(u2_col_in_461),
    .col_in_462(u2_col_in_462),
    .col_in_463(u2_col_in_463),
    .col_in_464(u2_col_in_464),
    .col_in_465(u2_col_in_465),
    .col_in_466(u2_col_in_466),
    .col_in_467(u2_col_in_467),
    .col_in_468(u2_col_in_468),
    .col_in_469(u2_col_in_469),
    .col_in_470(u2_col_in_470),
    .col_in_471(u2_col_in_471),
    .col_in_472(u2_col_in_472),
    .col_in_473(u2_col_in_473),
    .col_in_474(u2_col_in_474),
    .col_in_475(u2_col_in_475),
    .col_in_476(u2_col_in_476),
    .col_in_477(u2_col_in_477),
    .col_in_478(u2_col_in_478),
    .col_in_479(u2_col_in_479),
    .col_in_480(u2_col_in_480),
    .col_in_481(u2_col_in_481),
    .col_in_482(u2_col_in_482),
    .col_in_483(u2_col_in_483),
    .col_in_484(u2_col_in_484),
    .col_in_485(u2_col_in_485),
    .col_in_486(u2_col_in_486),
    .col_in_487(u2_col_in_487),
    .col_in_488(u2_col_in_488),
    .col_in_489(u2_col_in_489),
    .col_in_490(u2_col_in_490),
    .col_in_491(u2_col_in_491),
    .col_in_492(u2_col_in_492),
    .col_in_493(u2_col_in_493),
    .col_in_494(u2_col_in_494),
    .col_in_495(u2_col_in_495),
    .col_in_496(u2_col_in_496),
    .col_in_497(u2_col_in_497),
    .col_in_498(u2_col_in_498),
    .col_in_499(u2_col_in_499),
    .col_in_500(u2_col_in_500),
    .col_in_501(u2_col_in_501),
    .col_in_502(u2_col_in_502),
    .col_in_503(u2_col_in_503),
    .col_in_504(u2_col_in_504),
    .col_in_505(u2_col_in_505),
    .col_in_506(u2_col_in_506),
    .col_in_507(u2_col_in_507),
    .col_in_508(u2_col_in_508),
    .col_in_509(u2_col_in_509),
    .col_in_510(u2_col_in_510),
    .col_in_511(u2_col_in_511),
    .col_in_512(u2_col_in_512),
    .col_in_513(u2_col_in_513),
    .col_in_514(u2_col_in_514),
    .col_in_515(u2_col_in_515),
    .col_in_516(u2_col_in_516),
    .col_in_517(u2_col_in_517),
    .col_in_518(u2_col_in_518),
    .col_in_519(u2_col_in_519),
    .col_in_520(u2_col_in_520),
    .col_in_521(u2_col_in_521),
    .col_in_522(u2_col_in_522),
    .col_in_523(u2_col_in_523),
    .col_in_524(u2_col_in_524),
    .col_in_525(u2_col_in_525),
    .col_in_526(u2_col_in_526),
    .col_in_527(u2_col_in_527),
    .col_in_528(u2_col_in_528),
    .col_in_529(u2_col_in_529),
    .col_in_530(u2_col_in_530),
    .col_in_531(u2_col_in_531),
    .col_in_532(u2_col_in_532),
    .col_in_533(u2_col_in_533),
    .col_in_534(u2_col_in_534),
    .col_in_535(u2_col_in_535),
    .col_in_536(u2_col_in_536),
    .col_in_537(u2_col_in_537),
    .col_in_538(u2_col_in_538),
    .col_in_539(u2_col_in_539),
    .col_in_540(u2_col_in_540),
    .col_in_541(u2_col_in_541),
    .col_in_542(u2_col_in_542),
    .col_in_543(u2_col_in_543),
    .col_in_544(u2_col_in_544),
    .col_in_545(u2_col_in_545),
    .col_in_546(u2_col_in_546),
    .col_in_547(u2_col_in_547),
    .col_in_548(u2_col_in_548),
    .col_in_549(u2_col_in_549),
    .col_in_550(u2_col_in_550),
    .col_in_551(u2_col_in_551),
    .col_in_552(u2_col_in_552),
    .col_in_553(u2_col_in_553),
    .col_in_554(u2_col_in_554),
    .col_in_555(u2_col_in_555),
    .col_in_556(u2_col_in_556),
    .col_in_557(u2_col_in_557),
    .col_in_558(u2_col_in_558),
    .col_in_559(u2_col_in_559),
    .col_in_560(u2_col_in_560),
    .col_in_561(u2_col_in_561),
    .col_in_562(u2_col_in_562),
    .col_in_563(u2_col_in_563),
    .col_in_564(u2_col_in_564),
    .col_in_565(u2_col_in_565),
    .col_in_566(u2_col_in_566),
    .col_in_567(u2_col_in_567),
    .col_in_568(u2_col_in_568),
    .col_in_569(u2_col_in_569),
    .col_in_570(u2_col_in_570),
    .col_in_571(u2_col_in_571),
    .col_in_572(u2_col_in_572),
    .col_in_573(u2_col_in_573),
    .col_in_574(u2_col_in_574),
    .col_in_575(u2_col_in_575),
    .col_in_576(u2_col_in_576),
    .col_in_577(u2_col_in_577),
    .col_in_578(u2_col_in_578),
    .col_in_579(u2_col_in_579),
    .col_in_580(u2_col_in_580),
    .col_in_581(u2_col_in_581),
    .col_in_582(u2_col_in_582),
    .col_in_583(u2_col_in_583),
    .col_in_584(u2_col_in_584),
    .col_in_585(u2_col_in_585),
    .col_in_586(u2_col_in_586),
    .col_in_587(u2_col_in_587),
    .col_in_588(u2_col_in_588),
    .col_in_589(u2_col_in_589),
    .col_in_590(u2_col_in_590),
    .col_in_591(u2_col_in_591),
    .col_in_592(u2_col_in_592),
    .col_in_593(u2_col_in_593),
    .col_in_594(u2_col_in_594),
    .col_in_595(u2_col_in_595),
    .col_in_596(u2_col_in_596),
    .col_in_597(u2_col_in_597),
    .col_in_598(u2_col_in_598),
    .col_in_599(u2_col_in_599),
    .col_in_600(u2_col_in_600),
    .col_in_601(u2_col_in_601),
    .col_in_602(u2_col_in_602),
    .col_in_603(u2_col_in_603),
    .col_in_604(u2_col_in_604),
    .col_in_605(u2_col_in_605),
    .col_in_606(u2_col_in_606),
    .col_in_607(u2_col_in_607),
    .col_in_608(u2_col_in_608),
    .col_in_609(u2_col_in_609),
    .col_in_610(u2_col_in_610),
    .col_in_611(u2_col_in_611),
    .col_in_612(u2_col_in_612),
    .col_in_613(u2_col_in_613),
    .col_in_614(u2_col_in_614),
    .col_in_615(u2_col_in_615),
    .col_in_616(u2_col_in_616),
    .col_in_617(u2_col_in_617),
    .col_in_618(u2_col_in_618),
    .col_in_619(u2_col_in_619),
    .col_in_620(u2_col_in_620),
    .col_in_621(u2_col_in_621),
    .col_in_622(u2_col_in_622),
    .col_in_623(u2_col_in_623),
    .col_in_624(u2_col_in_624),
    .col_in_625(u2_col_in_625),
    .col_in_626(u2_col_in_626),
    .col_in_627(u2_col_in_627),
    .col_in_628(u2_col_in_628),
    .col_in_629(u2_col_in_629),
    .col_in_630(u2_col_in_630),
    .col_in_631(u2_col_in_631),
    .col_in_632(u2_col_in_632),
    .col_in_633(u2_col_in_633),
    .col_in_634(u2_col_in_634),
    .col_in_635(u2_col_in_635),
    .col_in_636(u2_col_in_636),
    .col_in_637(u2_col_in_637),
    .col_in_638(u2_col_in_638),
    .col_in_639(u2_col_in_639),
    .col_in_640(u2_col_in_640),
    .col_in_641(u2_col_in_641),
    .col_in_642(u2_col_in_642),
    .col_in_643(u2_col_in_643),
    .col_in_644(u2_col_in_644),
    .col_in_645(u2_col_in_645),
    .col_in_646(u2_col_in_646),
    .col_in_647(u2_col_in_647),
    .col_in_648(u2_col_in_648),
    .col_in_649(u2_col_in_649),
    .col_in_650(u2_col_in_650),
    .col_in_651(u2_col_in_651),
    .col_in_652(u2_col_in_652),
    .col_in_653(u2_col_in_653),
    .col_in_654(u2_col_in_654),
    .col_in_655(u2_col_in_655),
    .col_in_656(u2_col_in_656),
    .col_in_657(u2_col_in_657),
    .col_in_658(u2_col_in_658),
    .col_in_659(u2_col_in_659),
    .col_in_660(u2_col_in_660),
    .col_in_661(u2_col_in_661),
    .col_in_662(u2_col_in_662),
    .col_in_663(u2_col_in_663),
    .col_in_664(u2_col_in_664),
    .col_in_665(u2_col_in_665),
    .col_in_666(u2_col_in_666),
    .col_in_667(u2_col_in_667),
    .col_in_668(u2_col_in_668),
    .col_in_669(u2_col_in_669),
    .col_in_670(u2_col_in_670),
    .col_in_671(u2_col_in_671),
    .col_in_672(u2_col_in_672),
    .col_in_673(u2_col_in_673),
    .col_in_674(u2_col_in_674),
    .col_in_675(u2_col_in_675),
    .col_in_676(u2_col_in_676),
    .col_in_677(u2_col_in_677),
    .col_in_678(u2_col_in_678),
    .col_in_679(u2_col_in_679),
    .col_in_680(u2_col_in_680),
    .col_in_681(u2_col_in_681),
    .col_in_682(u2_col_in_682),
    .col_in_683(u2_col_in_683),
    .col_in_684(u2_col_in_684),
    .col_in_685(u2_col_in_685),
    .col_in_686(u2_col_in_686),
    .col_in_687(u2_col_in_687),
    .col_in_688(u2_col_in_688),
    .col_in_689(u2_col_in_689),
    .col_in_690(u2_col_in_690),
    .col_in_691(u2_col_in_691),
    .col_in_692(u2_col_in_692),
    .col_in_693(u2_col_in_693),
    .col_in_694(u2_col_in_694),
    .col_in_695(u2_col_in_695),
    .col_in_696(u2_col_in_696),
    .col_in_697(u2_col_in_697),
    .col_in_698(u2_col_in_698),
    .col_in_699(u2_col_in_699),
    .col_in_700(u2_col_in_700),
    .col_in_701(u2_col_in_701),
    .col_in_702(u2_col_in_702),
    .col_in_703(u2_col_in_703),
    .col_in_704(u2_col_in_704),
    .col_in_705(u2_col_in_705),
    .col_in_706(u2_col_in_706),
    .col_in_707(u2_col_in_707),
    .col_in_708(u2_col_in_708),
    .col_in_709(u2_col_in_709),
    .col_in_710(u2_col_in_710),
    .col_in_711(u2_col_in_711),
    .col_in_712(u2_col_in_712),
    .col_in_713(u2_col_in_713),
    .col_in_714(u2_col_in_714),
    .col_in_715(u2_col_in_715),
    .col_in_716(u2_col_in_716),
    .col_in_717(u2_col_in_717),
    .col_in_718(u2_col_in_718),
    .col_in_719(u2_col_in_719),
    .col_in_720(u2_col_in_720),
    .col_in_721(u2_col_in_721),
    .col_in_722(u2_col_in_722),
    .col_in_723(u2_col_in_723),
    .col_in_724(u2_col_in_724),
    .col_in_725(u2_col_in_725),
    .col_in_726(u2_col_in_726),
    .col_in_727(u2_col_in_727),
    .col_in_728(u2_col_in_728),
    .col_in_729(u2_col_in_729),
    .col_in_730(u2_col_in_730),
    .col_in_731(u2_col_in_731),
    .col_in_732(u2_col_in_732),
    .col_in_733(u2_col_in_733),
    .col_in_734(u2_col_in_734),
    .col_in_735(u2_col_in_735),
    .col_in_736(u2_col_in_736),
    .col_in_737(u2_col_in_737),
    .col_in_738(u2_col_in_738),
    .col_in_739(u2_col_in_739),
    .col_in_740(u2_col_in_740),
    .col_in_741(u2_col_in_741),
    .col_in_742(u2_col_in_742),
    .col_in_743(u2_col_in_743),
    .col_in_744(u2_col_in_744),
    .col_in_745(u2_col_in_745),
    .col_in_746(u2_col_in_746),
    .col_in_747(u2_col_in_747),
    .col_in_748(u2_col_in_748),
    .col_in_749(u2_col_in_749),
    .col_in_750(u2_col_in_750),
    .col_in_751(u2_col_in_751),
    .col_in_752(u2_col_in_752),
    .col_in_753(u2_col_in_753),
    .col_in_754(u2_col_in_754),
    .col_in_755(u2_col_in_755),
    .col_in_756(u2_col_in_756),
    .col_in_757(u2_col_in_757),
    .col_in_758(u2_col_in_758),
    .col_in_759(u2_col_in_759),
    .col_in_760(u2_col_in_760),
    .col_in_761(u2_col_in_761),
    .col_in_762(u2_col_in_762),
    .col_in_763(u2_col_in_763),
    .col_in_764(u2_col_in_764),
    .col_in_765(u2_col_in_765),
    .col_in_766(u2_col_in_766),
    .col_in_767(u2_col_in_767),
    .col_in_768(u2_col_in_768),
    .col_in_769(u2_col_in_769),
    .col_in_770(u2_col_in_770),
    .col_in_771(u2_col_in_771),
    .col_in_772(u2_col_in_772),
    .col_in_773(u2_col_in_773),
    .col_in_774(u2_col_in_774),
    .col_in_775(u2_col_in_775),
    .col_in_776(u2_col_in_776),
    .col_in_777(u2_col_in_777),
    .col_in_778(u2_col_in_778),
    .col_in_779(u2_col_in_779),
    .col_in_780(u2_col_in_780),
    .col_in_781(u2_col_in_781),
    .col_in_782(u2_col_in_782),
    .col_in_783(u2_col_in_783),
    .col_in_784(u2_col_in_784),
    .col_in_785(u2_col_in_785),
    .col_in_786(u2_col_in_786),
    .col_in_787(u2_col_in_787),
    .col_in_788(u2_col_in_788),
    .col_in_789(u2_col_in_789),
    .col_in_790(u2_col_in_790),
    .col_in_791(u2_col_in_791),
    .col_in_792(u2_col_in_792),
    .col_in_793(u2_col_in_793),
    .col_in_794(u2_col_in_794),
    .col_in_795(u2_col_in_795),
    .col_in_796(u2_col_in_796),
    .col_in_797(u2_col_in_797),
    .col_in_798(u2_col_in_798),
    .col_in_799(u2_col_in_799),
    .col_in_800(u2_col_in_800),
    .col_in_801(u2_col_in_801),
    .col_in_802(u2_col_in_802),
    .col_in_803(u2_col_in_803),
    .col_in_804(u2_col_in_804),
    .col_in_805(u2_col_in_805),
    .col_in_806(u2_col_in_806),
    .col_in_807(u2_col_in_807),
    .col_in_808(u2_col_in_808),
    .col_in_809(u2_col_in_809),
    .col_in_810(u2_col_in_810),
    .col_in_811(u2_col_in_811),
    .col_in_812(u2_col_in_812),
    .col_in_813(u2_col_in_813),
    .col_in_814(u2_col_in_814),
    .col_in_815(u2_col_in_815),
    .col_in_816(u2_col_in_816),
    .col_in_817(u2_col_in_817),
    .col_in_818(u2_col_in_818),
    .col_in_819(u2_col_in_819),
    .col_in_820(u2_col_in_820),
    .col_in_821(u2_col_in_821),
    .col_in_822(u2_col_in_822),
    .col_in_823(u2_col_in_823),
    .col_in_824(u2_col_in_824),
    .col_in_825(u2_col_in_825),
    .col_in_826(u2_col_in_826),
    .col_in_827(u2_col_in_827),
    .col_in_828(u2_col_in_828),
    .col_in_829(u2_col_in_829),
    .col_in_830(u2_col_in_830),
    .col_in_831(u2_col_in_831),
    .col_in_832(u2_col_in_832),
    .col_in_833(u2_col_in_833),
    .col_in_834(u2_col_in_834),
    .col_in_835(u2_col_in_835),
    .col_in_836(u2_col_in_836),
    .col_in_837(u2_col_in_837),
    .col_in_838(u2_col_in_838),
    .col_in_839(u2_col_in_839),
    .col_in_840(u2_col_in_840),
    .col_in_841(u2_col_in_841),
    .col_in_842(u2_col_in_842),
    .col_in_843(u2_col_in_843),
    .col_in_844(u2_col_in_844),
    .col_in_845(u2_col_in_845),
    .col_in_846(u2_col_in_846),
    .col_in_847(u2_col_in_847),
    .col_in_848(u2_col_in_848),
    .col_in_849(u2_col_in_849),
    .col_in_850(u2_col_in_850),
    .col_in_851(u2_col_in_851),
    .col_in_852(u2_col_in_852),
    .col_in_853(u2_col_in_853),
    .col_in_854(u2_col_in_854),
    .col_in_855(u2_col_in_855),
    .col_in_856(u2_col_in_856),
    .col_in_857(u2_col_in_857),
    .col_in_858(u2_col_in_858),
    .col_in_859(u2_col_in_859),
    .col_in_860(u2_col_in_860),
    .col_in_861(u2_col_in_861),
    .col_in_862(u2_col_in_862),
    .col_in_863(u2_col_in_863),
    .col_in_864(u2_col_in_864),
    .col_in_865(u2_col_in_865),
    .col_in_866(u2_col_in_866),
    .col_in_867(u2_col_in_867),
    .col_in_868(u2_col_in_868),
    .col_in_869(u2_col_in_869),
    .col_in_870(u2_col_in_870),
    .col_in_871(u2_col_in_871),
    .col_in_872(u2_col_in_872),
    .col_in_873(u2_col_in_873),
    .col_in_874(u2_col_in_874),
    .col_in_875(u2_col_in_875),
    .col_in_876(u2_col_in_876),
    .col_in_877(u2_col_in_877),
    .col_in_878(u2_col_in_878),
    .col_in_879(u2_col_in_879),
    .col_in_880(u2_col_in_880),
    .col_in_881(u2_col_in_881),
    .col_in_882(u2_col_in_882),
    .col_in_883(u2_col_in_883),
    .col_in_884(u2_col_in_884),
    .col_in_885(u2_col_in_885),
    .col_in_886(u2_col_in_886),
    .col_in_887(u2_col_in_887),
    .col_in_888(u2_col_in_888),
    .col_in_889(u2_col_in_889),
    .col_in_890(u2_col_in_890),
    .col_in_891(u2_col_in_891),
    .col_in_892(u2_col_in_892),
    .col_in_893(u2_col_in_893),
    .col_in_894(u2_col_in_894),
    .col_in_895(u2_col_in_895),
    .col_in_896(u2_col_in_896),
    .col_in_897(u2_col_in_897),
    .col_in_898(u2_col_in_898),
    .col_in_899(u2_col_in_899),
    .col_in_900(u2_col_in_900),
    .col_in_901(u2_col_in_901),
    .col_in_902(u2_col_in_902),
    .col_in_903(u2_col_in_903),
    .col_in_904(u2_col_in_904),
    .col_in_905(u2_col_in_905),
    .col_in_906(u2_col_in_906),
    .col_in_907(u2_col_in_907),
    .col_in_908(u2_col_in_908),
    .col_in_909(u2_col_in_909),
    .col_in_910(u2_col_in_910),
    .col_in_911(u2_col_in_911),
    .col_in_912(u2_col_in_912),
    .col_in_913(u2_col_in_913),
    .col_in_914(u2_col_in_914),
    .col_in_915(u2_col_in_915),
    .col_in_916(u2_col_in_916),
    .col_in_917(u2_col_in_917),
    .col_in_918(u2_col_in_918),
    .col_in_919(u2_col_in_919),
    .col_in_920(u2_col_in_920),
    .col_in_921(u2_col_in_921),
    .col_in_922(u2_col_in_922),
    .col_in_923(u2_col_in_923),
    .col_in_924(u2_col_in_924),
    .col_in_925(u2_col_in_925),
    .col_in_926(u2_col_in_926),
    .col_in_927(u2_col_in_927),
    .col_in_928(u2_col_in_928),
    .col_in_929(u2_col_in_929),
    .col_in_930(u2_col_in_930),
    .col_in_931(u2_col_in_931),
    .col_in_932(u2_col_in_932),
    .col_in_933(u2_col_in_933),
    .col_in_934(u2_col_in_934),
    .col_in_935(u2_col_in_935),
    .col_in_936(u2_col_in_936),
    .col_in_937(u2_col_in_937),
    .col_in_938(u2_col_in_938),
    .col_in_939(u2_col_in_939),
    .col_in_940(u2_col_in_940),
    .col_in_941(u2_col_in_941),
    .col_in_942(u2_col_in_942),
    .col_in_943(u2_col_in_943),
    .col_in_944(u2_col_in_944),
    .col_in_945(u2_col_in_945),
    .col_in_946(u2_col_in_946),
    .col_in_947(u2_col_in_947),
    .col_in_948(u2_col_in_948),
    .col_in_949(u2_col_in_949),
    .col_in_950(u2_col_in_950),
    .col_in_951(u2_col_in_951),
    .col_in_952(u2_col_in_952),
    .col_in_953(u2_col_in_953),
    .col_in_954(u2_col_in_954),
    .col_in_955(u2_col_in_955),
    .col_in_956(u2_col_in_956),
    .col_in_957(u2_col_in_957),
    .col_in_958(u2_col_in_958),
    .col_in_959(u2_col_in_959),
    .col_in_960(u2_col_in_960),
    .col_in_961(u2_col_in_961),
    .col_in_962(u2_col_in_962),
    .col_in_963(u2_col_in_963),
    .col_in_964(u2_col_in_964),
    .col_in_965(u2_col_in_965),
    .col_in_966(u2_col_in_966),
    .col_in_967(u2_col_in_967),
    .col_in_968(u2_col_in_968),
    .col_in_969(u2_col_in_969),
    .col_in_970(u2_col_in_970),
    .col_in_971(u2_col_in_971),
    .col_in_972(u2_col_in_972),
    .col_in_973(u2_col_in_973),
    .col_in_974(u2_col_in_974),
    .col_in_975(u2_col_in_975),
    .col_in_976(u2_col_in_976),
    .col_in_977(u2_col_in_977),
    .col_in_978(u2_col_in_978),
    .col_in_979(u2_col_in_979),
    .col_in_980(u2_col_in_980),
    .col_in_981(u2_col_in_981),
    .col_in_982(u2_col_in_982),
    .col_in_983(u2_col_in_983),
    .col_in_984(u2_col_in_984),
    .col_in_985(u2_col_in_985),
    .col_in_986(u2_col_in_986),
    .col_in_987(u2_col_in_987),
    .col_in_988(u2_col_in_988),
    .col_in_989(u2_col_in_989),
    .col_in_990(u2_col_in_990),
    .col_in_991(u2_col_in_991),
    .col_in_992(u2_col_in_992),
    .col_in_993(u2_col_in_993),
    .col_in_994(u2_col_in_994),
    .col_in_995(u2_col_in_995),
    .col_in_996(u2_col_in_996),
    .col_in_997(u2_col_in_997),
    .col_in_998(u2_col_in_998),
    .col_in_999(u2_col_in_999),
    .col_in_1000(u2_col_in_1000),
    .col_in_1001(u2_col_in_1001),
    .col_in_1002(u2_col_in_1002),
    .col_in_1003(u2_col_in_1003),
    .col_in_1004(u2_col_in_1004),
    .col_in_1005(u2_col_in_1005),
    .col_in_1006(u2_col_in_1006),
    .col_in_1007(u2_col_in_1007),
    .col_in_1008(u2_col_in_1008),
    .col_in_1009(u2_col_in_1009),
    .col_in_1010(u2_col_in_1010),
    .col_in_1011(u2_col_in_1011),
    .col_in_1012(u2_col_in_1012),
    .col_in_1013(u2_col_in_1013),
    .col_in_1014(u2_col_in_1014),
    .col_in_1015(u2_col_in_1015),
    .col_in_1016(u2_col_in_1016),
    .col_in_1017(u2_col_in_1017),
    .col_in_1018(u2_col_in_1018),
    .col_in_1019(u2_col_in_1019),
    .col_in_1020(u2_col_in_1020),
    .col_in_1021(u2_col_in_1021),
    .col_in_1022(u2_col_in_1022),
    .col_in_1023(u2_col_in_1023),
    .col_in_1024(u2_col_in_1024),
    .col_in_1025(u2_col_in_1025),
    .col_in_1026(u2_col_in_1026),
    .col_in_1027(u2_col_in_1027),
    .col_in_1028(u2_col_in_1028),
    .col_in_1029(u2_col_in_1029),

    .col_out_0(u2_col_out_0),
    .col_out_1(u2_col_out_1),
    .col_out_2(u2_col_out_2),
    .col_out_3(u2_col_out_3),
    .col_out_4(u2_col_out_4),
    .col_out_5(u2_col_out_5),
    .col_out_6(u2_col_out_6),
    .col_out_7(u2_col_out_7),
    .col_out_8(u2_col_out_8),
    .col_out_9(u2_col_out_9),
    .col_out_10(u2_col_out_10),
    .col_out_11(u2_col_out_11),
    .col_out_12(u2_col_out_12),
    .col_out_13(u2_col_out_13),
    .col_out_14(u2_col_out_14),
    .col_out_15(u2_col_out_15),
    .col_out_16(u2_col_out_16),
    .col_out_17(u2_col_out_17),
    .col_out_18(u2_col_out_18),
    .col_out_19(u2_col_out_19),
    .col_out_20(u2_col_out_20),
    .col_out_21(u2_col_out_21),
    .col_out_22(u2_col_out_22),
    .col_out_23(u2_col_out_23),
    .col_out_24(u2_col_out_24),
    .col_out_25(u2_col_out_25),
    .col_out_26(u2_col_out_26),
    .col_out_27(u2_col_out_27),
    .col_out_28(u2_col_out_28),
    .col_out_29(u2_col_out_29),
    .col_out_30(u2_col_out_30),
    .col_out_31(u2_col_out_31),
    .col_out_32(u2_col_out_32),
    .col_out_33(u2_col_out_33),
    .col_out_34(u2_col_out_34),
    .col_out_35(u2_col_out_35),
    .col_out_36(u2_col_out_36),
    .col_out_37(u2_col_out_37),
    .col_out_38(u2_col_out_38),
    .col_out_39(u2_col_out_39),
    .col_out_40(u2_col_out_40),
    .col_out_41(u2_col_out_41),
    .col_out_42(u2_col_out_42),
    .col_out_43(u2_col_out_43),
    .col_out_44(u2_col_out_44),
    .col_out_45(u2_col_out_45),
    .col_out_46(u2_col_out_46),
    .col_out_47(u2_col_out_47),
    .col_out_48(u2_col_out_48),
    .col_out_49(u2_col_out_49),
    .col_out_50(u2_col_out_50),
    .col_out_51(u2_col_out_51),
    .col_out_52(u2_col_out_52),
    .col_out_53(u2_col_out_53),
    .col_out_54(u2_col_out_54),
    .col_out_55(u2_col_out_55),
    .col_out_56(u2_col_out_56),
    .col_out_57(u2_col_out_57),
    .col_out_58(u2_col_out_58),
    .col_out_59(u2_col_out_59),
    .col_out_60(u2_col_out_60),
    .col_out_61(u2_col_out_61),
    .col_out_62(u2_col_out_62),
    .col_out_63(u2_col_out_63),
    .col_out_64(u2_col_out_64),
    .col_out_65(u2_col_out_65),
    .col_out_66(u2_col_out_66),
    .col_out_67(u2_col_out_67),
    .col_out_68(u2_col_out_68),
    .col_out_69(u2_col_out_69),
    .col_out_70(u2_col_out_70),
    .col_out_71(u2_col_out_71),
    .col_out_72(u2_col_out_72),
    .col_out_73(u2_col_out_73),
    .col_out_74(u2_col_out_74),
    .col_out_75(u2_col_out_75),
    .col_out_76(u2_col_out_76),
    .col_out_77(u2_col_out_77),
    .col_out_78(u2_col_out_78),
    .col_out_79(u2_col_out_79),
    .col_out_80(u2_col_out_80),
    .col_out_81(u2_col_out_81),
    .col_out_82(u2_col_out_82),
    .col_out_83(u2_col_out_83),
    .col_out_84(u2_col_out_84),
    .col_out_85(u2_col_out_85),
    .col_out_86(u2_col_out_86),
    .col_out_87(u2_col_out_87),
    .col_out_88(u2_col_out_88),
    .col_out_89(u2_col_out_89),
    .col_out_90(u2_col_out_90),
    .col_out_91(u2_col_out_91),
    .col_out_92(u2_col_out_92),
    .col_out_93(u2_col_out_93),
    .col_out_94(u2_col_out_94),
    .col_out_95(u2_col_out_95),
    .col_out_96(u2_col_out_96),
    .col_out_97(u2_col_out_97),
    .col_out_98(u2_col_out_98),
    .col_out_99(u2_col_out_99),
    .col_out_100(u2_col_out_100),
    .col_out_101(u2_col_out_101),
    .col_out_102(u2_col_out_102),
    .col_out_103(u2_col_out_103),
    .col_out_104(u2_col_out_104),
    .col_out_105(u2_col_out_105),
    .col_out_106(u2_col_out_106),
    .col_out_107(u2_col_out_107),
    .col_out_108(u2_col_out_108),
    .col_out_109(u2_col_out_109),
    .col_out_110(u2_col_out_110),
    .col_out_111(u2_col_out_111),
    .col_out_112(u2_col_out_112),
    .col_out_113(u2_col_out_113),
    .col_out_114(u2_col_out_114),
    .col_out_115(u2_col_out_115),
    .col_out_116(u2_col_out_116),
    .col_out_117(u2_col_out_117),
    .col_out_118(u2_col_out_118),
    .col_out_119(u2_col_out_119),
    .col_out_120(u2_col_out_120),
    .col_out_121(u2_col_out_121),
    .col_out_122(u2_col_out_122),
    .col_out_123(u2_col_out_123),
    .col_out_124(u2_col_out_124),
    .col_out_125(u2_col_out_125),
    .col_out_126(u2_col_out_126),
    .col_out_127(u2_col_out_127),
    .col_out_128(u2_col_out_128),
    .col_out_129(u2_col_out_129),
    .col_out_130(u2_col_out_130),
    .col_out_131(u2_col_out_131),
    .col_out_132(u2_col_out_132),
    .col_out_133(u2_col_out_133),
    .col_out_134(u2_col_out_134),
    .col_out_135(u2_col_out_135),
    .col_out_136(u2_col_out_136),
    .col_out_137(u2_col_out_137),
    .col_out_138(u2_col_out_138),
    .col_out_139(u2_col_out_139),
    .col_out_140(u2_col_out_140),
    .col_out_141(u2_col_out_141),
    .col_out_142(u2_col_out_142),
    .col_out_143(u2_col_out_143),
    .col_out_144(u2_col_out_144),
    .col_out_145(u2_col_out_145),
    .col_out_146(u2_col_out_146),
    .col_out_147(u2_col_out_147),
    .col_out_148(u2_col_out_148),
    .col_out_149(u2_col_out_149),
    .col_out_150(u2_col_out_150),
    .col_out_151(u2_col_out_151),
    .col_out_152(u2_col_out_152),
    .col_out_153(u2_col_out_153),
    .col_out_154(u2_col_out_154),
    .col_out_155(u2_col_out_155),
    .col_out_156(u2_col_out_156),
    .col_out_157(u2_col_out_157),
    .col_out_158(u2_col_out_158),
    .col_out_159(u2_col_out_159),
    .col_out_160(u2_col_out_160),
    .col_out_161(u2_col_out_161),
    .col_out_162(u2_col_out_162),
    .col_out_163(u2_col_out_163),
    .col_out_164(u2_col_out_164),
    .col_out_165(u2_col_out_165),
    .col_out_166(u2_col_out_166),
    .col_out_167(u2_col_out_167),
    .col_out_168(u2_col_out_168),
    .col_out_169(u2_col_out_169),
    .col_out_170(u2_col_out_170),
    .col_out_171(u2_col_out_171),
    .col_out_172(u2_col_out_172),
    .col_out_173(u2_col_out_173),
    .col_out_174(u2_col_out_174),
    .col_out_175(u2_col_out_175),
    .col_out_176(u2_col_out_176),
    .col_out_177(u2_col_out_177),
    .col_out_178(u2_col_out_178),
    .col_out_179(u2_col_out_179),
    .col_out_180(u2_col_out_180),
    .col_out_181(u2_col_out_181),
    .col_out_182(u2_col_out_182),
    .col_out_183(u2_col_out_183),
    .col_out_184(u2_col_out_184),
    .col_out_185(u2_col_out_185),
    .col_out_186(u2_col_out_186),
    .col_out_187(u2_col_out_187),
    .col_out_188(u2_col_out_188),
    .col_out_189(u2_col_out_189),
    .col_out_190(u2_col_out_190),
    .col_out_191(u2_col_out_191),
    .col_out_192(u2_col_out_192),
    .col_out_193(u2_col_out_193),
    .col_out_194(u2_col_out_194),
    .col_out_195(u2_col_out_195),
    .col_out_196(u2_col_out_196),
    .col_out_197(u2_col_out_197),
    .col_out_198(u2_col_out_198),
    .col_out_199(u2_col_out_199),
    .col_out_200(u2_col_out_200),
    .col_out_201(u2_col_out_201),
    .col_out_202(u2_col_out_202),
    .col_out_203(u2_col_out_203),
    .col_out_204(u2_col_out_204),
    .col_out_205(u2_col_out_205),
    .col_out_206(u2_col_out_206),
    .col_out_207(u2_col_out_207),
    .col_out_208(u2_col_out_208),
    .col_out_209(u2_col_out_209),
    .col_out_210(u2_col_out_210),
    .col_out_211(u2_col_out_211),
    .col_out_212(u2_col_out_212),
    .col_out_213(u2_col_out_213),
    .col_out_214(u2_col_out_214),
    .col_out_215(u2_col_out_215),
    .col_out_216(u2_col_out_216),
    .col_out_217(u2_col_out_217),
    .col_out_218(u2_col_out_218),
    .col_out_219(u2_col_out_219),
    .col_out_220(u2_col_out_220),
    .col_out_221(u2_col_out_221),
    .col_out_222(u2_col_out_222),
    .col_out_223(u2_col_out_223),
    .col_out_224(u2_col_out_224),
    .col_out_225(u2_col_out_225),
    .col_out_226(u2_col_out_226),
    .col_out_227(u2_col_out_227),
    .col_out_228(u2_col_out_228),
    .col_out_229(u2_col_out_229),
    .col_out_230(u2_col_out_230),
    .col_out_231(u2_col_out_231),
    .col_out_232(u2_col_out_232),
    .col_out_233(u2_col_out_233),
    .col_out_234(u2_col_out_234),
    .col_out_235(u2_col_out_235),
    .col_out_236(u2_col_out_236),
    .col_out_237(u2_col_out_237),
    .col_out_238(u2_col_out_238),
    .col_out_239(u2_col_out_239),
    .col_out_240(u2_col_out_240),
    .col_out_241(u2_col_out_241),
    .col_out_242(u2_col_out_242),
    .col_out_243(u2_col_out_243),
    .col_out_244(u2_col_out_244),
    .col_out_245(u2_col_out_245),
    .col_out_246(u2_col_out_246),
    .col_out_247(u2_col_out_247),
    .col_out_248(u2_col_out_248),
    .col_out_249(u2_col_out_249),
    .col_out_250(u2_col_out_250),
    .col_out_251(u2_col_out_251),
    .col_out_252(u2_col_out_252),
    .col_out_253(u2_col_out_253),
    .col_out_254(u2_col_out_254),
    .col_out_255(u2_col_out_255),
    .col_out_256(u2_col_out_256),
    .col_out_257(u2_col_out_257),
    .col_out_258(u2_col_out_258),
    .col_out_259(u2_col_out_259),
    .col_out_260(u2_col_out_260),
    .col_out_261(u2_col_out_261),
    .col_out_262(u2_col_out_262),
    .col_out_263(u2_col_out_263),
    .col_out_264(u2_col_out_264),
    .col_out_265(u2_col_out_265),
    .col_out_266(u2_col_out_266),
    .col_out_267(u2_col_out_267),
    .col_out_268(u2_col_out_268),
    .col_out_269(u2_col_out_269),
    .col_out_270(u2_col_out_270),
    .col_out_271(u2_col_out_271),
    .col_out_272(u2_col_out_272),
    .col_out_273(u2_col_out_273),
    .col_out_274(u2_col_out_274),
    .col_out_275(u2_col_out_275),
    .col_out_276(u2_col_out_276),
    .col_out_277(u2_col_out_277),
    .col_out_278(u2_col_out_278),
    .col_out_279(u2_col_out_279),
    .col_out_280(u2_col_out_280),
    .col_out_281(u2_col_out_281),
    .col_out_282(u2_col_out_282),
    .col_out_283(u2_col_out_283),
    .col_out_284(u2_col_out_284),
    .col_out_285(u2_col_out_285),
    .col_out_286(u2_col_out_286),
    .col_out_287(u2_col_out_287),
    .col_out_288(u2_col_out_288),
    .col_out_289(u2_col_out_289),
    .col_out_290(u2_col_out_290),
    .col_out_291(u2_col_out_291),
    .col_out_292(u2_col_out_292),
    .col_out_293(u2_col_out_293),
    .col_out_294(u2_col_out_294),
    .col_out_295(u2_col_out_295),
    .col_out_296(u2_col_out_296),
    .col_out_297(u2_col_out_297),
    .col_out_298(u2_col_out_298),
    .col_out_299(u2_col_out_299),
    .col_out_300(u2_col_out_300),
    .col_out_301(u2_col_out_301),
    .col_out_302(u2_col_out_302),
    .col_out_303(u2_col_out_303),
    .col_out_304(u2_col_out_304),
    .col_out_305(u2_col_out_305),
    .col_out_306(u2_col_out_306),
    .col_out_307(u2_col_out_307),
    .col_out_308(u2_col_out_308),
    .col_out_309(u2_col_out_309),
    .col_out_310(u2_col_out_310),
    .col_out_311(u2_col_out_311),
    .col_out_312(u2_col_out_312),
    .col_out_313(u2_col_out_313),
    .col_out_314(u2_col_out_314),
    .col_out_315(u2_col_out_315),
    .col_out_316(u2_col_out_316),
    .col_out_317(u2_col_out_317),
    .col_out_318(u2_col_out_318),
    .col_out_319(u2_col_out_319),
    .col_out_320(u2_col_out_320),
    .col_out_321(u2_col_out_321),
    .col_out_322(u2_col_out_322),
    .col_out_323(u2_col_out_323),
    .col_out_324(u2_col_out_324),
    .col_out_325(u2_col_out_325),
    .col_out_326(u2_col_out_326),
    .col_out_327(u2_col_out_327),
    .col_out_328(u2_col_out_328),
    .col_out_329(u2_col_out_329),
    .col_out_330(u2_col_out_330),
    .col_out_331(u2_col_out_331),
    .col_out_332(u2_col_out_332),
    .col_out_333(u2_col_out_333),
    .col_out_334(u2_col_out_334),
    .col_out_335(u2_col_out_335),
    .col_out_336(u2_col_out_336),
    .col_out_337(u2_col_out_337),
    .col_out_338(u2_col_out_338),
    .col_out_339(u2_col_out_339),
    .col_out_340(u2_col_out_340),
    .col_out_341(u2_col_out_341),
    .col_out_342(u2_col_out_342),
    .col_out_343(u2_col_out_343),
    .col_out_344(u2_col_out_344),
    .col_out_345(u2_col_out_345),
    .col_out_346(u2_col_out_346),
    .col_out_347(u2_col_out_347),
    .col_out_348(u2_col_out_348),
    .col_out_349(u2_col_out_349),
    .col_out_350(u2_col_out_350),
    .col_out_351(u2_col_out_351),
    .col_out_352(u2_col_out_352),
    .col_out_353(u2_col_out_353),
    .col_out_354(u2_col_out_354),
    .col_out_355(u2_col_out_355),
    .col_out_356(u2_col_out_356),
    .col_out_357(u2_col_out_357),
    .col_out_358(u2_col_out_358),
    .col_out_359(u2_col_out_359),
    .col_out_360(u2_col_out_360),
    .col_out_361(u2_col_out_361),
    .col_out_362(u2_col_out_362),
    .col_out_363(u2_col_out_363),
    .col_out_364(u2_col_out_364),
    .col_out_365(u2_col_out_365),
    .col_out_366(u2_col_out_366),
    .col_out_367(u2_col_out_367),
    .col_out_368(u2_col_out_368),
    .col_out_369(u2_col_out_369),
    .col_out_370(u2_col_out_370),
    .col_out_371(u2_col_out_371),
    .col_out_372(u2_col_out_372),
    .col_out_373(u2_col_out_373),
    .col_out_374(u2_col_out_374),
    .col_out_375(u2_col_out_375),
    .col_out_376(u2_col_out_376),
    .col_out_377(u2_col_out_377),
    .col_out_378(u2_col_out_378),
    .col_out_379(u2_col_out_379),
    .col_out_380(u2_col_out_380),
    .col_out_381(u2_col_out_381),
    .col_out_382(u2_col_out_382),
    .col_out_383(u2_col_out_383),
    .col_out_384(u2_col_out_384),
    .col_out_385(u2_col_out_385),
    .col_out_386(u2_col_out_386),
    .col_out_387(u2_col_out_387),
    .col_out_388(u2_col_out_388),
    .col_out_389(u2_col_out_389),
    .col_out_390(u2_col_out_390),
    .col_out_391(u2_col_out_391),
    .col_out_392(u2_col_out_392),
    .col_out_393(u2_col_out_393),
    .col_out_394(u2_col_out_394),
    .col_out_395(u2_col_out_395),
    .col_out_396(u2_col_out_396),
    .col_out_397(u2_col_out_397),
    .col_out_398(u2_col_out_398),
    .col_out_399(u2_col_out_399),
    .col_out_400(u2_col_out_400),
    .col_out_401(u2_col_out_401),
    .col_out_402(u2_col_out_402),
    .col_out_403(u2_col_out_403),
    .col_out_404(u2_col_out_404),
    .col_out_405(u2_col_out_405),
    .col_out_406(u2_col_out_406),
    .col_out_407(u2_col_out_407),
    .col_out_408(u2_col_out_408),
    .col_out_409(u2_col_out_409),
    .col_out_410(u2_col_out_410),
    .col_out_411(u2_col_out_411),
    .col_out_412(u2_col_out_412),
    .col_out_413(u2_col_out_413),
    .col_out_414(u2_col_out_414),
    .col_out_415(u2_col_out_415),
    .col_out_416(u2_col_out_416),
    .col_out_417(u2_col_out_417),
    .col_out_418(u2_col_out_418),
    .col_out_419(u2_col_out_419),
    .col_out_420(u2_col_out_420),
    .col_out_421(u2_col_out_421),
    .col_out_422(u2_col_out_422),
    .col_out_423(u2_col_out_423),
    .col_out_424(u2_col_out_424),
    .col_out_425(u2_col_out_425),
    .col_out_426(u2_col_out_426),
    .col_out_427(u2_col_out_427),
    .col_out_428(u2_col_out_428),
    .col_out_429(u2_col_out_429),
    .col_out_430(u2_col_out_430),
    .col_out_431(u2_col_out_431),
    .col_out_432(u2_col_out_432),
    .col_out_433(u2_col_out_433),
    .col_out_434(u2_col_out_434),
    .col_out_435(u2_col_out_435),
    .col_out_436(u2_col_out_436),
    .col_out_437(u2_col_out_437),
    .col_out_438(u2_col_out_438),
    .col_out_439(u2_col_out_439),
    .col_out_440(u2_col_out_440),
    .col_out_441(u2_col_out_441),
    .col_out_442(u2_col_out_442),
    .col_out_443(u2_col_out_443),
    .col_out_444(u2_col_out_444),
    .col_out_445(u2_col_out_445),
    .col_out_446(u2_col_out_446),
    .col_out_447(u2_col_out_447),
    .col_out_448(u2_col_out_448),
    .col_out_449(u2_col_out_449),
    .col_out_450(u2_col_out_450),
    .col_out_451(u2_col_out_451),
    .col_out_452(u2_col_out_452),
    .col_out_453(u2_col_out_453),
    .col_out_454(u2_col_out_454),
    .col_out_455(u2_col_out_455),
    .col_out_456(u2_col_out_456),
    .col_out_457(u2_col_out_457),
    .col_out_458(u2_col_out_458),
    .col_out_459(u2_col_out_459),
    .col_out_460(u2_col_out_460),
    .col_out_461(u2_col_out_461),
    .col_out_462(u2_col_out_462),
    .col_out_463(u2_col_out_463),
    .col_out_464(u2_col_out_464),
    .col_out_465(u2_col_out_465),
    .col_out_466(u2_col_out_466),
    .col_out_467(u2_col_out_467),
    .col_out_468(u2_col_out_468),
    .col_out_469(u2_col_out_469),
    .col_out_470(u2_col_out_470),
    .col_out_471(u2_col_out_471),
    .col_out_472(u2_col_out_472),
    .col_out_473(u2_col_out_473),
    .col_out_474(u2_col_out_474),
    .col_out_475(u2_col_out_475),
    .col_out_476(u2_col_out_476),
    .col_out_477(u2_col_out_477),
    .col_out_478(u2_col_out_478),
    .col_out_479(u2_col_out_479),
    .col_out_480(u2_col_out_480),
    .col_out_481(u2_col_out_481),
    .col_out_482(u2_col_out_482),
    .col_out_483(u2_col_out_483),
    .col_out_484(u2_col_out_484),
    .col_out_485(u2_col_out_485),
    .col_out_486(u2_col_out_486),
    .col_out_487(u2_col_out_487),
    .col_out_488(u2_col_out_488),
    .col_out_489(u2_col_out_489),
    .col_out_490(u2_col_out_490),
    .col_out_491(u2_col_out_491),
    .col_out_492(u2_col_out_492),
    .col_out_493(u2_col_out_493),
    .col_out_494(u2_col_out_494),
    .col_out_495(u2_col_out_495),
    .col_out_496(u2_col_out_496),
    .col_out_497(u2_col_out_497),
    .col_out_498(u2_col_out_498),
    .col_out_499(u2_col_out_499),
    .col_out_500(u2_col_out_500),
    .col_out_501(u2_col_out_501),
    .col_out_502(u2_col_out_502),
    .col_out_503(u2_col_out_503),
    .col_out_504(u2_col_out_504),
    .col_out_505(u2_col_out_505),
    .col_out_506(u2_col_out_506),
    .col_out_507(u2_col_out_507),
    .col_out_508(u2_col_out_508),
    .col_out_509(u2_col_out_509),
    .col_out_510(u2_col_out_510),
    .col_out_511(u2_col_out_511),
    .col_out_512(u2_col_out_512),
    .col_out_513(u2_col_out_513),
    .col_out_514(u2_col_out_514),
    .col_out_515(u2_col_out_515),
    .col_out_516(u2_col_out_516),
    .col_out_517(u2_col_out_517),
    .col_out_518(u2_col_out_518),
    .col_out_519(u2_col_out_519),
    .col_out_520(u2_col_out_520),
    .col_out_521(u2_col_out_521),
    .col_out_522(u2_col_out_522),
    .col_out_523(u2_col_out_523),
    .col_out_524(u2_col_out_524),
    .col_out_525(u2_col_out_525),
    .col_out_526(u2_col_out_526),
    .col_out_527(u2_col_out_527),
    .col_out_528(u2_col_out_528),
    .col_out_529(u2_col_out_529),
    .col_out_530(u2_col_out_530),
    .col_out_531(u2_col_out_531),
    .col_out_532(u2_col_out_532),
    .col_out_533(u2_col_out_533),
    .col_out_534(u2_col_out_534),
    .col_out_535(u2_col_out_535),
    .col_out_536(u2_col_out_536),
    .col_out_537(u2_col_out_537),
    .col_out_538(u2_col_out_538),
    .col_out_539(u2_col_out_539),
    .col_out_540(u2_col_out_540),
    .col_out_541(u2_col_out_541),
    .col_out_542(u2_col_out_542),
    .col_out_543(u2_col_out_543),
    .col_out_544(u2_col_out_544),
    .col_out_545(u2_col_out_545),
    .col_out_546(u2_col_out_546),
    .col_out_547(u2_col_out_547),
    .col_out_548(u2_col_out_548),
    .col_out_549(u2_col_out_549),
    .col_out_550(u2_col_out_550),
    .col_out_551(u2_col_out_551),
    .col_out_552(u2_col_out_552),
    .col_out_553(u2_col_out_553),
    .col_out_554(u2_col_out_554),
    .col_out_555(u2_col_out_555),
    .col_out_556(u2_col_out_556),
    .col_out_557(u2_col_out_557),
    .col_out_558(u2_col_out_558),
    .col_out_559(u2_col_out_559),
    .col_out_560(u2_col_out_560),
    .col_out_561(u2_col_out_561),
    .col_out_562(u2_col_out_562),
    .col_out_563(u2_col_out_563),
    .col_out_564(u2_col_out_564),
    .col_out_565(u2_col_out_565),
    .col_out_566(u2_col_out_566),
    .col_out_567(u2_col_out_567),
    .col_out_568(u2_col_out_568),
    .col_out_569(u2_col_out_569),
    .col_out_570(u2_col_out_570),
    .col_out_571(u2_col_out_571),
    .col_out_572(u2_col_out_572),
    .col_out_573(u2_col_out_573),
    .col_out_574(u2_col_out_574),
    .col_out_575(u2_col_out_575),
    .col_out_576(u2_col_out_576),
    .col_out_577(u2_col_out_577),
    .col_out_578(u2_col_out_578),
    .col_out_579(u2_col_out_579),
    .col_out_580(u2_col_out_580),
    .col_out_581(u2_col_out_581),
    .col_out_582(u2_col_out_582),
    .col_out_583(u2_col_out_583),
    .col_out_584(u2_col_out_584),
    .col_out_585(u2_col_out_585),
    .col_out_586(u2_col_out_586),
    .col_out_587(u2_col_out_587),
    .col_out_588(u2_col_out_588),
    .col_out_589(u2_col_out_589),
    .col_out_590(u2_col_out_590),
    .col_out_591(u2_col_out_591),
    .col_out_592(u2_col_out_592),
    .col_out_593(u2_col_out_593),
    .col_out_594(u2_col_out_594),
    .col_out_595(u2_col_out_595),
    .col_out_596(u2_col_out_596),
    .col_out_597(u2_col_out_597),
    .col_out_598(u2_col_out_598),
    .col_out_599(u2_col_out_599),
    .col_out_600(u2_col_out_600),
    .col_out_601(u2_col_out_601),
    .col_out_602(u2_col_out_602),
    .col_out_603(u2_col_out_603),
    .col_out_604(u2_col_out_604),
    .col_out_605(u2_col_out_605),
    .col_out_606(u2_col_out_606),
    .col_out_607(u2_col_out_607),
    .col_out_608(u2_col_out_608),
    .col_out_609(u2_col_out_609),
    .col_out_610(u2_col_out_610),
    .col_out_611(u2_col_out_611),
    .col_out_612(u2_col_out_612),
    .col_out_613(u2_col_out_613),
    .col_out_614(u2_col_out_614),
    .col_out_615(u2_col_out_615),
    .col_out_616(u2_col_out_616),
    .col_out_617(u2_col_out_617),
    .col_out_618(u2_col_out_618),
    .col_out_619(u2_col_out_619),
    .col_out_620(u2_col_out_620),
    .col_out_621(u2_col_out_621),
    .col_out_622(u2_col_out_622),
    .col_out_623(u2_col_out_623),
    .col_out_624(u2_col_out_624),
    .col_out_625(u2_col_out_625),
    .col_out_626(u2_col_out_626),
    .col_out_627(u2_col_out_627),
    .col_out_628(u2_col_out_628),
    .col_out_629(u2_col_out_629),
    .col_out_630(u2_col_out_630),
    .col_out_631(u2_col_out_631),
    .col_out_632(u2_col_out_632),
    .col_out_633(u2_col_out_633),
    .col_out_634(u2_col_out_634),
    .col_out_635(u2_col_out_635),
    .col_out_636(u2_col_out_636),
    .col_out_637(u2_col_out_637),
    .col_out_638(u2_col_out_638),
    .col_out_639(u2_col_out_639),
    .col_out_640(u2_col_out_640),
    .col_out_641(u2_col_out_641),
    .col_out_642(u2_col_out_642),
    .col_out_643(u2_col_out_643),
    .col_out_644(u2_col_out_644),
    .col_out_645(u2_col_out_645),
    .col_out_646(u2_col_out_646),
    .col_out_647(u2_col_out_647),
    .col_out_648(u2_col_out_648),
    .col_out_649(u2_col_out_649),
    .col_out_650(u2_col_out_650),
    .col_out_651(u2_col_out_651),
    .col_out_652(u2_col_out_652),
    .col_out_653(u2_col_out_653),
    .col_out_654(u2_col_out_654),
    .col_out_655(u2_col_out_655),
    .col_out_656(u2_col_out_656),
    .col_out_657(u2_col_out_657),
    .col_out_658(u2_col_out_658),
    .col_out_659(u2_col_out_659),
    .col_out_660(u2_col_out_660),
    .col_out_661(u2_col_out_661),
    .col_out_662(u2_col_out_662),
    .col_out_663(u2_col_out_663),
    .col_out_664(u2_col_out_664),
    .col_out_665(u2_col_out_665),
    .col_out_666(u2_col_out_666),
    .col_out_667(u2_col_out_667),
    .col_out_668(u2_col_out_668),
    .col_out_669(u2_col_out_669),
    .col_out_670(u2_col_out_670),
    .col_out_671(u2_col_out_671),
    .col_out_672(u2_col_out_672),
    .col_out_673(u2_col_out_673),
    .col_out_674(u2_col_out_674),
    .col_out_675(u2_col_out_675),
    .col_out_676(u2_col_out_676),
    .col_out_677(u2_col_out_677),
    .col_out_678(u2_col_out_678),
    .col_out_679(u2_col_out_679),
    .col_out_680(u2_col_out_680),
    .col_out_681(u2_col_out_681),
    .col_out_682(u2_col_out_682),
    .col_out_683(u2_col_out_683),
    .col_out_684(u2_col_out_684),
    .col_out_685(u2_col_out_685),
    .col_out_686(u2_col_out_686),
    .col_out_687(u2_col_out_687),
    .col_out_688(u2_col_out_688),
    .col_out_689(u2_col_out_689),
    .col_out_690(u2_col_out_690),
    .col_out_691(u2_col_out_691),
    .col_out_692(u2_col_out_692),
    .col_out_693(u2_col_out_693),
    .col_out_694(u2_col_out_694),
    .col_out_695(u2_col_out_695),
    .col_out_696(u2_col_out_696),
    .col_out_697(u2_col_out_697),
    .col_out_698(u2_col_out_698),
    .col_out_699(u2_col_out_699),
    .col_out_700(u2_col_out_700),
    .col_out_701(u2_col_out_701),
    .col_out_702(u2_col_out_702),
    .col_out_703(u2_col_out_703),
    .col_out_704(u2_col_out_704),
    .col_out_705(u2_col_out_705),
    .col_out_706(u2_col_out_706),
    .col_out_707(u2_col_out_707),
    .col_out_708(u2_col_out_708),
    .col_out_709(u2_col_out_709),
    .col_out_710(u2_col_out_710),
    .col_out_711(u2_col_out_711),
    .col_out_712(u2_col_out_712),
    .col_out_713(u2_col_out_713),
    .col_out_714(u2_col_out_714),
    .col_out_715(u2_col_out_715),
    .col_out_716(u2_col_out_716),
    .col_out_717(u2_col_out_717),
    .col_out_718(u2_col_out_718),
    .col_out_719(u2_col_out_719),
    .col_out_720(u2_col_out_720),
    .col_out_721(u2_col_out_721),
    .col_out_722(u2_col_out_722),
    .col_out_723(u2_col_out_723),
    .col_out_724(u2_col_out_724),
    .col_out_725(u2_col_out_725),
    .col_out_726(u2_col_out_726),
    .col_out_727(u2_col_out_727),
    .col_out_728(u2_col_out_728),
    .col_out_729(u2_col_out_729),
    .col_out_730(u2_col_out_730),
    .col_out_731(u2_col_out_731),
    .col_out_732(u2_col_out_732),
    .col_out_733(u2_col_out_733),
    .col_out_734(u2_col_out_734),
    .col_out_735(u2_col_out_735),
    .col_out_736(u2_col_out_736),
    .col_out_737(u2_col_out_737),
    .col_out_738(u2_col_out_738),
    .col_out_739(u2_col_out_739),
    .col_out_740(u2_col_out_740),
    .col_out_741(u2_col_out_741),
    .col_out_742(u2_col_out_742),
    .col_out_743(u2_col_out_743),
    .col_out_744(u2_col_out_744),
    .col_out_745(u2_col_out_745),
    .col_out_746(u2_col_out_746),
    .col_out_747(u2_col_out_747),
    .col_out_748(u2_col_out_748),
    .col_out_749(u2_col_out_749),
    .col_out_750(u2_col_out_750),
    .col_out_751(u2_col_out_751),
    .col_out_752(u2_col_out_752),
    .col_out_753(u2_col_out_753),
    .col_out_754(u2_col_out_754),
    .col_out_755(u2_col_out_755),
    .col_out_756(u2_col_out_756),
    .col_out_757(u2_col_out_757),
    .col_out_758(u2_col_out_758),
    .col_out_759(u2_col_out_759),
    .col_out_760(u2_col_out_760),
    .col_out_761(u2_col_out_761),
    .col_out_762(u2_col_out_762),
    .col_out_763(u2_col_out_763),
    .col_out_764(u2_col_out_764),
    .col_out_765(u2_col_out_765),
    .col_out_766(u2_col_out_766),
    .col_out_767(u2_col_out_767),
    .col_out_768(u2_col_out_768),
    .col_out_769(u2_col_out_769),
    .col_out_770(u2_col_out_770),
    .col_out_771(u2_col_out_771),
    .col_out_772(u2_col_out_772),
    .col_out_773(u2_col_out_773),
    .col_out_774(u2_col_out_774),
    .col_out_775(u2_col_out_775),
    .col_out_776(u2_col_out_776),
    .col_out_777(u2_col_out_777),
    .col_out_778(u2_col_out_778),
    .col_out_779(u2_col_out_779),
    .col_out_780(u2_col_out_780),
    .col_out_781(u2_col_out_781),
    .col_out_782(u2_col_out_782),
    .col_out_783(u2_col_out_783),
    .col_out_784(u2_col_out_784),
    .col_out_785(u2_col_out_785),
    .col_out_786(u2_col_out_786),
    .col_out_787(u2_col_out_787),
    .col_out_788(u2_col_out_788),
    .col_out_789(u2_col_out_789),
    .col_out_790(u2_col_out_790),
    .col_out_791(u2_col_out_791),
    .col_out_792(u2_col_out_792),
    .col_out_793(u2_col_out_793),
    .col_out_794(u2_col_out_794),
    .col_out_795(u2_col_out_795),
    .col_out_796(u2_col_out_796),
    .col_out_797(u2_col_out_797),
    .col_out_798(u2_col_out_798),
    .col_out_799(u2_col_out_799),
    .col_out_800(u2_col_out_800),
    .col_out_801(u2_col_out_801),
    .col_out_802(u2_col_out_802),
    .col_out_803(u2_col_out_803),
    .col_out_804(u2_col_out_804),
    .col_out_805(u2_col_out_805),
    .col_out_806(u2_col_out_806),
    .col_out_807(u2_col_out_807),
    .col_out_808(u2_col_out_808),
    .col_out_809(u2_col_out_809),
    .col_out_810(u2_col_out_810),
    .col_out_811(u2_col_out_811),
    .col_out_812(u2_col_out_812),
    .col_out_813(u2_col_out_813),
    .col_out_814(u2_col_out_814),
    .col_out_815(u2_col_out_815),
    .col_out_816(u2_col_out_816),
    .col_out_817(u2_col_out_817),
    .col_out_818(u2_col_out_818),
    .col_out_819(u2_col_out_819),
    .col_out_820(u2_col_out_820),
    .col_out_821(u2_col_out_821),
    .col_out_822(u2_col_out_822),
    .col_out_823(u2_col_out_823),
    .col_out_824(u2_col_out_824),
    .col_out_825(u2_col_out_825),
    .col_out_826(u2_col_out_826),
    .col_out_827(u2_col_out_827),
    .col_out_828(u2_col_out_828),
    .col_out_829(u2_col_out_829),
    .col_out_830(u2_col_out_830),
    .col_out_831(u2_col_out_831),
    .col_out_832(u2_col_out_832),
    .col_out_833(u2_col_out_833),
    .col_out_834(u2_col_out_834),
    .col_out_835(u2_col_out_835),
    .col_out_836(u2_col_out_836),
    .col_out_837(u2_col_out_837),
    .col_out_838(u2_col_out_838),
    .col_out_839(u2_col_out_839),
    .col_out_840(u2_col_out_840),
    .col_out_841(u2_col_out_841),
    .col_out_842(u2_col_out_842),
    .col_out_843(u2_col_out_843),
    .col_out_844(u2_col_out_844),
    .col_out_845(u2_col_out_845),
    .col_out_846(u2_col_out_846),
    .col_out_847(u2_col_out_847),
    .col_out_848(u2_col_out_848),
    .col_out_849(u2_col_out_849),
    .col_out_850(u2_col_out_850),
    .col_out_851(u2_col_out_851),
    .col_out_852(u2_col_out_852),
    .col_out_853(u2_col_out_853),
    .col_out_854(u2_col_out_854),
    .col_out_855(u2_col_out_855),
    .col_out_856(u2_col_out_856),
    .col_out_857(u2_col_out_857),
    .col_out_858(u2_col_out_858),
    .col_out_859(u2_col_out_859),
    .col_out_860(u2_col_out_860),
    .col_out_861(u2_col_out_861),
    .col_out_862(u2_col_out_862),
    .col_out_863(u2_col_out_863),
    .col_out_864(u2_col_out_864),
    .col_out_865(u2_col_out_865),
    .col_out_866(u2_col_out_866),
    .col_out_867(u2_col_out_867),
    .col_out_868(u2_col_out_868),
    .col_out_869(u2_col_out_869),
    .col_out_870(u2_col_out_870),
    .col_out_871(u2_col_out_871),
    .col_out_872(u2_col_out_872),
    .col_out_873(u2_col_out_873),
    .col_out_874(u2_col_out_874),
    .col_out_875(u2_col_out_875),
    .col_out_876(u2_col_out_876),
    .col_out_877(u2_col_out_877),
    .col_out_878(u2_col_out_878),
    .col_out_879(u2_col_out_879),
    .col_out_880(u2_col_out_880),
    .col_out_881(u2_col_out_881),
    .col_out_882(u2_col_out_882),
    .col_out_883(u2_col_out_883),
    .col_out_884(u2_col_out_884),
    .col_out_885(u2_col_out_885),
    .col_out_886(u2_col_out_886),
    .col_out_887(u2_col_out_887),
    .col_out_888(u2_col_out_888),
    .col_out_889(u2_col_out_889),
    .col_out_890(u2_col_out_890),
    .col_out_891(u2_col_out_891),
    .col_out_892(u2_col_out_892),
    .col_out_893(u2_col_out_893),
    .col_out_894(u2_col_out_894),
    .col_out_895(u2_col_out_895),
    .col_out_896(u2_col_out_896),
    .col_out_897(u2_col_out_897),
    .col_out_898(u2_col_out_898),
    .col_out_899(u2_col_out_899),
    .col_out_900(u2_col_out_900),
    .col_out_901(u2_col_out_901),
    .col_out_902(u2_col_out_902),
    .col_out_903(u2_col_out_903),
    .col_out_904(u2_col_out_904),
    .col_out_905(u2_col_out_905),
    .col_out_906(u2_col_out_906),
    .col_out_907(u2_col_out_907),
    .col_out_908(u2_col_out_908),
    .col_out_909(u2_col_out_909),
    .col_out_910(u2_col_out_910),
    .col_out_911(u2_col_out_911),
    .col_out_912(u2_col_out_912),
    .col_out_913(u2_col_out_913),
    .col_out_914(u2_col_out_914),
    .col_out_915(u2_col_out_915),
    .col_out_916(u2_col_out_916),
    .col_out_917(u2_col_out_917),
    .col_out_918(u2_col_out_918),
    .col_out_919(u2_col_out_919),
    .col_out_920(u2_col_out_920),
    .col_out_921(u2_col_out_921),
    .col_out_922(u2_col_out_922),
    .col_out_923(u2_col_out_923),
    .col_out_924(u2_col_out_924),
    .col_out_925(u2_col_out_925),
    .col_out_926(u2_col_out_926),
    .col_out_927(u2_col_out_927),
    .col_out_928(u2_col_out_928),
    .col_out_929(u2_col_out_929),
    .col_out_930(u2_col_out_930),
    .col_out_931(u2_col_out_931),
    .col_out_932(u2_col_out_932),
    .col_out_933(u2_col_out_933),
    .col_out_934(u2_col_out_934),
    .col_out_935(u2_col_out_935),
    .col_out_936(u2_col_out_936),
    .col_out_937(u2_col_out_937),
    .col_out_938(u2_col_out_938),
    .col_out_939(u2_col_out_939),
    .col_out_940(u2_col_out_940),
    .col_out_941(u2_col_out_941),
    .col_out_942(u2_col_out_942),
    .col_out_943(u2_col_out_943),
    .col_out_944(u2_col_out_944),
    .col_out_945(u2_col_out_945),
    .col_out_946(u2_col_out_946),
    .col_out_947(u2_col_out_947),
    .col_out_948(u2_col_out_948),
    .col_out_949(u2_col_out_949),
    .col_out_950(u2_col_out_950),
    .col_out_951(u2_col_out_951),
    .col_out_952(u2_col_out_952),
    .col_out_953(u2_col_out_953),
    .col_out_954(u2_col_out_954),
    .col_out_955(u2_col_out_955),
    .col_out_956(u2_col_out_956),
    .col_out_957(u2_col_out_957),
    .col_out_958(u2_col_out_958),
    .col_out_959(u2_col_out_959),
    .col_out_960(u2_col_out_960),
    .col_out_961(u2_col_out_961),
    .col_out_962(u2_col_out_962),
    .col_out_963(u2_col_out_963),
    .col_out_964(u2_col_out_964),
    .col_out_965(u2_col_out_965),
    .col_out_966(u2_col_out_966),
    .col_out_967(u2_col_out_967),
    .col_out_968(u2_col_out_968),
    .col_out_969(u2_col_out_969),
    .col_out_970(u2_col_out_970),
    .col_out_971(u2_col_out_971),
    .col_out_972(u2_col_out_972),
    .col_out_973(u2_col_out_973),
    .col_out_974(u2_col_out_974),
    .col_out_975(u2_col_out_975),
    .col_out_976(u2_col_out_976),
    .col_out_977(u2_col_out_977),
    .col_out_978(u2_col_out_978),
    .col_out_979(u2_col_out_979),
    .col_out_980(u2_col_out_980),
    .col_out_981(u2_col_out_981),
    .col_out_982(u2_col_out_982),
    .col_out_983(u2_col_out_983),
    .col_out_984(u2_col_out_984),
    .col_out_985(u2_col_out_985),
    .col_out_986(u2_col_out_986),
    .col_out_987(u2_col_out_987),
    .col_out_988(u2_col_out_988),
    .col_out_989(u2_col_out_989),
    .col_out_990(u2_col_out_990),
    .col_out_991(u2_col_out_991),
    .col_out_992(u2_col_out_992),
    .col_out_993(u2_col_out_993),
    .col_out_994(u2_col_out_994),
    .col_out_995(u2_col_out_995),
    .col_out_996(u2_col_out_996),
    .col_out_997(u2_col_out_997),
    .col_out_998(u2_col_out_998),
    .col_out_999(u2_col_out_999),
    .col_out_1000(u2_col_out_1000),
    .col_out_1001(u2_col_out_1001),
    .col_out_1002(u2_col_out_1002),
    .col_out_1003(u2_col_out_1003),
    .col_out_1004(u2_col_out_1004),
    .col_out_1005(u2_col_out_1005),
    .col_out_1006(u2_col_out_1006),
    .col_out_1007(u2_col_out_1007),
    .col_out_1008(u2_col_out_1008),
    .col_out_1009(u2_col_out_1009),
    .col_out_1010(u2_col_out_1010),
    .col_out_1011(u2_col_out_1011),
    .col_out_1012(u2_col_out_1012),
    .col_out_1013(u2_col_out_1013),
    .col_out_1014(u2_col_out_1014),
    .col_out_1015(u2_col_out_1015),
    .col_out_1016(u2_col_out_1016),
    .col_out_1017(u2_col_out_1017),
    .col_out_1018(u2_col_out_1018),
    .col_out_1019(u2_col_out_1019),
    .col_out_1020(u2_col_out_1020),
    .col_out_1021(u2_col_out_1021),
    .col_out_1022(u2_col_out_1022),
    .col_out_1023(u2_col_out_1023),
    .col_out_1024(u2_col_out_1024),
    .col_out_1025(u2_col_out_1025),
    .col_out_1026(u2_col_out_1026),
    .col_out_1027(u2_col_out_1027),
    .col_out_1028(u2_col_out_1028),
    .col_out_1029(u2_col_out_1029),
    .col_out_1030(u2_col_out_1030),
    .col_out_1031(u2_col_out_1031),
    .col_out_1032(u2_col_out_1032)
);


//*****************************************************
//**************输出赋值******************************
//*****************************************************
assign col_out_0 = u2_col_out_0;
assign col_out_1 = u2_col_out_1;
assign col_out_2 = u2_col_out_2;
assign col_out_3 = u2_col_out_3;
assign col_out_4 = u2_col_out_4;
assign col_out_5 = u2_col_out_5;
assign col_out_6 = u2_col_out_6;
assign col_out_7 = u2_col_out_7;
assign col_out_8 = u2_col_out_8;
assign col_out_9 = u2_col_out_9;
assign col_out_10 = u2_col_out_10;
assign col_out_11 = u2_col_out_11;
assign col_out_12 = u2_col_out_12;
assign col_out_13 = u2_col_out_13;
assign col_out_14 = u2_col_out_14;
assign col_out_15 = u2_col_out_15;
assign col_out_16 = u2_col_out_16;
assign col_out_17 = u2_col_out_17;
assign col_out_18 = u2_col_out_18;
assign col_out_19 = u2_col_out_19;
assign col_out_20 = u2_col_out_20;
assign col_out_21 = u2_col_out_21;
assign col_out_22 = u2_col_out_22;
assign col_out_23 = u2_col_out_23;
assign col_out_24 = u2_col_out_24;
assign col_out_25 = u2_col_out_25;
assign col_out_26 = u2_col_out_26;
assign col_out_27 = u2_col_out_27;
assign col_out_28 = u2_col_out_28;
assign col_out_29 = u2_col_out_29;
assign col_out_30 = u2_col_out_30;
assign col_out_31 = u2_col_out_31;
assign col_out_32 = u2_col_out_32;
assign col_out_33 = u2_col_out_33;
assign col_out_34 = u2_col_out_34;
assign col_out_35 = u2_col_out_35;
assign col_out_36 = u2_col_out_36;
assign col_out_37 = u2_col_out_37;
assign col_out_38 = u2_col_out_38;
assign col_out_39 = u2_col_out_39;
assign col_out_40 = u2_col_out_40;
assign col_out_41 = u2_col_out_41;
assign col_out_42 = u2_col_out_42;
assign col_out_43 = u2_col_out_43;
assign col_out_44 = u2_col_out_44;
assign col_out_45 = u2_col_out_45;
assign col_out_46 = u2_col_out_46;
assign col_out_47 = u2_col_out_47;
assign col_out_48 = u2_col_out_48;
assign col_out_49 = u2_col_out_49;
assign col_out_50 = u2_col_out_50;
assign col_out_51 = u2_col_out_51;
assign col_out_52 = u2_col_out_52;
assign col_out_53 = u2_col_out_53;
assign col_out_54 = u2_col_out_54;
assign col_out_55 = u2_col_out_55;
assign col_out_56 = u2_col_out_56;
assign col_out_57 = u2_col_out_57;
assign col_out_58 = u2_col_out_58;
assign col_out_59 = u2_col_out_59;
assign col_out_60 = u2_col_out_60;
assign col_out_61 = u2_col_out_61;
assign col_out_62 = u2_col_out_62;
assign col_out_63 = u2_col_out_63;
assign col_out_64 = u2_col_out_64;
assign col_out_65 = u2_col_out_65;
assign col_out_66 = u2_col_out_66;
assign col_out_67 = u2_col_out_67;
assign col_out_68 = u2_col_out_68;
assign col_out_69 = u2_col_out_69;
assign col_out_70 = u2_col_out_70;
assign col_out_71 = u2_col_out_71;
assign col_out_72 = u2_col_out_72;
assign col_out_73 = u2_col_out_73;
assign col_out_74 = u2_col_out_74;
assign col_out_75 = u2_col_out_75;
assign col_out_76 = u2_col_out_76;
assign col_out_77 = u2_col_out_77;
assign col_out_78 = u2_col_out_78;
assign col_out_79 = u2_col_out_79;
assign col_out_80 = u2_col_out_80;
assign col_out_81 = u2_col_out_81;
assign col_out_82 = u2_col_out_82;
assign col_out_83 = u2_col_out_83;
assign col_out_84 = u2_col_out_84;
assign col_out_85 = u2_col_out_85;
assign col_out_86 = u2_col_out_86;
assign col_out_87 = u2_col_out_87;
assign col_out_88 = u2_col_out_88;
assign col_out_89 = u2_col_out_89;
assign col_out_90 = u2_col_out_90;
assign col_out_91 = u2_col_out_91;
assign col_out_92 = u2_col_out_92;
assign col_out_93 = u2_col_out_93;
assign col_out_94 = u2_col_out_94;
assign col_out_95 = u2_col_out_95;
assign col_out_96 = u2_col_out_96;
assign col_out_97 = u2_col_out_97;
assign col_out_98 = u2_col_out_98;
assign col_out_99 = u2_col_out_99;
assign col_out_100 = u2_col_out_100;
assign col_out_101 = u2_col_out_101;
assign col_out_102 = u2_col_out_102;
assign col_out_103 = u2_col_out_103;
assign col_out_104 = u2_col_out_104;
assign col_out_105 = u2_col_out_105;
assign col_out_106 = u2_col_out_106;
assign col_out_107 = u2_col_out_107;
assign col_out_108 = u2_col_out_108;
assign col_out_109 = u2_col_out_109;
assign col_out_110 = u2_col_out_110;
assign col_out_111 = u2_col_out_111;
assign col_out_112 = u2_col_out_112;
assign col_out_113 = u2_col_out_113;
assign col_out_114 = u2_col_out_114;
assign col_out_115 = u2_col_out_115;
assign col_out_116 = u2_col_out_116;
assign col_out_117 = u2_col_out_117;
assign col_out_118 = u2_col_out_118;
assign col_out_119 = u2_col_out_119;
assign col_out_120 = u2_col_out_120;
assign col_out_121 = u2_col_out_121;
assign col_out_122 = u2_col_out_122;
assign col_out_123 = u2_col_out_123;
assign col_out_124 = u2_col_out_124;
assign col_out_125 = u2_col_out_125;
assign col_out_126 = u2_col_out_126;
assign col_out_127 = u2_col_out_127;
assign col_out_128 = u2_col_out_128;
assign col_out_129 = u2_col_out_129;
assign col_out_130 = u2_col_out_130;
assign col_out_131 = u2_col_out_131;
assign col_out_132 = u2_col_out_132;
assign col_out_133 = u2_col_out_133;
assign col_out_134 = u2_col_out_134;
assign col_out_135 = u2_col_out_135;
assign col_out_136 = u2_col_out_136;
assign col_out_137 = u2_col_out_137;
assign col_out_138 = u2_col_out_138;
assign col_out_139 = u2_col_out_139;
assign col_out_140 = u2_col_out_140;
assign col_out_141 = u2_col_out_141;
assign col_out_142 = u2_col_out_142;
assign col_out_143 = u2_col_out_143;
assign col_out_144 = u2_col_out_144;
assign col_out_145 = u2_col_out_145;
assign col_out_146 = u2_col_out_146;
assign col_out_147 = u2_col_out_147;
assign col_out_148 = u2_col_out_148;
assign col_out_149 = u2_col_out_149;
assign col_out_150 = u2_col_out_150;
assign col_out_151 = u2_col_out_151;
assign col_out_152 = u2_col_out_152;
assign col_out_153 = u2_col_out_153;
assign col_out_154 = u2_col_out_154;
assign col_out_155 = u2_col_out_155;
assign col_out_156 = u2_col_out_156;
assign col_out_157 = u2_col_out_157;
assign col_out_158 = u2_col_out_158;
assign col_out_159 = u2_col_out_159;
assign col_out_160 = u2_col_out_160;
assign col_out_161 = u2_col_out_161;
assign col_out_162 = u2_col_out_162;
assign col_out_163 = u2_col_out_163;
assign col_out_164 = u2_col_out_164;
assign col_out_165 = u2_col_out_165;
assign col_out_166 = u2_col_out_166;
assign col_out_167 = u2_col_out_167;
assign col_out_168 = u2_col_out_168;
assign col_out_169 = u2_col_out_169;
assign col_out_170 = u2_col_out_170;
assign col_out_171 = u2_col_out_171;
assign col_out_172 = u2_col_out_172;
assign col_out_173 = u2_col_out_173;
assign col_out_174 = u2_col_out_174;
assign col_out_175 = u2_col_out_175;
assign col_out_176 = u2_col_out_176;
assign col_out_177 = u2_col_out_177;
assign col_out_178 = u2_col_out_178;
assign col_out_179 = u2_col_out_179;
assign col_out_180 = u2_col_out_180;
assign col_out_181 = u2_col_out_181;
assign col_out_182 = u2_col_out_182;
assign col_out_183 = u2_col_out_183;
assign col_out_184 = u2_col_out_184;
assign col_out_185 = u2_col_out_185;
assign col_out_186 = u2_col_out_186;
assign col_out_187 = u2_col_out_187;
assign col_out_188 = u2_col_out_188;
assign col_out_189 = u2_col_out_189;
assign col_out_190 = u2_col_out_190;
assign col_out_191 = u2_col_out_191;
assign col_out_192 = u2_col_out_192;
assign col_out_193 = u2_col_out_193;
assign col_out_194 = u2_col_out_194;
assign col_out_195 = u2_col_out_195;
assign col_out_196 = u2_col_out_196;
assign col_out_197 = u2_col_out_197;
assign col_out_198 = u2_col_out_198;
assign col_out_199 = u2_col_out_199;
assign col_out_200 = u2_col_out_200;
assign col_out_201 = u2_col_out_201;
assign col_out_202 = u2_col_out_202;
assign col_out_203 = u2_col_out_203;
assign col_out_204 = u2_col_out_204;
assign col_out_205 = u2_col_out_205;
assign col_out_206 = u2_col_out_206;
assign col_out_207 = u2_col_out_207;
assign col_out_208 = u2_col_out_208;
assign col_out_209 = u2_col_out_209;
assign col_out_210 = u2_col_out_210;
assign col_out_211 = u2_col_out_211;
assign col_out_212 = u2_col_out_212;
assign col_out_213 = u2_col_out_213;
assign col_out_214 = u2_col_out_214;
assign col_out_215 = u2_col_out_215;
assign col_out_216 = u2_col_out_216;
assign col_out_217 = u2_col_out_217;
assign col_out_218 = u2_col_out_218;
assign col_out_219 = u2_col_out_219;
assign col_out_220 = u2_col_out_220;
assign col_out_221 = u2_col_out_221;
assign col_out_222 = u2_col_out_222;
assign col_out_223 = u2_col_out_223;
assign col_out_224 = u2_col_out_224;
assign col_out_225 = u2_col_out_225;
assign col_out_226 = u2_col_out_226;
assign col_out_227 = u2_col_out_227;
assign col_out_228 = u2_col_out_228;
assign col_out_229 = u2_col_out_229;
assign col_out_230 = u2_col_out_230;
assign col_out_231 = u2_col_out_231;
assign col_out_232 = u2_col_out_232;
assign col_out_233 = u2_col_out_233;
assign col_out_234 = u2_col_out_234;
assign col_out_235 = u2_col_out_235;
assign col_out_236 = u2_col_out_236;
assign col_out_237 = u2_col_out_237;
assign col_out_238 = u2_col_out_238;
assign col_out_239 = u2_col_out_239;
assign col_out_240 = u2_col_out_240;
assign col_out_241 = u2_col_out_241;
assign col_out_242 = u2_col_out_242;
assign col_out_243 = u2_col_out_243;
assign col_out_244 = u2_col_out_244;
assign col_out_245 = u2_col_out_245;
assign col_out_246 = u2_col_out_246;
assign col_out_247 = u2_col_out_247;
assign col_out_248 = u2_col_out_248;
assign col_out_249 = u2_col_out_249;
assign col_out_250 = u2_col_out_250;
assign col_out_251 = u2_col_out_251;
assign col_out_252 = u2_col_out_252;
assign col_out_253 = u2_col_out_253;
assign col_out_254 = u2_col_out_254;
assign col_out_255 = u2_col_out_255;
assign col_out_256 = u2_col_out_256;
assign col_out_257 = u2_col_out_257;
assign col_out_258 = u2_col_out_258;
assign col_out_259 = u2_col_out_259;
assign col_out_260 = u2_col_out_260;
assign col_out_261 = u2_col_out_261;
assign col_out_262 = u2_col_out_262;
assign col_out_263 = u2_col_out_263;
assign col_out_264 = u2_col_out_264;
assign col_out_265 = u2_col_out_265;
assign col_out_266 = u2_col_out_266;
assign col_out_267 = u2_col_out_267;
assign col_out_268 = u2_col_out_268;
assign col_out_269 = u2_col_out_269;
assign col_out_270 = u2_col_out_270;
assign col_out_271 = u2_col_out_271;
assign col_out_272 = u2_col_out_272;
assign col_out_273 = u2_col_out_273;
assign col_out_274 = u2_col_out_274;
assign col_out_275 = u2_col_out_275;
assign col_out_276 = u2_col_out_276;
assign col_out_277 = u2_col_out_277;
assign col_out_278 = u2_col_out_278;
assign col_out_279 = u2_col_out_279;
assign col_out_280 = u2_col_out_280;
assign col_out_281 = u2_col_out_281;
assign col_out_282 = u2_col_out_282;
assign col_out_283 = u2_col_out_283;
assign col_out_284 = u2_col_out_284;
assign col_out_285 = u2_col_out_285;
assign col_out_286 = u2_col_out_286;
assign col_out_287 = u2_col_out_287;
assign col_out_288 = u2_col_out_288;
assign col_out_289 = u2_col_out_289;
assign col_out_290 = u2_col_out_290;
assign col_out_291 = u2_col_out_291;
assign col_out_292 = u2_col_out_292;
assign col_out_293 = u2_col_out_293;
assign col_out_294 = u2_col_out_294;
assign col_out_295 = u2_col_out_295;
assign col_out_296 = u2_col_out_296;
assign col_out_297 = u2_col_out_297;
assign col_out_298 = u2_col_out_298;
assign col_out_299 = u2_col_out_299;
assign col_out_300 = u2_col_out_300;
assign col_out_301 = u2_col_out_301;
assign col_out_302 = u2_col_out_302;
assign col_out_303 = u2_col_out_303;
assign col_out_304 = u2_col_out_304;
assign col_out_305 = u2_col_out_305;
assign col_out_306 = u2_col_out_306;
assign col_out_307 = u2_col_out_307;
assign col_out_308 = u2_col_out_308;
assign col_out_309 = u2_col_out_309;
assign col_out_310 = u2_col_out_310;
assign col_out_311 = u2_col_out_311;
assign col_out_312 = u2_col_out_312;
assign col_out_313 = u2_col_out_313;
assign col_out_314 = u2_col_out_314;
assign col_out_315 = u2_col_out_315;
assign col_out_316 = u2_col_out_316;
assign col_out_317 = u2_col_out_317;
assign col_out_318 = u2_col_out_318;
assign col_out_319 = u2_col_out_319;
assign col_out_320 = u2_col_out_320;
assign col_out_321 = u2_col_out_321;
assign col_out_322 = u2_col_out_322;
assign col_out_323 = u2_col_out_323;
assign col_out_324 = u2_col_out_324;
assign col_out_325 = u2_col_out_325;
assign col_out_326 = u2_col_out_326;
assign col_out_327 = u2_col_out_327;
assign col_out_328 = u2_col_out_328;
assign col_out_329 = u2_col_out_329;
assign col_out_330 = u2_col_out_330;
assign col_out_331 = u2_col_out_331;
assign col_out_332 = u2_col_out_332;
assign col_out_333 = u2_col_out_333;
assign col_out_334 = u2_col_out_334;
assign col_out_335 = u2_col_out_335;
assign col_out_336 = u2_col_out_336;
assign col_out_337 = u2_col_out_337;
assign col_out_338 = u2_col_out_338;
assign col_out_339 = u2_col_out_339;
assign col_out_340 = u2_col_out_340;
assign col_out_341 = u2_col_out_341;
assign col_out_342 = u2_col_out_342;
assign col_out_343 = u2_col_out_343;
assign col_out_344 = u2_col_out_344;
assign col_out_345 = u2_col_out_345;
assign col_out_346 = u2_col_out_346;
assign col_out_347 = u2_col_out_347;
assign col_out_348 = u2_col_out_348;
assign col_out_349 = u2_col_out_349;
assign col_out_350 = u2_col_out_350;
assign col_out_351 = u2_col_out_351;
assign col_out_352 = u2_col_out_352;
assign col_out_353 = u2_col_out_353;
assign col_out_354 = u2_col_out_354;
assign col_out_355 = u2_col_out_355;
assign col_out_356 = u2_col_out_356;
assign col_out_357 = u2_col_out_357;
assign col_out_358 = u2_col_out_358;
assign col_out_359 = u2_col_out_359;
assign col_out_360 = u2_col_out_360;
assign col_out_361 = u2_col_out_361;
assign col_out_362 = u2_col_out_362;
assign col_out_363 = u2_col_out_363;
assign col_out_364 = u2_col_out_364;
assign col_out_365 = u2_col_out_365;
assign col_out_366 = u2_col_out_366;
assign col_out_367 = u2_col_out_367;
assign col_out_368 = u2_col_out_368;
assign col_out_369 = u2_col_out_369;
assign col_out_370 = u2_col_out_370;
assign col_out_371 = u2_col_out_371;
assign col_out_372 = u2_col_out_372;
assign col_out_373 = u2_col_out_373;
assign col_out_374 = u2_col_out_374;
assign col_out_375 = u2_col_out_375;
assign col_out_376 = u2_col_out_376;
assign col_out_377 = u2_col_out_377;
assign col_out_378 = u2_col_out_378;
assign col_out_379 = u2_col_out_379;
assign col_out_380 = u2_col_out_380;
assign col_out_381 = u2_col_out_381;
assign col_out_382 = u2_col_out_382;
assign col_out_383 = u2_col_out_383;
assign col_out_384 = u2_col_out_384;
assign col_out_385 = u2_col_out_385;
assign col_out_386 = u2_col_out_386;
assign col_out_387 = u2_col_out_387;
assign col_out_388 = u2_col_out_388;
assign col_out_389 = u2_col_out_389;
assign col_out_390 = u2_col_out_390;
assign col_out_391 = u2_col_out_391;
assign col_out_392 = u2_col_out_392;
assign col_out_393 = u2_col_out_393;
assign col_out_394 = u2_col_out_394;
assign col_out_395 = u2_col_out_395;
assign col_out_396 = u2_col_out_396;
assign col_out_397 = u2_col_out_397;
assign col_out_398 = u2_col_out_398;
assign col_out_399 = u2_col_out_399;
assign col_out_400 = u2_col_out_400;
assign col_out_401 = u2_col_out_401;
assign col_out_402 = u2_col_out_402;
assign col_out_403 = u2_col_out_403;
assign col_out_404 = u2_col_out_404;
assign col_out_405 = u2_col_out_405;
assign col_out_406 = u2_col_out_406;
assign col_out_407 = u2_col_out_407;
assign col_out_408 = u2_col_out_408;
assign col_out_409 = u2_col_out_409;
assign col_out_410 = u2_col_out_410;
assign col_out_411 = u2_col_out_411;
assign col_out_412 = u2_col_out_412;
assign col_out_413 = u2_col_out_413;
assign col_out_414 = u2_col_out_414;
assign col_out_415 = u2_col_out_415;
assign col_out_416 = u2_col_out_416;
assign col_out_417 = u2_col_out_417;
assign col_out_418 = u2_col_out_418;
assign col_out_419 = u2_col_out_419;
assign col_out_420 = u2_col_out_420;
assign col_out_421 = u2_col_out_421;
assign col_out_422 = u2_col_out_422;
assign col_out_423 = u2_col_out_423;
assign col_out_424 = u2_col_out_424;
assign col_out_425 = u2_col_out_425;
assign col_out_426 = u2_col_out_426;
assign col_out_427 = u2_col_out_427;
assign col_out_428 = u2_col_out_428;
assign col_out_429 = u2_col_out_429;
assign col_out_430 = u2_col_out_430;
assign col_out_431 = u2_col_out_431;
assign col_out_432 = u2_col_out_432;
assign col_out_433 = u2_col_out_433;
assign col_out_434 = u2_col_out_434;
assign col_out_435 = u2_col_out_435;
assign col_out_436 = u2_col_out_436;
assign col_out_437 = u2_col_out_437;
assign col_out_438 = u2_col_out_438;
assign col_out_439 = u2_col_out_439;
assign col_out_440 = u2_col_out_440;
assign col_out_441 = u2_col_out_441;
assign col_out_442 = u2_col_out_442;
assign col_out_443 = u2_col_out_443;
assign col_out_444 = u2_col_out_444;
assign col_out_445 = u2_col_out_445;
assign col_out_446 = u2_col_out_446;
assign col_out_447 = u2_col_out_447;
assign col_out_448 = u2_col_out_448;
assign col_out_449 = u2_col_out_449;
assign col_out_450 = u2_col_out_450;
assign col_out_451 = u2_col_out_451;
assign col_out_452 = u2_col_out_452;
assign col_out_453 = u2_col_out_453;
assign col_out_454 = u2_col_out_454;
assign col_out_455 = u2_col_out_455;
assign col_out_456 = u2_col_out_456;
assign col_out_457 = u2_col_out_457;
assign col_out_458 = u2_col_out_458;
assign col_out_459 = u2_col_out_459;
assign col_out_460 = u2_col_out_460;
assign col_out_461 = u2_col_out_461;
assign col_out_462 = u2_col_out_462;
assign col_out_463 = u2_col_out_463;
assign col_out_464 = u2_col_out_464;
assign col_out_465 = u2_col_out_465;
assign col_out_466 = u2_col_out_466;
assign col_out_467 = u2_col_out_467;
assign col_out_468 = u2_col_out_468;
assign col_out_469 = u2_col_out_469;
assign col_out_470 = u2_col_out_470;
assign col_out_471 = u2_col_out_471;
assign col_out_472 = u2_col_out_472;
assign col_out_473 = u2_col_out_473;
assign col_out_474 = u2_col_out_474;
assign col_out_475 = u2_col_out_475;
assign col_out_476 = u2_col_out_476;
assign col_out_477 = u2_col_out_477;
assign col_out_478 = u2_col_out_478;
assign col_out_479 = u2_col_out_479;
assign col_out_480 = u2_col_out_480;
assign col_out_481 = u2_col_out_481;
assign col_out_482 = u2_col_out_482;
assign col_out_483 = u2_col_out_483;
assign col_out_484 = u2_col_out_484;
assign col_out_485 = u2_col_out_485;
assign col_out_486 = u2_col_out_486;
assign col_out_487 = u2_col_out_487;
assign col_out_488 = u2_col_out_488;
assign col_out_489 = u2_col_out_489;
assign col_out_490 = u2_col_out_490;
assign col_out_491 = u2_col_out_491;
assign col_out_492 = u2_col_out_492;
assign col_out_493 = u2_col_out_493;
assign col_out_494 = u2_col_out_494;
assign col_out_495 = u2_col_out_495;
assign col_out_496 = u2_col_out_496;
assign col_out_497 = u2_col_out_497;
assign col_out_498 = u2_col_out_498;
assign col_out_499 = u2_col_out_499;
assign col_out_500 = u2_col_out_500;
assign col_out_501 = u2_col_out_501;
assign col_out_502 = u2_col_out_502;
assign col_out_503 = u2_col_out_503;
assign col_out_504 = u2_col_out_504;
assign col_out_505 = u2_col_out_505;
assign col_out_506 = u2_col_out_506;
assign col_out_507 = u2_col_out_507;
assign col_out_508 = u2_col_out_508;
assign col_out_509 = u2_col_out_509;
assign col_out_510 = u2_col_out_510;
assign col_out_511 = u2_col_out_511;
assign col_out_512 = u2_col_out_512;
assign col_out_513 = u2_col_out_513;
assign col_out_514 = u2_col_out_514;
assign col_out_515 = u2_col_out_515;
assign col_out_516 = u2_col_out_516;
assign col_out_517 = u2_col_out_517;
assign col_out_518 = u2_col_out_518;
assign col_out_519 = u2_col_out_519;
assign col_out_520 = u2_col_out_520;
assign col_out_521 = u2_col_out_521;
assign col_out_522 = u2_col_out_522;
assign col_out_523 = u2_col_out_523;
assign col_out_524 = u2_col_out_524;
assign col_out_525 = u2_col_out_525;
assign col_out_526 = u2_col_out_526;
assign col_out_527 = u2_col_out_527;
assign col_out_528 = u2_col_out_528;
assign col_out_529 = u2_col_out_529;
assign col_out_530 = u2_col_out_530;
assign col_out_531 = u2_col_out_531;
assign col_out_532 = u2_col_out_532;
assign col_out_533 = u2_col_out_533;
assign col_out_534 = u2_col_out_534;
assign col_out_535 = u2_col_out_535;
assign col_out_536 = u2_col_out_536;
assign col_out_537 = u2_col_out_537;
assign col_out_538 = u2_col_out_538;
assign col_out_539 = u2_col_out_539;
assign col_out_540 = u2_col_out_540;
assign col_out_541 = u2_col_out_541;
assign col_out_542 = u2_col_out_542;
assign col_out_543 = u2_col_out_543;
assign col_out_544 = u2_col_out_544;
assign col_out_545 = u2_col_out_545;
assign col_out_546 = u2_col_out_546;
assign col_out_547 = u2_col_out_547;
assign col_out_548 = u2_col_out_548;
assign col_out_549 = u2_col_out_549;
assign col_out_550 = u2_col_out_550;
assign col_out_551 = u2_col_out_551;
assign col_out_552 = u2_col_out_552;
assign col_out_553 = u2_col_out_553;
assign col_out_554 = u2_col_out_554;
assign col_out_555 = u2_col_out_555;
assign col_out_556 = u2_col_out_556;
assign col_out_557 = u2_col_out_557;
assign col_out_558 = u2_col_out_558;
assign col_out_559 = u2_col_out_559;
assign col_out_560 = u2_col_out_560;
assign col_out_561 = u2_col_out_561;
assign col_out_562 = u2_col_out_562;
assign col_out_563 = u2_col_out_563;
assign col_out_564 = u2_col_out_564;
assign col_out_565 = u2_col_out_565;
assign col_out_566 = u2_col_out_566;
assign col_out_567 = u2_col_out_567;
assign col_out_568 = u2_col_out_568;
assign col_out_569 = u2_col_out_569;
assign col_out_570 = u2_col_out_570;
assign col_out_571 = u2_col_out_571;
assign col_out_572 = u2_col_out_572;
assign col_out_573 = u2_col_out_573;
assign col_out_574 = u2_col_out_574;
assign col_out_575 = u2_col_out_575;
assign col_out_576 = u2_col_out_576;
assign col_out_577 = u2_col_out_577;
assign col_out_578 = u2_col_out_578;
assign col_out_579 = u2_col_out_579;
assign col_out_580 = u2_col_out_580;
assign col_out_581 = u2_col_out_581;
assign col_out_582 = u2_col_out_582;
assign col_out_583 = u2_col_out_583;
assign col_out_584 = u2_col_out_584;
assign col_out_585 = u2_col_out_585;
assign col_out_586 = u2_col_out_586;
assign col_out_587 = u2_col_out_587;
assign col_out_588 = u2_col_out_588;
assign col_out_589 = u2_col_out_589;
assign col_out_590 = u2_col_out_590;
assign col_out_591 = u2_col_out_591;
assign col_out_592 = u2_col_out_592;
assign col_out_593 = u2_col_out_593;
assign col_out_594 = u2_col_out_594;
assign col_out_595 = u2_col_out_595;
assign col_out_596 = u2_col_out_596;
assign col_out_597 = u2_col_out_597;
assign col_out_598 = u2_col_out_598;
assign col_out_599 = u2_col_out_599;
assign col_out_600 = u2_col_out_600;
assign col_out_601 = u2_col_out_601;
assign col_out_602 = u2_col_out_602;
assign col_out_603 = u2_col_out_603;
assign col_out_604 = u2_col_out_604;
assign col_out_605 = u2_col_out_605;
assign col_out_606 = u2_col_out_606;
assign col_out_607 = u2_col_out_607;
assign col_out_608 = u2_col_out_608;
assign col_out_609 = u2_col_out_609;
assign col_out_610 = u2_col_out_610;
assign col_out_611 = u2_col_out_611;
assign col_out_612 = u2_col_out_612;
assign col_out_613 = u2_col_out_613;
assign col_out_614 = u2_col_out_614;
assign col_out_615 = u2_col_out_615;
assign col_out_616 = u2_col_out_616;
assign col_out_617 = u2_col_out_617;
assign col_out_618 = u2_col_out_618;
assign col_out_619 = u2_col_out_619;
assign col_out_620 = u2_col_out_620;
assign col_out_621 = u2_col_out_621;
assign col_out_622 = u2_col_out_622;
assign col_out_623 = u2_col_out_623;
assign col_out_624 = u2_col_out_624;
assign col_out_625 = u2_col_out_625;
assign col_out_626 = u2_col_out_626;
assign col_out_627 = u2_col_out_627;
assign col_out_628 = u2_col_out_628;
assign col_out_629 = u2_col_out_629;
assign col_out_630 = u2_col_out_630;
assign col_out_631 = u2_col_out_631;
assign col_out_632 = u2_col_out_632;
assign col_out_633 = u2_col_out_633;
assign col_out_634 = u2_col_out_634;
assign col_out_635 = u2_col_out_635;
assign col_out_636 = u2_col_out_636;
assign col_out_637 = u2_col_out_637;
assign col_out_638 = u2_col_out_638;
assign col_out_639 = u2_col_out_639;
assign col_out_640 = u2_col_out_640;
assign col_out_641 = u2_col_out_641;
assign col_out_642 = u2_col_out_642;
assign col_out_643 = u2_col_out_643;
assign col_out_644 = u2_col_out_644;
assign col_out_645 = u2_col_out_645;
assign col_out_646 = u2_col_out_646;
assign col_out_647 = u2_col_out_647;
assign col_out_648 = u2_col_out_648;
assign col_out_649 = u2_col_out_649;
assign col_out_650 = u2_col_out_650;
assign col_out_651 = u2_col_out_651;
assign col_out_652 = u2_col_out_652;
assign col_out_653 = u2_col_out_653;
assign col_out_654 = u2_col_out_654;
assign col_out_655 = u2_col_out_655;
assign col_out_656 = u2_col_out_656;
assign col_out_657 = u2_col_out_657;
assign col_out_658 = u2_col_out_658;
assign col_out_659 = u2_col_out_659;
assign col_out_660 = u2_col_out_660;
assign col_out_661 = u2_col_out_661;
assign col_out_662 = u2_col_out_662;
assign col_out_663 = u2_col_out_663;
assign col_out_664 = u2_col_out_664;
assign col_out_665 = u2_col_out_665;
assign col_out_666 = u2_col_out_666;
assign col_out_667 = u2_col_out_667;
assign col_out_668 = u2_col_out_668;
assign col_out_669 = u2_col_out_669;
assign col_out_670 = u2_col_out_670;
assign col_out_671 = u2_col_out_671;
assign col_out_672 = u2_col_out_672;
assign col_out_673 = u2_col_out_673;
assign col_out_674 = u2_col_out_674;
assign col_out_675 = u2_col_out_675;
assign col_out_676 = u2_col_out_676;
assign col_out_677 = u2_col_out_677;
assign col_out_678 = u2_col_out_678;
assign col_out_679 = u2_col_out_679;
assign col_out_680 = u2_col_out_680;
assign col_out_681 = u2_col_out_681;
assign col_out_682 = u2_col_out_682;
assign col_out_683 = u2_col_out_683;
assign col_out_684 = u2_col_out_684;
assign col_out_685 = u2_col_out_685;
assign col_out_686 = u2_col_out_686;
assign col_out_687 = u2_col_out_687;
assign col_out_688 = u2_col_out_688;
assign col_out_689 = u2_col_out_689;
assign col_out_690 = u2_col_out_690;
assign col_out_691 = u2_col_out_691;
assign col_out_692 = u2_col_out_692;
assign col_out_693 = u2_col_out_693;
assign col_out_694 = u2_col_out_694;
assign col_out_695 = u2_col_out_695;
assign col_out_696 = u2_col_out_696;
assign col_out_697 = u2_col_out_697;
assign col_out_698 = u2_col_out_698;
assign col_out_699 = u2_col_out_699;
assign col_out_700 = u2_col_out_700;
assign col_out_701 = u2_col_out_701;
assign col_out_702 = u2_col_out_702;
assign col_out_703 = u2_col_out_703;
assign col_out_704 = u2_col_out_704;
assign col_out_705 = u2_col_out_705;
assign col_out_706 = u2_col_out_706;
assign col_out_707 = u2_col_out_707;
assign col_out_708 = u2_col_out_708;
assign col_out_709 = u2_col_out_709;
assign col_out_710 = u2_col_out_710;
assign col_out_711 = u2_col_out_711;
assign col_out_712 = u2_col_out_712;
assign col_out_713 = u2_col_out_713;
assign col_out_714 = u2_col_out_714;
assign col_out_715 = u2_col_out_715;
assign col_out_716 = u2_col_out_716;
assign col_out_717 = u2_col_out_717;
assign col_out_718 = u2_col_out_718;
assign col_out_719 = u2_col_out_719;
assign col_out_720 = u2_col_out_720;
assign col_out_721 = u2_col_out_721;
assign col_out_722 = u2_col_out_722;
assign col_out_723 = u2_col_out_723;
assign col_out_724 = u2_col_out_724;
assign col_out_725 = u2_col_out_725;
assign col_out_726 = u2_col_out_726;
assign col_out_727 = u2_col_out_727;
assign col_out_728 = u2_col_out_728;
assign col_out_729 = u2_col_out_729;
assign col_out_730 = u2_col_out_730;
assign col_out_731 = u2_col_out_731;
assign col_out_732 = u2_col_out_732;
assign col_out_733 = u2_col_out_733;
assign col_out_734 = u2_col_out_734;
assign col_out_735 = u2_col_out_735;
assign col_out_736 = u2_col_out_736;
assign col_out_737 = u2_col_out_737;
assign col_out_738 = u2_col_out_738;
assign col_out_739 = u2_col_out_739;
assign col_out_740 = u2_col_out_740;
assign col_out_741 = u2_col_out_741;
assign col_out_742 = u2_col_out_742;
assign col_out_743 = u2_col_out_743;
assign col_out_744 = u2_col_out_744;
assign col_out_745 = u2_col_out_745;
assign col_out_746 = u2_col_out_746;
assign col_out_747 = u2_col_out_747;
assign col_out_748 = u2_col_out_748;
assign col_out_749 = u2_col_out_749;
assign col_out_750 = u2_col_out_750;
assign col_out_751 = u2_col_out_751;
assign col_out_752 = u2_col_out_752;
assign col_out_753 = u2_col_out_753;
assign col_out_754 = u2_col_out_754;
assign col_out_755 = u2_col_out_755;
assign col_out_756 = u2_col_out_756;
assign col_out_757 = u2_col_out_757;
assign col_out_758 = u2_col_out_758;
assign col_out_759 = u2_col_out_759;
assign col_out_760 = u2_col_out_760;
assign col_out_761 = u2_col_out_761;
assign col_out_762 = u2_col_out_762;
assign col_out_763 = u2_col_out_763;
assign col_out_764 = u2_col_out_764;
assign col_out_765 = u2_col_out_765;
assign col_out_766 = u2_col_out_766;
assign col_out_767 = u2_col_out_767;
assign col_out_768 = u2_col_out_768;
assign col_out_769 = u2_col_out_769;
assign col_out_770 = u2_col_out_770;
assign col_out_771 = u2_col_out_771;
assign col_out_772 = u2_col_out_772;
assign col_out_773 = u2_col_out_773;
assign col_out_774 = u2_col_out_774;
assign col_out_775 = u2_col_out_775;
assign col_out_776 = u2_col_out_776;
assign col_out_777 = u2_col_out_777;
assign col_out_778 = u2_col_out_778;
assign col_out_779 = u2_col_out_779;
assign col_out_780 = u2_col_out_780;
assign col_out_781 = u2_col_out_781;
assign col_out_782 = u2_col_out_782;
assign col_out_783 = u2_col_out_783;
assign col_out_784 = u2_col_out_784;
assign col_out_785 = u2_col_out_785;
assign col_out_786 = u2_col_out_786;
assign col_out_787 = u2_col_out_787;
assign col_out_788 = u2_col_out_788;
assign col_out_789 = u2_col_out_789;
assign col_out_790 = u2_col_out_790;
assign col_out_791 = u2_col_out_791;
assign col_out_792 = u2_col_out_792;
assign col_out_793 = u2_col_out_793;
assign col_out_794 = u2_col_out_794;
assign col_out_795 = u2_col_out_795;
assign col_out_796 = u2_col_out_796;
assign col_out_797 = u2_col_out_797;
assign col_out_798 = u2_col_out_798;
assign col_out_799 = u2_col_out_799;
assign col_out_800 = u2_col_out_800;
assign col_out_801 = u2_col_out_801;
assign col_out_802 = u2_col_out_802;
assign col_out_803 = u2_col_out_803;
assign col_out_804 = u2_col_out_804;
assign col_out_805 = u2_col_out_805;
assign col_out_806 = u2_col_out_806;
assign col_out_807 = u2_col_out_807;
assign col_out_808 = u2_col_out_808;
assign col_out_809 = u2_col_out_809;
assign col_out_810 = u2_col_out_810;
assign col_out_811 = u2_col_out_811;
assign col_out_812 = u2_col_out_812;
assign col_out_813 = u2_col_out_813;
assign col_out_814 = u2_col_out_814;
assign col_out_815 = u2_col_out_815;
assign col_out_816 = u2_col_out_816;
assign col_out_817 = u2_col_out_817;
assign col_out_818 = u2_col_out_818;
assign col_out_819 = u2_col_out_819;
assign col_out_820 = u2_col_out_820;
assign col_out_821 = u2_col_out_821;
assign col_out_822 = u2_col_out_822;
assign col_out_823 = u2_col_out_823;
assign col_out_824 = u2_col_out_824;
assign col_out_825 = u2_col_out_825;
assign col_out_826 = u2_col_out_826;
assign col_out_827 = u2_col_out_827;
assign col_out_828 = u2_col_out_828;
assign col_out_829 = u2_col_out_829;
assign col_out_830 = u2_col_out_830;
assign col_out_831 = u2_col_out_831;
assign col_out_832 = u2_col_out_832;
assign col_out_833 = u2_col_out_833;
assign col_out_834 = u2_col_out_834;
assign col_out_835 = u2_col_out_835;
assign col_out_836 = u2_col_out_836;
assign col_out_837 = u2_col_out_837;
assign col_out_838 = u2_col_out_838;
assign col_out_839 = u2_col_out_839;
assign col_out_840 = u2_col_out_840;
assign col_out_841 = u2_col_out_841;
assign col_out_842 = u2_col_out_842;
assign col_out_843 = u2_col_out_843;
assign col_out_844 = u2_col_out_844;
assign col_out_845 = u2_col_out_845;
assign col_out_846 = u2_col_out_846;
assign col_out_847 = u2_col_out_847;
assign col_out_848 = u2_col_out_848;
assign col_out_849 = u2_col_out_849;
assign col_out_850 = u2_col_out_850;
assign col_out_851 = u2_col_out_851;
assign col_out_852 = u2_col_out_852;
assign col_out_853 = u2_col_out_853;
assign col_out_854 = u2_col_out_854;
assign col_out_855 = u2_col_out_855;
assign col_out_856 = u2_col_out_856;
assign col_out_857 = u2_col_out_857;
assign col_out_858 = u2_col_out_858;
assign col_out_859 = u2_col_out_859;
assign col_out_860 = u2_col_out_860;
assign col_out_861 = u2_col_out_861;
assign col_out_862 = u2_col_out_862;
assign col_out_863 = u2_col_out_863;
assign col_out_864 = u2_col_out_864;
assign col_out_865 = u2_col_out_865;
assign col_out_866 = u2_col_out_866;
assign col_out_867 = u2_col_out_867;
assign col_out_868 = u2_col_out_868;
assign col_out_869 = u2_col_out_869;
assign col_out_870 = u2_col_out_870;
assign col_out_871 = u2_col_out_871;
assign col_out_872 = u2_col_out_872;
assign col_out_873 = u2_col_out_873;
assign col_out_874 = u2_col_out_874;
assign col_out_875 = u2_col_out_875;
assign col_out_876 = u2_col_out_876;
assign col_out_877 = u2_col_out_877;
assign col_out_878 = u2_col_out_878;
assign col_out_879 = u2_col_out_879;
assign col_out_880 = u2_col_out_880;
assign col_out_881 = u2_col_out_881;
assign col_out_882 = u2_col_out_882;
assign col_out_883 = u2_col_out_883;
assign col_out_884 = u2_col_out_884;
assign col_out_885 = u2_col_out_885;
assign col_out_886 = u2_col_out_886;
assign col_out_887 = u2_col_out_887;
assign col_out_888 = u2_col_out_888;
assign col_out_889 = u2_col_out_889;
assign col_out_890 = u2_col_out_890;
assign col_out_891 = u2_col_out_891;
assign col_out_892 = u2_col_out_892;
assign col_out_893 = u2_col_out_893;
assign col_out_894 = u2_col_out_894;
assign col_out_895 = u2_col_out_895;
assign col_out_896 = u2_col_out_896;
assign col_out_897 = u2_col_out_897;
assign col_out_898 = u2_col_out_898;
assign col_out_899 = u2_col_out_899;
assign col_out_900 = u2_col_out_900;
assign col_out_901 = u2_col_out_901;
assign col_out_902 = u2_col_out_902;
assign col_out_903 = u2_col_out_903;
assign col_out_904 = u2_col_out_904;
assign col_out_905 = u2_col_out_905;
assign col_out_906 = u2_col_out_906;
assign col_out_907 = u2_col_out_907;
assign col_out_908 = u2_col_out_908;
assign col_out_909 = u2_col_out_909;
assign col_out_910 = u2_col_out_910;
assign col_out_911 = u2_col_out_911;
assign col_out_912 = u2_col_out_912;
assign col_out_913 = u2_col_out_913;
assign col_out_914 = u2_col_out_914;
assign col_out_915 = u2_col_out_915;
assign col_out_916 = u2_col_out_916;
assign col_out_917 = u2_col_out_917;
assign col_out_918 = u2_col_out_918;
assign col_out_919 = u2_col_out_919;
assign col_out_920 = u2_col_out_920;
assign col_out_921 = u2_col_out_921;
assign col_out_922 = u2_col_out_922;
assign col_out_923 = u2_col_out_923;
assign col_out_924 = u2_col_out_924;
assign col_out_925 = u2_col_out_925;
assign col_out_926 = u2_col_out_926;
assign col_out_927 = u2_col_out_927;
assign col_out_928 = u2_col_out_928;
assign col_out_929 = u2_col_out_929;
assign col_out_930 = u2_col_out_930;
assign col_out_931 = u2_col_out_931;
assign col_out_932 = u2_col_out_932;
assign col_out_933 = u2_col_out_933;
assign col_out_934 = u2_col_out_934;
assign col_out_935 = u2_col_out_935;
assign col_out_936 = u2_col_out_936;
assign col_out_937 = u2_col_out_937;
assign col_out_938 = u2_col_out_938;
assign col_out_939 = u2_col_out_939;
assign col_out_940 = u2_col_out_940;
assign col_out_941 = u2_col_out_941;
assign col_out_942 = u2_col_out_942;
assign col_out_943 = u2_col_out_943;
assign col_out_944 = u2_col_out_944;
assign col_out_945 = u2_col_out_945;
assign col_out_946 = u2_col_out_946;
assign col_out_947 = u2_col_out_947;
assign col_out_948 = u2_col_out_948;
assign col_out_949 = u2_col_out_949;
assign col_out_950 = u2_col_out_950;
assign col_out_951 = u2_col_out_951;
assign col_out_952 = u2_col_out_952;
assign col_out_953 = u2_col_out_953;
assign col_out_954 = u2_col_out_954;
assign col_out_955 = u2_col_out_955;
assign col_out_956 = u2_col_out_956;
assign col_out_957 = u2_col_out_957;
assign col_out_958 = u2_col_out_958;
assign col_out_959 = u2_col_out_959;
assign col_out_960 = u2_col_out_960;
assign col_out_961 = u2_col_out_961;
assign col_out_962 = u2_col_out_962;
assign col_out_963 = u2_col_out_963;
assign col_out_964 = u2_col_out_964;
assign col_out_965 = u2_col_out_965;
assign col_out_966 = u2_col_out_966;
assign col_out_967 = u2_col_out_967;
assign col_out_968 = u2_col_out_968;
assign col_out_969 = u2_col_out_969;
assign col_out_970 = u2_col_out_970;
assign col_out_971 = u2_col_out_971;
assign col_out_972 = u2_col_out_972;
assign col_out_973 = u2_col_out_973;
assign col_out_974 = u2_col_out_974;
assign col_out_975 = u2_col_out_975;
assign col_out_976 = u2_col_out_976;
assign col_out_977 = u2_col_out_977;
assign col_out_978 = u2_col_out_978;
assign col_out_979 = u2_col_out_979;
assign col_out_980 = u2_col_out_980;
assign col_out_981 = u2_col_out_981;
assign col_out_982 = u2_col_out_982;
assign col_out_983 = u2_col_out_983;
assign col_out_984 = u2_col_out_984;
assign col_out_985 = u2_col_out_985;
assign col_out_986 = u2_col_out_986;
assign col_out_987 = u2_col_out_987;
assign col_out_988 = u2_col_out_988;
assign col_out_989 = u2_col_out_989;
assign col_out_990 = u2_col_out_990;
assign col_out_991 = u2_col_out_991;
assign col_out_992 = u2_col_out_992;
assign col_out_993 = u2_col_out_993;
assign col_out_994 = u2_col_out_994;
assign col_out_995 = u2_col_out_995;
assign col_out_996 = u2_col_out_996;
assign col_out_997 = u2_col_out_997;
assign col_out_998 = u2_col_out_998;
assign col_out_999 = u2_col_out_999;
assign col_out_1000 = u2_col_out_1000;
assign col_out_1001 = u2_col_out_1001;
assign col_out_1002 = u2_col_out_1002;
assign col_out_1003 = u2_col_out_1003;
assign col_out_1004 = u2_col_out_1004;
assign col_out_1005 = u2_col_out_1005;
assign col_out_1006 = u2_col_out_1006;
assign col_out_1007 = u2_col_out_1007;
assign col_out_1008 = u2_col_out_1008;
assign col_out_1009 = u2_col_out_1009;
assign col_out_1010 = u2_col_out_1010;
assign col_out_1011 = u2_col_out_1011;
assign col_out_1012 = u2_col_out_1012;
assign col_out_1013 = u2_col_out_1013;
assign col_out_1014 = u2_col_out_1014;
assign col_out_1015 = u2_col_out_1015;
assign col_out_1016 = u2_col_out_1016;
assign col_out_1017 = u2_col_out_1017;
assign col_out_1018 = u2_col_out_1018;
assign col_out_1019 = u2_col_out_1019;
assign col_out_1020 = u2_col_out_1020;
assign col_out_1021 = u2_col_out_1021;
assign col_out_1022 = u2_col_out_1022;
assign col_out_1023 = u2_col_out_1023;
assign col_out_1024 = u2_col_out_1024;
assign col_out_1025 = u2_col_out_1025;
assign col_out_1026 = u2_col_out_1026;
assign col_out_1027 = u2_col_out_1027;
assign col_out_1028 = u2_col_out_1028;
assign col_out_1029 = u2_col_out_1029;
assign col_out_1030 = u2_col_out_1030;
assign col_out_1031 = u2_col_out_1031;
assign col_out_1032 = u2_col_out_1032;

endmodule
module xpb_5_490
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5bbe32117faaac629ffd1a7080dc934d3df98065fafbe98e460c86137e7e43859784e038c6a3e2603f64b2a610eee8275c4c00098377fe249d90c09cac923cf0bd3ecd1a72b414604289892459294f4a673d49f33d0dc1611769e4d3bc8198117918004fbc2660d7c49f057c54c2a9865e6717387c601b9ccf3b9d11ca482ea1;
    5'b00010 : xpb = 1024'h6cf1ecd3d6723fc74f4bd09f15edf490a7cfd9b208032a50e3c52d149f9da032bc142f8c3214631df6b26053e7fbf84547dd82ce43d2bfd8a8241db1e520530062e658635d72b7b72790fa61976da63da759a4ded9555b1794737acbed88d90c3286e75c783c922027e2419b1b52ce36df44f8ea874da095807bf1f0badf6d7;
    5'b00011 : xpb = 1024'h628d50debd11d05f14f1d77a723b729648767e011b7c1c335448d8e4c8781d88c346233189c528921ecfd8ab4f6ea7abb0c9d83667b52a2228130277cae44220c36d32a0a88b3fdbb50298ca72a029ae41b2e4412aa3171290b11c807b5a25a23c406ec583aa29f9c71d29960677d669cc5b66c724d4f5a627435c30d5f62578;
    5'b00100 : xpb = 1024'hd9e3d9a7ace47f8e9e97a13e2bdbe9214f9fb364100654a1c78a5a293f3b406578285f186428c63bed64c0a7cff7f08a8fbb059c87a57fb150483b63ca40a600c5ccb0c6bae56f6e4f21f4c32edb4c7b4eb349bdb2aab62f28e6f597db11b218650dceb8f07924404fc4833636a59c6dbe89f1d50e9b412b00f7e3e175bedae;
    5'b00101 : xpb = 1024'h695c6fabfa78f45b89e69484639a51df52f37b9c3bfc4ed862852bb61271f78bef07662a4ce66ec3fe3afeb08dee67300547b0634bf2561fb2954452e9364750c99b9826de626b57277ba8708c1704121c287e8f18386cc409f8542d3a32b332ff68dd3b4b2df31bc99b4dafb82d034d3a4fb655cd49cfaf7f4b1b4fe1a41c4f;
    5'b00110 : xpb = 1024'h146d5c67b8356bf55ede371dd41c9ddb1f76f8d1618097ef2ab4f873dded8e098343c8ea4963d2959e41720fbb7f3e8cfd798886acb783f89f86c5915af60f90128b3092a1858272576b2ef24c648f2b8f60cee9c8c001146bd5a7063c89a8b249794b61568b5b66077a6c4d151f86aa49dceeabf95e8e1c08173d5d2309e485;
    5'b00111 : xpb = 1024'h702b8e7937e01857fedb518e54f931285d7079375c7c817d70c17e875c6bd18f1ac8a9231007b4f5dda624b5cc6e26b459c58890302f821d3d17862e07884c80cfc9fdad143996d299f4b816a58dde75f69e18dd05cdc275833f8bd9f90b40c3c2914bb112b1bc3dcc1971c969e23030a84405e475bea9b8d752da6eed521326;
    5'b01000 : xpb = 1024'h1b3c7b34f59c8ff1d3d2f427c57b7d2429f3f66c8200ca9438f14b4527e7680caf050be30c8518c77dac9814f9fefe1151f760b390f4aff62a09076c794814c018b99618d75cadedc9e43e9865db698f69d66937b65556c5e51cdeb2fb6236430ca1b9d71e0f248809f89066c6d4b38db7d13e3aa1d36825601efc7c2eb7db5c;
    5'b01001 : xpb = 1024'h76faad4675473c5473d00e984658107167ed76d27cfcb4227efdd158a665ab924689ec1bd328fb27bd114abb0aede638ae4360bd146cae1ac799c80925da51b0d5f863334a10c24e0c6dc7bcbf04b8d9d113b32af3631826fc86c386b7e3ce5485b9ba26da35855fce9795e31b975d14163855731e3383c22f5a998df90009fd;
    5'b01010 : xpb = 1024'h220b9a023303b3ee48c7b131b6da5c6d3470f407a280fd39472d9e1671e1420fdac64edbcfa65ef95d17be1a387ebd95a67538e07531dbf3b48b4947979a19f01ee7fb9f0d33d9693c5d4e3e7f5243f3444c0385a3eaac775e64165fba3ac3d3cfca284ce592edaa0c76b4807889e07125c58dc94a48422eb826bb9b3a65d233;
    5'b01011 : xpb = 1024'h7dc9cc13b2ae6050e8c4cba237b6efba726a746d9d7ce6c78d3a2429f05f8595724b2f14964a41599c7c70c0496da5bd02c138e9f8a9da18521c09e4442c56e0dc26c8b97fe7edc97ee6d762d87b933dab894d78e0f86dd875cdfb3376bc5be548e2289ca1b94e81d115b9fccd4c89f7842ca501c6a85dcb876258ad04ae00d4;
    5'b01100 : xpb = 1024'h28dab8cf706ad7eabdbc6e3ba8393bb63eedf1a2c3012fde5569f0e7bbdb1c13068791d492c7a52b3c82e41f76fe7d19faf3110d596f07f13f0d8b22b5ec1f2025166125430b04e4aed65de498c91e571ec19dd391800228d7ab4e0c7913516492f296c2ad16b6cc0ef4d89a2a3f0d5493b9dd57f2bd1c38102e7aba4613c90a;
    5'b01101 : xpb = 1024'h8498eae0f015844d5db988ac2915cf037ce77208bdfd196c9b7676fb3a595f989e0c720d596b878b7be796c587ed6541573f1116dce70615dc9e4bbf627e5c10e2552e3fb5bf1944f15fe708f1f26da185fee7c6ce8dc389ef1532e03594e9760c0a9712693d17a3d393de167f01b6daf220f4906f1d37d4df6a17cc105bf7ab;
    5'b01110 : xpb = 1024'h2fa9d79cadd1fbe732b12b4599981aff496aef3de381628363a643b905d4f6163248d4cd55e8eb5d1bee0a24b57e3c9e4f70e93a3dac33eec98fccfdd43e24502b44c6ab78e23060214f6d8ab23ff8baf93738217f1557da50f285b937ebdef5561b0538749a7fee1172fcb3dbf43a3801ae2ce69b31f641683639d951c1bfe1;
    5'b01111 : xpb = 1024'h8b6809ae2d7ca849d2ae45b61a74ae4c87646fa3de7d4c11a9b2c9cc8453399bc9cdb5061c8ccdbd5b52bccac66d24c5abbce943c124321367208d9a80d06140e88393c5eb9644c063d8f6af0b69480560748214bc23193b685c6a8cf46d7706cf33058830c0e0c5d612023030b6e3be6015441f179211de3771d6eb1c09ee82;
    5'b10000 : xpb = 1024'h3678f669eb391fe3a7a5e84f8af6fa4853e7ecd90401952871e2968a4fced0195e0a17c6190a318efb593029f3fdfc22a3eec16721e95fec54120ed8f290298031732c31aeb95bdb93c87d30cbb6d31ed3acd26f6caaad8bca39bd65f6c46c86194373ae3c1e491013f120cd8da9671b6fa27c7543a6d04ac03df8f85d6fb6b8;
    5'b10001 : xpb = 1024'h9237287b6ae3cc4647a302c00bd38d9591e16d3efefd7eb6b7ef1c9dce4d139ef58ef7fedfae13ef3abde2d004ece44a003ac170a5615e10f1a2cf759f226670eeb1f94c216d703bd652065524e022693aea1c62a9b86eece1a3a239b3460497925b73fdf844a9e7d8902649e26c10a1ce0993adc006ebe78f79960a27b7e559;
    5'b10010 : xpb = 1024'h3d48153728a043e01c9aa5597c55d9915e64ea742481c7cd801ee95b99c8aa1c89cb5abedc2b77c0dac4562f327dbba6f86c999406268be9de9450b410e22eb037a191b7e490875706418cd6e52dad82ae226cbd5a40033d4380f512b59cfa16dc6be22403a21232166f44e73f5e93fedd96cc03ec1baa541845b817691dad8f;
    5'b10011 : xpb = 1024'h99064748a84af042bc97bfc9fd326cde9c5e6ada1f7db15bc62b6f6f1846eda221503af7a2cf5a211a2908d5436ca3ce54b8999d899e8a0e7c251150bd746ba0f4e05ed257449bb748cb15fb3e56fccd155fb6b0974dc49e5aead9e6721e92285583e273bfc87309db0e4a6394213d853bfde33c687bc5f0e78155293365dc30;
    5'b10100 : xpb = 1024'h44173404660767dc918f62636db4b8da68e1e80f4501fa728e5b3c2ce3c2841fb58c9db79f4cbdf2ba2f7c3470fd7b2b4cea71c0ea63b7e76916928f2f3433e03dcff73e1a67b2d278ba9c7cfea487e68898070b47d558eebcc82cbf747587a79f945099cb25db5418ed6900f113c0e24b8b1b929490845d704d773674cba466;
    5'b10101 : xpb = 1024'h9fd56615e5b2143f318c7cd3ee914c27a6db68753ffde400d467c2406240c7a54d117df065f0a052f9942eda81ec6352a93671ca6ddbb60c06a7532bdbc670d0fb0ec4588d1bc732bb4425a157cdd730efd550fe84e31a4fd432119330f71fb918ac50e9874c3c2bdd8c6e7d45d66a68a9f232cb10f09ffa3f8914483f13d307;
    5'b10110 : xpb = 1024'h4ae652d1a36e8bd906841f6d5f139823735ee5aa65822d179c978efe2dbc5e22e14de0b0626e0424999aa239af7d3aafa16849edcea0e3e4f398d46a4d86391043fe5cc4503ede4deb33ac23181b624a630da159356aaea0360f646c334e153862bcbf0f92a9a4761b6b8d1aa2c8edc5b97f6b213d055e66c855365580799b3d;
    5'b10111 : xpb = 1024'ha6a484e32319383ba68139dddff02b70b1586610607e16a5e2a41511ac3aa1a878d2c0e92911e684d8ff54dfc06c22d6fdb449f75218e20991299506fa187601013d29dec2f2f2ae2dbd35477144b194ca4aeb4c727870014d79493fefcfad49dbd4bf5f4ed0054de00a9296f78b974c17e68259b9657a039790d3674ac1c9de;
    5'b11000 : xpb = 1024'h51b5719ee0d5afd57b78dc775072776c7ddbe34586025fbcaad3e1cf77b638260d0f23a9258f4a567905c83eedfcfa33f5e6221ab2de0fe27e1b16456bd83e404a2cc24a861609c95dacbbc931923cae3d833ba723000451af569c18f226a2c925e52d855a2d6d981de9b134547e1aa92773baafe57a3870205cf5748c279214;
    5'b11001 : xpb = 1024'had73a3b060805c381b75f6e7d14f0ab9bbd563ab80fe494af0e067e2f6347baba49403e1ec332cb6b86a7ae4feebe25b5232222436560e071babd6e2186a7b31076b8f64f8ca1e29a03644ed8abb8bf8a4c0859a600dc5b2c6c080ecaea83ada9efd2dd51653ce6fe288b6b0a940c42f85dad1e861da540cef989286566fc0b5;
    5'b11010 : xpb = 1024'h5884906c1e3cd3d1f06d998141d156b58858e0e0a6829261b91034a0c1b0122938d066a1e8b090885870ee442c7cb9b84a63fa47971b3be0089d58208a2a4370505b27d0bbed3544d025cb6f4b09171217f8d5f510955a03289dd3c5b0ff3059e90d9bfb21b136ba2067d54e0633478c95680a3e8def12797864b49397d588eb;
    5'b11011 : xpb = 1024'h3957d27dbf94b6bc5653c1ab253a2b154dc5e15cc06db788140015e8d2ba8a6cd0cc961e52df459f87761a35a0d91154295d26af7e069b8f58ed95efbea0baf994ac03c7f104c60001551f10b56a22b8b31264fc11cee538a7b269eb35625d9331e0a212d0e9f045e46f3eb6325cae9a4f54294ba03d0e60130d6a0d93b5121;
    5'b11100 : xpb = 1024'h5f53af395ba3f7ce6562568b333035fe92d5de7bc702c506c74c87720ba9ec2c6491a99aabd1d6ba37dc14496afc793c9ee1d2747b5867dd931f99fba87c48a056898d56f1c460c0429edb15647ff175f26e7042fe2aafb4a1e50b726fd7bdeaac360a70e934ffdc22e5f967b7e87470035c59cd3663ec82d06c73b2a3837fc2;
    5'b11101 : xpb = 1024'ha649bf519606f683a59f924a3b281fa5f595bb0ec870e1d8f7c542fd72582a9f8ce0c5aa84f3a8bd7e287a8988d50999713aa97dc1d95b680111b3a1a3c10df9f7925c2b4e777db728e619724cd7c8f65a6c09daeb2440503c25e4b722eb369f6467896f492682660c5180514daf7cd12e992236278aaef593895bfe4e947f8;
    5'b11110 : xpb = 1024'h6622ce06990b1bcada571395248f15479d52dc16e782f7abd588da4355a3c62f9052ec936ef31cec17473a4ea97c38c0f35faaa15f9593db1da1dbd6c6ce4dd05cb7f2dd279b8c3bb517eabb7df6cbd9cce40a90ebc005661b2c431f2eb04b7b6f5e78e6b0b8c8fe25641d81699da1537150a95bded8c68c287432d1af317699;
    5'b11111 : xpb = 1024'h1133bac256c79364af4eb62e9511614369d6594c0d0740c29db8a701211f5cad248f4f536b7080bdb74dadadd70d101deb9182c4c05ac1b40a935d15388e160fa5a78b48eabea356e507713d3e4456f3401c5aeb9c4799b67d0995f8310740fab96ee70cbc16314863433c1ec69024b080dde1b20aed84f8b14054def0973ecf;
    endcase
end

endmodule

module xpb_5_240
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6586e6a987c1f9be121243fdf5fda8920596c0b2d5c930de41bb8bc132473ce47e64b164a8e343836694e4c7dadc83e33f69720854f5489cbf2aed07899ee3026136a41a089dfd63ed9efec60944711136c9b37922fa2540343574d307a031e3fb3fd7504be91f87fbb429f195425001b69f75fcca7e9f816cd39333e31c5475;
    5'b00010 : xpb = 1024'h1a6087fd4d95beb3591f1024dba109d299b77e34d61ac145059a5e2cb18bccc0f980e55087a008782dcb8a48d25af6fc1ab8bc2a8737c0edcdb69ab0d86b51534e1e138561aafd82c8a3fae979ad1df1798e6d59b96e1d6fb2de57ab5515c135c7781c76e709468270a86d0432b479da1e650d1744b1e1d29337ab633d56427f;
    5'b00011 : xpb = 1024'h7fe76ea6d557b8716b315422d19eb2649f4e3ee7abe3f2234755e9ede3d309a577e596b530834bfb94606f10ad377adf5a222e32dc2d098a8ce187b8620a3455af54b79f6a48fae6b642f9af82f18f02b05820d2dc6842afe713cc7e5cb5f319c2b7f3c732f2660a6c5c96f5c7f6c9dbd50483140f308154000b3e97207296f4;
    5'b00100 : xpb = 1024'h34c10ffa9b2b7d66b23e2049b74213a5336efc69ac35828a0b34bc5963179981f301caa10f4010f05b971491a4b5edf8357178550e6f81db9b6d3561b0d6a2a69c3c270ac355fb059147f5d2f35a3be2f31cdab372dc3adf65bcaf56aa2b826b8ef038edce128d04e150da086568f3b43cca1a2e8963c3a5266f56c67aac84fe;
    5'b00101 : xpb = 1024'h9a47f6a422ed7724c4506447ad3fbc373905bd1c81feb3684cf0481a955ed66671667c05b8235473c22bf9597f9271db74daea5d6364ca785a9822693a7585a8fd72cb24cbf3f8697ee6f498fc9eacf429e68e2c95d6601f99f22429b1cbb44f8a30103e19fbac8cdd0503f9faab43b5f369902b53e263269342e9fa5dc8d973;
    5'b00110 : xpb = 1024'h4f2197f7e8c13c1a0b5d306e92e31d77cd267a9e825043cf10cf1a8614a36642ec82aff196e0196889629eda7710e4f4502a347f95a742c96923d0128941f3f9ea5a3a902500f88859ebf0bc6d0759d46cab480d2c4a584f189b0701ff4143a156685564b51bd38751f9470c981d6d8e5b2f2745ce15a577b9a70229b802c77d;
    5'b00111 : xpb = 1024'h3fb394bae95010f5269fc9578867eb86147382082a1d435d4adecf193e7f61f679ee3dd759cde5d5099445b6e8f580d2b797ea1c7e9bb1a77af7dbbd80e624ad741a9fb7e0df8a734f0ecdfdd7006b4af7001edc2be507e9743e9da4cb6d2f322a09a8b503bfa81c6ed8a1f358f9766c2f4be604848e7c8e00b1a59123cb587;
    5'b01000 : xpb = 1024'h69821ff53656facd647c40936e84274a66ddf8d3586b0514166978b2c62f3303e60395421e8021e0b72e2923496bdbf06ae2f0aa1cdf03b736da6ac361ad454d38784e1586abf60b228feba5e6b477c5e639b566e5b875becb795ead545704d71de071db9c251a09c2a1b410cad1e7687994345d12c7874a4cdead8cf55909fc;
    5'b01001 : xpb = 1024'h1e5bc148fc2abfc2ab890cba5427888afafeb65558bc957ada484b1e4573c2e0611fc92dfd3ce6d57e64cea440ea4f0946323acc4f217c084566186cb079b39e255fbd80dfb8f629fd94e7c9571d24a628fe6f477c2c6dee4a224185a1cc9428ea18b702374541043795f72368441140e159cb778cfac99b7342c5bc4f92f806;
    5'b01010 : xpb = 1024'h83e2a7f283ecb980bd9b50b84a25311d009577082e85c6591c03d6df77baffc4df847a92a6202a58e4f9b36c1bc6d2ec859bacd4a416c4a5049105743a1896a08696619ae856f38deb33e68f606195b75fc822c09f26932e7e57b658a96cc60ce5588e52832e608c334a2114fd86614297f941745779691ce01658f032af4c7b;
    5'b01011 : xpb = 1024'h38bc494649c07e7604a81cdf2fc8925d94b6348a2ed756bfdfe2a94af6ff8fa15aa0ae7e84dcef4dac3058ed1345460560eaf6f6d6593cf6131cb31d88e504f1737dd1064163f3acc638e2b2d0ca4297a28cdca1359a8b5dfd009930f6e2555eb190d3791e4e8786a83e64279af88b1affbed88ed1acab6e067a711f8ce93a85;
    5'b01100 : xpb = 1024'h9e432fefd182783416ba60dd25c63aef9a4cf53d04a0879e219e350c2946cc85d9055fe32dc032d112c53db4ee21c9e8a05468ff2b4e8592d247a0251283e7f3d4b475204a01f110b3d7e178da0eb3a8d956901a5894b09e31360e03fe828742acd0aac96a37a70ea3f28e19303adb1cb65e4e8b9c2b4aef734e045370058efa;
    5'b01101 : xpb = 1024'h531cd14397563d295dc72d040b699c302e6db2bf04f21804e57d0777a88b5c62542193cf0c7cf7c5d9fbe335e5a03d017ba3b3215d90fde3e0d34dce61505644c19be48ba30ef12f8edcdd9c4a7760891c1b49faef08a8cdafdef0dc4bf816947908eff00557ce0918e6d12bcdad04f51e23e5a6165e8d4099b21c82ca3f7d04;
    5'b01110 : xpb = 1024'h7f672975d2a021ea4d3f92af10cfd70c28e70410543a86ba95bd9e327cfec3ecf3dc7baeb39bcbaa13288b6dd1eb01a56f2fd438fd37634ef5efb77b01cc495ae8353f6fc1bf14e69e1d9bfbae00d695ee003db857ca0fd2e87d3b4996da5e645413516a077f5038ddb143e6b1f2ecd85e97cc09091cf91c01634b224796b0e;
    5'b01111 : xpb = 1024'h6d7d5940e4ebfbdcb6e63d28e70aa602c82530f3db0cd949eb1765a45a1729234da2791f941d003e07c76d7eb7fb33fd965c6f4be4c8bed1ae89e87f39bba7980fb9f81104b9eeb25780d885c4247e7a95a9b754a876c63d62bd4887a10dd7ca40810c66ec61148b898f3e3000617ecf3c88f2bd5b106f132ce9c7e60795bf83;
    5'b10000 : xpb = 1024'h2256fa94aabfc0d1fdf3094fccae07435c45ee75db5e69b0aef6380fd95bb8ffc8bead0b72d9c532cefe12ffaf79a71671abb96e170b3722bd159628888815e8fca1677c5dc6eed13285d4a9348d2b5ad86e71353eeabe6ce1662b5fee83671c0cb9518d87813b85fe8381429dd3a8a7a44e89d7d543b164534de01561cfad8d;
    5'b10001 : xpb = 1024'h87dde13e3281ba9010054d4dc2abafd561dcaf28b1279a8ef0b1c3d10ba2f5e447235e701bbd08b63592f7c78a562af9b1152b766c007fbf7c4083301226f8eb5dd80b966664ec352024d36f3dd19c6c0f3824ae61e4e3ad159ba032f623990007f928ddd36a5b0dfa37ab343315f8a95aedffd49fc250e5c021734944ec0202;
    5'b10010 : xpb = 1024'h3cb78291f8557f8557121974a84f1115f5fd6caab1792af5b490963c8ae785c0c23f925bfa79cdaafcc99d4881d49e128c6475989e42f8108acc30d960f3673c4abf7b01bf71ec53fb29cf92ae3a494c51fcde8ef858dbdc9444830b43992851d4316e046e8a82086f2bee46d0882281c2b396ef19f59336e6858b789f25f00c;
    5'b10011 : xpb = 1024'ha23e693b8017794369245d729e4cb9a7fb942d5d87425bd3f64c21fdbd2ec2a540a443c0a35d112e635e82105cb121f5cbcde7a0f33840ad49f71de0ea924a3eabf61f1bc80fe9b7e8c8ce58b77eba5d88c692081b53011cc879f7de4b395a35cf714554ba73a1906ae0183865ca728379530cebe47432b853591eac82424481;
    5'b10100 : xpb = 1024'h57180a8f45eb3e38b031299983f01ae88fb4eadf8793ec3aba2af4693c735281bbc077ac8219d6232a952791542f950ea71d31c3257ab8fe5882cb8a395eb88f98dd8e87211ce9d6c3cdca7c27e7673dcb8b4be8b1c6f94c4722dab698aee9879ba98a7b5593c88adfd45b4b033c9c5be118a4065ea7750979bd36dbdc7c328b;
    5'b10101 : xpb = 1024'hbf1abe30bbf032df73df5c069937c2923d5a86187e57ca17e09c6d4bbb7e25e36dcab9860d69b17f1cbcd124bae0827826c7be557bd314f670e7933882b26e085c4fdf27a29e9f59ed2c69f9850141e0e5005c9483af17bc5cbbd8ee62478d967e1cfa1f0b3ef8554c89e5da0aec63448de3b20d8dab75aa0214f0b36b62095;
    5'b10110 : xpb = 1024'h7178928c9380fcec095039be5f9124bb296c69145daead7fbfc55295edff1f42b5415cfd09b9de9b5860b1da268a8c0ac1d5ededacb279ec2639663b11ca09e2e6fba20c82c7e7598c71c565a194852f4519b9426b3516bbfa013261edc4aabd6321a6f23c9d0f0d507cc84f35f11635ff7db11da35956dc0cf4e23f19d2750a;
    5'b10111 : xpb = 1024'h265233e05954c1e1505d05e5453485fbbd8d26965e003de683a425016d43af1f305d90e8e876a3901f97575b1e08ff239d25380fdef4f23d34c513e460967833d3e31177dbd4e7786776c18911fd320f87de732301a90eeb78aa153a3b3a3a0f2f59ec18d7bd3607c5710b61d363400e674348381d8c992d3358fa6e740c6314;
    5'b11000 : xpb = 1024'h8bd91a89e116bb9f626f49e33b322e8dc323e74933c96ec4c55fb0c29f8aec03aec2424d9159e713862c3c22f8e58306dc8eaa1833ea3ad9f3f000ebea355b363519b591e472e4dc5515c04f1b41a320bea8269c24a3342bacdf8a0d42da6bf32a99c36923a6558fc125355368a590101de2be34e80b38aea02c8da25728b789;
    5'b11001 : xpb = 1024'h40b2bbdda6ea8094a97c160a20d58fce5744a4cb341aff2b893e832e1ecf7be029de76397016ac084d62e1a3f063f61fb7ddf43a662cb32b027bae953901c987220124fd3d7fe4fb301abc728baa5001016ce07cbb172c5b2b886ce5904ffb44f6d2088fbec67c8a361978660617b9e885a8554f623e7affc690a5d1b162a593;
    5'b11010 : xpb = 1024'ha639a2872eac7a52bb8e5a0816d338605cdb657e09e43009cafa0eef5116b8c4a843279e18f9ef8bb3f7c66bcb407a02f7476642bb21fbc7c1a69b9cc2a0ac898337c917461de25f1db9bb3894eec112383693f5de11519b5fbde1b897f02d28f211dfe00aaf9c1231cda2579b5a09ea3c47cb4c2cbd1a8133643905947efa08;
    5'b11011 : xpb = 1024'h5b1343daf4803f48029b262efc7699a0f0fc23000a35c0708ed8e15ad05b48a1235f5b89f7b6b4807b2e6becc2beed1bd296b064ed647418d0324946116d1ada701f38829f2ae27df8beb75c05576df27afb4dd6748549cade66c490e565bc7abe4a2506a5cfc30ca6c1e56a38cc33c2a40d6266a6f05cd259c85134eeb8e812;
    5'b11100 : xpb = 1024'hfece52eba54043d49a7f255e219fae1851ce0820a8750d752b7b3c64f9fd87d9e7b8f75d67379754265116dba3d6034ade5fa871fa6ec69debdf6ef6039892b5d06a7edf837e29cd3c3b37f75c01ad2bdc007b70af941fa5d0fa76932db4bcc8a826a2d40efea071bb6287cd63e5d9b0bd2f98121239f23802c696448f2d61c;
    5'b11101 : xpb = 1024'h7573cbd84215fdfb5bba3653d817a3738ab3a134e05081b594733f8781e715621ce040da7f56bcf8a8f9f6359519e417ed4f6c8f749c35069de8e3f6e9d86c2dbe3d4c0800d5e000c162b2457f048be3f489bb302df3673a91451c3c3a7b7db085c2417d8cd9098f176a526e6b80ad9cc2726f7deba23ea4ecfffc982c0f2a91;
    5'b11110 : xpb = 1024'h2a4d6d2c07e9c2f0a2c7027abdbb04b41ed45eb6e0a2121c585211f3012ba53e97fc74c65e1381ed70309bb68c985730c89eb6b1a6dead57ac7491a038a4da7eab24bb7359e2e01f9c67ae68ef6d38c4374e7510c4675f6a0fedff1487f10d0251fa86a427f930898c5e958108f2d7752a38069865d580f6136414c78649189b;
    5'b11111 : xpb = 1024'h8fd453d58fabbcaeb4d94678b3b8ad46246b1f69b66b42fa9a0d9db43372e2231661262b06f6c570d6c5807e6774db14080828b9fbd3f5f46b9f7ea7c243bd810c5b5f8d6280dd838a06ad2ef8b1a9d56e182889e76184aa442373e78f913ee64d3a5df473e250118812bf729e352776e0d77c95305420778037a7fb69656d10;
    endcase
end

endmodule

module xpb_5_315
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h69a2842ba3dd031a663c124b38b6de8cbec15239805b01865eef0204a0a77273ed94db2d815c63341ca1ec9b9bf2b13894679a1477bda6956c26d4def2ef51a30ea7a442b7ec8e132b55817b8d079d917dd8ee73bcaa52607ef3fedbc7bc25c1f6f3842d2b10c750ddeb858c4884227b30ad73cc9077d2bf4a29c7f040166fcc;
    5'b00010 : xpb = 1024'h2297c30185cbd16c0172acbf611375c80c0ca1422b3e629540014ab38e4c37dfd7e138e2389247d999e599f0548751a6c4b50c42ccc87cdf27ae6a5fab0c2e94a90013d6c0481ee144110054813376f207ace34eecce77b0485b6bbcd54da8f1bedf7630a55896143517243999381ecd128108b6d0a4484e4de414dbf74a792d;
    5'b00011 : xpb = 1024'h8c3a472d29a8d48667aebf0a99ca5454cacdf37bab99641b9ef04cb82ef3aa53c576140fb9eeab0db687868bf07a02df591ca6574486237493d53f3e9dfb8037b7a7b8197834acf46f6681d00e3b14838585d1c2a978ca10c74f6a989d09ceb3b5d2fa5dd0695d651302a9c5e1bc4148432e7c83611c1b0d980ddccc3760e8f9;
    5'b00100 : xpb = 1024'h452f86030b97a2d802e5597ec226eb9018194284567cc52a800295671c986fbfafc271c471248fb333cb33e0a90ea34d896a18859990f9be4f5cd4bf56185d29520027ad80903dc2882200a90266ede40f59c69dd99cef6090b6d779aa9b51e37dbeec614ab12c286a2e487332703d9a2502116da148909c9bc829b7ee94f25a;
    5'b00101 : xpb = 1024'haed20a2eaf74a5f269216bc9faddca1cd6da94bdd6d7c6b0def1976bbd3fe2339d574cf1f280f2e7506d207c450154861dd1b29a114ea053bb83a99e4907aecc60a7cbf0387ccbd5b37782248f6e8b758d32b511964741c10faad655725777a574b2708e75c1f3794819cdff7af4601555af853a31c0635be5f1f1a82eab6226;
    5'b00110 : xpb = 1024'h67c74904916374440458063e233a61582425e3c681bb27bfc003e01aaae4a79f87a3aaa6a9b6d78ccdb0cdd0fd95f4f44e1f24c86659769d770b3f1f01248bbdfb003b8440d85ca3cc3300fd839a64d61706a9ecc66b6710d91243367fe8fad53c9e6291f009c23c9f456caccba85c6737831a2471ecd8eae9ac3e93e5df6b87;
    5'b00111 : xpb = 1024'h20bc87da735242959f8ea0b24b96f893717132cf2c9e88cea11628c998896d0b71f0085b60ecbc324af47b25b62a95627e6c96f6bb644ce73292d49fb94168af9558ab184933ed71e4ee7fd677c63e36a0da9ec7f68f8c60a279b0178d7a7e05048a54956a5190fff6710b5a1c5c58b91956af0eb2194e79ed668b7f9d1374e8;
    5'b01000 : xpb = 1024'h8a5f0c06172f45b005cab2fd844dd72030328508acf98a5500052ace3930df7f5f84e388e2491f66679667c1521d469b12d4310b3321f37c9eb9a97eac30ba52a4004f5b01207b851044015204cddbc81eb38d3bb339dec1216daef35536a3c6fb7dd8c295625850d45c90e664e07b344a0422db429121393790536fdd29e4b4;
    5'b01001 : xpb = 1024'h43544adbf91e1401a1014d71acaa6e5b7d7dd41157dceb63e117737d26d5a4eb49d1413d997f040be4da15160ab1e7094321a339882cc9c65a413eff644d97443e58beef097c0c5328ff802af8f9b528a8878216e35e0410ead51bd462c826f6c369cac60faa27142b882f93b59477862bd7b7c582bd96c83b4aa05b945dee15;
    5'b01010 : xpb = 1024'hacf6cf079cfb171c073d5fbce5614ce83c3f264ad837ecea40067581c77d175f37661c6b1adb6740017c01b1a6a49841d7893d4dffea705bc66813de573ce8e74d006331c1689a66545501a6860152ba2660708aa008567169c91ab02a844cb8ba5d4ef33abaee650973b51ffe189a015c852b92133569878574684bd4745de1;
    5'b01011 : xpb = 1024'h65ec0ddd7ee9e56da273fa310dbde423898a7553831b4df92118be30b521dccb21b27a1fd2114be57ebfaf065f3938b007d6af7c54f546a581efa95f0f59c5d8e758d2c5c9c42b346d10807f7a2d2c1ab0346565d02c7bc1333087913815cfe8824940f6b502bd28609f53cd4ecc96533e58c07c5361df16892eb5378ba86742;
    5'b01100 : xpb = 1024'h1ee14cb360d8b3bf3daa94a5361a7b5ed6d5c45c2dfeaf08022b06dfa2c6a2370bfed7d48947308afc035c5b17cdd91e382421aaaa001cef3d773edfc776a2ca81b14259d21fbc0285cbff586e59057b3a085a410050a110fc97f47245a753184a3532fa2f4a8bebb7caf27a9f8092a5202c5566938e54a58ce9022342dc70a3;
    5'b01101 : xpb = 1024'h8883d0df04b5b6d9a3e6a6f06ed159eb95971695ae59b08e611a08e4436e14aaf993b3020aa393bf18a548f6b3c08a56cc8bbbbf21bdc384a99e13beba65f46d9058e69c8a0c4a15b12180d3fb60a30cb7e148b4bcfaf3717b8bf34e0d6378da4128b7275a5b533c95b67806e804b52050d9c93324062764d712ca1382f2e06f;
    5'b01110 : xpb = 1024'h41790fb4e6a4852b3f1d4164972df126e2e2659e593d119d422c51933112da16e3e010b6c1d9786495e8f64b6c552ac4fcd92ded76c899ce6525a93f7282d15f2ab156309267dae3c9dcffacef8c7c6d41b53d8fed1f18c144f3602f1af4fc0a0914a92ad4a321ffece216b438b8b17232ad5e1d64329cf3dacd16ff3a26e9d0;
    5'b01111 : xpb = 1024'hab1b93e08a818845a55953afcfe4cfb3a1a3b7d7d9981323a11b5397d1ba4c8ad174ebe44335db98b28ae2e70847dbfd9140c801ee864063d14c7e1e657223023958fa734a5468f6f53281287c9419febf8e2c03a9c96b21c3e75f0ae2b121cc00082d57ffb3e950cacd9c40813cd3ed635ad1e9f4aa6fb324f6deef7a3d599c;
    5'b10000 : xpb = 1024'h6410d2b66c705697408fee23f84166eeeeef06e0847b7432822d9c46bf5f11f6bbc14998fa6bc03e2fce903bc0dc7c6bc18e3a30439116ad8cd4139f1d8efff3d3b16a0752aff9c50dee000170bff35f496220ded9ed90718d4ecbebf042a4fbc7f41f5b79fbb81421f93aedd1f0d03f452e66d434d6e54228b12bdb317162fd;
    5'b10001 : xpb = 1024'h1d06118c4e5f24e8dbc68898209dfe2a3c3a55e92f5ed541633fe4f5ad03d762a60da74db1a1a4e3ad123d9079711cd9f1dbac5e989becf7485ba91fd5abdce56e09d99b5b0b8a9326a97eda64ebccbfd33615ba0a11b5c156b638ccfdd4282b8fe0115ef44386d77924d99b22a4cc912701fbbe75035ad12c6b78c6e8a56c5e;
    5'b10010 : xpb = 1024'h86a895b7f23c280342029ae35954dcb6fafba822afb9d6c7c22ee6fa4dab49d693a2827b32fe0817c9b42a2c1563ce12864346731059938cb4827dfec89b2e887cb17dde12f818a651ff0055f1f36a51510f042dc6bc0821d5aa37a8c5904ded86d3958c1f544e2857105f276b28ef0c57af6f8b057b2d90769540b728bbdc2a;
    5'b10011 : xpb = 1024'h3f9dd48dd42af654dd39355781b173f24846f72b5a9d37d6a3412fa93b500f427deee02fea33ecbd46f7d780cdf86e80b690b8a1656469d6700a137f80b80b7a1709ed721b53a9746aba7f2ee61f43b1dae2f908f6e02d719f11a489d321d11d4ebf878f999c1cebae3bfdd4bbdceb5e3983047545a7a31f7a4f8da2dfefe58b;
    5'b10100 : xpb = 1024'ha94058b97807f96f437547a2ba68527f07084964daf8395d023031addbf781b66b83bb5d6b904ff16399c41c69eb1fb94af852b5dd22106bdc30e85e73a75d1d25b191b4d3403787961000aa7326e14358bbe77cb38a7fd21e05a3659addf6df45b30bbcc4ace43c8c27836104610dd96a307841d61f75dec479559320065557;
    5'b10101 : xpb = 1024'h6235978f59f6c7c0deabe216e2c4e9ba5453986d85db9a6be3427a5cc99c472255d0191222c63496e0dd7171227fc0277b45c4e4322ce6b597b87ddf2bc43a0ec00a0148db9bc855aecb7f836752baa3e28fdc57e3aea521e76d1046a86f7a0f0d9efdc03ef4b2ffe353220e55150a2b4c040d2c164beb6dc833a27ed73a5eb8;
    5'b10110 : xpb = 1024'h1b2ad6653be5961279e27c8b0b2180f5a19ee77630befb7ac454c30bb7410c8e401c76c6d9fc193c5e211ec5db146095ab9337128737bcff5340135fe3e117005a6270dce3f75923c786fe5c5b7e94046c63d13313d2ca71b0d47d27b600fd3ed58aefc3b93c81c33a7ec0bba5c9067d2dd7a216567860fccbedef6a8e6e6819;
    5'b10111 : xpb = 1024'h84cd5a90dfc2992ce01e8ed643d85f82606039afb119fd012343c51057e87f022db151f45b587c707ac30b61770711ce3ffad126fef56394bf66e83ed6d068a3690a151f9be3e736f2dc7fd7e8863195ea3cbfa6d07d1cd22fc87c037dbd2300cc7e73f0e44d4914186a4647ee4d28f85e8515e2e6f033bc1617b75ace84d7e5;
    5'b11000 : xpb = 1024'h3dc29966c1b1677e7b55294a6c34f6bdadab88b85bfd5e1004560dbf458d446e17fdafa9128e6115f806b8b62f9bb23c70484355540039de7aee7dbf8eed4595036284b3a43f78050b97feb0dcb20af67410b48200a14221f92fe8e48b4ea630946a65f45e9517d76f95e4f53f01254a4058aacd271ca94b19d2044685b8e146;
    5'b11001 : xpb = 1024'ha7651d92658e6a98e1913b95a4ebd54a6c6cdaf1dc585f9663450fc3e634b6e205928ad693eac44a14a8a551cb8e637504afdd69cbbde073e715529e81dc9738120a28f65c2c061836ed802c69b9a887f1e9a2f5bd4b94827823e7c0530acbf28b5dea2189a5df284d816a81878547c571061e99b7947c0a63fbcc36c5cf5112;
    5'b11010 : xpb = 1024'h605a5c68477d38ea7cc7d609cd486c85b9b829fa873bc0a544575872d3d97c4defdee88b4b20a8ef91ec52a6842303e334fd4f9820c8b6bda29ce81f39f97429ac62988a648796e64fa8ff055de581e87bbd97d0ed6fb9d2418b54a1609c4f225349dc2503edadeba4ad092ed839441752d9b383f7c0f19967b619227d035a73;
    5'b11011 : xpb = 1024'h194f9b3e296c073c17fe707df5a503c107037903321f21b42569a121c17e41b9da2b464002568d950f2ffffb3cb7a451654ac1c675d38d075e247d9ff216511b46bb081e6ce327b468647dde52115b4905918cac1d93df220af2c1826e2dd2521b35ce287e357caefbd8a7dc28ed406934ad486e37ed67286b70660e343763d4;
    5'b11100 : xpb = 1024'h82f21f69cd490a567e3a82c92e5be24dc5c4cb3cb27a233a8458a3266225b42dc7c0216d83b2f0c92bd1ec96d8aa5589f9b25bdaed91339cca4b527ee505a2be5562ac6124cfb5c793b9ff59df18f8da836a7b1fda3e318289e6c05e35e9f81412295255a94643ffd9c42d68717162e4655abc3ac86539e7b59a2dfe744dd3a0;
    5'b11101 : xpb = 1024'h3be75e3faf37d8a819711d3d56b8798913101a455d5d8449656aebd54fca7999b20c7f223ae8d56ea91599eb913ef5f829ffce09429c09e685d2e7ff9d227fafefbb1bf52d2b4695ac757e32d344d23b0d3e6ffb0a6256d2534e2d3f437b7b43da154459238e12c330efcc15c2255f36472e51250891af76b9547aea2b81dd01;
    5'b11110 : xpb = 1024'ha589e26b5314dbc27fad2f888f6f5815d1d16c7eddb885cfc459edd9f071ec0d9fa15a4fbc4538a2c5b786872d31a730be67681dba59b07bf1f9bcde9011d152fe62c037e517d4a8d7caffae604c6fcc8b175e6ec70ca932d2422c1b0b37a105d108c8864e9eda140edb51a20aa981b177dbc4f199098236037e42da6b984ccd;
    5'b11111 : xpb = 1024'h5e7f21413503aa141ae3c9fcb7cbef511f1cbb87889be6dea56c3688de16b17989edb804737b1d4842fb33dbe5c6479eeeb4da4c0f6486c5ad81525f482eae4498bb2fcbed736576f0867e875478492d14eb5349f730ce829ba998fc18c9243598f4ba89c8e6a8d76606f04f5b5d7e0359af59dbd935f7c507388fc622cc562e;
    endcase
end

endmodule

module xpb_5_760
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h41db9df5eab3b59cfe7e9b972bbc42f9d6a3203330b22a3912098363ba4bbe51b30976cff9437132ce827e5eef8addcf7434a9e1522bc7f11821b45b8daee419e3796a061bd8b204ef01d839efbe362018dae1cdffe3eca04e22c60f9f01d373a802e508f970787aab79be7b7e17a814942b1169ede311890ed56b5e4b65305e;
    5'b00010 : xpb = 1024'h83b73bebd5676b39fcfd372e577885f3ad46406661645472241306c774977ca36612ed9ff286e2659d04fcbddf15bb9ee86953c2a4578fe2304368b71b5dc833c6f2d40c37b16409de03b073df7c6c4031b5c39bffc7d9409c458c1f3e03a6e75005ca11f2e0f0f556f37cf6fc2f5029285622d3dbc623121daad6bc96ca60bc;
    5'b00011 : xpb = 1024'h14e5948bfe2cec0e30765aee72da819c12735d68bc9ede33b83fd0d57be08ded15d3e6f721a3d509cc293bd5eb4288a3f883d5bdd3d0878797c5ddb46e3a379c361d0963a3f918c9ba6b860b365ede2f568babd1732598d034dbc03422dad7c8c9011cf13b8870e27bad54938276d2146da7555b795dd76ae610c716594d2aaf;
    5'b00100 : xpb = 1024'h56c13281e8e0a1ab2ef4f6859e96c495e9167d9bed51086cca495439362c4c3ec8dd5dc71ae7463c9aabba34dacd66736cb87f9f25fc4f78afe7920ffbe91bb619967369bfd1cacea96d5e45261d144f6f668d9f7309857082fe8643c1dcab3c710401fa34f8e95d2727130f008e7a2901d266c56740e8f3f4e63274a4b25b0d;
    5'b00101 : xpb = 1024'h989cd077d39457482d73921cca53078fbfb99dcf1e0332a5dc52d79cf0780a907be6d497142ab76f692e3893ca584442e0ed298078281769c809466b8997ffcffd0fdd6fdbaa7cd3986f367f15db4a6f88416f6d72ed7210d1214c5360de7eb01906e7032e6961d7d2a0d18a7ea6223d95fd782f5523fa7d03bb9dd2f0178b6b;
    5'b00110 : xpb = 1024'h29cb2917fc59d81c60ecb5dce5b5033824e6bad1793dbc67707fa1aaf7c11bda2ba7cdee4347aa13985277abd6851147f107ab7ba7a10f0f2f8bbb68dc746f386c3a12c747f2319374d70c166cbdbc5ead1757a2e64b31a069b7806845b5af91920239e27710e1c4f75aa92704eda428db4eaab6f2bbaed5cc218e2cb29a555e;
    5'b00111 : xpb = 1024'h6ba6c70de70d8db95f6b517411714631fb89db04a9efe6a08289250eb20cda2bdeb144be3c8b1b4666d4f60ac60fef17653c555cf9ccd70047ad6fc46a2353524fb37ccd63cae39863d8e4505c7bf27ec5f23970e62f1e40b7da4677e4b783053a051eeb70815a3fa2d467a283054c3d6f79bc20e09ec05edaf6f98afdff85bc;
    5'b01000 : xpb = 1024'had826503d1c143565de9ed0b3d2d892bd22cfb37daa210d99492a8726c58987d91babb8e35ce8c7935577469b59acce6d970ff3e4bf89ef15fcf241ff7d2376c332ce6d37fa3959d52dabc8a4c3a289edecd1b3ee6130ae105fd0c8783b95678e20803f469f1d2ba4e4e261e011cf45203a4cd8ace81d1e7e9cc64e94964b61a;
    5'b01001 : xpb = 1024'h3eb0bda3fa86c42a916310cb588f84d4375a183a35dc9a9b28bf728073a1a9c7417bb4e564eb7f1d647bb381c1c799ebe98b81397b719696c751991d4aaea6d4a2571c2aebeb4a5d2f429221a31c9a8e03a303745970ca709e93409c6890875a5b0356d3b29952a77307fdba8764763d48f600126c198640b23255430be7800d;
    5'b01010 : xpb = 1024'h808c5b99e53a79c78fe1ac62844bc7ce0dfd386d668ec4d43ac8f5e42ded6818f4852bb55e2ef05032fe31e0b15277bb5dc02b1acd9d5e87df734d78d85d8aee85d0863107c3fc621e446a5b92dad0ae1c7de5425954b710ecb606ac07925ace03063bdcac09cb221e81bc36057c1e51dd21117c59fc97c9c107c0a1574cb06b;
    5'b01011 : xpb = 1024'h11bab43a0dfffa9bc35ad0229fadc376732a556fc1c94e95cef5bff235367962a446250c8d4be2f4622270f8bd7f44c06ddaad15fd16562d46f5c2762b39fa56f4fabb88740bb121faac3ff2e9bd429d4153cd77ccb276a0854c3ac0ec698baf7c018ebbf4b14b0f433b93d28bc3a03d22724403f7944c22896db0fb19cf7a5e;
    5'b01100 : xpb = 1024'h5396522ff8b3b038c1d96bb9cb6a067049cd75a2f27b78cee0ff4355ef8237b4574f9bdc868f542730a4ef57ad0a228fe20f56f74f421e1e5f1776d1b8e8de70d874258e8fe46326e9ae182cd97b78bd5a2eaf45cc966340d36f00d08b6b5f23240473c4ee21c389eeb5524e09db4851b69d556de5775dab98431c596534aabc;
    5'b01101 : xpb = 1024'h9571f025e36765d5c0580750f726496a207095d6232da307f308c6b9a9cdf6060a5912ac7fd2c559ff276db69c95005f564400d8a16de60f77392b2d4697c28abbed8f94abbd152bd8aff066c939aedd73099113cc7a4fe12191c6e02a6d3296cc0758cde7923c049a2f10c987f2f0664ac866d7d35a6f34a71887b7b099db1a;
    5'b01110 : xpb = 1024'h26a048c60c2ce6a9f3d12b1112884512859db2d87e682cc9873590c7b117074fba1a0c03aeefb7fe2e4baccea8c1cd64665e82d3d0e6ddb4debba02a997431f32b17c4ec1804c9ebb517c5fe201c20cc97df79493fd80f70ba27faf50f4463784502abad3039bbf1bee8e8660e3a72519019995f70f2238d6f7e7811731ca50d;
    5'b01111 : xpb = 1024'h687be6bbf6e09c46f24fc6a83e44880c5c40d30baf1a5702993f142b6b62c5a16d2382d3a8332930fcce2b2d984cab33da932cb52312a5a5f6dd54862723160d0e912ef233dd7bf0a4199e380fda56ecb0ba5b173fbbfc11084ac104ae4636ebed0590b629aa346c6a62a6e18c521a662444aac95ed535167e53e36fbe81d56b;
    5'b10000 : xpb = 1024'haa5784b1e19451e3f0ce623f6a00cb0632e3f33edfcc813bab48978f25ae83f3202cf9a3a1769a63cb50a98c87d789034ec7d696753e6d970eff08e1b4d1fa26f20a98f84fb62df5931b7671ff988d0cc9953ce53f9fe8b1566d87144d480a5f950875bf231aace715dc655d0a69c27ab86fbc334cb8469f8d294ece09e705c9;
    5'b10001 : xpb = 1024'h3b85dd520a59d2b8244785ff8562c6ae981110413b070afd3f75619d2cf7953ccfedf2fad0938d07fa74e8a4940456085ee25891a4b7653c76817ddf07ae698f6134ce4fbbfde2b56f834c09567afefbee6b251ab2fda840ef03bb29321f3b410e03c89e6bc22cd43a963cf990b14465fdc0eebaea4ffaf8558f3f27cc69cfbc;
    5'b10010 : xpb = 1024'h7d617b47f50d885522c62196b11f09a86eb430746bb93536517ee500e743538e82f769cac9d6fe3ac8f76703838f33d7d3170272f6e32d2d8ea3323a955d4da944ae3855d7d694ba5e8524434639351c074606e8b2e194e13d268138d1210eb4b606ada76532a54ee60ffb750ec8ec7a91ec0024d8330c816464aa8617cf001a;
    5'b10011 : xpb = 1024'he8fd3e81dd30929563f4556cc810550d3e14d76c6f3bef7e5abaf0eee8c64d832b86321f8f3f0def81ba61b8fbc00dce331846e265c24d2f625a737e839bd11b3d86dad441e497a3aecf9da9d1ba70b2c1bef1e263f5470d5bcb54db5f83f962f020086adda253c0ac9d31195106e65d73d32ac75cac0da2cca9adfda51ca0d;
    5'b10100 : xpb = 1024'h506b71de0886bec654bde0edf83d484aaa846da9f7a5e930f7b53272a8d82329e5c1d9f1f2376211c69e247a7f46deac57662e4f7887ecc40e475b9375e8a12b9751d7b35ff6fb7f29eed2148cd9dd2b44f6d0ec2623411123df7b5d54fa1309d704e58fa74a9db6b643918d1328167a6b68441663add2633ba0063e25b6fa6b;
    5'b10101 : xpb = 1024'h92470fd3f33a7463533c7c8523f98b4481278ddd2858136a09beb5d66323e17b98cb50c1eb7ad3449520a2d96ed1bc7bcb9ad830cab3b4b526690fef039785457acb41b97bcfad8418f0aa4e7c98134b5dd1b2ba26072db17202416cf3fbe67d7f07ca98a0bb163161bd5008913fbe8eff9355805190e3ec4a75719c711c2ac9;
    5'b10110 : xpb = 1024'h237568741bfff53786b5a0453f5b86ece654aadf83929d2b9deb7fe46a6cf2c5488c4a191a97c5e8c444e1f17afe8980dbb55a2bfa2cac5a8deb84ec5673f4ade9f57710e8176243f5587fe5d37a853a82a79aef9964ed410a987581d8d3175ef8031d77e962961e867727a51787407a44e48807ef28984512db61f6339ef4bc;
    5'b10111 : xpb = 1024'h6551066a06b3aad485343bdc6b17c9e6bcf7cb12b444c764aff5034824b8b116fb95c0e913db371b92c760506a8967504fea040d4c58744ba60d3947e422d8c7cd6ee11703f01448e45a581fc338bb5a9b827cbd9948d9e158bb3b9177d4ead2a0060280e2d30e9931f0e620959ee88ed90f9971dd0ba9ce21b0cd547f04251a;
    5'b11000 : xpb = 1024'ha72ca45ff167607183b2d77396d40ce0939aeb45e4f6f19dc1fe86abdf046f68ae9f37b90d1ea84e6149deaf5a14451fc41eadee9e843c3cbe2eeda371d1bce1b0e84b1d1fc8c64dd35c3059b2f6f17ab45d5e8b992cc681a6de01a116d6be464808e789dc438713dd6aa49c13b690a36d3aaadbcaeebb57308638b2ca695578;
    5'b11001 : xpb = 1024'h385afd001a2ce145b72bfb33b2360888f8c8084840317b5f562b50b9e64d80b25e6031103c3b9af2906e1dc766411224d4392fe9cdfd33e225b162a0c4ae2c4a201280748c107b0dafc405f109d96369d93346c10c8a86113f7435b5fbadef27c1043a6924eb070102247c3899fe128eb28bdd6368866faff8ec290c8cec1f6b;
    5'b11010 : xpb = 1024'h7a369af604e096e2b5aa96caddf24b82cf6b287b70e3a5986834d41da0993f041169a7e0357f0c255ef09c2655cbeff4486dd9cb2028fbd33dd316fc525d1064038bea7aa7e92d129ec5de2af9979989f20e288f0c6e72b18d96fbc59aafc29b69071f721e5b7f7bad9e3ab41815baa346b6eecd5669813907c1946ad8514fc9;
    5'b11011 : xpb = 1024'hb64f3962da617b6e923ba8af954472b3498457dcc1e2f59fc619e2ba7e2504dc12aa137649bfec98e14db3e61f8bcf958885bc64fa1f378a5558bf9a5397fcc72b61fd21430e1d27b2db3c2507a0b7916e410c47fcc3241262d2fda7f86f37ce20272516702ff68d25812509e5d3c8e8c082154f4013591d02784c49ad419bc;
    5'b11100 : xpb = 1024'h4d40918c1859cd53e7a2562225108a250b3b65b0fcd059930e6b218f622e0e9f743418075ddf6ffc5c97599d51839ac8ccbd05a7a1cdbb69bd77405532e863e6562f89d8300993d76a2f8bfc403841992fbef2927fb01ee1744ff5ea1e88c6f08a05575a607377e37dd1d0cc1c74e4a3203332bee1e4471adefcf022e6394a1a;
    5'b11101 : xpb = 1024'h8f1c2f82030d82f0e620f1b950cccd1ee1de85e42d8283cc2074a4f31c79ccf1273d8ed75722e12f2b19d7fc410e789840f1af88f3f9835ad598f4b0c097480039a8f3de4be245dc593164362ff677b94899d4607f940b81c272bbf9bd8a9a6432083c6359e3f05e294b8f479a8c8cb7b45e4428cfc758a3edd25b81319e7a78;
    5'b11110 : xpb = 1024'h204a88222bd303c5199a15796c2ec8c7470ba2e688bd0d8db4a16f0123c2de3ad6fe882e863fd3d35a3e17144d3b459d510c318423727b003d1b69ae1373b768a8d32935b829fa9c359939cd86d8e9a86d6fbc95f2f1cb115b08f00ea261cb45ab038f42a28b704b4e0566e420d40ea2f9af76b06d5f0cfcb6384bdaf421446b;
    5'b11111 : xpb = 1024'h622626181686b9621818b11097eb0bc11daec319b96f37c6c6aaf264de0e9c8c8a07fefe7f83450628c095733cc6236cc540db65759e42f1553d1e09a1229b828c4c933bd402aca1249b120776971fc8864a9e63f2d5b7b1a92bb61e41639eb95306744b9bfbe8c5f97f255f9eebb6b78dda881a5b421e85c50db7393f8674c9;
    endcase
end

endmodule

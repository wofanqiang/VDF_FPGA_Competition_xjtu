module xpb_5_395
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h389c38ac4f875f4055cde347473bcc32eabc832c4e077550bfdfc6649c424f407bdc8eb3c2966fc722e55d14587b81f22927ae55e4ec2a3ab4f8d01c262655b9d0b0d2ee457b86e5388a7ba5c5117423fc01600c65339ee42e253dc4846dd824322b341f07eebb74e82cf177f656510dac9fdabf082bc77383c282750c382d1e;
    5'b00010 : xpb = 1024'h713871589f0ebe80ab9bc68e8e779865d57906589c0eeaa17fbf8cc938849e80f7b91d67852cdf8e45caba28b0f703e4524f5cabc9d8547569f1a0384c4cab73a161a5dc8af70dca7114f74b8a22e847f802c018ca673dc85c4a7b8908dbb0486456683e0fdd76e9d059e2efecaca21b593fb57e10578ee7078504ea18705a3c;
    5'b00011 : xpb = 1024'ha9d4aa04ee961dc10169a9d5d5b36498c0358984ea165ff23f9f532dd4c6edc17395ac1b47c34f5568b0173d097285d67b770b01aec47eb01eea70547273012d721278cad07294afa99f72f14f345c6bf40420252f9adcac8a6fb94d8d49886c96819c5d17cc325eb886d467e302f32905df903d1883565a8b47875f24a8875a;
    5'b00100 : xpb = 1024'h31c39d5b7c2f48388c3215460c94e97a397c098062a634cb81a2603cbe068ff9ec29bd564033408dec37350a7e8ff6fe4084917170fdd89f234401125dc6e235ce74170a665d1e4fcf8febf47b6a0c5efc00869908484e8003086517578cbdfe99a53e526ef1f54619f3df00e1891e0d63a58c19d063c09dc89a8ecfa7fe4e0d;
    5'b00101 : xpb = 1024'h6a5fd607cbb6a778e1fff88d53d0b5ad24388cacb0adaa1c418226a15a48df3a68064c0a02c9b0550f1c921ed70b78f069ac3fc755ea02d9d83cd12e83ed37ef9f24e9f8abd8a535081a679a407b8082f801e6a56d7bed64312da2dbdbfa9622cbd0727176e0b0bb0220d078d7df6f1b104566d8d88f88114c5d1144b4367b2b;
    5'b00110 : xpb = 1024'ha2fc0eb41b3e06b937cddbd49b0c81e00ef50fd8feb51f6d0161ed05f68b2e7ae3e2dabdc560201c3201ef332f86fae292d3ee1d3ad62d148d35a14aaa138da96fd5bce6f1542c1a40a4e340058cf4a6f40346b1d2af8c485f52e0a060686e46fdfba6907ecf6c2fea4dc1f0ce35c028bce54197e0bb4f84d01f93b9c06ea849;
    5'b00111 : xpb = 1024'h2aeb020aa8d73130c2964744d1ee06c1883b8fd47744f4464364fa14dfcad0b35c76ebf8bdd01154b5890d00a4a46c0a57e1748cfd0f8703918f320895676eb1cc375b26873eb5ba66955c4331c2a499fbffad25ab5cfe1bd7eb8c6a2aaba3d9011f4885d5f52f174bbacc89ccbbeb0d1aab3d74989bb9c80d729b2a43c46efc;
    5'b01000 : xpb = 1024'h63873ab6f85e907118642a8c1929d2f472f81300c54c69970344c0797c0d1ff3d8537aac8066811bd86e6a14fd1fedfc810922e2e1fbb13e46880224bb8dc46b9ce82e14ccba3c9f9f1fd7e8f6d418bdf8010d3210909d000610ca2eaf197bfd334a7ca4dde3ea8c33e7be01c3123c1ac74b1833a0c7813b91351d9f4ffc9c1a;
    5'b01001 : xpb = 1024'h9c23736347e5efb16e320dd360659f275db4962d1353dee7c32486de184f6f345430096042fcf0e2fb53c729559b6feeaa30d138c6e7db78fb80d240e1b41a256d9901031235c384d7aa538ebbe58ce1f4026d3e75c43be4343607f3338754216575b0c3e5d2a6011c14af79b9688d2873eaf2f2a8f348af14f7a0145c34c938;
    5'b01010 : xpb = 1024'h241266b9d57f1a28f8fa794397472408d6fb16288be3b3c1052793ed018f116cccc41a9b3b6ce21b7edae4f6cab8e1166f3e57a889213567ffda62fecd07fb2dc9fa9f42a8204d24fd9acc91e81b3cd4fbfed3b24e71adb7acceb3bcfdca89b3689952b93cf868e87d81ba12b7eeb80cd1b0eecf60d3b2f2524aa784df8a8feb;
    5'b01011 : xpb = 1024'h5cae9f66250679694ec85c8ade82f03bc1b79954d9eb2911c5075a519dd160ad48a0a94efe0351e2a1c0420b23346308986605fe6e0d5fa2b4d3331af32e50e79aab7230ed9bd40a36254837ad2cb0f8f80033beb3a54c9bdaf3f181823861d79ac486d844e7245d65aeab8aae45091a7e50c98e68ff7a65d60d29f9ebc2bd09;
    5'b01100 : xpb = 1024'h954ad812748dd8a9a4963fd225bebc6eac741c8127f29e6284e720b63a13afedc47d3802c099c1a9c4a59f1f7bafe4fac18db45452f989dd69cc03371954a6a16b5c451f33175aef6eafc3dd723e251cf40193cb18d8eb8009192f4606a639fbccefbaf74cd5dfd24ddb9d02a49b5a282af0a44d712b41d959cfac6ef7faea27;
    5'b01101 : xpb = 1024'h1d39cb69022703212f5eab425ca0415025ba9c7ca082733bc6ea2dc5235352263d11493db909b2e2482cbcecf0cd5622869b3ac41532e3cc6e2593f504a887a9c7bde35ec901e48f94a03ce09e73d50ffbfdfa3ef1865d5381b1db0fd0e96f8dd0135ceca3fba2b9af48a79ba321850c88b6a02a290bac1c9722b3df7b50b0da;
    5'b01110 : xpb = 1024'h55d6041551ae6261852c8e89a3dc0d8310771fa8ee89e88c86c9f429bf95a166b8edd7f17ba022a96b121a014948d814afc2e919fa1f0e07231e64112acedd63986eb64d0e7d6b74cd2ab88663854933f7ff5a4b56b9fc37afd718d4555747b2023e910babea5e2e977599139977d61a35567ae9313773901ae536548788ddf8;
    5'b01111 : xpb = 1024'h8e723cc1a135c1a1dafa71d0eb17d9b5fb33a2d53c915ddd46a9ba8e5bd7f0a734ca66a53e3692708df77715a1c45a06d8ea976fdf0b3841d817342d50f5331d691f893b53f8f25a05b5342c2896bd57f400ba57bbed9b1bddfc5698d9c51fd63469c52ab3d919a37fa28a8b8fce2727e1f655a839633b039ea7b8c993c10b16;
    5'b10000 : xpb = 1024'h166130182eceec1965c2dd4121f95e97747a22d0b52132b688acc79d451792dfad5e77e036a683a9117e94e316e1cb2e9df81ddfa1449230dc70c4eb3c491425c581277ae9e37bfa2ba5ad2f54cc6d4afbfd20cb949b0cef56950262a4085568378d67200afedc8ae10f95248e54520c3fbc5184f143a546dbfac03a1716d1c9;
    5'b10001 : xpb = 1024'h4efd68c47e564b59bb90c08869352aca5f36a5fd0328a807488c8e01e159e220293b0693f93cf3703463f1f76f5d4d20c71fcc358630bc6b91699507626f69df9631fa692f5f02df643028d519dde16ef7fe80d7f9ceabd384ba402728762d8c69b89b3f12ed97ffc93c869c84aaa319ec5c2c43f96f6cba5fbd42af234efee7;
    5'b10010 : xpb = 1024'h8799a170cdddaa9a115ea3cfb070f6fd49f3292951301d58086c54667d9c3160a5179547bbd3633757494f0bc7d8cf12f0477a8b6b1ce6a6466265238895bf9966e2cd5774da89c49cbaa47adeef5592f3ffe0e45f024ab7b2df7debace405b09be3cf5e1adc5374b16978147b00f42798fc0703019b342de37fc5242f872c05;
    5'b10011 : xpb = 1024'hf8894c75b76d5119c270f3fe7527bdec339a924c9bff2314a6f617566dbd3991daba682b443546fdad06cd93cf6403ab55500fb2d5640954abbf5e173e9a0a1c3446b970ac51364c2ab1d7e0b250585fbfc475837afbc8b2b7829b577273b429f0771537202165c12d682ad79871f0bf6c202dfb97b9e7120d2cc94b2dcf2b8;
    5'b10100 : xpb = 1024'h4824cd73aafe3451f1f4f2872e8e4811adf62c5117c767820a4f27da031e22d99988353676d9c436fdb5c9ed9571c22cde7caf5112426acfffb4c5fd9a0ff65b93f53e8550409a49fb359923d03679a9f7fda7649ce35b6f599d6779fb951366d132a57279f0d1d0fb0374256fdd7019a361dd9ec1a765e4a4954f09bf151fd6;
    5'b10101 : xpb = 1024'h80c1061ffa85939247c2d5ce75ca144498b2af7d65cedcd2ca2eee3e9f60721a1564c3ea397033fe209b2701eded441f07a45da6f72e950ab4ad9619c0364c1564a6117395bc212f33c014c99547edcdf3ff07710216fa5387c2a53e8002eb8b035dd99181df8d45e330659d6633c1275001b85dc9d32d582857d17ecb4d4cf4;
    5'b10110 : xpb = 1024'h8aff976881ebe09d28b413eacab992611f92f78de5eb1ac0c31fb4d88a014528df8d52531e02536a42244cf630ab546ccb1e416b967eef9b90726d7ab8a2d1dc107afb32ba6aacf59b08dccc17d9dc0fbfb6de4dac46c27005b51084a46211d06817b86d905502d449d703664b9ec0badc7b43a81b3979b65aad8ef4ea313a7;
    5'b10111 : xpb = 1024'h414c3222d7a61d4a28592485f3e76558fcb5b2a52c6626fccc11c1b224e2639309d563d8f47694fdc707a1e3bb863738f5d9926c9e5419346dfff6f3d1b082d791b882a1712231b4923b0972868f11e4f7fccdf13ff80b0b2e808eccceb3f94138acafa5e0f40ba22cca61ae5b103d195a678ef989df5f0ee96d5b645adb40c5;
    5'b11000 : xpb = 1024'h79e86acf272d7c8a7e2707cd3b23318be77235d17a6d9c4d8bf18816c124b2d385b1f28cb70d04c4e9ecfef81401b92b1f0140c28340436f22f8c70ff7d6d8916269558fb69db899cac585184ba08608f3fe2dfda52ba9ef5ca5cc915321d1656ad7e3c4e8e2c71714f7532651668e27070769b8920b26826d2fddd967136de3;
    5'b11001 : xpb = 1024'h1d75e25b4c6a70208ef733d7204b66d60b8b5ccf2fd7126cdf49525aa64550bfe4603c7af7cf5fd6d741cc5891f2a52e40ec73245799d5e275257cde32ab999becaf3cf4c884239f0b5fe1b77d635fbfbfa94717dd91bc2d53e785b1d6506f76dfb85ba400889fe76645dbf4fecb90b64cd659549eb90c5aa82e549ea693496;
    5'b11010 : xpb = 1024'h3a7396d2044e06425ebd5684b94082a04b7538f94104e6778dd45b8a46a6a44c7a22927b721365c4905979d9e19aac450d3675882a65c798dc4b27ea09510f538f7bc6bd9203c91f294079c13ce7aa1ff7fbf47de30cbaa70363b61fa1d2df1ba026b9d947f745735e914f3746430a19116d4054521758392e4567bef6a161b4;
    5'b11011 : xpb = 1024'h730fcf7e53d56582b48b39cc007c4ed33631bc258f0c5bc84db421eee2e8f38cf5ff212f34a9d58bb33ed6ee3a162e37365e23de0f51f1d39143f8062f77650d602c99abd77f500461caf56701f91e43f3fd548a4840598b3188f3e42640b73fd251edf84fe600e846be40af3c995b26be0d1b135a431facb207ea3402d98ed2;
    5'b11100 : xpb = 1024'habac082aa35cc4c30a591d1347b81b0620ee3f51dd13d1190d93e8537f2b42cd71dbafe2f7404552d62434029291b0295f85d233f43e1c0e463cc822559dbac730dd6c9a1cfad6e99a55710cc70a9267effeb496ad73f86f5fae31a8aaae8f64047d221757d4bc5d2eeb322732efac346aacf5d2626ee72035ca6ca90f11bbf0;
    5'b11101 : xpb = 1024'h339afb8130f5ef3a952188837e999fe79a34bf4d55a3a5f24f96f562686ae505ea6fc11defb0368b59ab51d007af2151249358a3b67775fd4a9658e040f19bcf8d3f0ad9b2e56089c045ea0ff340425af7fb1b0a86216a42d846dd7274f1c4f607a0c40caefa7f4490583cc03175d718c872f1af1a4f5163731d7419926782a3;
    5'b11110 : xpb = 1024'h6c37342d807d4e7aeaef6bcac5d56c1a84f14279a3ab1b430f76bbc704ad3446664c4fd1b246a6527c90aee4602aa3434dbb06f99b63a037ff8f28fc6717f1895defddc7f860e76ef8d065b5b851b67ef3fc7b16eb550927066c1b36f95f9d1a39cbf82bb6e93ab978852e3827cc28267512cc6e227b18d6f6dff68e9e9fafc1;
    5'b11111 : xpb = 1024'ha4d36cd9d004adbb40bd4f120d11384d6fadc5a5f1b29093cf56822ba0ef8386e228de8574dd16199f760bf8b8a6253576e2b54f804fca72b487f9188d3e47432ea0b0b63ddc6e54315ae15b7d632aa2effddb235088a80b349158fb7dcd753e6bf72c4abed7f62e60b21fb01e22793421b2a72d2aa6e04a7aa27903aad7dcdf;
    endcase
end

endmodule

module xpb_5_1015
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7cea60f163ebe675c2bf399b02e5a8ad3acc9a15a2021f8db25369a33f4ee4982ba99767f2eb404b0dcd51424d913d00fead2ff4c515d299a9b5567cc2399495d6c157022fe2811186afcb2b1c94ada07d4544b3c3c296dd9493915b76d8d92a4c93861b84c00d2fdc193a81339793785c4599ce06930d8451ab809a9d08c6b8;
    5'b00010 : xpb = 1024'h49277c8d05e99822ba78fb5ef5710a09042330fa6e8c9ea3e6ca19f0cb9b1c28540ab1571bb002077c3c633db7c46937994038036778d4e7a2cb6d9b49a0b47a39337955b03404ddfac593b3a04d971006858fcefaff00aa739a90bc33870fc26a1f7a0d58b721d231728e236f5f00c769b154b9bcdabdd85ce78630b12f2705;
    5'b00011 : xpb = 1024'h15649828a7e749cfb232bd22e7fc6b64cd79c7df3b171dba1b40ca3e57e753b87c6bcb464474c3c3eaab753921f7956e33d3401209dbd7359be184b9d107d45e9ba59ba9308588aa6edb5c3c2406807f8fc5daea323b6a7752a1901cf035465a87ab6dff2cae367486cbe1c5ab266e16771d0fa573226e2c68238bc6c5558752;
    5'b00100 : xpb = 1024'h924ef91a0bd3304574f1f6bdeae21412084661f4dd193d47cd9433e197363850a81562ae3760040ef878c67b6f88d26f32807006cef1a9cf4596db36934168f47266f2ab606809bbf58b2767409b2e200d0b1f9df5fe0154e7352178670e1f84d43ef41ab16e43a462e51c46debe018ed362a97379b57bb0b9cf0c61625e4e0a;
    5'b00101 : xpb = 1024'h5e8c14b5add0e1f26cabb881dd6d756dd19cf8d9a9a3bc5e020ae42f23826fe0d0767c9d6024c5cb66e7d876d9bbfea5cd1378157154ac1d3eacf2551aa888d8d4d914fee0b98d8869a0efefc454178f964b6ab92d3a6b21c63c20d923bc561cf1cae80c85655846b83e6fe91a856edde0ce645f2ffd2c04c50b11f77684ae57;
    5'b00110 : xpb = 1024'h2ac930514fce939f64657a45cff8d6c99af38fbe762e3b743681947cafcea770f8d7968c88e98787d556ea7243ef2adc67a6802413b7ae6b37c30973a20fa8bd374b3752610b1154ddb6b878480d00ff1f8bb5d46476d4eea5432039e06a8cb50f56dbfe595c6ce90d97c38b564cdc2cee3a1f4ae644dc58d047178d8aab0ea4;
    5'b00111 : xpb = 1024'ha7b39142b3ba7a152724b3e0d2de7f76d5c029d418305b01e8d4fe1fef1d8c0924812df47bd4c7d2e3243bb4918067dd6653b018d8cd8104e1785ff064493d530e0c8e5490ed9266646683a364a1ae9f9cd0fa8828396bcc39d6b195574365df5bea6219de1c7a18e9b0fe0c89e46fa54a7fb918ecd7e9dd21f2982827b3d55c;
    5'b01000 : xpb = 1024'h73f0acde55b82bc21ede75a4c569e0d29f16c0b8e4bada181d4bae6d7b69c3994ce247e3a499898f51934daffbb3941400e6b8277b308352da8e770eebb05d37707eb0a8113f1632d87c4c2be85a980f261145a35f75d59918ddb0f613f19c777976560bb2138ebb3f0a51aec5abdcf457eb7404a31f9a312d2e9dbe3bda35a9;
    5'b01001 : xpb = 1024'h402dc879f7b5dd6f16983768b7f5422e686d579db145592e51c25ebb07b5fb29754361d2cd5e4b4bc0025fab65e6c04a9b79c0361d9385a0d3a48e2d73177d1bd2f0d2fb919099ff4c9214b46c13817eaf5190be96b23f65f7e4b056d09fd30f970249fd860aa35d9463a55101734a4365572ef059674a85386aa354500095f6;
    5'b01010 : xpb = 1024'hc6ae41599b38f1c0e51f92caa80a38a31c3ee827dcfd84486390f08940232b99da47bc1f6230d082e7171a6d019ec81360cc844bff687eeccbaa54bfa7e9d003562f54f11e21dcbc0a7dd3cefcc6aee3891dbd9cdeea932d6ebafb78d4e09a7b48e3def5a01b7ffe9bcf8f33d3ab79272c2e9dc0faefad943a6a8ea6426f643;
    5'b01011 : xpb = 1024'h89554506fd9f7591d11132c7ad664c376c9088981fd1f7d2388c78abd3511751c94e1329e90e4d533c3ec2e91dab298234b9f839850c5a88766ffbc8bcb831960c244c5141c49edd4757a8680c61188eb5d7208d91b140106b7f41130426e2d20121c40adec1c52fc5d6337470d24b0acf0883aa1642085d95522985012fbcfb;
    5'b01100 : xpb = 1024'h559260a29f9d273ec8caf48b9ff1ad9335e71f7cec5c76e86d0328f95f9d4ee1f1af2d1911d30f0faaadd4e487de55b8cf4d0048276f5cd66f8612e7441f517a6e966ea4c21622a9bb6d70f0901a01fe3f176ba8c8eda9dd4a864073c0d5196a1eadb7fcb2b8d9d21b2f8716ac99b859dc743e95cc89b8b1a08e2f1b15561d48;
    5'b01101 : xpb = 1024'h21cf7c3e419ad8ebc084b64f927d0eeeff3db661b8e6f5fea179d946ebe986721a1047083a97d0cc191ce6dff21181ef69e00856c9d25f24689c2a05cb86715ed10890f84267a6762f83397913d2eb6dc857b6c4002a13aa298d3fd47d8350023c39abee86afee747088dab8e86125a8e9dff98182d16905abca34b1297c7d95;
    5'b01110 : xpb = 1024'h9eb9dd2fa586bf618343efea9562b79c3a0a50775ae9158c53cd42ea2b386b0a45b9de702d83111726ea38223fa2bef0688d384b8ee831be125180828dc005f4a7c9e7fa724a2787b63304a43067990e459cfb77c3ecaa87be20d12ff45c292c88cd320a0b6ffba44ca2153a1bf8b9214625934f89647689fd75b54bc685444d;
    5'b01111 : xpb = 1024'h6af6f8cb4784710e7afdb1ae87ee18f80360e75c277394a28843f337b784a29a6e1af85f5647d2d395594a1da9d5eb270320405a314b340c0b6797a1152725d90a3c0a4df29bab542a48cd2cb420827dcedd4692fb2914549d27d090b10a5fc4a65925fbdf671046a1fb68dc57c0267053914e3b3fac26de08b1bae1daaba49a;
    5'b10000 : xpb = 1024'h37341466e98222bb72b773727a797a53ccb77e40f3fe13b8bcbaa38543d0da2a967c124e7f0c949003c85c191409175d9db34868d3ae365a047daebf9c8e45bd6cae2ca172ed2f209e5e95b537d96bed581d91ae32657e217c2ecff16db8965cc3e519edb35e24e8f754bc7e938793bf60fd0926f5f3d73213edc077eed204e7;
    5'b10001 : xpb = 1024'h37130028b7fd4686a7135366d04dbaf960e1525c08892cef13153d2d01d11babedd2c3da7d1564c72376e147e3c439438465077761138a7fd93c5de23f565a1cf204ef4f33eb2ed12745e3dbb92555ce15ddcc969a1e7ee5b35cf522a66ccf4e1710ddf8755398b4cae1020cf4f010e6e68c412ac3b87861f29c60e02f86534;
    5'b10010 : xpb = 1024'h805b90f3ef6bbade2d306ed16fea845cd0daaf3b628ab25ca384bd760f6bf652ea86c3a59abc96978004bf56cbcd809536f3806c3b270b41a7491c5ae62efa37a5e1a5f7232133fe99242968d82702fd5ea3217d2d647ecbefc960ada13fa61f2e0493fb0c1546bb28c74aa202e69486caae5de0b2ce950a70d546a8a0012bec;
    5'b10011 : xpb = 1024'h4c98ac8f91696c8b24ea30956275e5b89a3146202f153172d7fb6dc39bb82de312e7dd94c3815853ee73d1523600accbd186887add8a0d8fa05f33796d961a1c0853c84aa372b7cb0d39f1f15bdfec6ce7e36c9864a0e898ced0600e5deddcb74b9087ece00c5b5d7e209e443eae01d5d81a18cc6916455e7c114c3eb4278c39;
    5'b10100 : xpb = 1024'h18d5c82b33671e381ca3f259550147146387dd04fb9fb0890c721e11280465733b48f783ec461a105ce2e34da033d9026c1990897fed0fdd99754a97f4fd3a006ac5ea9e23c43b97814fba79df98d5dc7123b7b39bdd5265add75f6f1a9c134f691c7bdeb4036fffd379f1e67a756f24e585d3b81f5df5b2874d51d4c84dec86;
    5'b10101 : xpb = 1024'h95c0291c975304addf632bf457e6efc19e54771a9da1d016bec587b467534a0b66f28eebdf315a5b6ab0348fedc516036ac6c07e4502e277432aa114b736ce96418741a053a6bca907ff85a4fc2d837cee68fc675f9fe943426af0ca9174ec79b5b001fa38c37d2faf932c67ae0d029d41cb6d8625f10336d8f8d26f6556b33e;
    5'b10110 : xpb = 1024'h61fd44b83950b65ad71cedb84a72511d67ab0dff6a2c4f2cf33c3801f39f819b8f53a8db07f61c17d91f468b57f8423a0559c88ce765e4c53c40b8333e9dee7aa3f963f3d3f840757c154e2d7fe66cec77a9478296dc53102171f02b4e232311d33bf5ec0cba91d204ec8009e9d46fec4f372871dc38b38ae434d805797d138b;
    5'b10111 : xpb = 1024'h2e3a6053db4e6807ced6af7c3cfdb2793101a4e436b6ce4327b2e84f7febb92bb7b4c2ca30baddd4478e5886c22b6e709fecd09b89c8e7133556cf51c6050e5f066b86475449c441f02b16b6039f565c00e9929dce18bcdd0078ef8c0ad159a9f0c7e9dde0b1a6745a45d3ac259bdd3b5ca2e35d928063deef70dd9b8da373d8;
    5'b11000 : xpb = 1024'hab24c1453f3a4e7d9195e9173fe35b266bce3ef9d8b8edd0da0651f2bf3a9dc3e35e5a3223a61e1f555ba9c90fbcab719e9a00904edeb9acdf0c25ce883ea2f4dd2cdd49842c455376dae1e1203403fc7e2ed75191db53ba950c80e781aa32d43d5b6ff96571b3a4365f0e2d593370b3b8e87d2b99137163411c5e362aac3a90;
    5'b11001 : xpb = 1024'h7761dce0e138002a894faadb326ebc823524d5dea5436ce70e7d02404b86d5540bbf74214c6adfdbc3cabbc479efd7a8392d089ef141bbfad8223ced0fa5c2d93f9eff9d047dc91feaf0aa69a3eced6c076f226cc917bd87741380483e58696c5ae763eb3968c8468bb861cf94fade02c65438174f5b21b74c5863cc3ed29add;
    5'b11010 : xpb = 1024'h439ef87c8335b1d781096c9f24fa1dddfe7b6cc371cdebfd42f3b28dd7d30ce434208e10752fa1983239cdbfe42303ded3c010ad93a4be48d138540b970ce2bda21121f084cf4cec5f0672f227a5d6db90af6d8800542754531a7fa8fb06a004787357dd0d5fdce8e111b571d0c24b51d3bff30305a2d20b5794696252f8fb2a;
    5'b11011 : xpb = 1024'hfdc14182533638478c32e6317857f39c7d203a83e586b13776a62db641f44745c81a7ff9df46354a0a8dfbb4e5630156e5318bc3607c096ca4e6b2a1e7402a2048344440520d0b8d31c3b7aab5ec04b19efb8a33790912132217f09b7b4d69c95ff4bcee156f18b366b09140c89b8a0e12badeebbea825f62d06ef8671f5b77;
    5'b11100 : xpb = 1024'h8cc67509891f49fa3b8267fe1a6b27e7029e9dbde05a8aa129bdcc7ea36e290c882b3f6790dfa39fae7630fd9be76d166d0048b0fb1d93307403c1a6e0ad9737db449b46350351ca59cc06a5c7f36deb9734fd56fb5327fec6b510652e8dafc6e292d1ea6616febb1284439540214c193d7147bcc27d8fe3b47bef930428222f;
    5'b11101 : xpb = 1024'h590390a52b1cfba7333c29c20cf68942cbf534a2ace509b75e347ccc2fba609cb08c5956b9a4655c1ce542f9061a994d079350bf9d80957e6d19d8c56814b71c3db6bd99b554d596cde1cf2e4bac575b20754872328f91cba5bc0fc5eb3be65f001ec5dc3a0e135d67dd97377be8b9684add02a878c54037bfb7f529184e827c;
    5'b11110 : xpb = 1024'h2540ac40cd1aad542af5eb85ff81ea9e954bcb87796f88cd92ab2d19bc06982cd8ed7345e26927188b5454f4704dc583a22658ce3fe397cc662fefe3ef7bd700a028dfed35a6596341f797b6cf6540caa9b5938d69cbfb9884c30f26a7ea1cf71daab9ce0e0527ffbd36ead9b7b026b75848bd942f0cf08bcaf3fabf2c74e2c9;
    5'b11111 : xpb = 1024'ha22b0d32310693c9edb525210267934bd018659d1b71a85b44fe96bcfb557cc504970aadd55467639921a636bddf0284a0d388c304f96a660fe54660b1b56b9676ea36ef6588da74c8a762e1ebf9ee6b26fad8412d8e92761956a0821ec2f6216a3e3fe992c5352f9950255aeb47ba2fb48e5762359ffe101c9f7b59c97da981;
    endcase
end

endmodule

module xpb_5_205
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9c0f8ddf46cf47d59f7cc6e8d51171de1c2e4712488c4f37b65370f9f0d4e4ca88befad793c2549fbc56a32c232fb1a2905d746324f0a2d89286b110b0874c7b1a3723780cd02968ebc1d41a0b30cfcd68f35a0cb668c8eba0bc840b348fe819b16fff78b3bd7a9c40187b30099a1368fe05b22404a5a344eebf73cd85f81021;
    5'b00010 : xpb = 1024'h8771d668cbb05ae273f415fa99c89c6ac6e68af3bba0fdf7eeca289e2ea71c8d0e3578365d5e2ab0d94f07116301527abca0c0e0272e7565746e22c3263c2444c01f12416a0f558cc4e9a5917d85db69dde1ba80e04b64c68bec761baef52da133d86cc7b6b1fcaaf9710f811b6400a8ad318565b8ffe959970f6c96830db9d7;
    5'b00011 : xpb = 1024'h72d41ef250916def486b650c5e7fc6f7719eced52eb5acb82740e0426c79544f93abf59526fa00c1f6476af6a2d2f352e8e40d5d296c47f2565594759bf0fc0e6607010ac74e81b09e117708efdae70652d01af50a2e00a1771c682c295a7328b640da16b9a67eb9b2c9a3d22d2dede85c5d58a76d5a2f6e3f5f655f8023638d;
    5'b00100 : xpb = 1024'h5e36677bd57280fc1ce2b41e2336f1841c5712b6a1ca5b785fb797e6aa4b8c12192272f3f095d6d3133fcedbe2a4942b152759da2baa1a7f383d062811a5d3d80beeefd4248dadd477394880622ff2a2c7be7b6934109c7c624c5a3ca3bfb8b038a94765bc9b00c86c2238233ef7db280b892be921b47582e7af5e287d390d43;
    5'b00101 : xpb = 1024'h4998b0055a539408f15a032fe7ee1c10c70f569814df0a38982e4f8ae81dc3d49e98f052ba31ace4303832c122763503416aa6572de7ed0c1a2477da875aaba1b1d6de9d81ccd9f8506119f7d484fe3f3cacdbdd5df338574d7c4c4d1e24fe37bb11b4b4bf8f82d7257acc7450c1c867bab4ff2ad60ebb978fff56f17a4eb6f9;
    5'b00110 : xpb = 1024'h34faf88edf34a715c5d15241aca5469d71c79a7987f3b8f8d0a5072f25effb97240f6db183cd82f54d3096a66247d5db6dadf2d43025bf98fc0be98cfd0f836b57becd66df0c061c2988eb6f46da09dbb19b3c5187d5d43238ac3e5d988a43bf3d7a2203c28404e5ded360c5628bb5a769e0d26c8a6901ac384f4fba776460af;
    5'b00111 : xpb = 1024'h205d41186415ba229a48a153715c712a1c7fde5afb0867b9091bbed363c23359a985eb104d6959066a28fa8ba21976b399f13f5132639225ddf35b3f72c45b34fda6bc303c4b324002b0bce6b92f157826899cc5b1b8700d23dc306e12ef8946bfe28f52c57886f4982bf5167455a2e7190ca5ae3ec347c0e09f4883747a0a65;
    5'b01000 : xpb = 1024'hbbf89a1e8f6cd2f6ebff06536139bb6c738223c6e1d167941927677a1946b1c2efc686f17052f1787215e70e1eb178bc6348bce34a164b2bfdaccf1e87932fea38eaaf9998a5e63dbd88e5e2b8421149b77fd39db9b0be80f0c227e8d54cece424afca1c86d090351848967861f9026c83878eff31d8dd588ef414c718fb41b;
    5'b01001 : xpb = 1024'ha7cf17812fc615050e3cb74e0b250d94e366694eb6a965b0f7e5e77192694fe6b7bb6346aac783b74378019d051ac92e569200315992078b52617e0299007f79bdc5ce71a65a87ccc79a627836b4f0e2046b57469203d4d3afc8a689c1e4b6e7f3bafc1a7c2a839f919d04978fb9a38fc63e2b13f7c3311a77aeb519f787c43c;
    5'b01010 : xpb = 1024'h9331600ab4a72811e2b4065fcfdc38218e1ead3029be1471305c9f15d03b87a93d31e0a5746359c86070658244ec6a0682d54cae5bcfda183448efb50eb5574363adbd3b0399b3f0a0c233efa909fc7e7959b7babbe670ae9af8989a3c49fc6f762369697f1f05ae4af598e8a18390cf7569fe55ac1d772f1ffeade2f49d6df2;
    5'b01011 : xpb = 1024'h7e93a89439883b1eb72b5571949362ae38d6f1119cd2c33168d356ba0e0dbf6bc2a85e043dff2fd97d68c96784be0adeaf18992b5e0daca516306167846a2f0d0995ac0460d8e01479ea05671b5f081aee48182ee5c90c8986288aaab6af41f6f88bd6b8821387bd044e2d39b34d7e0f2495d1976077bd43c84ea6abf1b317a8;
    5'b01100 : xpb = 1024'h69f5f11dbe694e2b8ba2a483594a8d3ae38f34f30fe771f1a14a0e5e4bdff72e481edb63079b05ea9a612d4cc48fabb6db5be5a8604b7f31f817d319fa1f06d6af7d9acdbe180c385311d6de8db413b7633678a30faba86471587cbb3114877e7af44407850809cbbda6c18ac5176b4ed3c1a4d914d20358709e9f74eec8c15e;
    5'b01101 : xpb = 1024'h555839a7434a61386019f3951e01b7c78e4778d482fc20b1d9c0c60289b22ef0cd9558c1d136dbfbb759913204614c8f079f3225628951bed9ff44cc6fd3dea0556589971b57385c2c39a85600091f53d824d917398e443f5c886ecbab79cd05fd5cb15687fc8bda76ff55dbd6e1588e82ed781ac92c496d18ee983debde6b14;
    5'b01110 : xpb = 1024'h40ba8230c82b7445349142a6e2b8e25438ffbcb5f610cf7212377da6c78466b3530bd6209ad2b20cd451f5174432ed6733e27ea264c7244bbbe6b67ee588b669fb4d786078966480056179cd725e2af04d13398b6370e01a47b860dc25df128d7fc51ea58af10de93057ea2ce8ab45ce32194b5c7d868f81c13e9106e8f414ca;
    5'b01111 : xpb = 1024'h2c1ccaba4d0c8752090891b8a7700ce0e3b8009769257e324aae354b05569e75d882537f646e881df14a58fc84048e3f6025cb1f6704f6d89dce28315b3d8e33a1356729d5d590a3de894b44e4b3368cc20199ff8d537bf532e852eca0445815022d8bf48de58ff7e9b07e7dfa75330de1451e9e31e0d596698e89cfe609be80;
    5'b10000 : xpb = 1024'h177f1343d1ed9a5edd7fe0ca6c27376d8e704478dc3a2cf28324ecef4328d6385df8d0de2e0a5e2f0e42bce1c3d62f178c69179c6942c9657fb599e3d0f265fd471d55f33314bcc7b7b11cbc5708422936effa73b73617d01e1844fd1aa99d9c8495f94390da1206a30912cf0c3f204d9070f1dfe63b1bab11de8298e31f6836;
    5'b10001 : xpb = 1024'h2e15bcd56cead6bb1f72fdc30de61fa3928885a4f4edbb2bb9ba49380fb0dfae36f4e3cf7a634402b3b20c703a7cfefb8ac64196b809bf2619d0b9646a73dc6ed0544bc9053e8eb90d8ee33c95d4dc5abde5ae7e118b3ab0948370d950ee32406fe669293ce94155c61a7201e090d8d3f9cc5219a9561bfba2e7b61e03511ec;
    5'b10010 : xpb = 1024'h9ef0e9ac9d9df5415173f6c505efd3d85556cf6c97db2aea71ef158d71cff2c56c2e49148b6888dfe791c3f326d781924909d87c90713ecaf423bca6f72e8a42073c68349d2412547c9ac24dd48e1d9314d1b4f497817c96aa04bb18c99ecb3db86e660b478c0eb19c7a225027a320f63da277459f3b0504a8edef2f662d220d;
    5'b10011 : xpb = 1024'h8a533236227f084e25eb45d6caa6fe65000f134e0aefd9aaaa65cd31afa22a87f1a4c67355045ef1048a27d866a9226a754d24f992af1157d60b2e596ce3620bad2456fdfa633e7855c293c546e3292f89c01568c16418719534ad29440410c53ad6d35a4a8090c055d2b6a1396d0e35ecce4a8753954b19513de7f86342cbc3;
    5'b10100 : xpb = 1024'h75b57abfa7601b5afa6294e88f5e28f1aac7572f7e04886ae2dc84d5ed74624a771b43d21ea0350221828bbda67ac342a190717694ece3e4b7f2a00be29839d5530c45c757a26a9c2eea653cb93834cbfeae75dceb46b44c80649f39be69564cbd3f40a94d7512cf0f2b4af24b36fb759bfa1dc907ef912df98de0c160587579;
    5'b10101 : xpb = 1024'h6117c3492c412e67ced9e3fa5415537e557f9b10f119372b1b533c7a2b469a0cfc91c130e83c0b133e7aefa2e64c641acdd3bdf3972ab67199da11be584d119ef8f43490b4e196c0081236b42b8d4068739cd651152950276b94914a38ce9bd43fa7adf8506994ddc883df435d00e8b54b25f10abc49d742a1ddd98a5d6e1f2f;
    5'b10110 : xpb = 1024'h4c7a0bd2b1224174a351330c18cc7e0b0037def2642de5eb53c9f41e6918d1cf82083e8fb1d7e1245b735388261e04f2fa170a70996888fe7bc18370ce01e9689edc235a1220c2e3e13a082b9de24c04e88b36c53f0bec0256c4835ab333e15bc2101b47535e16ec81dc73946ecad5f4fa51c44c70a41d574a2dd2535a83c8e5;
    5'b10111 : xpb = 1024'h37dc545c3603548177c8821ddd83a897aaf022d3d74294ab8c40abc2a6eb0992077ebbee7b73b735786bb76d65efa5cb265a56ed9ba65b8b5da8f52343b6c13244c412236f5fef07ba61d9a3103757a15d79973968ee87dd41f4756b2d9926e344788896565298fb3b3507e58094c334a97d978e24fe636bf27dcb1c5799729b;
    5'b11000 : xpb = 1024'h233e9ce5bae4678e4c3fd12fa23ad32455a866b54a57436bc4b76366e4bd41548cf5394d450f8d4695641b52a5c146a3529da36a9de42e183f9066d5b96b98fbeaac00eccc9f1b2b9389ab1a828c633dd267f7ad92d123b82d24677ba7fe6c6ac6e0f5e559471b09f48d9c36925eb07458a96acfd958a9809acdc3e554af1c51;
    5'b11001 : xpb = 1024'hea0e56f3fc57a9b20b7204166f1fdb10060aa96bd6bf22bfd2e1b0b228f7917126bb6ac0eab6357b25c7f37e592e77b7ee0efe7a02200a52177d8882f2070c59093efb629de474f6cb17c91f4e16eda47565821bcb3bf931854598c2263b1f2494963345c3b9d18ade63087a4289db407d53e118db2ef95431dbcae51c4c607;
    5'b11010 : xpb = 1024'haab0734e8694c270c033e72a3c036f8f1c8ef1a905f84163b3818c0513645de19b2ab183a26db7f76eb3226408c2991e0f3e644ac512a37db3fe8998dfa7bd40aacb132e36ae70b8587350ac00123ea7b049b22e731c887eb910dd9756f39a0bfab962ad0ff917b4edfeabb7adc2b11d05daf035925892da31dd307bd7bcd628;
    5'b11011 : xpb = 1024'h9612bbd80b75d57d94ab363c00ba9a1bc747358a790cf023ebf843a9513695a420a12ee26c098e088bab8649489439f63b81b0c7c750760a95e5fb4b555c950a50b301f793ed9cdc319b222372674a44253812a29cff2459a440cfa7d158df937d21cffc12ed99c3a7574008bf8c9e5cb506c37746b2d8eeda2d2944d4d27fde;
    5'b11100 : xpb = 1024'h817504619056e88a6922854dc571c4a871ff796bec219ee4246efb4d8f08cd66a617ac4135a56419a8a3ea2e8865dace67c4fd44c98e489777cd6cfdcb116cd3f69af0c0f12cc9000ac2f39ae4bc55e09a267316c6e1c0348f70c1b84bbe251aff8a3d4b15e21bd260afd459d1568b9c643296b8fb0d1f03827d220dd1e82994;
    5'b11101 : xpb = 1024'h6cd74ceb1537fb973d99d45f8a28ef351cb7bd4d5f364da45ce5b2f1ccdb05292b8e299fff413a2ac59c4e13c8377ba6940849c1cbcc1b2459b4deb040c6449d9c82df8a4e6bf523e3eac5125711617d0f14d38af0c45c0f7aa0b3c8c6236aa281f2aa9a18d69de11a0868aae32078dc135e69faaf6765182acd1ad6cefdd34a;
    5'b11110 : xpb = 1024'h583995749a190ea4121123714ee019c1c770012ed24afc64955c6a960aad3cebb104a6fec8dd103be294b1f908091c7ec04b963ece09edb13b9c5062b67b1c67426ace53abab2147bd129689c9666d19840333ff1aa6f7ea65d0a5d94088b02a045b17e91bcb1fefd360fcfbf4ea661bc28a3d3c63c1ab2cd31d139fcc137d00;
    5'b11111 : xpb = 1024'h439bddfe1efa21b0e68872831397444e72284510455fab24cdd3223a487f74ae367b245d9278e64cff8d15de47dabd56ec8ee2bbd047c03e1d83c2152c2ff430e852bd1d08ea4d6b963a68013bbb78b5f8f19473448993c5510097e9baedf5b186c385381ebfa1fe8cb9914d06b4535b71b6107e181bf1417b6d0c68c92926b6;
    endcase
end

endmodule

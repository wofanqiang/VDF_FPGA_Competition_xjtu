module xpb_5_550
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hab9aa9d9f1185787bb57f5b6c31958667e20f0359e7f881bc9df1aeec01a0f5312ac40520413fb90c1c867729c5879e927e4fe891fa5e8c62a7ca623d5b671e9bc25ed23b2919a63d480f5f1621d78459676f07af4556a8d9665e99e0b688d67295813138c56087c72d44823853854f805300946e6a9c8fd7ad66c35ed2ed027;
    5'b00010 : xpb = 1024'ha6880e5e20427a46abaa739675d8697b8acbdd3a67876fc015e17c87cd31719e2210032b3e017892e4328f9e5552e307ebafd52c1c990140a45a0ce9709a6f2203fca598b59237829667e9402b5f2c5a38e8e75d5c24a80a773f41415ca6783c23a893fd67e3186b5ee8a96812a083c6bb8633ab7d0834caaf3d5d67517b39e3;
    5'b00011 : xpb = 1024'ha17572e24f6c9d059bfcf17628977a909776ca3f308f576461e3de20da48d3e93173c60477eef595069cb7ca0e4d4c26af7aabcf198c19bb1e3773af0b7e6c5a4bd35e0db892d4a1584edc8ef4a0e06edb5ade3fc3f3e587581898e4ade463111df914e74370285a4afd0aaca008b29571dc5e101366a097e3a44e98b5c7a39f;
    5'b00100 : xpb = 1024'h9c62d7667e96bfc48c4f6f55db568ba5a421b743f9973f08ade63fb9e760363440d788ddb1dc72972906dff5c747b54573458272167f32359814da74a662699293aa1682bb9371c01a35cfddbde294837dccd5222bc3230438f1f087ff224de6184995d11efd384937116bf12d70e16428328874a9c50c65180b3fca1a140d5b;
    5'b00101 : xpb = 1024'h97503beaadc0e2837ca1ed358e159cbab0cca448c29f26acf9e8a152f477987f503b4bb6ebc9ef994b71082180421e643710591513724ab011f2413a414666cadb80cef7be940ededc1cc32c87244898203ecc049392608119cb482b506038bb129a16bafa8a48382325cd35bad91032de88b2d9402378324c7230fb7e607717;
    5'b00110 : xpb = 1024'h923da06edceb05426cf46b1540d4adcfbd77914d8ba70e5145eb02ec018efaca5f9f0e9025b76c9b6ddb304d393c8782fadb2fb81065632a8bcfa7ffdc2a64032357876cc194abfd9e03b67b5065fcacc2b0c2e6fb619dfdfaa49fcea19e23900cea97a4d61758270f3a2e7a48413f0194dedd3dd681e3ff80d9222ce2ace0d3;
    5'b00111 : xpb = 1024'h8d2b04f30c1528015d46e8f4f393bee4ca227e5254aef5f591ed64850ea65d156f02d1695fa4e99d90455878f236f0a1bea6065b0d587ba505ad0ec5770e613b6b2e3fe1c495491c5feaa9ca19a7b0c16522b9c96330db7adb7df771f2dc0e65073b188eb1a46815fb4e8fbed5a96dd04b3507a26ce04fccb540135e46f94a8f;
    5'b01000 : xpb = 1024'h881869773b3f4ac04d9966d4a652cff9d6cd6b571db6dd99ddefc61e1bbdbf607e6694429992669fb2af80a4ab3159c08270dcfe0a4b941f7f8a758b11f25e73b304f856c795e63b21d19d18e2e964d60794b0abcb0018f7bc574f154419f93a018b99788d317804e762f10363119c9f018b3207033ebb99e9a7048fab45b44b;
    5'b01001 : xpb = 1024'h8305cdfb6a696d7f3debe4b45911e10ee378585be6bec53e29f227b728d521ab8dca571bd37fe3a1d519a8d0642bc2df463bb3a1073eac99f967dc50acd65babfadbb0cbca968359e3b89067ac2b18eaaa06a78e32cf56749d30a6b89557e40efbdc1a6268be87f3d3775247f079cb6db7e15c6b999d27671e0df5c10f921e07;
    5'b01010 : xpb = 1024'h7df3327f9993903e2e3e62940bd0f223f0234560afc6ace275f4895035ec83f69d2e19f50d6d60a3f783d0fc1d262bfe0a068a440431c5147345431647ba58e442b26940cd972078a59f83b6756cccff4c789e709a9e93f17e09fe5be695cee3f62c9b4c444b97e2bf8bb38c7de1fa3c6e3786d02ffb93345274e6f273de87c3;
    5'b01011 : xpb = 1024'h78e09703c8bdb2fd1e90e073be900338fcce326578ce9486c1f6eae94303e641ac91dcce475adda619edf927d620951ccdd160e70124dd8eed22a9dbe29e561c8a8921b5d097bd97678677053eae8113eeea9553026dd16e5ee355ff37d3b9b8f07d1c361fd8a7d1aba014d10b4a290b248db134c659ff0186dbd823d82af17f;
    5'b01100 : xpb = 1024'h73cdfb87f7e7d5bc0ee35e53714f144e09791f6a41d67c2b0df94c82501b488cbbf59fa781485aa83c5821538f1afe3b919c3789fe17f609670010a17d825354d25fda2ad3985ab6296d6a5407f03528915c8c356a3d0eeb3fbcada28911a48deacd9d1ffb65b7c097b4761598b257d9dae3db995cb86acebb42c9553c775b3b;
    5'b01101 : xpb = 1024'h6ebb600c2711f87aff35dc33240e256316240c6f0ade63cf59fbae1b5d32aad7cb596280bb35d7aa5ec2497f4815675a55670e2cfb0b0e83e0dd77671866508d1a36929fd698f7d4eb545da2d131e93d33ce8317d20c4c6820960545da4f8f62e51e1e09d6f2c7af83c8d75a261a86a8913a05fdf316d69befa9ba86a0c3c4f7;
    5'b01110 : xpb = 1024'h69a8c490563c1b39ef885a12d6cd367822cef973d3e64b73a5fe0fb46a4a0d22dabd2559f52354ac812c71ab010fd0791931e4cff7fe26fe5abade2cb34a4dc5620d4b14d99994f3ad3b50f19a739d51d64079fa39db89e5016f5ce92b8d7a37df6e9ef3b27fd79e6fdd389eb382b57747903062897542692410abb805102eb3;
    5'b01111 : xpb = 1024'h6496291485663df8dfdad7f2898c478d2f79e6789cee3317f200714d77616f6dea20e8332f10d1aea39699d6ba0a3997dcfcbb72f4f13f78d49844f24e2e4afda9e40389dc9a32126f22444063b5516678b270dca1aac761e248b48c7ccb650cd9bf1fdd8e0ce78d5bf199e340eae445fde65ac71fd3ae3658779ce9695c986f;
    5'b10000 : xpb = 1024'h5f838d98b49060b7d02d55d23c4b58a23c24d37d65f61abc3e02d2e68478d1b8f984ab0c68fe4eb0c600c2027304a2b6a0c79215f1e457f34e75abb7e9124835f1babbfedf9acf313109378f2cf7057b1b2467bf097a04dec3220c2fce094fe1d40fa0c76999f77c4805fb27ce531314b43c852bb6321a038cde8e1acda9022b;
    5'b10001 : xpb = 1024'h5a70f21ce3ba8376c07fd3b1ef0a69b748cfc0822efe02608a05347f9190340408e86de5a2ebcbb2e86aea2e2bff0bd5649268b8eed7706dc853127d83f6456e39917473e29b6c4ff2f02addf638b98fbd965ea17149425ba3fb63d31f473ab6ce6021b14527076b341a5c6c5bbb41e36a92af904c9085d0c1457f4c31f56be7;
    5'b10010 : xpb = 1024'h555e56a112e4a635b0d25191a1c97acc557aad86f805ea04d60796189ea7964f184c30bedcd948b50ad51259e4f974f4285d3f5bebca88e8423079431eda42a681682ce8e59c096eb4d71e2cbf7a6da460085583d9187fd884d4bb767085258bc8b0a29b20b4175a202ebdb0e92370b220e8d9f4e2eef19df5ac707d9641d5a3;
    5'b10011 : xpb = 1024'h504bbb25420ec8f4a124cf7154888be162259a8bc10dd1a92209f7b1abbef89a27aff39816c6c5b72d3f3a859df3de12ec2815fee8bda162bc0de008b9be3fdec93ee55de89ca68d76be117b88bc21b9027a4c6640e7bd5565ae1319c1c31060c3012384fc4127490c431ef5768b9f80d73f0459794d5d6b2a1361aefa8e3f5f;
    5'b10100 : xpb = 1024'h4b391fa97138ebb391774d5107479cf66ed087908a15b94d6e0c594ab8d65ae53713b67150b442b94fa962b156ee4731aff2eca1e5b0b9dd35eb46ce54a23d1711159dd2eb9d43ac38a504ca51fdd5cda4ec4348a8b6fad246876abd1300fb35bd51a46ed7ce3737f857803a03f3ce4f8d952ebe0fabc9385e7a52e05edaa91b;
    5'b10101 : xpb = 1024'h4626842da0630e7281c9cb30ba06ae0b7b7b7495531da0f1ba0ebae3c5edbd304677794a8aa1bfbb72138add0fe8b05073bdc344e2a3d257afc8ad93ef863a4f58ec5647ee9de0cafa8bf8191b3f89e2475e3a2b1086384f2760c260643ee60ab7a22558b35b4726e46be17e915bfd1e43eb5922a60a350592e14411c32712d7;
    5'b10110 : xpb = 1024'h4113e8b1cf8d3131721c49106cc5bf208826619a1c25889606111c7cd3051f7b55db3c23c48f3cbd947db308c8e3196f378899e7df96ead229a614598a6a3787a0c30ebcf19e7de9bc72eb67e4813df6e9d0310d785575cc083a1a03b57cd0dfb1f2a6428ee85715d08042c31ec42becfa4183873c68a0d2c748354327737c93;
    5'b10111 : xpb = 1024'h3c014d35feb753f0626ec6f01f84d03594d14e9ee52d703a52137e15e01c81c6653efefcfe7cb9bfb6e7db3481dd828dfb53708adc8a034ca3837b1f254e34bfe899c731f49f1b087e59deb6adc2f20b8c4227efe024b348e91371a706babbb4ac43272c6a756704bc94a407ac2c5abbb097adebd2c70c9ffbaf26748bbfe64f;
    5'b11000 : xpb = 1024'h36eeb1ba2de176af52c144cfd243e14aa17c3ba3ae3557de9e15dfaeed33e41174a2c1d6386a36c1d95203603ad7ebacbf1e472dd97d1bc71d60e1e4c03231f830707fa6f79fb8274040d2057704a6202eb41ed247f3f0c5c9ecc94a57f8a689a693a816460276f3a8a9054c3994898a66edd8506925786d301617a5f00c500b;
    5'b11001 : xpb = 1024'h31dc163e5d0b996e4313c2af8502f25fae2728a8773d3f82ea184147fa4b465c840684af7257b3c3fbbc2b8bf3d254cb82e91dd0d6703441973e48aa5b162f307847381bfaa055460227c55440465a34d12615b4afc32e42aac620eda936915ea0e42900218f86e294bd6690c6fcb8591d4402b4ff83e43a647d08d75458b9c7;
    5'b11010 : xpb = 1024'h2cc97ac28c35bc2d3366408f37c20374bad215ad40452727361aa2e10762a8a7936a4788ac4530c61e2653b7acccbdea46b3f473d3634cbc111baf6ff5fa2c68c01df090fda0f264c40eb8a309880e4973980c9717926bbf8b9f7890fa747c339b34a9e9fd1c96d180d1c7d55464e727d39a2d1995e2500798e3fa08b8a52383;
    5'b11011 : xpb = 1024'h27b6df46bb5fdeec23b8be6eea811489c77d02b2094d0ecb821d047a147a0af2a2ce0a61e632adc840907be365c727090a7ecb16d05665368af9163590de29a107f4a90600a18f8385f5abf1d2c9c25e160a03797f61a93c6c78d0344bb2670895852ad3d8a9a6c06ce62919e1cd15f689f0577e2c40bbd4cd4aeb3a1cf18d3f;
    5'b11100 : xpb = 1024'h22a443caea8a01ab140b3c4e9d40259ed427efb6d254f66fce1f661321916d3db231cd3b20202aca62faa40f1ec19027ce49a1b9cd497db104d67cfb2bc226d94fcb617b03a22ca247dc9f409c0b7672b87bfa5be730e6b94d5227d79cf051dd8fd5abbdb436b6af58fa8a5e6f3544c5404681e2c29f27a201b1dc6b813df6fb;
    5'b11101 : xpb = 1024'h1d91a84f19b4246a045dba2e4fff36b3e0d2dcbb9b5cde141a21c7ac2ea8cf88c19590145a0da7cc8564cc3ad7bbf9469214785cca3c962b7eb3e3c0c6a6241197a219f006a2c9c109c3928f654d2a875aedf13e4f0024362e2b7f7aee2e3cb28a262ca78fc3c69e450eeba2fc9d7393f69cac4758fd936f3618cd9ce58a60b7;
    5'b11110 : xpb = 1024'h187f0cd348de4728f4b0380e02be47c8ed7dc9c06464c5b8662429453bc031d3d0f952ed93fb24cea7cef46690b6626555df4effc72faea5f8914a86618a2149df78d26509a366dfcbaa85de2e8ede9bfd5fe820b6cf61b30f04d71e3f6c27878476ad916b50d68d31234ce78a05a262acf2d6abef5bff3c6a7fbece49d6ca73;
    5'b11111 : xpb = 1024'h136c7157780869e7e502b5edb57d58ddfa28b6c52d6cad5cb2268ade48d7941ee05d15c6cde8a1d0ca391c9249b0cb8419aa25a2c422c720726eb14bfc6e1e82274f8ada0ca403fe8d91792cf7d092b09fd1df031e9e9f2fefde2ec190aa125c7ec72e7b46dde67c1d37ae2c176dd1316349011085ba6b099ee6afffae23342f;
    endcase
end

endmodule

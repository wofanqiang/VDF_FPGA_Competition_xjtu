module compressor_array_6_4_1024
(
    input  [5:0] col_in_0,
    input  [5:0] col_in_1,
    input  [5:0] col_in_2,
    input  [5:0] col_in_3,
    input  [5:0] col_in_4,
    input  [5:0] col_in_5,
    input  [5:0] col_in_6,
    input  [5:0] col_in_7,
    input  [5:0] col_in_8,
    input  [5:0] col_in_9,
    input  [5:0] col_in_10,
    input  [5:0] col_in_11,
    input  [5:0] col_in_12,
    input  [5:0] col_in_13,
    input  [5:0] col_in_14,
    input  [5:0] col_in_15,
    input  [5:0] col_in_16,
    input  [5:0] col_in_17,
    input  [5:0] col_in_18,
    input  [5:0] col_in_19,
    input  [5:0] col_in_20,
    input  [5:0] col_in_21,
    input  [5:0] col_in_22,
    input  [5:0] col_in_23,
    input  [5:0] col_in_24,
    input  [5:0] col_in_25,
    input  [5:0] col_in_26,
    input  [5:0] col_in_27,
    input  [5:0] col_in_28,
    input  [5:0] col_in_29,
    input  [5:0] col_in_30,
    input  [5:0] col_in_31,
    input  [5:0] col_in_32,
    input  [5:0] col_in_33,
    input  [5:0] col_in_34,
    input  [5:0] col_in_35,
    input  [5:0] col_in_36,
    input  [5:0] col_in_37,
    input  [5:0] col_in_38,
    input  [5:0] col_in_39,
    input  [5:0] col_in_40,
    input  [5:0] col_in_41,
    input  [5:0] col_in_42,
    input  [5:0] col_in_43,
    input  [5:0] col_in_44,
    input  [5:0] col_in_45,
    input  [5:0] col_in_46,
    input  [5:0] col_in_47,
    input  [5:0] col_in_48,
    input  [5:0] col_in_49,
    input  [5:0] col_in_50,
    input  [5:0] col_in_51,
    input  [5:0] col_in_52,
    input  [5:0] col_in_53,
    input  [5:0] col_in_54,
    input  [5:0] col_in_55,
    input  [5:0] col_in_56,
    input  [5:0] col_in_57,
    input  [5:0] col_in_58,
    input  [5:0] col_in_59,
    input  [5:0] col_in_60,
    input  [5:0] col_in_61,
    input  [5:0] col_in_62,
    input  [5:0] col_in_63,
    input  [5:0] col_in_64,
    input  [5:0] col_in_65,
    input  [5:0] col_in_66,
    input  [5:0] col_in_67,
    input  [5:0] col_in_68,
    input  [5:0] col_in_69,
    input  [5:0] col_in_70,
    input  [5:0] col_in_71,
    input  [5:0] col_in_72,
    input  [5:0] col_in_73,
    input  [5:0] col_in_74,
    input  [5:0] col_in_75,
    input  [5:0] col_in_76,
    input  [5:0] col_in_77,
    input  [5:0] col_in_78,
    input  [5:0] col_in_79,
    input  [5:0] col_in_80,
    input  [5:0] col_in_81,
    input  [5:0] col_in_82,
    input  [5:0] col_in_83,
    input  [5:0] col_in_84,
    input  [5:0] col_in_85,
    input  [5:0] col_in_86,
    input  [5:0] col_in_87,
    input  [5:0] col_in_88,
    input  [5:0] col_in_89,
    input  [5:0] col_in_90,
    input  [5:0] col_in_91,
    input  [5:0] col_in_92,
    input  [5:0] col_in_93,
    input  [5:0] col_in_94,
    input  [5:0] col_in_95,
    input  [5:0] col_in_96,
    input  [5:0] col_in_97,
    input  [5:0] col_in_98,
    input  [5:0] col_in_99,
    input  [5:0] col_in_100,
    input  [5:0] col_in_101,
    input  [5:0] col_in_102,
    input  [5:0] col_in_103,
    input  [5:0] col_in_104,
    input  [5:0] col_in_105,
    input  [5:0] col_in_106,
    input  [5:0] col_in_107,
    input  [5:0] col_in_108,
    input  [5:0] col_in_109,
    input  [5:0] col_in_110,
    input  [5:0] col_in_111,
    input  [5:0] col_in_112,
    input  [5:0] col_in_113,
    input  [5:0] col_in_114,
    input  [5:0] col_in_115,
    input  [5:0] col_in_116,
    input  [5:0] col_in_117,
    input  [5:0] col_in_118,
    input  [5:0] col_in_119,
    input  [5:0] col_in_120,
    input  [5:0] col_in_121,
    input  [5:0] col_in_122,
    input  [5:0] col_in_123,
    input  [5:0] col_in_124,
    input  [5:0] col_in_125,
    input  [5:0] col_in_126,
    input  [5:0] col_in_127,
    input  [5:0] col_in_128,
    input  [5:0] col_in_129,
    input  [5:0] col_in_130,
    input  [5:0] col_in_131,
    input  [5:0] col_in_132,
    input  [5:0] col_in_133,
    input  [5:0] col_in_134,
    input  [5:0] col_in_135,
    input  [5:0] col_in_136,
    input  [5:0] col_in_137,
    input  [5:0] col_in_138,
    input  [5:0] col_in_139,
    input  [5:0] col_in_140,
    input  [5:0] col_in_141,
    input  [5:0] col_in_142,
    input  [5:0] col_in_143,
    input  [5:0] col_in_144,
    input  [5:0] col_in_145,
    input  [5:0] col_in_146,
    input  [5:0] col_in_147,
    input  [5:0] col_in_148,
    input  [5:0] col_in_149,
    input  [5:0] col_in_150,
    input  [5:0] col_in_151,
    input  [5:0] col_in_152,
    input  [5:0] col_in_153,
    input  [5:0] col_in_154,
    input  [5:0] col_in_155,
    input  [5:0] col_in_156,
    input  [5:0] col_in_157,
    input  [5:0] col_in_158,
    input  [5:0] col_in_159,
    input  [5:0] col_in_160,
    input  [5:0] col_in_161,
    input  [5:0] col_in_162,
    input  [5:0] col_in_163,
    input  [5:0] col_in_164,
    input  [5:0] col_in_165,
    input  [5:0] col_in_166,
    input  [5:0] col_in_167,
    input  [5:0] col_in_168,
    input  [5:0] col_in_169,
    input  [5:0] col_in_170,
    input  [5:0] col_in_171,
    input  [5:0] col_in_172,
    input  [5:0] col_in_173,
    input  [5:0] col_in_174,
    input  [5:0] col_in_175,
    input  [5:0] col_in_176,
    input  [5:0] col_in_177,
    input  [5:0] col_in_178,
    input  [5:0] col_in_179,
    input  [5:0] col_in_180,
    input  [5:0] col_in_181,
    input  [5:0] col_in_182,
    input  [5:0] col_in_183,
    input  [5:0] col_in_184,
    input  [5:0] col_in_185,
    input  [5:0] col_in_186,
    input  [5:0] col_in_187,
    input  [5:0] col_in_188,
    input  [5:0] col_in_189,
    input  [5:0] col_in_190,
    input  [5:0] col_in_191,
    input  [5:0] col_in_192,
    input  [5:0] col_in_193,
    input  [5:0] col_in_194,
    input  [5:0] col_in_195,
    input  [5:0] col_in_196,
    input  [5:0] col_in_197,
    input  [5:0] col_in_198,
    input  [5:0] col_in_199,
    input  [5:0] col_in_200,
    input  [5:0] col_in_201,
    input  [5:0] col_in_202,
    input  [5:0] col_in_203,
    input  [5:0] col_in_204,
    input  [5:0] col_in_205,
    input  [5:0] col_in_206,
    input  [5:0] col_in_207,
    input  [5:0] col_in_208,
    input  [5:0] col_in_209,
    input  [5:0] col_in_210,
    input  [5:0] col_in_211,
    input  [5:0] col_in_212,
    input  [5:0] col_in_213,
    input  [5:0] col_in_214,
    input  [5:0] col_in_215,
    input  [5:0] col_in_216,
    input  [5:0] col_in_217,
    input  [5:0] col_in_218,
    input  [5:0] col_in_219,
    input  [5:0] col_in_220,
    input  [5:0] col_in_221,
    input  [5:0] col_in_222,
    input  [5:0] col_in_223,
    input  [5:0] col_in_224,
    input  [5:0] col_in_225,
    input  [5:0] col_in_226,
    input  [5:0] col_in_227,
    input  [5:0] col_in_228,
    input  [5:0] col_in_229,
    input  [5:0] col_in_230,
    input  [5:0] col_in_231,
    input  [5:0] col_in_232,
    input  [5:0] col_in_233,
    input  [5:0] col_in_234,
    input  [5:0] col_in_235,
    input  [5:0] col_in_236,
    input  [5:0] col_in_237,
    input  [5:0] col_in_238,
    input  [5:0] col_in_239,
    input  [5:0] col_in_240,
    input  [5:0] col_in_241,
    input  [5:0] col_in_242,
    input  [5:0] col_in_243,
    input  [5:0] col_in_244,
    input  [5:0] col_in_245,
    input  [5:0] col_in_246,
    input  [5:0] col_in_247,
    input  [5:0] col_in_248,
    input  [5:0] col_in_249,
    input  [5:0] col_in_250,
    input  [5:0] col_in_251,
    input  [5:0] col_in_252,
    input  [5:0] col_in_253,
    input  [5:0] col_in_254,
    input  [5:0] col_in_255,
    input  [5:0] col_in_256,
    input  [5:0] col_in_257,
    input  [5:0] col_in_258,
    input  [5:0] col_in_259,
    input  [5:0] col_in_260,
    input  [5:0] col_in_261,
    input  [5:0] col_in_262,
    input  [5:0] col_in_263,
    input  [5:0] col_in_264,
    input  [5:0] col_in_265,
    input  [5:0] col_in_266,
    input  [5:0] col_in_267,
    input  [5:0] col_in_268,
    input  [5:0] col_in_269,
    input  [5:0] col_in_270,
    input  [5:0] col_in_271,
    input  [5:0] col_in_272,
    input  [5:0] col_in_273,
    input  [5:0] col_in_274,
    input  [5:0] col_in_275,
    input  [5:0] col_in_276,
    input  [5:0] col_in_277,
    input  [5:0] col_in_278,
    input  [5:0] col_in_279,
    input  [5:0] col_in_280,
    input  [5:0] col_in_281,
    input  [5:0] col_in_282,
    input  [5:0] col_in_283,
    input  [5:0] col_in_284,
    input  [5:0] col_in_285,
    input  [5:0] col_in_286,
    input  [5:0] col_in_287,
    input  [5:0] col_in_288,
    input  [5:0] col_in_289,
    input  [5:0] col_in_290,
    input  [5:0] col_in_291,
    input  [5:0] col_in_292,
    input  [5:0] col_in_293,
    input  [5:0] col_in_294,
    input  [5:0] col_in_295,
    input  [5:0] col_in_296,
    input  [5:0] col_in_297,
    input  [5:0] col_in_298,
    input  [5:0] col_in_299,
    input  [5:0] col_in_300,
    input  [5:0] col_in_301,
    input  [5:0] col_in_302,
    input  [5:0] col_in_303,
    input  [5:0] col_in_304,
    input  [5:0] col_in_305,
    input  [5:0] col_in_306,
    input  [5:0] col_in_307,
    input  [5:0] col_in_308,
    input  [5:0] col_in_309,
    input  [5:0] col_in_310,
    input  [5:0] col_in_311,
    input  [5:0] col_in_312,
    input  [5:0] col_in_313,
    input  [5:0] col_in_314,
    input  [5:0] col_in_315,
    input  [5:0] col_in_316,
    input  [5:0] col_in_317,
    input  [5:0] col_in_318,
    input  [5:0] col_in_319,
    input  [5:0] col_in_320,
    input  [5:0] col_in_321,
    input  [5:0] col_in_322,
    input  [5:0] col_in_323,
    input  [5:0] col_in_324,
    input  [5:0] col_in_325,
    input  [5:0] col_in_326,
    input  [5:0] col_in_327,
    input  [5:0] col_in_328,
    input  [5:0] col_in_329,
    input  [5:0] col_in_330,
    input  [5:0] col_in_331,
    input  [5:0] col_in_332,
    input  [5:0] col_in_333,
    input  [5:0] col_in_334,
    input  [5:0] col_in_335,
    input  [5:0] col_in_336,
    input  [5:0] col_in_337,
    input  [5:0] col_in_338,
    input  [5:0] col_in_339,
    input  [5:0] col_in_340,
    input  [5:0] col_in_341,
    input  [5:0] col_in_342,
    input  [5:0] col_in_343,
    input  [5:0] col_in_344,
    input  [5:0] col_in_345,
    input  [5:0] col_in_346,
    input  [5:0] col_in_347,
    input  [5:0] col_in_348,
    input  [5:0] col_in_349,
    input  [5:0] col_in_350,
    input  [5:0] col_in_351,
    input  [5:0] col_in_352,
    input  [5:0] col_in_353,
    input  [5:0] col_in_354,
    input  [5:0] col_in_355,
    input  [5:0] col_in_356,
    input  [5:0] col_in_357,
    input  [5:0] col_in_358,
    input  [5:0] col_in_359,
    input  [5:0] col_in_360,
    input  [5:0] col_in_361,
    input  [5:0] col_in_362,
    input  [5:0] col_in_363,
    input  [5:0] col_in_364,
    input  [5:0] col_in_365,
    input  [5:0] col_in_366,
    input  [5:0] col_in_367,
    input  [5:0] col_in_368,
    input  [5:0] col_in_369,
    input  [5:0] col_in_370,
    input  [5:0] col_in_371,
    input  [5:0] col_in_372,
    input  [5:0] col_in_373,
    input  [5:0] col_in_374,
    input  [5:0] col_in_375,
    input  [5:0] col_in_376,
    input  [5:0] col_in_377,
    input  [5:0] col_in_378,
    input  [5:0] col_in_379,
    input  [5:0] col_in_380,
    input  [5:0] col_in_381,
    input  [5:0] col_in_382,
    input  [5:0] col_in_383,
    input  [5:0] col_in_384,
    input  [5:0] col_in_385,
    input  [5:0] col_in_386,
    input  [5:0] col_in_387,
    input  [5:0] col_in_388,
    input  [5:0] col_in_389,
    input  [5:0] col_in_390,
    input  [5:0] col_in_391,
    input  [5:0] col_in_392,
    input  [5:0] col_in_393,
    input  [5:0] col_in_394,
    input  [5:0] col_in_395,
    input  [5:0] col_in_396,
    input  [5:0] col_in_397,
    input  [5:0] col_in_398,
    input  [5:0] col_in_399,
    input  [5:0] col_in_400,
    input  [5:0] col_in_401,
    input  [5:0] col_in_402,
    input  [5:0] col_in_403,
    input  [5:0] col_in_404,
    input  [5:0] col_in_405,
    input  [5:0] col_in_406,
    input  [5:0] col_in_407,
    input  [5:0] col_in_408,
    input  [5:0] col_in_409,
    input  [5:0] col_in_410,
    input  [5:0] col_in_411,
    input  [5:0] col_in_412,
    input  [5:0] col_in_413,
    input  [5:0] col_in_414,
    input  [5:0] col_in_415,
    input  [5:0] col_in_416,
    input  [5:0] col_in_417,
    input  [5:0] col_in_418,
    input  [5:0] col_in_419,
    input  [5:0] col_in_420,
    input  [5:0] col_in_421,
    input  [5:0] col_in_422,
    input  [5:0] col_in_423,
    input  [5:0] col_in_424,
    input  [5:0] col_in_425,
    input  [5:0] col_in_426,
    input  [5:0] col_in_427,
    input  [5:0] col_in_428,
    input  [5:0] col_in_429,
    input  [5:0] col_in_430,
    input  [5:0] col_in_431,
    input  [5:0] col_in_432,
    input  [5:0] col_in_433,
    input  [5:0] col_in_434,
    input  [5:0] col_in_435,
    input  [5:0] col_in_436,
    input  [5:0] col_in_437,
    input  [5:0] col_in_438,
    input  [5:0] col_in_439,
    input  [5:0] col_in_440,
    input  [5:0] col_in_441,
    input  [5:0] col_in_442,
    input  [5:0] col_in_443,
    input  [5:0] col_in_444,
    input  [5:0] col_in_445,
    input  [5:0] col_in_446,
    input  [5:0] col_in_447,
    input  [5:0] col_in_448,
    input  [5:0] col_in_449,
    input  [5:0] col_in_450,
    input  [5:0] col_in_451,
    input  [5:0] col_in_452,
    input  [5:0] col_in_453,
    input  [5:0] col_in_454,
    input  [5:0] col_in_455,
    input  [5:0] col_in_456,
    input  [5:0] col_in_457,
    input  [5:0] col_in_458,
    input  [5:0] col_in_459,
    input  [5:0] col_in_460,
    input  [5:0] col_in_461,
    input  [5:0] col_in_462,
    input  [5:0] col_in_463,
    input  [5:0] col_in_464,
    input  [5:0] col_in_465,
    input  [5:0] col_in_466,
    input  [5:0] col_in_467,
    input  [5:0] col_in_468,
    input  [5:0] col_in_469,
    input  [5:0] col_in_470,
    input  [5:0] col_in_471,
    input  [5:0] col_in_472,
    input  [5:0] col_in_473,
    input  [5:0] col_in_474,
    input  [5:0] col_in_475,
    input  [5:0] col_in_476,
    input  [5:0] col_in_477,
    input  [5:0] col_in_478,
    input  [5:0] col_in_479,
    input  [5:0] col_in_480,
    input  [5:0] col_in_481,
    input  [5:0] col_in_482,
    input  [5:0] col_in_483,
    input  [5:0] col_in_484,
    input  [5:0] col_in_485,
    input  [5:0] col_in_486,
    input  [5:0] col_in_487,
    input  [5:0] col_in_488,
    input  [5:0] col_in_489,
    input  [5:0] col_in_490,
    input  [5:0] col_in_491,
    input  [5:0] col_in_492,
    input  [5:0] col_in_493,
    input  [5:0] col_in_494,
    input  [5:0] col_in_495,
    input  [5:0] col_in_496,
    input  [5:0] col_in_497,
    input  [5:0] col_in_498,
    input  [5:0] col_in_499,
    input  [5:0] col_in_500,
    input  [5:0] col_in_501,
    input  [5:0] col_in_502,
    input  [5:0] col_in_503,
    input  [5:0] col_in_504,
    input  [5:0] col_in_505,
    input  [5:0] col_in_506,
    input  [5:0] col_in_507,
    input  [5:0] col_in_508,
    input  [5:0] col_in_509,
    input  [5:0] col_in_510,
    input  [5:0] col_in_511,
    input  [5:0] col_in_512,
    input  [5:0] col_in_513,
    input  [5:0] col_in_514,
    input  [5:0] col_in_515,
    input  [5:0] col_in_516,
    input  [5:0] col_in_517,
    input  [5:0] col_in_518,
    input  [5:0] col_in_519,
    input  [5:0] col_in_520,
    input  [5:0] col_in_521,
    input  [5:0] col_in_522,
    input  [5:0] col_in_523,
    input  [5:0] col_in_524,
    input  [5:0] col_in_525,
    input  [5:0] col_in_526,
    input  [5:0] col_in_527,
    input  [5:0] col_in_528,
    input  [5:0] col_in_529,
    input  [5:0] col_in_530,
    input  [5:0] col_in_531,
    input  [5:0] col_in_532,
    input  [5:0] col_in_533,
    input  [5:0] col_in_534,
    input  [5:0] col_in_535,
    input  [5:0] col_in_536,
    input  [5:0] col_in_537,
    input  [5:0] col_in_538,
    input  [5:0] col_in_539,
    input  [5:0] col_in_540,
    input  [5:0] col_in_541,
    input  [5:0] col_in_542,
    input  [5:0] col_in_543,
    input  [5:0] col_in_544,
    input  [5:0] col_in_545,
    input  [5:0] col_in_546,
    input  [5:0] col_in_547,
    input  [5:0] col_in_548,
    input  [5:0] col_in_549,
    input  [5:0] col_in_550,
    input  [5:0] col_in_551,
    input  [5:0] col_in_552,
    input  [5:0] col_in_553,
    input  [5:0] col_in_554,
    input  [5:0] col_in_555,
    input  [5:0] col_in_556,
    input  [5:0] col_in_557,
    input  [5:0] col_in_558,
    input  [5:0] col_in_559,
    input  [5:0] col_in_560,
    input  [5:0] col_in_561,
    input  [5:0] col_in_562,
    input  [5:0] col_in_563,
    input  [5:0] col_in_564,
    input  [5:0] col_in_565,
    input  [5:0] col_in_566,
    input  [5:0] col_in_567,
    input  [5:0] col_in_568,
    input  [5:0] col_in_569,
    input  [5:0] col_in_570,
    input  [5:0] col_in_571,
    input  [5:0] col_in_572,
    input  [5:0] col_in_573,
    input  [5:0] col_in_574,
    input  [5:0] col_in_575,
    input  [5:0] col_in_576,
    input  [5:0] col_in_577,
    input  [5:0] col_in_578,
    input  [5:0] col_in_579,
    input  [5:0] col_in_580,
    input  [5:0] col_in_581,
    input  [5:0] col_in_582,
    input  [5:0] col_in_583,
    input  [5:0] col_in_584,
    input  [5:0] col_in_585,
    input  [5:0] col_in_586,
    input  [5:0] col_in_587,
    input  [5:0] col_in_588,
    input  [5:0] col_in_589,
    input  [5:0] col_in_590,
    input  [5:0] col_in_591,
    input  [5:0] col_in_592,
    input  [5:0] col_in_593,
    input  [5:0] col_in_594,
    input  [5:0] col_in_595,
    input  [5:0] col_in_596,
    input  [5:0] col_in_597,
    input  [5:0] col_in_598,
    input  [5:0] col_in_599,
    input  [5:0] col_in_600,
    input  [5:0] col_in_601,
    input  [5:0] col_in_602,
    input  [5:0] col_in_603,
    input  [5:0] col_in_604,
    input  [5:0] col_in_605,
    input  [5:0] col_in_606,
    input  [5:0] col_in_607,
    input  [5:0] col_in_608,
    input  [5:0] col_in_609,
    input  [5:0] col_in_610,
    input  [5:0] col_in_611,
    input  [5:0] col_in_612,
    input  [5:0] col_in_613,
    input  [5:0] col_in_614,
    input  [5:0] col_in_615,
    input  [5:0] col_in_616,
    input  [5:0] col_in_617,
    input  [5:0] col_in_618,
    input  [5:0] col_in_619,
    input  [5:0] col_in_620,
    input  [5:0] col_in_621,
    input  [5:0] col_in_622,
    input  [5:0] col_in_623,
    input  [5:0] col_in_624,
    input  [5:0] col_in_625,
    input  [5:0] col_in_626,
    input  [5:0] col_in_627,
    input  [5:0] col_in_628,
    input  [5:0] col_in_629,
    input  [5:0] col_in_630,
    input  [5:0] col_in_631,
    input  [5:0] col_in_632,
    input  [5:0] col_in_633,
    input  [5:0] col_in_634,
    input  [5:0] col_in_635,
    input  [5:0] col_in_636,
    input  [5:0] col_in_637,
    input  [5:0] col_in_638,
    input  [5:0] col_in_639,
    input  [5:0] col_in_640,
    input  [5:0] col_in_641,
    input  [5:0] col_in_642,
    input  [5:0] col_in_643,
    input  [5:0] col_in_644,
    input  [5:0] col_in_645,
    input  [5:0] col_in_646,
    input  [5:0] col_in_647,
    input  [5:0] col_in_648,
    input  [5:0] col_in_649,
    input  [5:0] col_in_650,
    input  [5:0] col_in_651,
    input  [5:0] col_in_652,
    input  [5:0] col_in_653,
    input  [5:0] col_in_654,
    input  [5:0] col_in_655,
    input  [5:0] col_in_656,
    input  [5:0] col_in_657,
    input  [5:0] col_in_658,
    input  [5:0] col_in_659,
    input  [5:0] col_in_660,
    input  [5:0] col_in_661,
    input  [5:0] col_in_662,
    input  [5:0] col_in_663,
    input  [5:0] col_in_664,
    input  [5:0] col_in_665,
    input  [5:0] col_in_666,
    input  [5:0] col_in_667,
    input  [5:0] col_in_668,
    input  [5:0] col_in_669,
    input  [5:0] col_in_670,
    input  [5:0] col_in_671,
    input  [5:0] col_in_672,
    input  [5:0] col_in_673,
    input  [5:0] col_in_674,
    input  [5:0] col_in_675,
    input  [5:0] col_in_676,
    input  [5:0] col_in_677,
    input  [5:0] col_in_678,
    input  [5:0] col_in_679,
    input  [5:0] col_in_680,
    input  [5:0] col_in_681,
    input  [5:0] col_in_682,
    input  [5:0] col_in_683,
    input  [5:0] col_in_684,
    input  [5:0] col_in_685,
    input  [5:0] col_in_686,
    input  [5:0] col_in_687,
    input  [5:0] col_in_688,
    input  [5:0] col_in_689,
    input  [5:0] col_in_690,
    input  [5:0] col_in_691,
    input  [5:0] col_in_692,
    input  [5:0] col_in_693,
    input  [5:0] col_in_694,
    input  [5:0] col_in_695,
    input  [5:0] col_in_696,
    input  [5:0] col_in_697,
    input  [5:0] col_in_698,
    input  [5:0] col_in_699,
    input  [5:0] col_in_700,
    input  [5:0] col_in_701,
    input  [5:0] col_in_702,
    input  [5:0] col_in_703,
    input  [5:0] col_in_704,
    input  [5:0] col_in_705,
    input  [5:0] col_in_706,
    input  [5:0] col_in_707,
    input  [5:0] col_in_708,
    input  [5:0] col_in_709,
    input  [5:0] col_in_710,
    input  [5:0] col_in_711,
    input  [5:0] col_in_712,
    input  [5:0] col_in_713,
    input  [5:0] col_in_714,
    input  [5:0] col_in_715,
    input  [5:0] col_in_716,
    input  [5:0] col_in_717,
    input  [5:0] col_in_718,
    input  [5:0] col_in_719,
    input  [5:0] col_in_720,
    input  [5:0] col_in_721,
    input  [5:0] col_in_722,
    input  [5:0] col_in_723,
    input  [5:0] col_in_724,
    input  [5:0] col_in_725,
    input  [5:0] col_in_726,
    input  [5:0] col_in_727,
    input  [5:0] col_in_728,
    input  [5:0] col_in_729,
    input  [5:0] col_in_730,
    input  [5:0] col_in_731,
    input  [5:0] col_in_732,
    input  [5:0] col_in_733,
    input  [5:0] col_in_734,
    input  [5:0] col_in_735,
    input  [5:0] col_in_736,
    input  [5:0] col_in_737,
    input  [5:0] col_in_738,
    input  [5:0] col_in_739,
    input  [5:0] col_in_740,
    input  [5:0] col_in_741,
    input  [5:0] col_in_742,
    input  [5:0] col_in_743,
    input  [5:0] col_in_744,
    input  [5:0] col_in_745,
    input  [5:0] col_in_746,
    input  [5:0] col_in_747,
    input  [5:0] col_in_748,
    input  [5:0] col_in_749,
    input  [5:0] col_in_750,
    input  [5:0] col_in_751,
    input  [5:0] col_in_752,
    input  [5:0] col_in_753,
    input  [5:0] col_in_754,
    input  [5:0] col_in_755,
    input  [5:0] col_in_756,
    input  [5:0] col_in_757,
    input  [5:0] col_in_758,
    input  [5:0] col_in_759,
    input  [5:0] col_in_760,
    input  [5:0] col_in_761,
    input  [5:0] col_in_762,
    input  [5:0] col_in_763,
    input  [5:0] col_in_764,
    input  [5:0] col_in_765,
    input  [5:0] col_in_766,
    input  [5:0] col_in_767,
    input  [5:0] col_in_768,
    input  [5:0] col_in_769,
    input  [5:0] col_in_770,
    input  [5:0] col_in_771,
    input  [5:0] col_in_772,
    input  [5:0] col_in_773,
    input  [5:0] col_in_774,
    input  [5:0] col_in_775,
    input  [5:0] col_in_776,
    input  [5:0] col_in_777,
    input  [5:0] col_in_778,
    input  [5:0] col_in_779,
    input  [5:0] col_in_780,
    input  [5:0] col_in_781,
    input  [5:0] col_in_782,
    input  [5:0] col_in_783,
    input  [5:0] col_in_784,
    input  [5:0] col_in_785,
    input  [5:0] col_in_786,
    input  [5:0] col_in_787,
    input  [5:0] col_in_788,
    input  [5:0] col_in_789,
    input  [5:0] col_in_790,
    input  [5:0] col_in_791,
    input  [5:0] col_in_792,
    input  [5:0] col_in_793,
    input  [5:0] col_in_794,
    input  [5:0] col_in_795,
    input  [5:0] col_in_796,
    input  [5:0] col_in_797,
    input  [5:0] col_in_798,
    input  [5:0] col_in_799,
    input  [5:0] col_in_800,
    input  [5:0] col_in_801,
    input  [5:0] col_in_802,
    input  [5:0] col_in_803,
    input  [5:0] col_in_804,
    input  [5:0] col_in_805,
    input  [5:0] col_in_806,
    input  [5:0] col_in_807,
    input  [5:0] col_in_808,
    input  [5:0] col_in_809,
    input  [5:0] col_in_810,
    input  [5:0] col_in_811,
    input  [5:0] col_in_812,
    input  [5:0] col_in_813,
    input  [5:0] col_in_814,
    input  [5:0] col_in_815,
    input  [5:0] col_in_816,
    input  [5:0] col_in_817,
    input  [5:0] col_in_818,
    input  [5:0] col_in_819,
    input  [5:0] col_in_820,
    input  [5:0] col_in_821,
    input  [5:0] col_in_822,
    input  [5:0] col_in_823,
    input  [5:0] col_in_824,
    input  [5:0] col_in_825,
    input  [5:0] col_in_826,
    input  [5:0] col_in_827,
    input  [5:0] col_in_828,
    input  [5:0] col_in_829,
    input  [5:0] col_in_830,
    input  [5:0] col_in_831,
    input  [5:0] col_in_832,
    input  [5:0] col_in_833,
    input  [5:0] col_in_834,
    input  [5:0] col_in_835,
    input  [5:0] col_in_836,
    input  [5:0] col_in_837,
    input  [5:0] col_in_838,
    input  [5:0] col_in_839,
    input  [5:0] col_in_840,
    input  [5:0] col_in_841,
    input  [5:0] col_in_842,
    input  [5:0] col_in_843,
    input  [5:0] col_in_844,
    input  [5:0] col_in_845,
    input  [5:0] col_in_846,
    input  [5:0] col_in_847,
    input  [5:0] col_in_848,
    input  [5:0] col_in_849,
    input  [5:0] col_in_850,
    input  [5:0] col_in_851,
    input  [5:0] col_in_852,
    input  [5:0] col_in_853,
    input  [5:0] col_in_854,
    input  [5:0] col_in_855,
    input  [5:0] col_in_856,
    input  [5:0] col_in_857,
    input  [5:0] col_in_858,
    input  [5:0] col_in_859,
    input  [5:0] col_in_860,
    input  [5:0] col_in_861,
    input  [5:0] col_in_862,
    input  [5:0] col_in_863,
    input  [5:0] col_in_864,
    input  [5:0] col_in_865,
    input  [5:0] col_in_866,
    input  [5:0] col_in_867,
    input  [5:0] col_in_868,
    input  [5:0] col_in_869,
    input  [5:0] col_in_870,
    input  [5:0] col_in_871,
    input  [5:0] col_in_872,
    input  [5:0] col_in_873,
    input  [5:0] col_in_874,
    input  [5:0] col_in_875,
    input  [5:0] col_in_876,
    input  [5:0] col_in_877,
    input  [5:0] col_in_878,
    input  [5:0] col_in_879,
    input  [5:0] col_in_880,
    input  [5:0] col_in_881,
    input  [5:0] col_in_882,
    input  [5:0] col_in_883,
    input  [5:0] col_in_884,
    input  [5:0] col_in_885,
    input  [5:0] col_in_886,
    input  [5:0] col_in_887,
    input  [5:0] col_in_888,
    input  [5:0] col_in_889,
    input  [5:0] col_in_890,
    input  [5:0] col_in_891,
    input  [5:0] col_in_892,
    input  [5:0] col_in_893,
    input  [5:0] col_in_894,
    input  [5:0] col_in_895,
    input  [5:0] col_in_896,
    input  [5:0] col_in_897,
    input  [5:0] col_in_898,
    input  [5:0] col_in_899,
    input  [5:0] col_in_900,
    input  [5:0] col_in_901,
    input  [5:0] col_in_902,
    input  [5:0] col_in_903,
    input  [5:0] col_in_904,
    input  [5:0] col_in_905,
    input  [5:0] col_in_906,
    input  [5:0] col_in_907,
    input  [5:0] col_in_908,
    input  [5:0] col_in_909,
    input  [5:0] col_in_910,
    input  [5:0] col_in_911,
    input  [5:0] col_in_912,
    input  [5:0] col_in_913,
    input  [5:0] col_in_914,
    input  [5:0] col_in_915,
    input  [5:0] col_in_916,
    input  [5:0] col_in_917,
    input  [5:0] col_in_918,
    input  [5:0] col_in_919,
    input  [5:0] col_in_920,
    input  [5:0] col_in_921,
    input  [5:0] col_in_922,
    input  [5:0] col_in_923,
    input  [5:0] col_in_924,
    input  [5:0] col_in_925,
    input  [5:0] col_in_926,
    input  [5:0] col_in_927,
    input  [5:0] col_in_928,
    input  [5:0] col_in_929,
    input  [5:0] col_in_930,
    input  [5:0] col_in_931,
    input  [5:0] col_in_932,
    input  [5:0] col_in_933,
    input  [5:0] col_in_934,
    input  [5:0] col_in_935,
    input  [5:0] col_in_936,
    input  [5:0] col_in_937,
    input  [5:0] col_in_938,
    input  [5:0] col_in_939,
    input  [5:0] col_in_940,
    input  [5:0] col_in_941,
    input  [5:0] col_in_942,
    input  [5:0] col_in_943,
    input  [5:0] col_in_944,
    input  [5:0] col_in_945,
    input  [5:0] col_in_946,
    input  [5:0] col_in_947,
    input  [5:0] col_in_948,
    input  [5:0] col_in_949,
    input  [5:0] col_in_950,
    input  [5:0] col_in_951,
    input  [5:0] col_in_952,
    input  [5:0] col_in_953,
    input  [5:0] col_in_954,
    input  [5:0] col_in_955,
    input  [5:0] col_in_956,
    input  [5:0] col_in_957,
    input  [5:0] col_in_958,
    input  [5:0] col_in_959,
    input  [5:0] col_in_960,
    input  [5:0] col_in_961,
    input  [5:0] col_in_962,
    input  [5:0] col_in_963,
    input  [5:0] col_in_964,
    input  [5:0] col_in_965,
    input  [5:0] col_in_966,
    input  [5:0] col_in_967,
    input  [5:0] col_in_968,
    input  [5:0] col_in_969,
    input  [5:0] col_in_970,
    input  [5:0] col_in_971,
    input  [5:0] col_in_972,
    input  [5:0] col_in_973,
    input  [5:0] col_in_974,
    input  [5:0] col_in_975,
    input  [5:0] col_in_976,
    input  [5:0] col_in_977,
    input  [5:0] col_in_978,
    input  [5:0] col_in_979,
    input  [5:0] col_in_980,
    input  [5:0] col_in_981,
    input  [5:0] col_in_982,
    input  [5:0] col_in_983,
    input  [5:0] col_in_984,
    input  [5:0] col_in_985,
    input  [5:0] col_in_986,
    input  [5:0] col_in_987,
    input  [5:0] col_in_988,
    input  [5:0] col_in_989,
    input  [5:0] col_in_990,
    input  [5:0] col_in_991,
    input  [5:0] col_in_992,
    input  [5:0] col_in_993,
    input  [5:0] col_in_994,
    input  [5:0] col_in_995,
    input  [5:0] col_in_996,
    input  [5:0] col_in_997,
    input  [5:0] col_in_998,
    input  [5:0] col_in_999,
    input  [5:0] col_in_1000,
    input  [5:0] col_in_1001,
    input  [5:0] col_in_1002,
    input  [5:0] col_in_1003,
    input  [5:0] col_in_1004,
    input  [5:0] col_in_1005,
    input  [5:0] col_in_1006,
    input  [5:0] col_in_1007,
    input  [5:0] col_in_1008,
    input  [5:0] col_in_1009,
    input  [5:0] col_in_1010,
    input  [5:0] col_in_1011,
    input  [5:0] col_in_1012,
    input  [5:0] col_in_1013,
    input  [5:0] col_in_1014,
    input  [5:0] col_in_1015,
    input  [5:0] col_in_1016,
    input  [5:0] col_in_1017,
    input  [5:0] col_in_1018,
    input  [5:0] col_in_1019,
    input  [5:0] col_in_1020,
    input  [5:0] col_in_1021,
    input  [5:0] col_in_1022,
    input  [5:0] col_in_1023,

    output [3:0] col_out_0,
    output [3:0] col_out_1,
    output [3:0] col_out_2,
    output [3:0] col_out_3,
    output [3:0] col_out_4,
    output [3:0] col_out_5,
    output [3:0] col_out_6,
    output [3:0] col_out_7,
    output [3:0] col_out_8,
    output [3:0] col_out_9,
    output [3:0] col_out_10,
    output [3:0] col_out_11,
    output [3:0] col_out_12,
    output [3:0] col_out_13,
    output [3:0] col_out_14,
    output [3:0] col_out_15,
    output [3:0] col_out_16,
    output [3:0] col_out_17,
    output [3:0] col_out_18,
    output [3:0] col_out_19,
    output [3:0] col_out_20,
    output [3:0] col_out_21,
    output [3:0] col_out_22,
    output [3:0] col_out_23,
    output [3:0] col_out_24,
    output [3:0] col_out_25,
    output [3:0] col_out_26,
    output [3:0] col_out_27,
    output [3:0] col_out_28,
    output [3:0] col_out_29,
    output [3:0] col_out_30,
    output [3:0] col_out_31,
    output [3:0] col_out_32,
    output [3:0] col_out_33,
    output [3:0] col_out_34,
    output [3:0] col_out_35,
    output [3:0] col_out_36,
    output [3:0] col_out_37,
    output [3:0] col_out_38,
    output [3:0] col_out_39,
    output [3:0] col_out_40,
    output [3:0] col_out_41,
    output [3:0] col_out_42,
    output [3:0] col_out_43,
    output [3:0] col_out_44,
    output [3:0] col_out_45,
    output [3:0] col_out_46,
    output [3:0] col_out_47,
    output [3:0] col_out_48,
    output [3:0] col_out_49,
    output [3:0] col_out_50,
    output [3:0] col_out_51,
    output [3:0] col_out_52,
    output [3:0] col_out_53,
    output [3:0] col_out_54,
    output [3:0] col_out_55,
    output [3:0] col_out_56,
    output [3:0] col_out_57,
    output [3:0] col_out_58,
    output [3:0] col_out_59,
    output [3:0] col_out_60,
    output [3:0] col_out_61,
    output [3:0] col_out_62,
    output [3:0] col_out_63,
    output [3:0] col_out_64,
    output [3:0] col_out_65,
    output [3:0] col_out_66,
    output [3:0] col_out_67,
    output [3:0] col_out_68,
    output [3:0] col_out_69,
    output [3:0] col_out_70,
    output [3:0] col_out_71,
    output [3:0] col_out_72,
    output [3:0] col_out_73,
    output [3:0] col_out_74,
    output [3:0] col_out_75,
    output [3:0] col_out_76,
    output [3:0] col_out_77,
    output [3:0] col_out_78,
    output [3:0] col_out_79,
    output [3:0] col_out_80,
    output [3:0] col_out_81,
    output [3:0] col_out_82,
    output [3:0] col_out_83,
    output [3:0] col_out_84,
    output [3:0] col_out_85,
    output [3:0] col_out_86,
    output [3:0] col_out_87,
    output [3:0] col_out_88,
    output [3:0] col_out_89,
    output [3:0] col_out_90,
    output [3:0] col_out_91,
    output [3:0] col_out_92,
    output [3:0] col_out_93,
    output [3:0] col_out_94,
    output [3:0] col_out_95,
    output [3:0] col_out_96,
    output [3:0] col_out_97,
    output [3:0] col_out_98,
    output [3:0] col_out_99,
    output [3:0] col_out_100,
    output [3:0] col_out_101,
    output [3:0] col_out_102,
    output [3:0] col_out_103,
    output [3:0] col_out_104,
    output [3:0] col_out_105,
    output [3:0] col_out_106,
    output [3:0] col_out_107,
    output [3:0] col_out_108,
    output [3:0] col_out_109,
    output [3:0] col_out_110,
    output [3:0] col_out_111,
    output [3:0] col_out_112,
    output [3:0] col_out_113,
    output [3:0] col_out_114,
    output [3:0] col_out_115,
    output [3:0] col_out_116,
    output [3:0] col_out_117,
    output [3:0] col_out_118,
    output [3:0] col_out_119,
    output [3:0] col_out_120,
    output [3:0] col_out_121,
    output [3:0] col_out_122,
    output [3:0] col_out_123,
    output [3:0] col_out_124,
    output [3:0] col_out_125,
    output [3:0] col_out_126,
    output [3:0] col_out_127,
    output [3:0] col_out_128,
    output [3:0] col_out_129,
    output [3:0] col_out_130,
    output [3:0] col_out_131,
    output [3:0] col_out_132,
    output [3:0] col_out_133,
    output [3:0] col_out_134,
    output [3:0] col_out_135,
    output [3:0] col_out_136,
    output [3:0] col_out_137,
    output [3:0] col_out_138,
    output [3:0] col_out_139,
    output [3:0] col_out_140,
    output [3:0] col_out_141,
    output [3:0] col_out_142,
    output [3:0] col_out_143,
    output [3:0] col_out_144,
    output [3:0] col_out_145,
    output [3:0] col_out_146,
    output [3:0] col_out_147,
    output [3:0] col_out_148,
    output [3:0] col_out_149,
    output [3:0] col_out_150,
    output [3:0] col_out_151,
    output [3:0] col_out_152,
    output [3:0] col_out_153,
    output [3:0] col_out_154,
    output [3:0] col_out_155,
    output [3:0] col_out_156,
    output [3:0] col_out_157,
    output [3:0] col_out_158,
    output [3:0] col_out_159,
    output [3:0] col_out_160,
    output [3:0] col_out_161,
    output [3:0] col_out_162,
    output [3:0] col_out_163,
    output [3:0] col_out_164,
    output [3:0] col_out_165,
    output [3:0] col_out_166,
    output [3:0] col_out_167,
    output [3:0] col_out_168,
    output [3:0] col_out_169,
    output [3:0] col_out_170,
    output [3:0] col_out_171,
    output [3:0] col_out_172,
    output [3:0] col_out_173,
    output [3:0] col_out_174,
    output [3:0] col_out_175,
    output [3:0] col_out_176,
    output [3:0] col_out_177,
    output [3:0] col_out_178,
    output [3:0] col_out_179,
    output [3:0] col_out_180,
    output [3:0] col_out_181,
    output [3:0] col_out_182,
    output [3:0] col_out_183,
    output [3:0] col_out_184,
    output [3:0] col_out_185,
    output [3:0] col_out_186,
    output [3:0] col_out_187,
    output [3:0] col_out_188,
    output [3:0] col_out_189,
    output [3:0] col_out_190,
    output [3:0] col_out_191,
    output [3:0] col_out_192,
    output [3:0] col_out_193,
    output [3:0] col_out_194,
    output [3:0] col_out_195,
    output [3:0] col_out_196,
    output [3:0] col_out_197,
    output [3:0] col_out_198,
    output [3:0] col_out_199,
    output [3:0] col_out_200,
    output [3:0] col_out_201,
    output [3:0] col_out_202,
    output [3:0] col_out_203,
    output [3:0] col_out_204,
    output [3:0] col_out_205,
    output [3:0] col_out_206,
    output [3:0] col_out_207,
    output [3:0] col_out_208,
    output [3:0] col_out_209,
    output [3:0] col_out_210,
    output [3:0] col_out_211,
    output [3:0] col_out_212,
    output [3:0] col_out_213,
    output [3:0] col_out_214,
    output [3:0] col_out_215,
    output [3:0] col_out_216,
    output [3:0] col_out_217,
    output [3:0] col_out_218,
    output [3:0] col_out_219,
    output [3:0] col_out_220,
    output [3:0] col_out_221,
    output [3:0] col_out_222,
    output [3:0] col_out_223,
    output [3:0] col_out_224,
    output [3:0] col_out_225,
    output [3:0] col_out_226,
    output [3:0] col_out_227,
    output [3:0] col_out_228,
    output [3:0] col_out_229,
    output [3:0] col_out_230,
    output [3:0] col_out_231,
    output [3:0] col_out_232,
    output [3:0] col_out_233,
    output [3:0] col_out_234,
    output [3:0] col_out_235,
    output [3:0] col_out_236,
    output [3:0] col_out_237,
    output [3:0] col_out_238,
    output [3:0] col_out_239,
    output [3:0] col_out_240,
    output [3:0] col_out_241,
    output [3:0] col_out_242,
    output [3:0] col_out_243,
    output [3:0] col_out_244,
    output [3:0] col_out_245,
    output [3:0] col_out_246,
    output [3:0] col_out_247,
    output [3:0] col_out_248,
    output [3:0] col_out_249,
    output [3:0] col_out_250,
    output [3:0] col_out_251,
    output [3:0] col_out_252,
    output [3:0] col_out_253,
    output [3:0] col_out_254,
    output [3:0] col_out_255,
    output [3:0] col_out_256,
    output [3:0] col_out_257,
    output [3:0] col_out_258,
    output [3:0] col_out_259,
    output [3:0] col_out_260,
    output [3:0] col_out_261,
    output [3:0] col_out_262,
    output [3:0] col_out_263,
    output [3:0] col_out_264,
    output [3:0] col_out_265,
    output [3:0] col_out_266,
    output [3:0] col_out_267,
    output [3:0] col_out_268,
    output [3:0] col_out_269,
    output [3:0] col_out_270,
    output [3:0] col_out_271,
    output [3:0] col_out_272,
    output [3:0] col_out_273,
    output [3:0] col_out_274,
    output [3:0] col_out_275,
    output [3:0] col_out_276,
    output [3:0] col_out_277,
    output [3:0] col_out_278,
    output [3:0] col_out_279,
    output [3:0] col_out_280,
    output [3:0] col_out_281,
    output [3:0] col_out_282,
    output [3:0] col_out_283,
    output [3:0] col_out_284,
    output [3:0] col_out_285,
    output [3:0] col_out_286,
    output [3:0] col_out_287,
    output [3:0] col_out_288,
    output [3:0] col_out_289,
    output [3:0] col_out_290,
    output [3:0] col_out_291,
    output [3:0] col_out_292,
    output [3:0] col_out_293,
    output [3:0] col_out_294,
    output [3:0] col_out_295,
    output [3:0] col_out_296,
    output [3:0] col_out_297,
    output [3:0] col_out_298,
    output [3:0] col_out_299,
    output [3:0] col_out_300,
    output [3:0] col_out_301,
    output [3:0] col_out_302,
    output [3:0] col_out_303,
    output [3:0] col_out_304,
    output [3:0] col_out_305,
    output [3:0] col_out_306,
    output [3:0] col_out_307,
    output [3:0] col_out_308,
    output [3:0] col_out_309,
    output [3:0] col_out_310,
    output [3:0] col_out_311,
    output [3:0] col_out_312,
    output [3:0] col_out_313,
    output [3:0] col_out_314,
    output [3:0] col_out_315,
    output [3:0] col_out_316,
    output [3:0] col_out_317,
    output [3:0] col_out_318,
    output [3:0] col_out_319,
    output [3:0] col_out_320,
    output [3:0] col_out_321,
    output [3:0] col_out_322,
    output [3:0] col_out_323,
    output [3:0] col_out_324,
    output [3:0] col_out_325,
    output [3:0] col_out_326,
    output [3:0] col_out_327,
    output [3:0] col_out_328,
    output [3:0] col_out_329,
    output [3:0] col_out_330,
    output [3:0] col_out_331,
    output [3:0] col_out_332,
    output [3:0] col_out_333,
    output [3:0] col_out_334,
    output [3:0] col_out_335,
    output [3:0] col_out_336,
    output [3:0] col_out_337,
    output [3:0] col_out_338,
    output [3:0] col_out_339,
    output [3:0] col_out_340,
    output [3:0] col_out_341,
    output [3:0] col_out_342,
    output [3:0] col_out_343,
    output [3:0] col_out_344,
    output [3:0] col_out_345,
    output [3:0] col_out_346,
    output [3:0] col_out_347,
    output [3:0] col_out_348,
    output [3:0] col_out_349,
    output [3:0] col_out_350,
    output [3:0] col_out_351,
    output [3:0] col_out_352,
    output [3:0] col_out_353,
    output [3:0] col_out_354,
    output [3:0] col_out_355,
    output [3:0] col_out_356,
    output [3:0] col_out_357,
    output [3:0] col_out_358,
    output [3:0] col_out_359,
    output [3:0] col_out_360,
    output [3:0] col_out_361,
    output [3:0] col_out_362,
    output [3:0] col_out_363,
    output [3:0] col_out_364,
    output [3:0] col_out_365,
    output [3:0] col_out_366,
    output [3:0] col_out_367,
    output [3:0] col_out_368,
    output [3:0] col_out_369,
    output [3:0] col_out_370,
    output [3:0] col_out_371,
    output [3:0] col_out_372,
    output [3:0] col_out_373,
    output [3:0] col_out_374,
    output [3:0] col_out_375,
    output [3:0] col_out_376,
    output [3:0] col_out_377,
    output [3:0] col_out_378,
    output [3:0] col_out_379,
    output [3:0] col_out_380,
    output [3:0] col_out_381,
    output [3:0] col_out_382,
    output [3:0] col_out_383,
    output [3:0] col_out_384,
    output [3:0] col_out_385,
    output [3:0] col_out_386,
    output [3:0] col_out_387,
    output [3:0] col_out_388,
    output [3:0] col_out_389,
    output [3:0] col_out_390,
    output [3:0] col_out_391,
    output [3:0] col_out_392,
    output [3:0] col_out_393,
    output [3:0] col_out_394,
    output [3:0] col_out_395,
    output [3:0] col_out_396,
    output [3:0] col_out_397,
    output [3:0] col_out_398,
    output [3:0] col_out_399,
    output [3:0] col_out_400,
    output [3:0] col_out_401,
    output [3:0] col_out_402,
    output [3:0] col_out_403,
    output [3:0] col_out_404,
    output [3:0] col_out_405,
    output [3:0] col_out_406,
    output [3:0] col_out_407,
    output [3:0] col_out_408,
    output [3:0] col_out_409,
    output [3:0] col_out_410,
    output [3:0] col_out_411,
    output [3:0] col_out_412,
    output [3:0] col_out_413,
    output [3:0] col_out_414,
    output [3:0] col_out_415,
    output [3:0] col_out_416,
    output [3:0] col_out_417,
    output [3:0] col_out_418,
    output [3:0] col_out_419,
    output [3:0] col_out_420,
    output [3:0] col_out_421,
    output [3:0] col_out_422,
    output [3:0] col_out_423,
    output [3:0] col_out_424,
    output [3:0] col_out_425,
    output [3:0] col_out_426,
    output [3:0] col_out_427,
    output [3:0] col_out_428,
    output [3:0] col_out_429,
    output [3:0] col_out_430,
    output [3:0] col_out_431,
    output [3:0] col_out_432,
    output [3:0] col_out_433,
    output [3:0] col_out_434,
    output [3:0] col_out_435,
    output [3:0] col_out_436,
    output [3:0] col_out_437,
    output [3:0] col_out_438,
    output [3:0] col_out_439,
    output [3:0] col_out_440,
    output [3:0] col_out_441,
    output [3:0] col_out_442,
    output [3:0] col_out_443,
    output [3:0] col_out_444,
    output [3:0] col_out_445,
    output [3:0] col_out_446,
    output [3:0] col_out_447,
    output [3:0] col_out_448,
    output [3:0] col_out_449,
    output [3:0] col_out_450,
    output [3:0] col_out_451,
    output [3:0] col_out_452,
    output [3:0] col_out_453,
    output [3:0] col_out_454,
    output [3:0] col_out_455,
    output [3:0] col_out_456,
    output [3:0] col_out_457,
    output [3:0] col_out_458,
    output [3:0] col_out_459,
    output [3:0] col_out_460,
    output [3:0] col_out_461,
    output [3:0] col_out_462,
    output [3:0] col_out_463,
    output [3:0] col_out_464,
    output [3:0] col_out_465,
    output [3:0] col_out_466,
    output [3:0] col_out_467,
    output [3:0] col_out_468,
    output [3:0] col_out_469,
    output [3:0] col_out_470,
    output [3:0] col_out_471,
    output [3:0] col_out_472,
    output [3:0] col_out_473,
    output [3:0] col_out_474,
    output [3:0] col_out_475,
    output [3:0] col_out_476,
    output [3:0] col_out_477,
    output [3:0] col_out_478,
    output [3:0] col_out_479,
    output [3:0] col_out_480,
    output [3:0] col_out_481,
    output [3:0] col_out_482,
    output [3:0] col_out_483,
    output [3:0] col_out_484,
    output [3:0] col_out_485,
    output [3:0] col_out_486,
    output [3:0] col_out_487,
    output [3:0] col_out_488,
    output [3:0] col_out_489,
    output [3:0] col_out_490,
    output [3:0] col_out_491,
    output [3:0] col_out_492,
    output [3:0] col_out_493,
    output [3:0] col_out_494,
    output [3:0] col_out_495,
    output [3:0] col_out_496,
    output [3:0] col_out_497,
    output [3:0] col_out_498,
    output [3:0] col_out_499,
    output [3:0] col_out_500,
    output [3:0] col_out_501,
    output [3:0] col_out_502,
    output [3:0] col_out_503,
    output [3:0] col_out_504,
    output [3:0] col_out_505,
    output [3:0] col_out_506,
    output [3:0] col_out_507,
    output [3:0] col_out_508,
    output [3:0] col_out_509,
    output [3:0] col_out_510,
    output [3:0] col_out_511,
    output [3:0] col_out_512,
    output [3:0] col_out_513,
    output [3:0] col_out_514,
    output [3:0] col_out_515,
    output [3:0] col_out_516,
    output [3:0] col_out_517,
    output [3:0] col_out_518,
    output [3:0] col_out_519,
    output [3:0] col_out_520,
    output [3:0] col_out_521,
    output [3:0] col_out_522,
    output [3:0] col_out_523,
    output [3:0] col_out_524,
    output [3:0] col_out_525,
    output [3:0] col_out_526,
    output [3:0] col_out_527,
    output [3:0] col_out_528,
    output [3:0] col_out_529,
    output [3:0] col_out_530,
    output [3:0] col_out_531,
    output [3:0] col_out_532,
    output [3:0] col_out_533,
    output [3:0] col_out_534,
    output [3:0] col_out_535,
    output [3:0] col_out_536,
    output [3:0] col_out_537,
    output [3:0] col_out_538,
    output [3:0] col_out_539,
    output [3:0] col_out_540,
    output [3:0] col_out_541,
    output [3:0] col_out_542,
    output [3:0] col_out_543,
    output [3:0] col_out_544,
    output [3:0] col_out_545,
    output [3:0] col_out_546,
    output [3:0] col_out_547,
    output [3:0] col_out_548,
    output [3:0] col_out_549,
    output [3:0] col_out_550,
    output [3:0] col_out_551,
    output [3:0] col_out_552,
    output [3:0] col_out_553,
    output [3:0] col_out_554,
    output [3:0] col_out_555,
    output [3:0] col_out_556,
    output [3:0] col_out_557,
    output [3:0] col_out_558,
    output [3:0] col_out_559,
    output [3:0] col_out_560,
    output [3:0] col_out_561,
    output [3:0] col_out_562,
    output [3:0] col_out_563,
    output [3:0] col_out_564,
    output [3:0] col_out_565,
    output [3:0] col_out_566,
    output [3:0] col_out_567,
    output [3:0] col_out_568,
    output [3:0] col_out_569,
    output [3:0] col_out_570,
    output [3:0] col_out_571,
    output [3:0] col_out_572,
    output [3:0] col_out_573,
    output [3:0] col_out_574,
    output [3:0] col_out_575,
    output [3:0] col_out_576,
    output [3:0] col_out_577,
    output [3:0] col_out_578,
    output [3:0] col_out_579,
    output [3:0] col_out_580,
    output [3:0] col_out_581,
    output [3:0] col_out_582,
    output [3:0] col_out_583,
    output [3:0] col_out_584,
    output [3:0] col_out_585,
    output [3:0] col_out_586,
    output [3:0] col_out_587,
    output [3:0] col_out_588,
    output [3:0] col_out_589,
    output [3:0] col_out_590,
    output [3:0] col_out_591,
    output [3:0] col_out_592,
    output [3:0] col_out_593,
    output [3:0] col_out_594,
    output [3:0] col_out_595,
    output [3:0] col_out_596,
    output [3:0] col_out_597,
    output [3:0] col_out_598,
    output [3:0] col_out_599,
    output [3:0] col_out_600,
    output [3:0] col_out_601,
    output [3:0] col_out_602,
    output [3:0] col_out_603,
    output [3:0] col_out_604,
    output [3:0] col_out_605,
    output [3:0] col_out_606,
    output [3:0] col_out_607,
    output [3:0] col_out_608,
    output [3:0] col_out_609,
    output [3:0] col_out_610,
    output [3:0] col_out_611,
    output [3:0] col_out_612,
    output [3:0] col_out_613,
    output [3:0] col_out_614,
    output [3:0] col_out_615,
    output [3:0] col_out_616,
    output [3:0] col_out_617,
    output [3:0] col_out_618,
    output [3:0] col_out_619,
    output [3:0] col_out_620,
    output [3:0] col_out_621,
    output [3:0] col_out_622,
    output [3:0] col_out_623,
    output [3:0] col_out_624,
    output [3:0] col_out_625,
    output [3:0] col_out_626,
    output [3:0] col_out_627,
    output [3:0] col_out_628,
    output [3:0] col_out_629,
    output [3:0] col_out_630,
    output [3:0] col_out_631,
    output [3:0] col_out_632,
    output [3:0] col_out_633,
    output [3:0] col_out_634,
    output [3:0] col_out_635,
    output [3:0] col_out_636,
    output [3:0] col_out_637,
    output [3:0] col_out_638,
    output [3:0] col_out_639,
    output [3:0] col_out_640,
    output [3:0] col_out_641,
    output [3:0] col_out_642,
    output [3:0] col_out_643,
    output [3:0] col_out_644,
    output [3:0] col_out_645,
    output [3:0] col_out_646,
    output [3:0] col_out_647,
    output [3:0] col_out_648,
    output [3:0] col_out_649,
    output [3:0] col_out_650,
    output [3:0] col_out_651,
    output [3:0] col_out_652,
    output [3:0] col_out_653,
    output [3:0] col_out_654,
    output [3:0] col_out_655,
    output [3:0] col_out_656,
    output [3:0] col_out_657,
    output [3:0] col_out_658,
    output [3:0] col_out_659,
    output [3:0] col_out_660,
    output [3:0] col_out_661,
    output [3:0] col_out_662,
    output [3:0] col_out_663,
    output [3:0] col_out_664,
    output [3:0] col_out_665,
    output [3:0] col_out_666,
    output [3:0] col_out_667,
    output [3:0] col_out_668,
    output [3:0] col_out_669,
    output [3:0] col_out_670,
    output [3:0] col_out_671,
    output [3:0] col_out_672,
    output [3:0] col_out_673,
    output [3:0] col_out_674,
    output [3:0] col_out_675,
    output [3:0] col_out_676,
    output [3:0] col_out_677,
    output [3:0] col_out_678,
    output [3:0] col_out_679,
    output [3:0] col_out_680,
    output [3:0] col_out_681,
    output [3:0] col_out_682,
    output [3:0] col_out_683,
    output [3:0] col_out_684,
    output [3:0] col_out_685,
    output [3:0] col_out_686,
    output [3:0] col_out_687,
    output [3:0] col_out_688,
    output [3:0] col_out_689,
    output [3:0] col_out_690,
    output [3:0] col_out_691,
    output [3:0] col_out_692,
    output [3:0] col_out_693,
    output [3:0] col_out_694,
    output [3:0] col_out_695,
    output [3:0] col_out_696,
    output [3:0] col_out_697,
    output [3:0] col_out_698,
    output [3:0] col_out_699,
    output [3:0] col_out_700,
    output [3:0] col_out_701,
    output [3:0] col_out_702,
    output [3:0] col_out_703,
    output [3:0] col_out_704,
    output [3:0] col_out_705,
    output [3:0] col_out_706,
    output [3:0] col_out_707,
    output [3:0] col_out_708,
    output [3:0] col_out_709,
    output [3:0] col_out_710,
    output [3:0] col_out_711,
    output [3:0] col_out_712,
    output [3:0] col_out_713,
    output [3:0] col_out_714,
    output [3:0] col_out_715,
    output [3:0] col_out_716,
    output [3:0] col_out_717,
    output [3:0] col_out_718,
    output [3:0] col_out_719,
    output [3:0] col_out_720,
    output [3:0] col_out_721,
    output [3:0] col_out_722,
    output [3:0] col_out_723,
    output [3:0] col_out_724,
    output [3:0] col_out_725,
    output [3:0] col_out_726,
    output [3:0] col_out_727,
    output [3:0] col_out_728,
    output [3:0] col_out_729,
    output [3:0] col_out_730,
    output [3:0] col_out_731,
    output [3:0] col_out_732,
    output [3:0] col_out_733,
    output [3:0] col_out_734,
    output [3:0] col_out_735,
    output [3:0] col_out_736,
    output [3:0] col_out_737,
    output [3:0] col_out_738,
    output [3:0] col_out_739,
    output [3:0] col_out_740,
    output [3:0] col_out_741,
    output [3:0] col_out_742,
    output [3:0] col_out_743,
    output [3:0] col_out_744,
    output [3:0] col_out_745,
    output [3:0] col_out_746,
    output [3:0] col_out_747,
    output [3:0] col_out_748,
    output [3:0] col_out_749,
    output [3:0] col_out_750,
    output [3:0] col_out_751,
    output [3:0] col_out_752,
    output [3:0] col_out_753,
    output [3:0] col_out_754,
    output [3:0] col_out_755,
    output [3:0] col_out_756,
    output [3:0] col_out_757,
    output [3:0] col_out_758,
    output [3:0] col_out_759,
    output [3:0] col_out_760,
    output [3:0] col_out_761,
    output [3:0] col_out_762,
    output [3:0] col_out_763,
    output [3:0] col_out_764,
    output [3:0] col_out_765,
    output [3:0] col_out_766,
    output [3:0] col_out_767,
    output [3:0] col_out_768,
    output [3:0] col_out_769,
    output [3:0] col_out_770,
    output [3:0] col_out_771,
    output [3:0] col_out_772,
    output [3:0] col_out_773,
    output [3:0] col_out_774,
    output [3:0] col_out_775,
    output [3:0] col_out_776,
    output [3:0] col_out_777,
    output [3:0] col_out_778,
    output [3:0] col_out_779,
    output [3:0] col_out_780,
    output [3:0] col_out_781,
    output [3:0] col_out_782,
    output [3:0] col_out_783,
    output [3:0] col_out_784,
    output [3:0] col_out_785,
    output [3:0] col_out_786,
    output [3:0] col_out_787,
    output [3:0] col_out_788,
    output [3:0] col_out_789,
    output [3:0] col_out_790,
    output [3:0] col_out_791,
    output [3:0] col_out_792,
    output [3:0] col_out_793,
    output [3:0] col_out_794,
    output [3:0] col_out_795,
    output [3:0] col_out_796,
    output [3:0] col_out_797,
    output [3:0] col_out_798,
    output [3:0] col_out_799,
    output [3:0] col_out_800,
    output [3:0] col_out_801,
    output [3:0] col_out_802,
    output [3:0] col_out_803,
    output [3:0] col_out_804,
    output [3:0] col_out_805,
    output [3:0] col_out_806,
    output [3:0] col_out_807,
    output [3:0] col_out_808,
    output [3:0] col_out_809,
    output [3:0] col_out_810,
    output [3:0] col_out_811,
    output [3:0] col_out_812,
    output [3:0] col_out_813,
    output [3:0] col_out_814,
    output [3:0] col_out_815,
    output [3:0] col_out_816,
    output [3:0] col_out_817,
    output [3:0] col_out_818,
    output [3:0] col_out_819,
    output [3:0] col_out_820,
    output [3:0] col_out_821,
    output [3:0] col_out_822,
    output [3:0] col_out_823,
    output [3:0] col_out_824,
    output [3:0] col_out_825,
    output [3:0] col_out_826,
    output [3:0] col_out_827,
    output [3:0] col_out_828,
    output [3:0] col_out_829,
    output [3:0] col_out_830,
    output [3:0] col_out_831,
    output [3:0] col_out_832,
    output [3:0] col_out_833,
    output [3:0] col_out_834,
    output [3:0] col_out_835,
    output [3:0] col_out_836,
    output [3:0] col_out_837,
    output [3:0] col_out_838,
    output [3:0] col_out_839,
    output [3:0] col_out_840,
    output [3:0] col_out_841,
    output [3:0] col_out_842,
    output [3:0] col_out_843,
    output [3:0] col_out_844,
    output [3:0] col_out_845,
    output [3:0] col_out_846,
    output [3:0] col_out_847,
    output [3:0] col_out_848,
    output [3:0] col_out_849,
    output [3:0] col_out_850,
    output [3:0] col_out_851,
    output [3:0] col_out_852,
    output [3:0] col_out_853,
    output [3:0] col_out_854,
    output [3:0] col_out_855,
    output [3:0] col_out_856,
    output [3:0] col_out_857,
    output [3:0] col_out_858,
    output [3:0] col_out_859,
    output [3:0] col_out_860,
    output [3:0] col_out_861,
    output [3:0] col_out_862,
    output [3:0] col_out_863,
    output [3:0] col_out_864,
    output [3:0] col_out_865,
    output [3:0] col_out_866,
    output [3:0] col_out_867,
    output [3:0] col_out_868,
    output [3:0] col_out_869,
    output [3:0] col_out_870,
    output [3:0] col_out_871,
    output [3:0] col_out_872,
    output [3:0] col_out_873,
    output [3:0] col_out_874,
    output [3:0] col_out_875,
    output [3:0] col_out_876,
    output [3:0] col_out_877,
    output [3:0] col_out_878,
    output [3:0] col_out_879,
    output [3:0] col_out_880,
    output [3:0] col_out_881,
    output [3:0] col_out_882,
    output [3:0] col_out_883,
    output [3:0] col_out_884,
    output [3:0] col_out_885,
    output [3:0] col_out_886,
    output [3:0] col_out_887,
    output [3:0] col_out_888,
    output [3:0] col_out_889,
    output [3:0] col_out_890,
    output [3:0] col_out_891,
    output [3:0] col_out_892,
    output [3:0] col_out_893,
    output [3:0] col_out_894,
    output [3:0] col_out_895,
    output [3:0] col_out_896,
    output [3:0] col_out_897,
    output [3:0] col_out_898,
    output [3:0] col_out_899,
    output [3:0] col_out_900,
    output [3:0] col_out_901,
    output [3:0] col_out_902,
    output [3:0] col_out_903,
    output [3:0] col_out_904,
    output [3:0] col_out_905,
    output [3:0] col_out_906,
    output [3:0] col_out_907,
    output [3:0] col_out_908,
    output [3:0] col_out_909,
    output [3:0] col_out_910,
    output [3:0] col_out_911,
    output [3:0] col_out_912,
    output [3:0] col_out_913,
    output [3:0] col_out_914,
    output [3:0] col_out_915,
    output [3:0] col_out_916,
    output [3:0] col_out_917,
    output [3:0] col_out_918,
    output [3:0] col_out_919,
    output [3:0] col_out_920,
    output [3:0] col_out_921,
    output [3:0] col_out_922,
    output [3:0] col_out_923,
    output [3:0] col_out_924,
    output [3:0] col_out_925,
    output [3:0] col_out_926,
    output [3:0] col_out_927,
    output [3:0] col_out_928,
    output [3:0] col_out_929,
    output [3:0] col_out_930,
    output [3:0] col_out_931,
    output [3:0] col_out_932,
    output [3:0] col_out_933,
    output [3:0] col_out_934,
    output [3:0] col_out_935,
    output [3:0] col_out_936,
    output [3:0] col_out_937,
    output [3:0] col_out_938,
    output [3:0] col_out_939,
    output [3:0] col_out_940,
    output [3:0] col_out_941,
    output [3:0] col_out_942,
    output [3:0] col_out_943,
    output [3:0] col_out_944,
    output [3:0] col_out_945,
    output [3:0] col_out_946,
    output [3:0] col_out_947,
    output [3:0] col_out_948,
    output [3:0] col_out_949,
    output [3:0] col_out_950,
    output [3:0] col_out_951,
    output [3:0] col_out_952,
    output [3:0] col_out_953,
    output [3:0] col_out_954,
    output [3:0] col_out_955,
    output [3:0] col_out_956,
    output [3:0] col_out_957,
    output [3:0] col_out_958,
    output [3:0] col_out_959,
    output [3:0] col_out_960,
    output [3:0] col_out_961,
    output [3:0] col_out_962,
    output [3:0] col_out_963,
    output [3:0] col_out_964,
    output [3:0] col_out_965,
    output [3:0] col_out_966,
    output [3:0] col_out_967,
    output [3:0] col_out_968,
    output [3:0] col_out_969,
    output [3:0] col_out_970,
    output [3:0] col_out_971,
    output [3:0] col_out_972,
    output [3:0] col_out_973,
    output [3:0] col_out_974,
    output [3:0] col_out_975,
    output [3:0] col_out_976,
    output [3:0] col_out_977,
    output [3:0] col_out_978,
    output [3:0] col_out_979,
    output [3:0] col_out_980,
    output [3:0] col_out_981,
    output [3:0] col_out_982,
    output [3:0] col_out_983,
    output [3:0] col_out_984,
    output [3:0] col_out_985,
    output [3:0] col_out_986,
    output [3:0] col_out_987,
    output [3:0] col_out_988,
    output [3:0] col_out_989,
    output [3:0] col_out_990,
    output [3:0] col_out_991,
    output [3:0] col_out_992,
    output [3:0] col_out_993,
    output [3:0] col_out_994,
    output [3:0] col_out_995,
    output [3:0] col_out_996,
    output [3:0] col_out_997,
    output [3:0] col_out_998,
    output [3:0] col_out_999,
    output [3:0] col_out_1000,
    output [3:0] col_out_1001,
    output [3:0] col_out_1002,
    output [3:0] col_out_1003,
    output [3:0] col_out_1004,
    output [3:0] col_out_1005,
    output [3:0] col_out_1006,
    output [3:0] col_out_1007,
    output [3:0] col_out_1008,
    output [3:0] col_out_1009,
    output [3:0] col_out_1010,
    output [3:0] col_out_1011,
    output [3:0] col_out_1012,
    output [3:0] col_out_1013,
    output [3:0] col_out_1014,
    output [3:0] col_out_1015,
    output [3:0] col_out_1016,
    output [3:0] col_out_1017,
    output [3:0] col_out_1018,
    output [3:0] col_out_1019,
    output [3:0] col_out_1020,
    output [3:0] col_out_1021,
    output [3:0] col_out_1022,
    output [3:0] col_out_1023,
    output [3:0] col_out_1024
);



//--compressor_array input and output----------------------

wire [5:0] u_ca_in_0;
wire [5:0] u_ca_in_1;
wire [5:0] u_ca_in_2;
wire [5:0] u_ca_in_3;
wire [5:0] u_ca_in_4;
wire [5:0] u_ca_in_5;
wire [5:0] u_ca_in_6;
wire [5:0] u_ca_in_7;
wire [5:0] u_ca_in_8;
wire [5:0] u_ca_in_9;
wire [5:0] u_ca_in_10;
wire [5:0] u_ca_in_11;
wire [5:0] u_ca_in_12;
wire [5:0] u_ca_in_13;
wire [5:0] u_ca_in_14;
wire [5:0] u_ca_in_15;
wire [5:0] u_ca_in_16;
wire [5:0] u_ca_in_17;
wire [5:0] u_ca_in_18;
wire [5:0] u_ca_in_19;
wire [5:0] u_ca_in_20;
wire [5:0] u_ca_in_21;
wire [5:0] u_ca_in_22;
wire [5:0] u_ca_in_23;
wire [5:0] u_ca_in_24;
wire [5:0] u_ca_in_25;
wire [5:0] u_ca_in_26;
wire [5:0] u_ca_in_27;
wire [5:0] u_ca_in_28;
wire [5:0] u_ca_in_29;
wire [5:0] u_ca_in_30;
wire [5:0] u_ca_in_31;
wire [5:0] u_ca_in_32;
wire [5:0] u_ca_in_33;
wire [5:0] u_ca_in_34;
wire [5:0] u_ca_in_35;
wire [5:0] u_ca_in_36;
wire [5:0] u_ca_in_37;
wire [5:0] u_ca_in_38;
wire [5:0] u_ca_in_39;
wire [5:0] u_ca_in_40;
wire [5:0] u_ca_in_41;
wire [5:0] u_ca_in_42;
wire [5:0] u_ca_in_43;
wire [5:0] u_ca_in_44;
wire [5:0] u_ca_in_45;
wire [5:0] u_ca_in_46;
wire [5:0] u_ca_in_47;
wire [5:0] u_ca_in_48;
wire [5:0] u_ca_in_49;
wire [5:0] u_ca_in_50;
wire [5:0] u_ca_in_51;
wire [5:0] u_ca_in_52;
wire [5:0] u_ca_in_53;
wire [5:0] u_ca_in_54;
wire [5:0] u_ca_in_55;
wire [5:0] u_ca_in_56;
wire [5:0] u_ca_in_57;
wire [5:0] u_ca_in_58;
wire [5:0] u_ca_in_59;
wire [5:0] u_ca_in_60;
wire [5:0] u_ca_in_61;
wire [5:0] u_ca_in_62;
wire [5:0] u_ca_in_63;
wire [5:0] u_ca_in_64;
wire [5:0] u_ca_in_65;
wire [5:0] u_ca_in_66;
wire [5:0] u_ca_in_67;
wire [5:0] u_ca_in_68;
wire [5:0] u_ca_in_69;
wire [5:0] u_ca_in_70;
wire [5:0] u_ca_in_71;
wire [5:0] u_ca_in_72;
wire [5:0] u_ca_in_73;
wire [5:0] u_ca_in_74;
wire [5:0] u_ca_in_75;
wire [5:0] u_ca_in_76;
wire [5:0] u_ca_in_77;
wire [5:0] u_ca_in_78;
wire [5:0] u_ca_in_79;
wire [5:0] u_ca_in_80;
wire [5:0] u_ca_in_81;
wire [5:0] u_ca_in_82;
wire [5:0] u_ca_in_83;
wire [5:0] u_ca_in_84;
wire [5:0] u_ca_in_85;
wire [5:0] u_ca_in_86;
wire [5:0] u_ca_in_87;
wire [5:0] u_ca_in_88;
wire [5:0] u_ca_in_89;
wire [5:0] u_ca_in_90;
wire [5:0] u_ca_in_91;
wire [5:0] u_ca_in_92;
wire [5:0] u_ca_in_93;
wire [5:0] u_ca_in_94;
wire [5:0] u_ca_in_95;
wire [5:0] u_ca_in_96;
wire [5:0] u_ca_in_97;
wire [5:0] u_ca_in_98;
wire [5:0] u_ca_in_99;
wire [5:0] u_ca_in_100;
wire [5:0] u_ca_in_101;
wire [5:0] u_ca_in_102;
wire [5:0] u_ca_in_103;
wire [5:0] u_ca_in_104;
wire [5:0] u_ca_in_105;
wire [5:0] u_ca_in_106;
wire [5:0] u_ca_in_107;
wire [5:0] u_ca_in_108;
wire [5:0] u_ca_in_109;
wire [5:0] u_ca_in_110;
wire [5:0] u_ca_in_111;
wire [5:0] u_ca_in_112;
wire [5:0] u_ca_in_113;
wire [5:0] u_ca_in_114;
wire [5:0] u_ca_in_115;
wire [5:0] u_ca_in_116;
wire [5:0] u_ca_in_117;
wire [5:0] u_ca_in_118;
wire [5:0] u_ca_in_119;
wire [5:0] u_ca_in_120;
wire [5:0] u_ca_in_121;
wire [5:0] u_ca_in_122;
wire [5:0] u_ca_in_123;
wire [5:0] u_ca_in_124;
wire [5:0] u_ca_in_125;
wire [5:0] u_ca_in_126;
wire [5:0] u_ca_in_127;
wire [5:0] u_ca_in_128;
wire [5:0] u_ca_in_129;
wire [5:0] u_ca_in_130;
wire [5:0] u_ca_in_131;
wire [5:0] u_ca_in_132;
wire [5:0] u_ca_in_133;
wire [5:0] u_ca_in_134;
wire [5:0] u_ca_in_135;
wire [5:0] u_ca_in_136;
wire [5:0] u_ca_in_137;
wire [5:0] u_ca_in_138;
wire [5:0] u_ca_in_139;
wire [5:0] u_ca_in_140;
wire [5:0] u_ca_in_141;
wire [5:0] u_ca_in_142;
wire [5:0] u_ca_in_143;
wire [5:0] u_ca_in_144;
wire [5:0] u_ca_in_145;
wire [5:0] u_ca_in_146;
wire [5:0] u_ca_in_147;
wire [5:0] u_ca_in_148;
wire [5:0] u_ca_in_149;
wire [5:0] u_ca_in_150;
wire [5:0] u_ca_in_151;
wire [5:0] u_ca_in_152;
wire [5:0] u_ca_in_153;
wire [5:0] u_ca_in_154;
wire [5:0] u_ca_in_155;
wire [5:0] u_ca_in_156;
wire [5:0] u_ca_in_157;
wire [5:0] u_ca_in_158;
wire [5:0] u_ca_in_159;
wire [5:0] u_ca_in_160;
wire [5:0] u_ca_in_161;
wire [5:0] u_ca_in_162;
wire [5:0] u_ca_in_163;
wire [5:0] u_ca_in_164;
wire [5:0] u_ca_in_165;
wire [5:0] u_ca_in_166;
wire [5:0] u_ca_in_167;
wire [5:0] u_ca_in_168;
wire [5:0] u_ca_in_169;
wire [5:0] u_ca_in_170;
wire [5:0] u_ca_in_171;
wire [5:0] u_ca_in_172;
wire [5:0] u_ca_in_173;
wire [5:0] u_ca_in_174;
wire [5:0] u_ca_in_175;
wire [5:0] u_ca_in_176;
wire [5:0] u_ca_in_177;
wire [5:0] u_ca_in_178;
wire [5:0] u_ca_in_179;
wire [5:0] u_ca_in_180;
wire [5:0] u_ca_in_181;
wire [5:0] u_ca_in_182;
wire [5:0] u_ca_in_183;
wire [5:0] u_ca_in_184;
wire [5:0] u_ca_in_185;
wire [5:0] u_ca_in_186;
wire [5:0] u_ca_in_187;
wire [5:0] u_ca_in_188;
wire [5:0] u_ca_in_189;
wire [5:0] u_ca_in_190;
wire [5:0] u_ca_in_191;
wire [5:0] u_ca_in_192;
wire [5:0] u_ca_in_193;
wire [5:0] u_ca_in_194;
wire [5:0] u_ca_in_195;
wire [5:0] u_ca_in_196;
wire [5:0] u_ca_in_197;
wire [5:0] u_ca_in_198;
wire [5:0] u_ca_in_199;
wire [5:0] u_ca_in_200;
wire [5:0] u_ca_in_201;
wire [5:0] u_ca_in_202;
wire [5:0] u_ca_in_203;
wire [5:0] u_ca_in_204;
wire [5:0] u_ca_in_205;
wire [5:0] u_ca_in_206;
wire [5:0] u_ca_in_207;
wire [5:0] u_ca_in_208;
wire [5:0] u_ca_in_209;
wire [5:0] u_ca_in_210;
wire [5:0] u_ca_in_211;
wire [5:0] u_ca_in_212;
wire [5:0] u_ca_in_213;
wire [5:0] u_ca_in_214;
wire [5:0] u_ca_in_215;
wire [5:0] u_ca_in_216;
wire [5:0] u_ca_in_217;
wire [5:0] u_ca_in_218;
wire [5:0] u_ca_in_219;
wire [5:0] u_ca_in_220;
wire [5:0] u_ca_in_221;
wire [5:0] u_ca_in_222;
wire [5:0] u_ca_in_223;
wire [5:0] u_ca_in_224;
wire [5:0] u_ca_in_225;
wire [5:0] u_ca_in_226;
wire [5:0] u_ca_in_227;
wire [5:0] u_ca_in_228;
wire [5:0] u_ca_in_229;
wire [5:0] u_ca_in_230;
wire [5:0] u_ca_in_231;
wire [5:0] u_ca_in_232;
wire [5:0] u_ca_in_233;
wire [5:0] u_ca_in_234;
wire [5:0] u_ca_in_235;
wire [5:0] u_ca_in_236;
wire [5:0] u_ca_in_237;
wire [5:0] u_ca_in_238;
wire [5:0] u_ca_in_239;
wire [5:0] u_ca_in_240;
wire [5:0] u_ca_in_241;
wire [5:0] u_ca_in_242;
wire [5:0] u_ca_in_243;
wire [5:0] u_ca_in_244;
wire [5:0] u_ca_in_245;
wire [5:0] u_ca_in_246;
wire [5:0] u_ca_in_247;
wire [5:0] u_ca_in_248;
wire [5:0] u_ca_in_249;
wire [5:0] u_ca_in_250;
wire [5:0] u_ca_in_251;
wire [5:0] u_ca_in_252;
wire [5:0] u_ca_in_253;
wire [5:0] u_ca_in_254;
wire [5:0] u_ca_in_255;
wire [5:0] u_ca_in_256;
wire [5:0] u_ca_in_257;
wire [5:0] u_ca_in_258;
wire [5:0] u_ca_in_259;
wire [5:0] u_ca_in_260;
wire [5:0] u_ca_in_261;
wire [5:0] u_ca_in_262;
wire [5:0] u_ca_in_263;
wire [5:0] u_ca_in_264;
wire [5:0] u_ca_in_265;
wire [5:0] u_ca_in_266;
wire [5:0] u_ca_in_267;
wire [5:0] u_ca_in_268;
wire [5:0] u_ca_in_269;
wire [5:0] u_ca_in_270;
wire [5:0] u_ca_in_271;
wire [5:0] u_ca_in_272;
wire [5:0] u_ca_in_273;
wire [5:0] u_ca_in_274;
wire [5:0] u_ca_in_275;
wire [5:0] u_ca_in_276;
wire [5:0] u_ca_in_277;
wire [5:0] u_ca_in_278;
wire [5:0] u_ca_in_279;
wire [5:0] u_ca_in_280;
wire [5:0] u_ca_in_281;
wire [5:0] u_ca_in_282;
wire [5:0] u_ca_in_283;
wire [5:0] u_ca_in_284;
wire [5:0] u_ca_in_285;
wire [5:0] u_ca_in_286;
wire [5:0] u_ca_in_287;
wire [5:0] u_ca_in_288;
wire [5:0] u_ca_in_289;
wire [5:0] u_ca_in_290;
wire [5:0] u_ca_in_291;
wire [5:0] u_ca_in_292;
wire [5:0] u_ca_in_293;
wire [5:0] u_ca_in_294;
wire [5:0] u_ca_in_295;
wire [5:0] u_ca_in_296;
wire [5:0] u_ca_in_297;
wire [5:0] u_ca_in_298;
wire [5:0] u_ca_in_299;
wire [5:0] u_ca_in_300;
wire [5:0] u_ca_in_301;
wire [5:0] u_ca_in_302;
wire [5:0] u_ca_in_303;
wire [5:0] u_ca_in_304;
wire [5:0] u_ca_in_305;
wire [5:0] u_ca_in_306;
wire [5:0] u_ca_in_307;
wire [5:0] u_ca_in_308;
wire [5:0] u_ca_in_309;
wire [5:0] u_ca_in_310;
wire [5:0] u_ca_in_311;
wire [5:0] u_ca_in_312;
wire [5:0] u_ca_in_313;
wire [5:0] u_ca_in_314;
wire [5:0] u_ca_in_315;
wire [5:0] u_ca_in_316;
wire [5:0] u_ca_in_317;
wire [5:0] u_ca_in_318;
wire [5:0] u_ca_in_319;
wire [5:0] u_ca_in_320;
wire [5:0] u_ca_in_321;
wire [5:0] u_ca_in_322;
wire [5:0] u_ca_in_323;
wire [5:0] u_ca_in_324;
wire [5:0] u_ca_in_325;
wire [5:0] u_ca_in_326;
wire [5:0] u_ca_in_327;
wire [5:0] u_ca_in_328;
wire [5:0] u_ca_in_329;
wire [5:0] u_ca_in_330;
wire [5:0] u_ca_in_331;
wire [5:0] u_ca_in_332;
wire [5:0] u_ca_in_333;
wire [5:0] u_ca_in_334;
wire [5:0] u_ca_in_335;
wire [5:0] u_ca_in_336;
wire [5:0] u_ca_in_337;
wire [5:0] u_ca_in_338;
wire [5:0] u_ca_in_339;
wire [5:0] u_ca_in_340;
wire [5:0] u_ca_in_341;
wire [5:0] u_ca_in_342;
wire [5:0] u_ca_in_343;
wire [5:0] u_ca_in_344;
wire [5:0] u_ca_in_345;
wire [5:0] u_ca_in_346;
wire [5:0] u_ca_in_347;
wire [5:0] u_ca_in_348;
wire [5:0] u_ca_in_349;
wire [5:0] u_ca_in_350;
wire [5:0] u_ca_in_351;
wire [5:0] u_ca_in_352;
wire [5:0] u_ca_in_353;
wire [5:0] u_ca_in_354;
wire [5:0] u_ca_in_355;
wire [5:0] u_ca_in_356;
wire [5:0] u_ca_in_357;
wire [5:0] u_ca_in_358;
wire [5:0] u_ca_in_359;
wire [5:0] u_ca_in_360;
wire [5:0] u_ca_in_361;
wire [5:0] u_ca_in_362;
wire [5:0] u_ca_in_363;
wire [5:0] u_ca_in_364;
wire [5:0] u_ca_in_365;
wire [5:0] u_ca_in_366;
wire [5:0] u_ca_in_367;
wire [5:0] u_ca_in_368;
wire [5:0] u_ca_in_369;
wire [5:0] u_ca_in_370;
wire [5:0] u_ca_in_371;
wire [5:0] u_ca_in_372;
wire [5:0] u_ca_in_373;
wire [5:0] u_ca_in_374;
wire [5:0] u_ca_in_375;
wire [5:0] u_ca_in_376;
wire [5:0] u_ca_in_377;
wire [5:0] u_ca_in_378;
wire [5:0] u_ca_in_379;
wire [5:0] u_ca_in_380;
wire [5:0] u_ca_in_381;
wire [5:0] u_ca_in_382;
wire [5:0] u_ca_in_383;
wire [5:0] u_ca_in_384;
wire [5:0] u_ca_in_385;
wire [5:0] u_ca_in_386;
wire [5:0] u_ca_in_387;
wire [5:0] u_ca_in_388;
wire [5:0] u_ca_in_389;
wire [5:0] u_ca_in_390;
wire [5:0] u_ca_in_391;
wire [5:0] u_ca_in_392;
wire [5:0] u_ca_in_393;
wire [5:0] u_ca_in_394;
wire [5:0] u_ca_in_395;
wire [5:0] u_ca_in_396;
wire [5:0] u_ca_in_397;
wire [5:0] u_ca_in_398;
wire [5:0] u_ca_in_399;
wire [5:0] u_ca_in_400;
wire [5:0] u_ca_in_401;
wire [5:0] u_ca_in_402;
wire [5:0] u_ca_in_403;
wire [5:0] u_ca_in_404;
wire [5:0] u_ca_in_405;
wire [5:0] u_ca_in_406;
wire [5:0] u_ca_in_407;
wire [5:0] u_ca_in_408;
wire [5:0] u_ca_in_409;
wire [5:0] u_ca_in_410;
wire [5:0] u_ca_in_411;
wire [5:0] u_ca_in_412;
wire [5:0] u_ca_in_413;
wire [5:0] u_ca_in_414;
wire [5:0] u_ca_in_415;
wire [5:0] u_ca_in_416;
wire [5:0] u_ca_in_417;
wire [5:0] u_ca_in_418;
wire [5:0] u_ca_in_419;
wire [5:0] u_ca_in_420;
wire [5:0] u_ca_in_421;
wire [5:0] u_ca_in_422;
wire [5:0] u_ca_in_423;
wire [5:0] u_ca_in_424;
wire [5:0] u_ca_in_425;
wire [5:0] u_ca_in_426;
wire [5:0] u_ca_in_427;
wire [5:0] u_ca_in_428;
wire [5:0] u_ca_in_429;
wire [5:0] u_ca_in_430;
wire [5:0] u_ca_in_431;
wire [5:0] u_ca_in_432;
wire [5:0] u_ca_in_433;
wire [5:0] u_ca_in_434;
wire [5:0] u_ca_in_435;
wire [5:0] u_ca_in_436;
wire [5:0] u_ca_in_437;
wire [5:0] u_ca_in_438;
wire [5:0] u_ca_in_439;
wire [5:0] u_ca_in_440;
wire [5:0] u_ca_in_441;
wire [5:0] u_ca_in_442;
wire [5:0] u_ca_in_443;
wire [5:0] u_ca_in_444;
wire [5:0] u_ca_in_445;
wire [5:0] u_ca_in_446;
wire [5:0] u_ca_in_447;
wire [5:0] u_ca_in_448;
wire [5:0] u_ca_in_449;
wire [5:0] u_ca_in_450;
wire [5:0] u_ca_in_451;
wire [5:0] u_ca_in_452;
wire [5:0] u_ca_in_453;
wire [5:0] u_ca_in_454;
wire [5:0] u_ca_in_455;
wire [5:0] u_ca_in_456;
wire [5:0] u_ca_in_457;
wire [5:0] u_ca_in_458;
wire [5:0] u_ca_in_459;
wire [5:0] u_ca_in_460;
wire [5:0] u_ca_in_461;
wire [5:0] u_ca_in_462;
wire [5:0] u_ca_in_463;
wire [5:0] u_ca_in_464;
wire [5:0] u_ca_in_465;
wire [5:0] u_ca_in_466;
wire [5:0] u_ca_in_467;
wire [5:0] u_ca_in_468;
wire [5:0] u_ca_in_469;
wire [5:0] u_ca_in_470;
wire [5:0] u_ca_in_471;
wire [5:0] u_ca_in_472;
wire [5:0] u_ca_in_473;
wire [5:0] u_ca_in_474;
wire [5:0] u_ca_in_475;
wire [5:0] u_ca_in_476;
wire [5:0] u_ca_in_477;
wire [5:0] u_ca_in_478;
wire [5:0] u_ca_in_479;
wire [5:0] u_ca_in_480;
wire [5:0] u_ca_in_481;
wire [5:0] u_ca_in_482;
wire [5:0] u_ca_in_483;
wire [5:0] u_ca_in_484;
wire [5:0] u_ca_in_485;
wire [5:0] u_ca_in_486;
wire [5:0] u_ca_in_487;
wire [5:0] u_ca_in_488;
wire [5:0] u_ca_in_489;
wire [5:0] u_ca_in_490;
wire [5:0] u_ca_in_491;
wire [5:0] u_ca_in_492;
wire [5:0] u_ca_in_493;
wire [5:0] u_ca_in_494;
wire [5:0] u_ca_in_495;
wire [5:0] u_ca_in_496;
wire [5:0] u_ca_in_497;
wire [5:0] u_ca_in_498;
wire [5:0] u_ca_in_499;
wire [5:0] u_ca_in_500;
wire [5:0] u_ca_in_501;
wire [5:0] u_ca_in_502;
wire [5:0] u_ca_in_503;
wire [5:0] u_ca_in_504;
wire [5:0] u_ca_in_505;
wire [5:0] u_ca_in_506;
wire [5:0] u_ca_in_507;
wire [5:0] u_ca_in_508;
wire [5:0] u_ca_in_509;
wire [5:0] u_ca_in_510;
wire [5:0] u_ca_in_511;
wire [5:0] u_ca_in_512;
wire [5:0] u_ca_in_513;
wire [5:0] u_ca_in_514;
wire [5:0] u_ca_in_515;
wire [5:0] u_ca_in_516;
wire [5:0] u_ca_in_517;
wire [5:0] u_ca_in_518;
wire [5:0] u_ca_in_519;
wire [5:0] u_ca_in_520;
wire [5:0] u_ca_in_521;
wire [5:0] u_ca_in_522;
wire [5:0] u_ca_in_523;
wire [5:0] u_ca_in_524;
wire [5:0] u_ca_in_525;
wire [5:0] u_ca_in_526;
wire [5:0] u_ca_in_527;
wire [5:0] u_ca_in_528;
wire [5:0] u_ca_in_529;
wire [5:0] u_ca_in_530;
wire [5:0] u_ca_in_531;
wire [5:0] u_ca_in_532;
wire [5:0] u_ca_in_533;
wire [5:0] u_ca_in_534;
wire [5:0] u_ca_in_535;
wire [5:0] u_ca_in_536;
wire [5:0] u_ca_in_537;
wire [5:0] u_ca_in_538;
wire [5:0] u_ca_in_539;
wire [5:0] u_ca_in_540;
wire [5:0] u_ca_in_541;
wire [5:0] u_ca_in_542;
wire [5:0] u_ca_in_543;
wire [5:0] u_ca_in_544;
wire [5:0] u_ca_in_545;
wire [5:0] u_ca_in_546;
wire [5:0] u_ca_in_547;
wire [5:0] u_ca_in_548;
wire [5:0] u_ca_in_549;
wire [5:0] u_ca_in_550;
wire [5:0] u_ca_in_551;
wire [5:0] u_ca_in_552;
wire [5:0] u_ca_in_553;
wire [5:0] u_ca_in_554;
wire [5:0] u_ca_in_555;
wire [5:0] u_ca_in_556;
wire [5:0] u_ca_in_557;
wire [5:0] u_ca_in_558;
wire [5:0] u_ca_in_559;
wire [5:0] u_ca_in_560;
wire [5:0] u_ca_in_561;
wire [5:0] u_ca_in_562;
wire [5:0] u_ca_in_563;
wire [5:0] u_ca_in_564;
wire [5:0] u_ca_in_565;
wire [5:0] u_ca_in_566;
wire [5:0] u_ca_in_567;
wire [5:0] u_ca_in_568;
wire [5:0] u_ca_in_569;
wire [5:0] u_ca_in_570;
wire [5:0] u_ca_in_571;
wire [5:0] u_ca_in_572;
wire [5:0] u_ca_in_573;
wire [5:0] u_ca_in_574;
wire [5:0] u_ca_in_575;
wire [5:0] u_ca_in_576;
wire [5:0] u_ca_in_577;
wire [5:0] u_ca_in_578;
wire [5:0] u_ca_in_579;
wire [5:0] u_ca_in_580;
wire [5:0] u_ca_in_581;
wire [5:0] u_ca_in_582;
wire [5:0] u_ca_in_583;
wire [5:0] u_ca_in_584;
wire [5:0] u_ca_in_585;
wire [5:0] u_ca_in_586;
wire [5:0] u_ca_in_587;
wire [5:0] u_ca_in_588;
wire [5:0] u_ca_in_589;
wire [5:0] u_ca_in_590;
wire [5:0] u_ca_in_591;
wire [5:0] u_ca_in_592;
wire [5:0] u_ca_in_593;
wire [5:0] u_ca_in_594;
wire [5:0] u_ca_in_595;
wire [5:0] u_ca_in_596;
wire [5:0] u_ca_in_597;
wire [5:0] u_ca_in_598;
wire [5:0] u_ca_in_599;
wire [5:0] u_ca_in_600;
wire [5:0] u_ca_in_601;
wire [5:0] u_ca_in_602;
wire [5:0] u_ca_in_603;
wire [5:0] u_ca_in_604;
wire [5:0] u_ca_in_605;
wire [5:0] u_ca_in_606;
wire [5:0] u_ca_in_607;
wire [5:0] u_ca_in_608;
wire [5:0] u_ca_in_609;
wire [5:0] u_ca_in_610;
wire [5:0] u_ca_in_611;
wire [5:0] u_ca_in_612;
wire [5:0] u_ca_in_613;
wire [5:0] u_ca_in_614;
wire [5:0] u_ca_in_615;
wire [5:0] u_ca_in_616;
wire [5:0] u_ca_in_617;
wire [5:0] u_ca_in_618;
wire [5:0] u_ca_in_619;
wire [5:0] u_ca_in_620;
wire [5:0] u_ca_in_621;
wire [5:0] u_ca_in_622;
wire [5:0] u_ca_in_623;
wire [5:0] u_ca_in_624;
wire [5:0] u_ca_in_625;
wire [5:0] u_ca_in_626;
wire [5:0] u_ca_in_627;
wire [5:0] u_ca_in_628;
wire [5:0] u_ca_in_629;
wire [5:0] u_ca_in_630;
wire [5:0] u_ca_in_631;
wire [5:0] u_ca_in_632;
wire [5:0] u_ca_in_633;
wire [5:0] u_ca_in_634;
wire [5:0] u_ca_in_635;
wire [5:0] u_ca_in_636;
wire [5:0] u_ca_in_637;
wire [5:0] u_ca_in_638;
wire [5:0] u_ca_in_639;
wire [5:0] u_ca_in_640;
wire [5:0] u_ca_in_641;
wire [5:0] u_ca_in_642;
wire [5:0] u_ca_in_643;
wire [5:0] u_ca_in_644;
wire [5:0] u_ca_in_645;
wire [5:0] u_ca_in_646;
wire [5:0] u_ca_in_647;
wire [5:0] u_ca_in_648;
wire [5:0] u_ca_in_649;
wire [5:0] u_ca_in_650;
wire [5:0] u_ca_in_651;
wire [5:0] u_ca_in_652;
wire [5:0] u_ca_in_653;
wire [5:0] u_ca_in_654;
wire [5:0] u_ca_in_655;
wire [5:0] u_ca_in_656;
wire [5:0] u_ca_in_657;
wire [5:0] u_ca_in_658;
wire [5:0] u_ca_in_659;
wire [5:0] u_ca_in_660;
wire [5:0] u_ca_in_661;
wire [5:0] u_ca_in_662;
wire [5:0] u_ca_in_663;
wire [5:0] u_ca_in_664;
wire [5:0] u_ca_in_665;
wire [5:0] u_ca_in_666;
wire [5:0] u_ca_in_667;
wire [5:0] u_ca_in_668;
wire [5:0] u_ca_in_669;
wire [5:0] u_ca_in_670;
wire [5:0] u_ca_in_671;
wire [5:0] u_ca_in_672;
wire [5:0] u_ca_in_673;
wire [5:0] u_ca_in_674;
wire [5:0] u_ca_in_675;
wire [5:0] u_ca_in_676;
wire [5:0] u_ca_in_677;
wire [5:0] u_ca_in_678;
wire [5:0] u_ca_in_679;
wire [5:0] u_ca_in_680;
wire [5:0] u_ca_in_681;
wire [5:0] u_ca_in_682;
wire [5:0] u_ca_in_683;
wire [5:0] u_ca_in_684;
wire [5:0] u_ca_in_685;
wire [5:0] u_ca_in_686;
wire [5:0] u_ca_in_687;
wire [5:0] u_ca_in_688;
wire [5:0] u_ca_in_689;
wire [5:0] u_ca_in_690;
wire [5:0] u_ca_in_691;
wire [5:0] u_ca_in_692;
wire [5:0] u_ca_in_693;
wire [5:0] u_ca_in_694;
wire [5:0] u_ca_in_695;
wire [5:0] u_ca_in_696;
wire [5:0] u_ca_in_697;
wire [5:0] u_ca_in_698;
wire [5:0] u_ca_in_699;
wire [5:0] u_ca_in_700;
wire [5:0] u_ca_in_701;
wire [5:0] u_ca_in_702;
wire [5:0] u_ca_in_703;
wire [5:0] u_ca_in_704;
wire [5:0] u_ca_in_705;
wire [5:0] u_ca_in_706;
wire [5:0] u_ca_in_707;
wire [5:0] u_ca_in_708;
wire [5:0] u_ca_in_709;
wire [5:0] u_ca_in_710;
wire [5:0] u_ca_in_711;
wire [5:0] u_ca_in_712;
wire [5:0] u_ca_in_713;
wire [5:0] u_ca_in_714;
wire [5:0] u_ca_in_715;
wire [5:0] u_ca_in_716;
wire [5:0] u_ca_in_717;
wire [5:0] u_ca_in_718;
wire [5:0] u_ca_in_719;
wire [5:0] u_ca_in_720;
wire [5:0] u_ca_in_721;
wire [5:0] u_ca_in_722;
wire [5:0] u_ca_in_723;
wire [5:0] u_ca_in_724;
wire [5:0] u_ca_in_725;
wire [5:0] u_ca_in_726;
wire [5:0] u_ca_in_727;
wire [5:0] u_ca_in_728;
wire [5:0] u_ca_in_729;
wire [5:0] u_ca_in_730;
wire [5:0] u_ca_in_731;
wire [5:0] u_ca_in_732;
wire [5:0] u_ca_in_733;
wire [5:0] u_ca_in_734;
wire [5:0] u_ca_in_735;
wire [5:0] u_ca_in_736;
wire [5:0] u_ca_in_737;
wire [5:0] u_ca_in_738;
wire [5:0] u_ca_in_739;
wire [5:0] u_ca_in_740;
wire [5:0] u_ca_in_741;
wire [5:0] u_ca_in_742;
wire [5:0] u_ca_in_743;
wire [5:0] u_ca_in_744;
wire [5:0] u_ca_in_745;
wire [5:0] u_ca_in_746;
wire [5:0] u_ca_in_747;
wire [5:0] u_ca_in_748;
wire [5:0] u_ca_in_749;
wire [5:0] u_ca_in_750;
wire [5:0] u_ca_in_751;
wire [5:0] u_ca_in_752;
wire [5:0] u_ca_in_753;
wire [5:0] u_ca_in_754;
wire [5:0] u_ca_in_755;
wire [5:0] u_ca_in_756;
wire [5:0] u_ca_in_757;
wire [5:0] u_ca_in_758;
wire [5:0] u_ca_in_759;
wire [5:0] u_ca_in_760;
wire [5:0] u_ca_in_761;
wire [5:0] u_ca_in_762;
wire [5:0] u_ca_in_763;
wire [5:0] u_ca_in_764;
wire [5:0] u_ca_in_765;
wire [5:0] u_ca_in_766;
wire [5:0] u_ca_in_767;
wire [5:0] u_ca_in_768;
wire [5:0] u_ca_in_769;
wire [5:0] u_ca_in_770;
wire [5:0] u_ca_in_771;
wire [5:0] u_ca_in_772;
wire [5:0] u_ca_in_773;
wire [5:0] u_ca_in_774;
wire [5:0] u_ca_in_775;
wire [5:0] u_ca_in_776;
wire [5:0] u_ca_in_777;
wire [5:0] u_ca_in_778;
wire [5:0] u_ca_in_779;
wire [5:0] u_ca_in_780;
wire [5:0] u_ca_in_781;
wire [5:0] u_ca_in_782;
wire [5:0] u_ca_in_783;
wire [5:0] u_ca_in_784;
wire [5:0] u_ca_in_785;
wire [5:0] u_ca_in_786;
wire [5:0] u_ca_in_787;
wire [5:0] u_ca_in_788;
wire [5:0] u_ca_in_789;
wire [5:0] u_ca_in_790;
wire [5:0] u_ca_in_791;
wire [5:0] u_ca_in_792;
wire [5:0] u_ca_in_793;
wire [5:0] u_ca_in_794;
wire [5:0] u_ca_in_795;
wire [5:0] u_ca_in_796;
wire [5:0] u_ca_in_797;
wire [5:0] u_ca_in_798;
wire [5:0] u_ca_in_799;
wire [5:0] u_ca_in_800;
wire [5:0] u_ca_in_801;
wire [5:0] u_ca_in_802;
wire [5:0] u_ca_in_803;
wire [5:0] u_ca_in_804;
wire [5:0] u_ca_in_805;
wire [5:0] u_ca_in_806;
wire [5:0] u_ca_in_807;
wire [5:0] u_ca_in_808;
wire [5:0] u_ca_in_809;
wire [5:0] u_ca_in_810;
wire [5:0] u_ca_in_811;
wire [5:0] u_ca_in_812;
wire [5:0] u_ca_in_813;
wire [5:0] u_ca_in_814;
wire [5:0] u_ca_in_815;
wire [5:0] u_ca_in_816;
wire [5:0] u_ca_in_817;
wire [5:0] u_ca_in_818;
wire [5:0] u_ca_in_819;
wire [5:0] u_ca_in_820;
wire [5:0] u_ca_in_821;
wire [5:0] u_ca_in_822;
wire [5:0] u_ca_in_823;
wire [5:0] u_ca_in_824;
wire [5:0] u_ca_in_825;
wire [5:0] u_ca_in_826;
wire [5:0] u_ca_in_827;
wire [5:0] u_ca_in_828;
wire [5:0] u_ca_in_829;
wire [5:0] u_ca_in_830;
wire [5:0] u_ca_in_831;
wire [5:0] u_ca_in_832;
wire [5:0] u_ca_in_833;
wire [5:0] u_ca_in_834;
wire [5:0] u_ca_in_835;
wire [5:0] u_ca_in_836;
wire [5:0] u_ca_in_837;
wire [5:0] u_ca_in_838;
wire [5:0] u_ca_in_839;
wire [5:0] u_ca_in_840;
wire [5:0] u_ca_in_841;
wire [5:0] u_ca_in_842;
wire [5:0] u_ca_in_843;
wire [5:0] u_ca_in_844;
wire [5:0] u_ca_in_845;
wire [5:0] u_ca_in_846;
wire [5:0] u_ca_in_847;
wire [5:0] u_ca_in_848;
wire [5:0] u_ca_in_849;
wire [5:0] u_ca_in_850;
wire [5:0] u_ca_in_851;
wire [5:0] u_ca_in_852;
wire [5:0] u_ca_in_853;
wire [5:0] u_ca_in_854;
wire [5:0] u_ca_in_855;
wire [5:0] u_ca_in_856;
wire [5:0] u_ca_in_857;
wire [5:0] u_ca_in_858;
wire [5:0] u_ca_in_859;
wire [5:0] u_ca_in_860;
wire [5:0] u_ca_in_861;
wire [5:0] u_ca_in_862;
wire [5:0] u_ca_in_863;
wire [5:0] u_ca_in_864;
wire [5:0] u_ca_in_865;
wire [5:0] u_ca_in_866;
wire [5:0] u_ca_in_867;
wire [5:0] u_ca_in_868;
wire [5:0] u_ca_in_869;
wire [5:0] u_ca_in_870;
wire [5:0] u_ca_in_871;
wire [5:0] u_ca_in_872;
wire [5:0] u_ca_in_873;
wire [5:0] u_ca_in_874;
wire [5:0] u_ca_in_875;
wire [5:0] u_ca_in_876;
wire [5:0] u_ca_in_877;
wire [5:0] u_ca_in_878;
wire [5:0] u_ca_in_879;
wire [5:0] u_ca_in_880;
wire [5:0] u_ca_in_881;
wire [5:0] u_ca_in_882;
wire [5:0] u_ca_in_883;
wire [5:0] u_ca_in_884;
wire [5:0] u_ca_in_885;
wire [5:0] u_ca_in_886;
wire [5:0] u_ca_in_887;
wire [5:0] u_ca_in_888;
wire [5:0] u_ca_in_889;
wire [5:0] u_ca_in_890;
wire [5:0] u_ca_in_891;
wire [5:0] u_ca_in_892;
wire [5:0] u_ca_in_893;
wire [5:0] u_ca_in_894;
wire [5:0] u_ca_in_895;
wire [5:0] u_ca_in_896;
wire [5:0] u_ca_in_897;
wire [5:0] u_ca_in_898;
wire [5:0] u_ca_in_899;
wire [5:0] u_ca_in_900;
wire [5:0] u_ca_in_901;
wire [5:0] u_ca_in_902;
wire [5:0] u_ca_in_903;
wire [5:0] u_ca_in_904;
wire [5:0] u_ca_in_905;
wire [5:0] u_ca_in_906;
wire [5:0] u_ca_in_907;
wire [5:0] u_ca_in_908;
wire [5:0] u_ca_in_909;
wire [5:0] u_ca_in_910;
wire [5:0] u_ca_in_911;
wire [5:0] u_ca_in_912;
wire [5:0] u_ca_in_913;
wire [5:0] u_ca_in_914;
wire [5:0] u_ca_in_915;
wire [5:0] u_ca_in_916;
wire [5:0] u_ca_in_917;
wire [5:0] u_ca_in_918;
wire [5:0] u_ca_in_919;
wire [5:0] u_ca_in_920;
wire [5:0] u_ca_in_921;
wire [5:0] u_ca_in_922;
wire [5:0] u_ca_in_923;
wire [5:0] u_ca_in_924;
wire [5:0] u_ca_in_925;
wire [5:0] u_ca_in_926;
wire [5:0] u_ca_in_927;
wire [5:0] u_ca_in_928;
wire [5:0] u_ca_in_929;
wire [5:0] u_ca_in_930;
wire [5:0] u_ca_in_931;
wire [5:0] u_ca_in_932;
wire [5:0] u_ca_in_933;
wire [5:0] u_ca_in_934;
wire [5:0] u_ca_in_935;
wire [5:0] u_ca_in_936;
wire [5:0] u_ca_in_937;
wire [5:0] u_ca_in_938;
wire [5:0] u_ca_in_939;
wire [5:0] u_ca_in_940;
wire [5:0] u_ca_in_941;
wire [5:0] u_ca_in_942;
wire [5:0] u_ca_in_943;
wire [5:0] u_ca_in_944;
wire [5:0] u_ca_in_945;
wire [5:0] u_ca_in_946;
wire [5:0] u_ca_in_947;
wire [5:0] u_ca_in_948;
wire [5:0] u_ca_in_949;
wire [5:0] u_ca_in_950;
wire [5:0] u_ca_in_951;
wire [5:0] u_ca_in_952;
wire [5:0] u_ca_in_953;
wire [5:0] u_ca_in_954;
wire [5:0] u_ca_in_955;
wire [5:0] u_ca_in_956;
wire [5:0] u_ca_in_957;
wire [5:0] u_ca_in_958;
wire [5:0] u_ca_in_959;
wire [5:0] u_ca_in_960;
wire [5:0] u_ca_in_961;
wire [5:0] u_ca_in_962;
wire [5:0] u_ca_in_963;
wire [5:0] u_ca_in_964;
wire [5:0] u_ca_in_965;
wire [5:0] u_ca_in_966;
wire [5:0] u_ca_in_967;
wire [5:0] u_ca_in_968;
wire [5:0] u_ca_in_969;
wire [5:0] u_ca_in_970;
wire [5:0] u_ca_in_971;
wire [5:0] u_ca_in_972;
wire [5:0] u_ca_in_973;
wire [5:0] u_ca_in_974;
wire [5:0] u_ca_in_975;
wire [5:0] u_ca_in_976;
wire [5:0] u_ca_in_977;
wire [5:0] u_ca_in_978;
wire [5:0] u_ca_in_979;
wire [5:0] u_ca_in_980;
wire [5:0] u_ca_in_981;
wire [5:0] u_ca_in_982;
wire [5:0] u_ca_in_983;
wire [5:0] u_ca_in_984;
wire [5:0] u_ca_in_985;
wire [5:0] u_ca_in_986;
wire [5:0] u_ca_in_987;
wire [5:0] u_ca_in_988;
wire [5:0] u_ca_in_989;
wire [5:0] u_ca_in_990;
wire [5:0] u_ca_in_991;
wire [5:0] u_ca_in_992;
wire [5:0] u_ca_in_993;
wire [5:0] u_ca_in_994;
wire [5:0] u_ca_in_995;
wire [5:0] u_ca_in_996;
wire [5:0] u_ca_in_997;
wire [5:0] u_ca_in_998;
wire [5:0] u_ca_in_999;
wire [5:0] u_ca_in_1000;
wire [5:0] u_ca_in_1001;
wire [5:0] u_ca_in_1002;
wire [5:0] u_ca_in_1003;
wire [5:0] u_ca_in_1004;
wire [5:0] u_ca_in_1005;
wire [5:0] u_ca_in_1006;
wire [5:0] u_ca_in_1007;
wire [5:0] u_ca_in_1008;
wire [5:0] u_ca_in_1009;
wire [5:0] u_ca_in_1010;
wire [5:0] u_ca_in_1011;
wire [5:0] u_ca_in_1012;
wire [5:0] u_ca_in_1013;
wire [5:0] u_ca_in_1014;
wire [5:0] u_ca_in_1015;
wire [5:0] u_ca_in_1016;
wire [5:0] u_ca_in_1017;
wire [5:0] u_ca_in_1018;
wire [5:0] u_ca_in_1019;
wire [5:0] u_ca_in_1020;
wire [5:0] u_ca_in_1021;
wire [5:0] u_ca_in_1022;
wire [5:0] u_ca_in_1023;
wire [3:0] u_ca_out_0;
wire [3:0] u_ca_out_1;
wire [3:0] u_ca_out_2;
wire [3:0] u_ca_out_3;
wire [3:0] u_ca_out_4;
wire [3:0] u_ca_out_5;
wire [3:0] u_ca_out_6;
wire [3:0] u_ca_out_7;
wire [3:0] u_ca_out_8;
wire [3:0] u_ca_out_9;
wire [3:0] u_ca_out_10;
wire [3:0] u_ca_out_11;
wire [3:0] u_ca_out_12;
wire [3:0] u_ca_out_13;
wire [3:0] u_ca_out_14;
wire [3:0] u_ca_out_15;
wire [3:0] u_ca_out_16;
wire [3:0] u_ca_out_17;
wire [3:0] u_ca_out_18;
wire [3:0] u_ca_out_19;
wire [3:0] u_ca_out_20;
wire [3:0] u_ca_out_21;
wire [3:0] u_ca_out_22;
wire [3:0] u_ca_out_23;
wire [3:0] u_ca_out_24;
wire [3:0] u_ca_out_25;
wire [3:0] u_ca_out_26;
wire [3:0] u_ca_out_27;
wire [3:0] u_ca_out_28;
wire [3:0] u_ca_out_29;
wire [3:0] u_ca_out_30;
wire [3:0] u_ca_out_31;
wire [3:0] u_ca_out_32;
wire [3:0] u_ca_out_33;
wire [3:0] u_ca_out_34;
wire [3:0] u_ca_out_35;
wire [3:0] u_ca_out_36;
wire [3:0] u_ca_out_37;
wire [3:0] u_ca_out_38;
wire [3:0] u_ca_out_39;
wire [3:0] u_ca_out_40;
wire [3:0] u_ca_out_41;
wire [3:0] u_ca_out_42;
wire [3:0] u_ca_out_43;
wire [3:0] u_ca_out_44;
wire [3:0] u_ca_out_45;
wire [3:0] u_ca_out_46;
wire [3:0] u_ca_out_47;
wire [3:0] u_ca_out_48;
wire [3:0] u_ca_out_49;
wire [3:0] u_ca_out_50;
wire [3:0] u_ca_out_51;
wire [3:0] u_ca_out_52;
wire [3:0] u_ca_out_53;
wire [3:0] u_ca_out_54;
wire [3:0] u_ca_out_55;
wire [3:0] u_ca_out_56;
wire [3:0] u_ca_out_57;
wire [3:0] u_ca_out_58;
wire [3:0] u_ca_out_59;
wire [3:0] u_ca_out_60;
wire [3:0] u_ca_out_61;
wire [3:0] u_ca_out_62;
wire [3:0] u_ca_out_63;
wire [3:0] u_ca_out_64;
wire [3:0] u_ca_out_65;
wire [3:0] u_ca_out_66;
wire [3:0] u_ca_out_67;
wire [3:0] u_ca_out_68;
wire [3:0] u_ca_out_69;
wire [3:0] u_ca_out_70;
wire [3:0] u_ca_out_71;
wire [3:0] u_ca_out_72;
wire [3:0] u_ca_out_73;
wire [3:0] u_ca_out_74;
wire [3:0] u_ca_out_75;
wire [3:0] u_ca_out_76;
wire [3:0] u_ca_out_77;
wire [3:0] u_ca_out_78;
wire [3:0] u_ca_out_79;
wire [3:0] u_ca_out_80;
wire [3:0] u_ca_out_81;
wire [3:0] u_ca_out_82;
wire [3:0] u_ca_out_83;
wire [3:0] u_ca_out_84;
wire [3:0] u_ca_out_85;
wire [3:0] u_ca_out_86;
wire [3:0] u_ca_out_87;
wire [3:0] u_ca_out_88;
wire [3:0] u_ca_out_89;
wire [3:0] u_ca_out_90;
wire [3:0] u_ca_out_91;
wire [3:0] u_ca_out_92;
wire [3:0] u_ca_out_93;
wire [3:0] u_ca_out_94;
wire [3:0] u_ca_out_95;
wire [3:0] u_ca_out_96;
wire [3:0] u_ca_out_97;
wire [3:0] u_ca_out_98;
wire [3:0] u_ca_out_99;
wire [3:0] u_ca_out_100;
wire [3:0] u_ca_out_101;
wire [3:0] u_ca_out_102;
wire [3:0] u_ca_out_103;
wire [3:0] u_ca_out_104;
wire [3:0] u_ca_out_105;
wire [3:0] u_ca_out_106;
wire [3:0] u_ca_out_107;
wire [3:0] u_ca_out_108;
wire [3:0] u_ca_out_109;
wire [3:0] u_ca_out_110;
wire [3:0] u_ca_out_111;
wire [3:0] u_ca_out_112;
wire [3:0] u_ca_out_113;
wire [3:0] u_ca_out_114;
wire [3:0] u_ca_out_115;
wire [3:0] u_ca_out_116;
wire [3:0] u_ca_out_117;
wire [3:0] u_ca_out_118;
wire [3:0] u_ca_out_119;
wire [3:0] u_ca_out_120;
wire [3:0] u_ca_out_121;
wire [3:0] u_ca_out_122;
wire [3:0] u_ca_out_123;
wire [3:0] u_ca_out_124;
wire [3:0] u_ca_out_125;
wire [3:0] u_ca_out_126;
wire [3:0] u_ca_out_127;
wire [3:0] u_ca_out_128;
wire [3:0] u_ca_out_129;
wire [3:0] u_ca_out_130;
wire [3:0] u_ca_out_131;
wire [3:0] u_ca_out_132;
wire [3:0] u_ca_out_133;
wire [3:0] u_ca_out_134;
wire [3:0] u_ca_out_135;
wire [3:0] u_ca_out_136;
wire [3:0] u_ca_out_137;
wire [3:0] u_ca_out_138;
wire [3:0] u_ca_out_139;
wire [3:0] u_ca_out_140;
wire [3:0] u_ca_out_141;
wire [3:0] u_ca_out_142;
wire [3:0] u_ca_out_143;
wire [3:0] u_ca_out_144;
wire [3:0] u_ca_out_145;
wire [3:0] u_ca_out_146;
wire [3:0] u_ca_out_147;
wire [3:0] u_ca_out_148;
wire [3:0] u_ca_out_149;
wire [3:0] u_ca_out_150;
wire [3:0] u_ca_out_151;
wire [3:0] u_ca_out_152;
wire [3:0] u_ca_out_153;
wire [3:0] u_ca_out_154;
wire [3:0] u_ca_out_155;
wire [3:0] u_ca_out_156;
wire [3:0] u_ca_out_157;
wire [3:0] u_ca_out_158;
wire [3:0] u_ca_out_159;
wire [3:0] u_ca_out_160;
wire [3:0] u_ca_out_161;
wire [3:0] u_ca_out_162;
wire [3:0] u_ca_out_163;
wire [3:0] u_ca_out_164;
wire [3:0] u_ca_out_165;
wire [3:0] u_ca_out_166;
wire [3:0] u_ca_out_167;
wire [3:0] u_ca_out_168;
wire [3:0] u_ca_out_169;
wire [3:0] u_ca_out_170;
wire [3:0] u_ca_out_171;
wire [3:0] u_ca_out_172;
wire [3:0] u_ca_out_173;
wire [3:0] u_ca_out_174;
wire [3:0] u_ca_out_175;
wire [3:0] u_ca_out_176;
wire [3:0] u_ca_out_177;
wire [3:0] u_ca_out_178;
wire [3:0] u_ca_out_179;
wire [3:0] u_ca_out_180;
wire [3:0] u_ca_out_181;
wire [3:0] u_ca_out_182;
wire [3:0] u_ca_out_183;
wire [3:0] u_ca_out_184;
wire [3:0] u_ca_out_185;
wire [3:0] u_ca_out_186;
wire [3:0] u_ca_out_187;
wire [3:0] u_ca_out_188;
wire [3:0] u_ca_out_189;
wire [3:0] u_ca_out_190;
wire [3:0] u_ca_out_191;
wire [3:0] u_ca_out_192;
wire [3:0] u_ca_out_193;
wire [3:0] u_ca_out_194;
wire [3:0] u_ca_out_195;
wire [3:0] u_ca_out_196;
wire [3:0] u_ca_out_197;
wire [3:0] u_ca_out_198;
wire [3:0] u_ca_out_199;
wire [3:0] u_ca_out_200;
wire [3:0] u_ca_out_201;
wire [3:0] u_ca_out_202;
wire [3:0] u_ca_out_203;
wire [3:0] u_ca_out_204;
wire [3:0] u_ca_out_205;
wire [3:0] u_ca_out_206;
wire [3:0] u_ca_out_207;
wire [3:0] u_ca_out_208;
wire [3:0] u_ca_out_209;
wire [3:0] u_ca_out_210;
wire [3:0] u_ca_out_211;
wire [3:0] u_ca_out_212;
wire [3:0] u_ca_out_213;
wire [3:0] u_ca_out_214;
wire [3:0] u_ca_out_215;
wire [3:0] u_ca_out_216;
wire [3:0] u_ca_out_217;
wire [3:0] u_ca_out_218;
wire [3:0] u_ca_out_219;
wire [3:0] u_ca_out_220;
wire [3:0] u_ca_out_221;
wire [3:0] u_ca_out_222;
wire [3:0] u_ca_out_223;
wire [3:0] u_ca_out_224;
wire [3:0] u_ca_out_225;
wire [3:0] u_ca_out_226;
wire [3:0] u_ca_out_227;
wire [3:0] u_ca_out_228;
wire [3:0] u_ca_out_229;
wire [3:0] u_ca_out_230;
wire [3:0] u_ca_out_231;
wire [3:0] u_ca_out_232;
wire [3:0] u_ca_out_233;
wire [3:0] u_ca_out_234;
wire [3:0] u_ca_out_235;
wire [3:0] u_ca_out_236;
wire [3:0] u_ca_out_237;
wire [3:0] u_ca_out_238;
wire [3:0] u_ca_out_239;
wire [3:0] u_ca_out_240;
wire [3:0] u_ca_out_241;
wire [3:0] u_ca_out_242;
wire [3:0] u_ca_out_243;
wire [3:0] u_ca_out_244;
wire [3:0] u_ca_out_245;
wire [3:0] u_ca_out_246;
wire [3:0] u_ca_out_247;
wire [3:0] u_ca_out_248;
wire [3:0] u_ca_out_249;
wire [3:0] u_ca_out_250;
wire [3:0] u_ca_out_251;
wire [3:0] u_ca_out_252;
wire [3:0] u_ca_out_253;
wire [3:0] u_ca_out_254;
wire [3:0] u_ca_out_255;
wire [3:0] u_ca_out_256;
wire [3:0] u_ca_out_257;
wire [3:0] u_ca_out_258;
wire [3:0] u_ca_out_259;
wire [3:0] u_ca_out_260;
wire [3:0] u_ca_out_261;
wire [3:0] u_ca_out_262;
wire [3:0] u_ca_out_263;
wire [3:0] u_ca_out_264;
wire [3:0] u_ca_out_265;
wire [3:0] u_ca_out_266;
wire [3:0] u_ca_out_267;
wire [3:0] u_ca_out_268;
wire [3:0] u_ca_out_269;
wire [3:0] u_ca_out_270;
wire [3:0] u_ca_out_271;
wire [3:0] u_ca_out_272;
wire [3:0] u_ca_out_273;
wire [3:0] u_ca_out_274;
wire [3:0] u_ca_out_275;
wire [3:0] u_ca_out_276;
wire [3:0] u_ca_out_277;
wire [3:0] u_ca_out_278;
wire [3:0] u_ca_out_279;
wire [3:0] u_ca_out_280;
wire [3:0] u_ca_out_281;
wire [3:0] u_ca_out_282;
wire [3:0] u_ca_out_283;
wire [3:0] u_ca_out_284;
wire [3:0] u_ca_out_285;
wire [3:0] u_ca_out_286;
wire [3:0] u_ca_out_287;
wire [3:0] u_ca_out_288;
wire [3:0] u_ca_out_289;
wire [3:0] u_ca_out_290;
wire [3:0] u_ca_out_291;
wire [3:0] u_ca_out_292;
wire [3:0] u_ca_out_293;
wire [3:0] u_ca_out_294;
wire [3:0] u_ca_out_295;
wire [3:0] u_ca_out_296;
wire [3:0] u_ca_out_297;
wire [3:0] u_ca_out_298;
wire [3:0] u_ca_out_299;
wire [3:0] u_ca_out_300;
wire [3:0] u_ca_out_301;
wire [3:0] u_ca_out_302;
wire [3:0] u_ca_out_303;
wire [3:0] u_ca_out_304;
wire [3:0] u_ca_out_305;
wire [3:0] u_ca_out_306;
wire [3:0] u_ca_out_307;
wire [3:0] u_ca_out_308;
wire [3:0] u_ca_out_309;
wire [3:0] u_ca_out_310;
wire [3:0] u_ca_out_311;
wire [3:0] u_ca_out_312;
wire [3:0] u_ca_out_313;
wire [3:0] u_ca_out_314;
wire [3:0] u_ca_out_315;
wire [3:0] u_ca_out_316;
wire [3:0] u_ca_out_317;
wire [3:0] u_ca_out_318;
wire [3:0] u_ca_out_319;
wire [3:0] u_ca_out_320;
wire [3:0] u_ca_out_321;
wire [3:0] u_ca_out_322;
wire [3:0] u_ca_out_323;
wire [3:0] u_ca_out_324;
wire [3:0] u_ca_out_325;
wire [3:0] u_ca_out_326;
wire [3:0] u_ca_out_327;
wire [3:0] u_ca_out_328;
wire [3:0] u_ca_out_329;
wire [3:0] u_ca_out_330;
wire [3:0] u_ca_out_331;
wire [3:0] u_ca_out_332;
wire [3:0] u_ca_out_333;
wire [3:0] u_ca_out_334;
wire [3:0] u_ca_out_335;
wire [3:0] u_ca_out_336;
wire [3:0] u_ca_out_337;
wire [3:0] u_ca_out_338;
wire [3:0] u_ca_out_339;
wire [3:0] u_ca_out_340;
wire [3:0] u_ca_out_341;
wire [3:0] u_ca_out_342;
wire [3:0] u_ca_out_343;
wire [3:0] u_ca_out_344;
wire [3:0] u_ca_out_345;
wire [3:0] u_ca_out_346;
wire [3:0] u_ca_out_347;
wire [3:0] u_ca_out_348;
wire [3:0] u_ca_out_349;
wire [3:0] u_ca_out_350;
wire [3:0] u_ca_out_351;
wire [3:0] u_ca_out_352;
wire [3:0] u_ca_out_353;
wire [3:0] u_ca_out_354;
wire [3:0] u_ca_out_355;
wire [3:0] u_ca_out_356;
wire [3:0] u_ca_out_357;
wire [3:0] u_ca_out_358;
wire [3:0] u_ca_out_359;
wire [3:0] u_ca_out_360;
wire [3:0] u_ca_out_361;
wire [3:0] u_ca_out_362;
wire [3:0] u_ca_out_363;
wire [3:0] u_ca_out_364;
wire [3:0] u_ca_out_365;
wire [3:0] u_ca_out_366;
wire [3:0] u_ca_out_367;
wire [3:0] u_ca_out_368;
wire [3:0] u_ca_out_369;
wire [3:0] u_ca_out_370;
wire [3:0] u_ca_out_371;
wire [3:0] u_ca_out_372;
wire [3:0] u_ca_out_373;
wire [3:0] u_ca_out_374;
wire [3:0] u_ca_out_375;
wire [3:0] u_ca_out_376;
wire [3:0] u_ca_out_377;
wire [3:0] u_ca_out_378;
wire [3:0] u_ca_out_379;
wire [3:0] u_ca_out_380;
wire [3:0] u_ca_out_381;
wire [3:0] u_ca_out_382;
wire [3:0] u_ca_out_383;
wire [3:0] u_ca_out_384;
wire [3:0] u_ca_out_385;
wire [3:0] u_ca_out_386;
wire [3:0] u_ca_out_387;
wire [3:0] u_ca_out_388;
wire [3:0] u_ca_out_389;
wire [3:0] u_ca_out_390;
wire [3:0] u_ca_out_391;
wire [3:0] u_ca_out_392;
wire [3:0] u_ca_out_393;
wire [3:0] u_ca_out_394;
wire [3:0] u_ca_out_395;
wire [3:0] u_ca_out_396;
wire [3:0] u_ca_out_397;
wire [3:0] u_ca_out_398;
wire [3:0] u_ca_out_399;
wire [3:0] u_ca_out_400;
wire [3:0] u_ca_out_401;
wire [3:0] u_ca_out_402;
wire [3:0] u_ca_out_403;
wire [3:0] u_ca_out_404;
wire [3:0] u_ca_out_405;
wire [3:0] u_ca_out_406;
wire [3:0] u_ca_out_407;
wire [3:0] u_ca_out_408;
wire [3:0] u_ca_out_409;
wire [3:0] u_ca_out_410;
wire [3:0] u_ca_out_411;
wire [3:0] u_ca_out_412;
wire [3:0] u_ca_out_413;
wire [3:0] u_ca_out_414;
wire [3:0] u_ca_out_415;
wire [3:0] u_ca_out_416;
wire [3:0] u_ca_out_417;
wire [3:0] u_ca_out_418;
wire [3:0] u_ca_out_419;
wire [3:0] u_ca_out_420;
wire [3:0] u_ca_out_421;
wire [3:0] u_ca_out_422;
wire [3:0] u_ca_out_423;
wire [3:0] u_ca_out_424;
wire [3:0] u_ca_out_425;
wire [3:0] u_ca_out_426;
wire [3:0] u_ca_out_427;
wire [3:0] u_ca_out_428;
wire [3:0] u_ca_out_429;
wire [3:0] u_ca_out_430;
wire [3:0] u_ca_out_431;
wire [3:0] u_ca_out_432;
wire [3:0] u_ca_out_433;
wire [3:0] u_ca_out_434;
wire [3:0] u_ca_out_435;
wire [3:0] u_ca_out_436;
wire [3:0] u_ca_out_437;
wire [3:0] u_ca_out_438;
wire [3:0] u_ca_out_439;
wire [3:0] u_ca_out_440;
wire [3:0] u_ca_out_441;
wire [3:0] u_ca_out_442;
wire [3:0] u_ca_out_443;
wire [3:0] u_ca_out_444;
wire [3:0] u_ca_out_445;
wire [3:0] u_ca_out_446;
wire [3:0] u_ca_out_447;
wire [3:0] u_ca_out_448;
wire [3:0] u_ca_out_449;
wire [3:0] u_ca_out_450;
wire [3:0] u_ca_out_451;
wire [3:0] u_ca_out_452;
wire [3:0] u_ca_out_453;
wire [3:0] u_ca_out_454;
wire [3:0] u_ca_out_455;
wire [3:0] u_ca_out_456;
wire [3:0] u_ca_out_457;
wire [3:0] u_ca_out_458;
wire [3:0] u_ca_out_459;
wire [3:0] u_ca_out_460;
wire [3:0] u_ca_out_461;
wire [3:0] u_ca_out_462;
wire [3:0] u_ca_out_463;
wire [3:0] u_ca_out_464;
wire [3:0] u_ca_out_465;
wire [3:0] u_ca_out_466;
wire [3:0] u_ca_out_467;
wire [3:0] u_ca_out_468;
wire [3:0] u_ca_out_469;
wire [3:0] u_ca_out_470;
wire [3:0] u_ca_out_471;
wire [3:0] u_ca_out_472;
wire [3:0] u_ca_out_473;
wire [3:0] u_ca_out_474;
wire [3:0] u_ca_out_475;
wire [3:0] u_ca_out_476;
wire [3:0] u_ca_out_477;
wire [3:0] u_ca_out_478;
wire [3:0] u_ca_out_479;
wire [3:0] u_ca_out_480;
wire [3:0] u_ca_out_481;
wire [3:0] u_ca_out_482;
wire [3:0] u_ca_out_483;
wire [3:0] u_ca_out_484;
wire [3:0] u_ca_out_485;
wire [3:0] u_ca_out_486;
wire [3:0] u_ca_out_487;
wire [3:0] u_ca_out_488;
wire [3:0] u_ca_out_489;
wire [3:0] u_ca_out_490;
wire [3:0] u_ca_out_491;
wire [3:0] u_ca_out_492;
wire [3:0] u_ca_out_493;
wire [3:0] u_ca_out_494;
wire [3:0] u_ca_out_495;
wire [3:0] u_ca_out_496;
wire [3:0] u_ca_out_497;
wire [3:0] u_ca_out_498;
wire [3:0] u_ca_out_499;
wire [3:0] u_ca_out_500;
wire [3:0] u_ca_out_501;
wire [3:0] u_ca_out_502;
wire [3:0] u_ca_out_503;
wire [3:0] u_ca_out_504;
wire [3:0] u_ca_out_505;
wire [3:0] u_ca_out_506;
wire [3:0] u_ca_out_507;
wire [3:0] u_ca_out_508;
wire [3:0] u_ca_out_509;
wire [3:0] u_ca_out_510;
wire [3:0] u_ca_out_511;
wire [3:0] u_ca_out_512;
wire [3:0] u_ca_out_513;
wire [3:0] u_ca_out_514;
wire [3:0] u_ca_out_515;
wire [3:0] u_ca_out_516;
wire [3:0] u_ca_out_517;
wire [3:0] u_ca_out_518;
wire [3:0] u_ca_out_519;
wire [3:0] u_ca_out_520;
wire [3:0] u_ca_out_521;
wire [3:0] u_ca_out_522;
wire [3:0] u_ca_out_523;
wire [3:0] u_ca_out_524;
wire [3:0] u_ca_out_525;
wire [3:0] u_ca_out_526;
wire [3:0] u_ca_out_527;
wire [3:0] u_ca_out_528;
wire [3:0] u_ca_out_529;
wire [3:0] u_ca_out_530;
wire [3:0] u_ca_out_531;
wire [3:0] u_ca_out_532;
wire [3:0] u_ca_out_533;
wire [3:0] u_ca_out_534;
wire [3:0] u_ca_out_535;
wire [3:0] u_ca_out_536;
wire [3:0] u_ca_out_537;
wire [3:0] u_ca_out_538;
wire [3:0] u_ca_out_539;
wire [3:0] u_ca_out_540;
wire [3:0] u_ca_out_541;
wire [3:0] u_ca_out_542;
wire [3:0] u_ca_out_543;
wire [3:0] u_ca_out_544;
wire [3:0] u_ca_out_545;
wire [3:0] u_ca_out_546;
wire [3:0] u_ca_out_547;
wire [3:0] u_ca_out_548;
wire [3:0] u_ca_out_549;
wire [3:0] u_ca_out_550;
wire [3:0] u_ca_out_551;
wire [3:0] u_ca_out_552;
wire [3:0] u_ca_out_553;
wire [3:0] u_ca_out_554;
wire [3:0] u_ca_out_555;
wire [3:0] u_ca_out_556;
wire [3:0] u_ca_out_557;
wire [3:0] u_ca_out_558;
wire [3:0] u_ca_out_559;
wire [3:0] u_ca_out_560;
wire [3:0] u_ca_out_561;
wire [3:0] u_ca_out_562;
wire [3:0] u_ca_out_563;
wire [3:0] u_ca_out_564;
wire [3:0] u_ca_out_565;
wire [3:0] u_ca_out_566;
wire [3:0] u_ca_out_567;
wire [3:0] u_ca_out_568;
wire [3:0] u_ca_out_569;
wire [3:0] u_ca_out_570;
wire [3:0] u_ca_out_571;
wire [3:0] u_ca_out_572;
wire [3:0] u_ca_out_573;
wire [3:0] u_ca_out_574;
wire [3:0] u_ca_out_575;
wire [3:0] u_ca_out_576;
wire [3:0] u_ca_out_577;
wire [3:0] u_ca_out_578;
wire [3:0] u_ca_out_579;
wire [3:0] u_ca_out_580;
wire [3:0] u_ca_out_581;
wire [3:0] u_ca_out_582;
wire [3:0] u_ca_out_583;
wire [3:0] u_ca_out_584;
wire [3:0] u_ca_out_585;
wire [3:0] u_ca_out_586;
wire [3:0] u_ca_out_587;
wire [3:0] u_ca_out_588;
wire [3:0] u_ca_out_589;
wire [3:0] u_ca_out_590;
wire [3:0] u_ca_out_591;
wire [3:0] u_ca_out_592;
wire [3:0] u_ca_out_593;
wire [3:0] u_ca_out_594;
wire [3:0] u_ca_out_595;
wire [3:0] u_ca_out_596;
wire [3:0] u_ca_out_597;
wire [3:0] u_ca_out_598;
wire [3:0] u_ca_out_599;
wire [3:0] u_ca_out_600;
wire [3:0] u_ca_out_601;
wire [3:0] u_ca_out_602;
wire [3:0] u_ca_out_603;
wire [3:0] u_ca_out_604;
wire [3:0] u_ca_out_605;
wire [3:0] u_ca_out_606;
wire [3:0] u_ca_out_607;
wire [3:0] u_ca_out_608;
wire [3:0] u_ca_out_609;
wire [3:0] u_ca_out_610;
wire [3:0] u_ca_out_611;
wire [3:0] u_ca_out_612;
wire [3:0] u_ca_out_613;
wire [3:0] u_ca_out_614;
wire [3:0] u_ca_out_615;
wire [3:0] u_ca_out_616;
wire [3:0] u_ca_out_617;
wire [3:0] u_ca_out_618;
wire [3:0] u_ca_out_619;
wire [3:0] u_ca_out_620;
wire [3:0] u_ca_out_621;
wire [3:0] u_ca_out_622;
wire [3:0] u_ca_out_623;
wire [3:0] u_ca_out_624;
wire [3:0] u_ca_out_625;
wire [3:0] u_ca_out_626;
wire [3:0] u_ca_out_627;
wire [3:0] u_ca_out_628;
wire [3:0] u_ca_out_629;
wire [3:0] u_ca_out_630;
wire [3:0] u_ca_out_631;
wire [3:0] u_ca_out_632;
wire [3:0] u_ca_out_633;
wire [3:0] u_ca_out_634;
wire [3:0] u_ca_out_635;
wire [3:0] u_ca_out_636;
wire [3:0] u_ca_out_637;
wire [3:0] u_ca_out_638;
wire [3:0] u_ca_out_639;
wire [3:0] u_ca_out_640;
wire [3:0] u_ca_out_641;
wire [3:0] u_ca_out_642;
wire [3:0] u_ca_out_643;
wire [3:0] u_ca_out_644;
wire [3:0] u_ca_out_645;
wire [3:0] u_ca_out_646;
wire [3:0] u_ca_out_647;
wire [3:0] u_ca_out_648;
wire [3:0] u_ca_out_649;
wire [3:0] u_ca_out_650;
wire [3:0] u_ca_out_651;
wire [3:0] u_ca_out_652;
wire [3:0] u_ca_out_653;
wire [3:0] u_ca_out_654;
wire [3:0] u_ca_out_655;
wire [3:0] u_ca_out_656;
wire [3:0] u_ca_out_657;
wire [3:0] u_ca_out_658;
wire [3:0] u_ca_out_659;
wire [3:0] u_ca_out_660;
wire [3:0] u_ca_out_661;
wire [3:0] u_ca_out_662;
wire [3:0] u_ca_out_663;
wire [3:0] u_ca_out_664;
wire [3:0] u_ca_out_665;
wire [3:0] u_ca_out_666;
wire [3:0] u_ca_out_667;
wire [3:0] u_ca_out_668;
wire [3:0] u_ca_out_669;
wire [3:0] u_ca_out_670;
wire [3:0] u_ca_out_671;
wire [3:0] u_ca_out_672;
wire [3:0] u_ca_out_673;
wire [3:0] u_ca_out_674;
wire [3:0] u_ca_out_675;
wire [3:0] u_ca_out_676;
wire [3:0] u_ca_out_677;
wire [3:0] u_ca_out_678;
wire [3:0] u_ca_out_679;
wire [3:0] u_ca_out_680;
wire [3:0] u_ca_out_681;
wire [3:0] u_ca_out_682;
wire [3:0] u_ca_out_683;
wire [3:0] u_ca_out_684;
wire [3:0] u_ca_out_685;
wire [3:0] u_ca_out_686;
wire [3:0] u_ca_out_687;
wire [3:0] u_ca_out_688;
wire [3:0] u_ca_out_689;
wire [3:0] u_ca_out_690;
wire [3:0] u_ca_out_691;
wire [3:0] u_ca_out_692;
wire [3:0] u_ca_out_693;
wire [3:0] u_ca_out_694;
wire [3:0] u_ca_out_695;
wire [3:0] u_ca_out_696;
wire [3:0] u_ca_out_697;
wire [3:0] u_ca_out_698;
wire [3:0] u_ca_out_699;
wire [3:0] u_ca_out_700;
wire [3:0] u_ca_out_701;
wire [3:0] u_ca_out_702;
wire [3:0] u_ca_out_703;
wire [3:0] u_ca_out_704;
wire [3:0] u_ca_out_705;
wire [3:0] u_ca_out_706;
wire [3:0] u_ca_out_707;
wire [3:0] u_ca_out_708;
wire [3:0] u_ca_out_709;
wire [3:0] u_ca_out_710;
wire [3:0] u_ca_out_711;
wire [3:0] u_ca_out_712;
wire [3:0] u_ca_out_713;
wire [3:0] u_ca_out_714;
wire [3:0] u_ca_out_715;
wire [3:0] u_ca_out_716;
wire [3:0] u_ca_out_717;
wire [3:0] u_ca_out_718;
wire [3:0] u_ca_out_719;
wire [3:0] u_ca_out_720;
wire [3:0] u_ca_out_721;
wire [3:0] u_ca_out_722;
wire [3:0] u_ca_out_723;
wire [3:0] u_ca_out_724;
wire [3:0] u_ca_out_725;
wire [3:0] u_ca_out_726;
wire [3:0] u_ca_out_727;
wire [3:0] u_ca_out_728;
wire [3:0] u_ca_out_729;
wire [3:0] u_ca_out_730;
wire [3:0] u_ca_out_731;
wire [3:0] u_ca_out_732;
wire [3:0] u_ca_out_733;
wire [3:0] u_ca_out_734;
wire [3:0] u_ca_out_735;
wire [3:0] u_ca_out_736;
wire [3:0] u_ca_out_737;
wire [3:0] u_ca_out_738;
wire [3:0] u_ca_out_739;
wire [3:0] u_ca_out_740;
wire [3:0] u_ca_out_741;
wire [3:0] u_ca_out_742;
wire [3:0] u_ca_out_743;
wire [3:0] u_ca_out_744;
wire [3:0] u_ca_out_745;
wire [3:0] u_ca_out_746;
wire [3:0] u_ca_out_747;
wire [3:0] u_ca_out_748;
wire [3:0] u_ca_out_749;
wire [3:0] u_ca_out_750;
wire [3:0] u_ca_out_751;
wire [3:0] u_ca_out_752;
wire [3:0] u_ca_out_753;
wire [3:0] u_ca_out_754;
wire [3:0] u_ca_out_755;
wire [3:0] u_ca_out_756;
wire [3:0] u_ca_out_757;
wire [3:0] u_ca_out_758;
wire [3:0] u_ca_out_759;
wire [3:0] u_ca_out_760;
wire [3:0] u_ca_out_761;
wire [3:0] u_ca_out_762;
wire [3:0] u_ca_out_763;
wire [3:0] u_ca_out_764;
wire [3:0] u_ca_out_765;
wire [3:0] u_ca_out_766;
wire [3:0] u_ca_out_767;
wire [3:0] u_ca_out_768;
wire [3:0] u_ca_out_769;
wire [3:0] u_ca_out_770;
wire [3:0] u_ca_out_771;
wire [3:0] u_ca_out_772;
wire [3:0] u_ca_out_773;
wire [3:0] u_ca_out_774;
wire [3:0] u_ca_out_775;
wire [3:0] u_ca_out_776;
wire [3:0] u_ca_out_777;
wire [3:0] u_ca_out_778;
wire [3:0] u_ca_out_779;
wire [3:0] u_ca_out_780;
wire [3:0] u_ca_out_781;
wire [3:0] u_ca_out_782;
wire [3:0] u_ca_out_783;
wire [3:0] u_ca_out_784;
wire [3:0] u_ca_out_785;
wire [3:0] u_ca_out_786;
wire [3:0] u_ca_out_787;
wire [3:0] u_ca_out_788;
wire [3:0] u_ca_out_789;
wire [3:0] u_ca_out_790;
wire [3:0] u_ca_out_791;
wire [3:0] u_ca_out_792;
wire [3:0] u_ca_out_793;
wire [3:0] u_ca_out_794;
wire [3:0] u_ca_out_795;
wire [3:0] u_ca_out_796;
wire [3:0] u_ca_out_797;
wire [3:0] u_ca_out_798;
wire [3:0] u_ca_out_799;
wire [3:0] u_ca_out_800;
wire [3:0] u_ca_out_801;
wire [3:0] u_ca_out_802;
wire [3:0] u_ca_out_803;
wire [3:0] u_ca_out_804;
wire [3:0] u_ca_out_805;
wire [3:0] u_ca_out_806;
wire [3:0] u_ca_out_807;
wire [3:0] u_ca_out_808;
wire [3:0] u_ca_out_809;
wire [3:0] u_ca_out_810;
wire [3:0] u_ca_out_811;
wire [3:0] u_ca_out_812;
wire [3:0] u_ca_out_813;
wire [3:0] u_ca_out_814;
wire [3:0] u_ca_out_815;
wire [3:0] u_ca_out_816;
wire [3:0] u_ca_out_817;
wire [3:0] u_ca_out_818;
wire [3:0] u_ca_out_819;
wire [3:0] u_ca_out_820;
wire [3:0] u_ca_out_821;
wire [3:0] u_ca_out_822;
wire [3:0] u_ca_out_823;
wire [3:0] u_ca_out_824;
wire [3:0] u_ca_out_825;
wire [3:0] u_ca_out_826;
wire [3:0] u_ca_out_827;
wire [3:0] u_ca_out_828;
wire [3:0] u_ca_out_829;
wire [3:0] u_ca_out_830;
wire [3:0] u_ca_out_831;
wire [3:0] u_ca_out_832;
wire [3:0] u_ca_out_833;
wire [3:0] u_ca_out_834;
wire [3:0] u_ca_out_835;
wire [3:0] u_ca_out_836;
wire [3:0] u_ca_out_837;
wire [3:0] u_ca_out_838;
wire [3:0] u_ca_out_839;
wire [3:0] u_ca_out_840;
wire [3:0] u_ca_out_841;
wire [3:0] u_ca_out_842;
wire [3:0] u_ca_out_843;
wire [3:0] u_ca_out_844;
wire [3:0] u_ca_out_845;
wire [3:0] u_ca_out_846;
wire [3:0] u_ca_out_847;
wire [3:0] u_ca_out_848;
wire [3:0] u_ca_out_849;
wire [3:0] u_ca_out_850;
wire [3:0] u_ca_out_851;
wire [3:0] u_ca_out_852;
wire [3:0] u_ca_out_853;
wire [3:0] u_ca_out_854;
wire [3:0] u_ca_out_855;
wire [3:0] u_ca_out_856;
wire [3:0] u_ca_out_857;
wire [3:0] u_ca_out_858;
wire [3:0] u_ca_out_859;
wire [3:0] u_ca_out_860;
wire [3:0] u_ca_out_861;
wire [3:0] u_ca_out_862;
wire [3:0] u_ca_out_863;
wire [3:0] u_ca_out_864;
wire [3:0] u_ca_out_865;
wire [3:0] u_ca_out_866;
wire [3:0] u_ca_out_867;
wire [3:0] u_ca_out_868;
wire [3:0] u_ca_out_869;
wire [3:0] u_ca_out_870;
wire [3:0] u_ca_out_871;
wire [3:0] u_ca_out_872;
wire [3:0] u_ca_out_873;
wire [3:0] u_ca_out_874;
wire [3:0] u_ca_out_875;
wire [3:0] u_ca_out_876;
wire [3:0] u_ca_out_877;
wire [3:0] u_ca_out_878;
wire [3:0] u_ca_out_879;
wire [3:0] u_ca_out_880;
wire [3:0] u_ca_out_881;
wire [3:0] u_ca_out_882;
wire [3:0] u_ca_out_883;
wire [3:0] u_ca_out_884;
wire [3:0] u_ca_out_885;
wire [3:0] u_ca_out_886;
wire [3:0] u_ca_out_887;
wire [3:0] u_ca_out_888;
wire [3:0] u_ca_out_889;
wire [3:0] u_ca_out_890;
wire [3:0] u_ca_out_891;
wire [3:0] u_ca_out_892;
wire [3:0] u_ca_out_893;
wire [3:0] u_ca_out_894;
wire [3:0] u_ca_out_895;
wire [3:0] u_ca_out_896;
wire [3:0] u_ca_out_897;
wire [3:0] u_ca_out_898;
wire [3:0] u_ca_out_899;
wire [3:0] u_ca_out_900;
wire [3:0] u_ca_out_901;
wire [3:0] u_ca_out_902;
wire [3:0] u_ca_out_903;
wire [3:0] u_ca_out_904;
wire [3:0] u_ca_out_905;
wire [3:0] u_ca_out_906;
wire [3:0] u_ca_out_907;
wire [3:0] u_ca_out_908;
wire [3:0] u_ca_out_909;
wire [3:0] u_ca_out_910;
wire [3:0] u_ca_out_911;
wire [3:0] u_ca_out_912;
wire [3:0] u_ca_out_913;
wire [3:0] u_ca_out_914;
wire [3:0] u_ca_out_915;
wire [3:0] u_ca_out_916;
wire [3:0] u_ca_out_917;
wire [3:0] u_ca_out_918;
wire [3:0] u_ca_out_919;
wire [3:0] u_ca_out_920;
wire [3:0] u_ca_out_921;
wire [3:0] u_ca_out_922;
wire [3:0] u_ca_out_923;
wire [3:0] u_ca_out_924;
wire [3:0] u_ca_out_925;
wire [3:0] u_ca_out_926;
wire [3:0] u_ca_out_927;
wire [3:0] u_ca_out_928;
wire [3:0] u_ca_out_929;
wire [3:0] u_ca_out_930;
wire [3:0] u_ca_out_931;
wire [3:0] u_ca_out_932;
wire [3:0] u_ca_out_933;
wire [3:0] u_ca_out_934;
wire [3:0] u_ca_out_935;
wire [3:0] u_ca_out_936;
wire [3:0] u_ca_out_937;
wire [3:0] u_ca_out_938;
wire [3:0] u_ca_out_939;
wire [3:0] u_ca_out_940;
wire [3:0] u_ca_out_941;
wire [3:0] u_ca_out_942;
wire [3:0] u_ca_out_943;
wire [3:0] u_ca_out_944;
wire [3:0] u_ca_out_945;
wire [3:0] u_ca_out_946;
wire [3:0] u_ca_out_947;
wire [3:0] u_ca_out_948;
wire [3:0] u_ca_out_949;
wire [3:0] u_ca_out_950;
wire [3:0] u_ca_out_951;
wire [3:0] u_ca_out_952;
wire [3:0] u_ca_out_953;
wire [3:0] u_ca_out_954;
wire [3:0] u_ca_out_955;
wire [3:0] u_ca_out_956;
wire [3:0] u_ca_out_957;
wire [3:0] u_ca_out_958;
wire [3:0] u_ca_out_959;
wire [3:0] u_ca_out_960;
wire [3:0] u_ca_out_961;
wire [3:0] u_ca_out_962;
wire [3:0] u_ca_out_963;
wire [3:0] u_ca_out_964;
wire [3:0] u_ca_out_965;
wire [3:0] u_ca_out_966;
wire [3:0] u_ca_out_967;
wire [3:0] u_ca_out_968;
wire [3:0] u_ca_out_969;
wire [3:0] u_ca_out_970;
wire [3:0] u_ca_out_971;
wire [3:0] u_ca_out_972;
wire [3:0] u_ca_out_973;
wire [3:0] u_ca_out_974;
wire [3:0] u_ca_out_975;
wire [3:0] u_ca_out_976;
wire [3:0] u_ca_out_977;
wire [3:0] u_ca_out_978;
wire [3:0] u_ca_out_979;
wire [3:0] u_ca_out_980;
wire [3:0] u_ca_out_981;
wire [3:0] u_ca_out_982;
wire [3:0] u_ca_out_983;
wire [3:0] u_ca_out_984;
wire [3:0] u_ca_out_985;
wire [3:0] u_ca_out_986;
wire [3:0] u_ca_out_987;
wire [3:0] u_ca_out_988;
wire [3:0] u_ca_out_989;
wire [3:0] u_ca_out_990;
wire [3:0] u_ca_out_991;
wire [3:0] u_ca_out_992;
wire [3:0] u_ca_out_993;
wire [3:0] u_ca_out_994;
wire [3:0] u_ca_out_995;
wire [3:0] u_ca_out_996;
wire [3:0] u_ca_out_997;
wire [3:0] u_ca_out_998;
wire [3:0] u_ca_out_999;
wire [3:0] u_ca_out_1000;
wire [3:0] u_ca_out_1001;
wire [3:0] u_ca_out_1002;
wire [3:0] u_ca_out_1003;
wire [3:0] u_ca_out_1004;
wire [3:0] u_ca_out_1005;
wire [3:0] u_ca_out_1006;
wire [3:0] u_ca_out_1007;
wire [3:0] u_ca_out_1008;
wire [3:0] u_ca_out_1009;
wire [3:0] u_ca_out_1010;
wire [3:0] u_ca_out_1011;
wire [3:0] u_ca_out_1012;
wire [3:0] u_ca_out_1013;
wire [3:0] u_ca_out_1014;
wire [3:0] u_ca_out_1015;
wire [3:0] u_ca_out_1016;
wire [3:0] u_ca_out_1017;
wire [3:0] u_ca_out_1018;
wire [3:0] u_ca_out_1019;
wire [3:0] u_ca_out_1020;
wire [3:0] u_ca_out_1021;
wire [3:0] u_ca_out_1022;
wire [3:0] u_ca_out_1023;

assign u_ca_in_0 = col_in_0;
assign u_ca_in_1 = col_in_1;
assign u_ca_in_2 = col_in_2;
assign u_ca_in_3 = col_in_3;
assign u_ca_in_4 = col_in_4;
assign u_ca_in_5 = col_in_5;
assign u_ca_in_6 = col_in_6;
assign u_ca_in_7 = col_in_7;
assign u_ca_in_8 = col_in_8;
assign u_ca_in_9 = col_in_9;
assign u_ca_in_10 = col_in_10;
assign u_ca_in_11 = col_in_11;
assign u_ca_in_12 = col_in_12;
assign u_ca_in_13 = col_in_13;
assign u_ca_in_14 = col_in_14;
assign u_ca_in_15 = col_in_15;
assign u_ca_in_16 = col_in_16;
assign u_ca_in_17 = col_in_17;
assign u_ca_in_18 = col_in_18;
assign u_ca_in_19 = col_in_19;
assign u_ca_in_20 = col_in_20;
assign u_ca_in_21 = col_in_21;
assign u_ca_in_22 = col_in_22;
assign u_ca_in_23 = col_in_23;
assign u_ca_in_24 = col_in_24;
assign u_ca_in_25 = col_in_25;
assign u_ca_in_26 = col_in_26;
assign u_ca_in_27 = col_in_27;
assign u_ca_in_28 = col_in_28;
assign u_ca_in_29 = col_in_29;
assign u_ca_in_30 = col_in_30;
assign u_ca_in_31 = col_in_31;
assign u_ca_in_32 = col_in_32;
assign u_ca_in_33 = col_in_33;
assign u_ca_in_34 = col_in_34;
assign u_ca_in_35 = col_in_35;
assign u_ca_in_36 = col_in_36;
assign u_ca_in_37 = col_in_37;
assign u_ca_in_38 = col_in_38;
assign u_ca_in_39 = col_in_39;
assign u_ca_in_40 = col_in_40;
assign u_ca_in_41 = col_in_41;
assign u_ca_in_42 = col_in_42;
assign u_ca_in_43 = col_in_43;
assign u_ca_in_44 = col_in_44;
assign u_ca_in_45 = col_in_45;
assign u_ca_in_46 = col_in_46;
assign u_ca_in_47 = col_in_47;
assign u_ca_in_48 = col_in_48;
assign u_ca_in_49 = col_in_49;
assign u_ca_in_50 = col_in_50;
assign u_ca_in_51 = col_in_51;
assign u_ca_in_52 = col_in_52;
assign u_ca_in_53 = col_in_53;
assign u_ca_in_54 = col_in_54;
assign u_ca_in_55 = col_in_55;
assign u_ca_in_56 = col_in_56;
assign u_ca_in_57 = col_in_57;
assign u_ca_in_58 = col_in_58;
assign u_ca_in_59 = col_in_59;
assign u_ca_in_60 = col_in_60;
assign u_ca_in_61 = col_in_61;
assign u_ca_in_62 = col_in_62;
assign u_ca_in_63 = col_in_63;
assign u_ca_in_64 = col_in_64;
assign u_ca_in_65 = col_in_65;
assign u_ca_in_66 = col_in_66;
assign u_ca_in_67 = col_in_67;
assign u_ca_in_68 = col_in_68;
assign u_ca_in_69 = col_in_69;
assign u_ca_in_70 = col_in_70;
assign u_ca_in_71 = col_in_71;
assign u_ca_in_72 = col_in_72;
assign u_ca_in_73 = col_in_73;
assign u_ca_in_74 = col_in_74;
assign u_ca_in_75 = col_in_75;
assign u_ca_in_76 = col_in_76;
assign u_ca_in_77 = col_in_77;
assign u_ca_in_78 = col_in_78;
assign u_ca_in_79 = col_in_79;
assign u_ca_in_80 = col_in_80;
assign u_ca_in_81 = col_in_81;
assign u_ca_in_82 = col_in_82;
assign u_ca_in_83 = col_in_83;
assign u_ca_in_84 = col_in_84;
assign u_ca_in_85 = col_in_85;
assign u_ca_in_86 = col_in_86;
assign u_ca_in_87 = col_in_87;
assign u_ca_in_88 = col_in_88;
assign u_ca_in_89 = col_in_89;
assign u_ca_in_90 = col_in_90;
assign u_ca_in_91 = col_in_91;
assign u_ca_in_92 = col_in_92;
assign u_ca_in_93 = col_in_93;
assign u_ca_in_94 = col_in_94;
assign u_ca_in_95 = col_in_95;
assign u_ca_in_96 = col_in_96;
assign u_ca_in_97 = col_in_97;
assign u_ca_in_98 = col_in_98;
assign u_ca_in_99 = col_in_99;
assign u_ca_in_100 = col_in_100;
assign u_ca_in_101 = col_in_101;
assign u_ca_in_102 = col_in_102;
assign u_ca_in_103 = col_in_103;
assign u_ca_in_104 = col_in_104;
assign u_ca_in_105 = col_in_105;
assign u_ca_in_106 = col_in_106;
assign u_ca_in_107 = col_in_107;
assign u_ca_in_108 = col_in_108;
assign u_ca_in_109 = col_in_109;
assign u_ca_in_110 = col_in_110;
assign u_ca_in_111 = col_in_111;
assign u_ca_in_112 = col_in_112;
assign u_ca_in_113 = col_in_113;
assign u_ca_in_114 = col_in_114;
assign u_ca_in_115 = col_in_115;
assign u_ca_in_116 = col_in_116;
assign u_ca_in_117 = col_in_117;
assign u_ca_in_118 = col_in_118;
assign u_ca_in_119 = col_in_119;
assign u_ca_in_120 = col_in_120;
assign u_ca_in_121 = col_in_121;
assign u_ca_in_122 = col_in_122;
assign u_ca_in_123 = col_in_123;
assign u_ca_in_124 = col_in_124;
assign u_ca_in_125 = col_in_125;
assign u_ca_in_126 = col_in_126;
assign u_ca_in_127 = col_in_127;
assign u_ca_in_128 = col_in_128;
assign u_ca_in_129 = col_in_129;
assign u_ca_in_130 = col_in_130;
assign u_ca_in_131 = col_in_131;
assign u_ca_in_132 = col_in_132;
assign u_ca_in_133 = col_in_133;
assign u_ca_in_134 = col_in_134;
assign u_ca_in_135 = col_in_135;
assign u_ca_in_136 = col_in_136;
assign u_ca_in_137 = col_in_137;
assign u_ca_in_138 = col_in_138;
assign u_ca_in_139 = col_in_139;
assign u_ca_in_140 = col_in_140;
assign u_ca_in_141 = col_in_141;
assign u_ca_in_142 = col_in_142;
assign u_ca_in_143 = col_in_143;
assign u_ca_in_144 = col_in_144;
assign u_ca_in_145 = col_in_145;
assign u_ca_in_146 = col_in_146;
assign u_ca_in_147 = col_in_147;
assign u_ca_in_148 = col_in_148;
assign u_ca_in_149 = col_in_149;
assign u_ca_in_150 = col_in_150;
assign u_ca_in_151 = col_in_151;
assign u_ca_in_152 = col_in_152;
assign u_ca_in_153 = col_in_153;
assign u_ca_in_154 = col_in_154;
assign u_ca_in_155 = col_in_155;
assign u_ca_in_156 = col_in_156;
assign u_ca_in_157 = col_in_157;
assign u_ca_in_158 = col_in_158;
assign u_ca_in_159 = col_in_159;
assign u_ca_in_160 = col_in_160;
assign u_ca_in_161 = col_in_161;
assign u_ca_in_162 = col_in_162;
assign u_ca_in_163 = col_in_163;
assign u_ca_in_164 = col_in_164;
assign u_ca_in_165 = col_in_165;
assign u_ca_in_166 = col_in_166;
assign u_ca_in_167 = col_in_167;
assign u_ca_in_168 = col_in_168;
assign u_ca_in_169 = col_in_169;
assign u_ca_in_170 = col_in_170;
assign u_ca_in_171 = col_in_171;
assign u_ca_in_172 = col_in_172;
assign u_ca_in_173 = col_in_173;
assign u_ca_in_174 = col_in_174;
assign u_ca_in_175 = col_in_175;
assign u_ca_in_176 = col_in_176;
assign u_ca_in_177 = col_in_177;
assign u_ca_in_178 = col_in_178;
assign u_ca_in_179 = col_in_179;
assign u_ca_in_180 = col_in_180;
assign u_ca_in_181 = col_in_181;
assign u_ca_in_182 = col_in_182;
assign u_ca_in_183 = col_in_183;
assign u_ca_in_184 = col_in_184;
assign u_ca_in_185 = col_in_185;
assign u_ca_in_186 = col_in_186;
assign u_ca_in_187 = col_in_187;
assign u_ca_in_188 = col_in_188;
assign u_ca_in_189 = col_in_189;
assign u_ca_in_190 = col_in_190;
assign u_ca_in_191 = col_in_191;
assign u_ca_in_192 = col_in_192;
assign u_ca_in_193 = col_in_193;
assign u_ca_in_194 = col_in_194;
assign u_ca_in_195 = col_in_195;
assign u_ca_in_196 = col_in_196;
assign u_ca_in_197 = col_in_197;
assign u_ca_in_198 = col_in_198;
assign u_ca_in_199 = col_in_199;
assign u_ca_in_200 = col_in_200;
assign u_ca_in_201 = col_in_201;
assign u_ca_in_202 = col_in_202;
assign u_ca_in_203 = col_in_203;
assign u_ca_in_204 = col_in_204;
assign u_ca_in_205 = col_in_205;
assign u_ca_in_206 = col_in_206;
assign u_ca_in_207 = col_in_207;
assign u_ca_in_208 = col_in_208;
assign u_ca_in_209 = col_in_209;
assign u_ca_in_210 = col_in_210;
assign u_ca_in_211 = col_in_211;
assign u_ca_in_212 = col_in_212;
assign u_ca_in_213 = col_in_213;
assign u_ca_in_214 = col_in_214;
assign u_ca_in_215 = col_in_215;
assign u_ca_in_216 = col_in_216;
assign u_ca_in_217 = col_in_217;
assign u_ca_in_218 = col_in_218;
assign u_ca_in_219 = col_in_219;
assign u_ca_in_220 = col_in_220;
assign u_ca_in_221 = col_in_221;
assign u_ca_in_222 = col_in_222;
assign u_ca_in_223 = col_in_223;
assign u_ca_in_224 = col_in_224;
assign u_ca_in_225 = col_in_225;
assign u_ca_in_226 = col_in_226;
assign u_ca_in_227 = col_in_227;
assign u_ca_in_228 = col_in_228;
assign u_ca_in_229 = col_in_229;
assign u_ca_in_230 = col_in_230;
assign u_ca_in_231 = col_in_231;
assign u_ca_in_232 = col_in_232;
assign u_ca_in_233 = col_in_233;
assign u_ca_in_234 = col_in_234;
assign u_ca_in_235 = col_in_235;
assign u_ca_in_236 = col_in_236;
assign u_ca_in_237 = col_in_237;
assign u_ca_in_238 = col_in_238;
assign u_ca_in_239 = col_in_239;
assign u_ca_in_240 = col_in_240;
assign u_ca_in_241 = col_in_241;
assign u_ca_in_242 = col_in_242;
assign u_ca_in_243 = col_in_243;
assign u_ca_in_244 = col_in_244;
assign u_ca_in_245 = col_in_245;
assign u_ca_in_246 = col_in_246;
assign u_ca_in_247 = col_in_247;
assign u_ca_in_248 = col_in_248;
assign u_ca_in_249 = col_in_249;
assign u_ca_in_250 = col_in_250;
assign u_ca_in_251 = col_in_251;
assign u_ca_in_252 = col_in_252;
assign u_ca_in_253 = col_in_253;
assign u_ca_in_254 = col_in_254;
assign u_ca_in_255 = col_in_255;
assign u_ca_in_256 = col_in_256;
assign u_ca_in_257 = col_in_257;
assign u_ca_in_258 = col_in_258;
assign u_ca_in_259 = col_in_259;
assign u_ca_in_260 = col_in_260;
assign u_ca_in_261 = col_in_261;
assign u_ca_in_262 = col_in_262;
assign u_ca_in_263 = col_in_263;
assign u_ca_in_264 = col_in_264;
assign u_ca_in_265 = col_in_265;
assign u_ca_in_266 = col_in_266;
assign u_ca_in_267 = col_in_267;
assign u_ca_in_268 = col_in_268;
assign u_ca_in_269 = col_in_269;
assign u_ca_in_270 = col_in_270;
assign u_ca_in_271 = col_in_271;
assign u_ca_in_272 = col_in_272;
assign u_ca_in_273 = col_in_273;
assign u_ca_in_274 = col_in_274;
assign u_ca_in_275 = col_in_275;
assign u_ca_in_276 = col_in_276;
assign u_ca_in_277 = col_in_277;
assign u_ca_in_278 = col_in_278;
assign u_ca_in_279 = col_in_279;
assign u_ca_in_280 = col_in_280;
assign u_ca_in_281 = col_in_281;
assign u_ca_in_282 = col_in_282;
assign u_ca_in_283 = col_in_283;
assign u_ca_in_284 = col_in_284;
assign u_ca_in_285 = col_in_285;
assign u_ca_in_286 = col_in_286;
assign u_ca_in_287 = col_in_287;
assign u_ca_in_288 = col_in_288;
assign u_ca_in_289 = col_in_289;
assign u_ca_in_290 = col_in_290;
assign u_ca_in_291 = col_in_291;
assign u_ca_in_292 = col_in_292;
assign u_ca_in_293 = col_in_293;
assign u_ca_in_294 = col_in_294;
assign u_ca_in_295 = col_in_295;
assign u_ca_in_296 = col_in_296;
assign u_ca_in_297 = col_in_297;
assign u_ca_in_298 = col_in_298;
assign u_ca_in_299 = col_in_299;
assign u_ca_in_300 = col_in_300;
assign u_ca_in_301 = col_in_301;
assign u_ca_in_302 = col_in_302;
assign u_ca_in_303 = col_in_303;
assign u_ca_in_304 = col_in_304;
assign u_ca_in_305 = col_in_305;
assign u_ca_in_306 = col_in_306;
assign u_ca_in_307 = col_in_307;
assign u_ca_in_308 = col_in_308;
assign u_ca_in_309 = col_in_309;
assign u_ca_in_310 = col_in_310;
assign u_ca_in_311 = col_in_311;
assign u_ca_in_312 = col_in_312;
assign u_ca_in_313 = col_in_313;
assign u_ca_in_314 = col_in_314;
assign u_ca_in_315 = col_in_315;
assign u_ca_in_316 = col_in_316;
assign u_ca_in_317 = col_in_317;
assign u_ca_in_318 = col_in_318;
assign u_ca_in_319 = col_in_319;
assign u_ca_in_320 = col_in_320;
assign u_ca_in_321 = col_in_321;
assign u_ca_in_322 = col_in_322;
assign u_ca_in_323 = col_in_323;
assign u_ca_in_324 = col_in_324;
assign u_ca_in_325 = col_in_325;
assign u_ca_in_326 = col_in_326;
assign u_ca_in_327 = col_in_327;
assign u_ca_in_328 = col_in_328;
assign u_ca_in_329 = col_in_329;
assign u_ca_in_330 = col_in_330;
assign u_ca_in_331 = col_in_331;
assign u_ca_in_332 = col_in_332;
assign u_ca_in_333 = col_in_333;
assign u_ca_in_334 = col_in_334;
assign u_ca_in_335 = col_in_335;
assign u_ca_in_336 = col_in_336;
assign u_ca_in_337 = col_in_337;
assign u_ca_in_338 = col_in_338;
assign u_ca_in_339 = col_in_339;
assign u_ca_in_340 = col_in_340;
assign u_ca_in_341 = col_in_341;
assign u_ca_in_342 = col_in_342;
assign u_ca_in_343 = col_in_343;
assign u_ca_in_344 = col_in_344;
assign u_ca_in_345 = col_in_345;
assign u_ca_in_346 = col_in_346;
assign u_ca_in_347 = col_in_347;
assign u_ca_in_348 = col_in_348;
assign u_ca_in_349 = col_in_349;
assign u_ca_in_350 = col_in_350;
assign u_ca_in_351 = col_in_351;
assign u_ca_in_352 = col_in_352;
assign u_ca_in_353 = col_in_353;
assign u_ca_in_354 = col_in_354;
assign u_ca_in_355 = col_in_355;
assign u_ca_in_356 = col_in_356;
assign u_ca_in_357 = col_in_357;
assign u_ca_in_358 = col_in_358;
assign u_ca_in_359 = col_in_359;
assign u_ca_in_360 = col_in_360;
assign u_ca_in_361 = col_in_361;
assign u_ca_in_362 = col_in_362;
assign u_ca_in_363 = col_in_363;
assign u_ca_in_364 = col_in_364;
assign u_ca_in_365 = col_in_365;
assign u_ca_in_366 = col_in_366;
assign u_ca_in_367 = col_in_367;
assign u_ca_in_368 = col_in_368;
assign u_ca_in_369 = col_in_369;
assign u_ca_in_370 = col_in_370;
assign u_ca_in_371 = col_in_371;
assign u_ca_in_372 = col_in_372;
assign u_ca_in_373 = col_in_373;
assign u_ca_in_374 = col_in_374;
assign u_ca_in_375 = col_in_375;
assign u_ca_in_376 = col_in_376;
assign u_ca_in_377 = col_in_377;
assign u_ca_in_378 = col_in_378;
assign u_ca_in_379 = col_in_379;
assign u_ca_in_380 = col_in_380;
assign u_ca_in_381 = col_in_381;
assign u_ca_in_382 = col_in_382;
assign u_ca_in_383 = col_in_383;
assign u_ca_in_384 = col_in_384;
assign u_ca_in_385 = col_in_385;
assign u_ca_in_386 = col_in_386;
assign u_ca_in_387 = col_in_387;
assign u_ca_in_388 = col_in_388;
assign u_ca_in_389 = col_in_389;
assign u_ca_in_390 = col_in_390;
assign u_ca_in_391 = col_in_391;
assign u_ca_in_392 = col_in_392;
assign u_ca_in_393 = col_in_393;
assign u_ca_in_394 = col_in_394;
assign u_ca_in_395 = col_in_395;
assign u_ca_in_396 = col_in_396;
assign u_ca_in_397 = col_in_397;
assign u_ca_in_398 = col_in_398;
assign u_ca_in_399 = col_in_399;
assign u_ca_in_400 = col_in_400;
assign u_ca_in_401 = col_in_401;
assign u_ca_in_402 = col_in_402;
assign u_ca_in_403 = col_in_403;
assign u_ca_in_404 = col_in_404;
assign u_ca_in_405 = col_in_405;
assign u_ca_in_406 = col_in_406;
assign u_ca_in_407 = col_in_407;
assign u_ca_in_408 = col_in_408;
assign u_ca_in_409 = col_in_409;
assign u_ca_in_410 = col_in_410;
assign u_ca_in_411 = col_in_411;
assign u_ca_in_412 = col_in_412;
assign u_ca_in_413 = col_in_413;
assign u_ca_in_414 = col_in_414;
assign u_ca_in_415 = col_in_415;
assign u_ca_in_416 = col_in_416;
assign u_ca_in_417 = col_in_417;
assign u_ca_in_418 = col_in_418;
assign u_ca_in_419 = col_in_419;
assign u_ca_in_420 = col_in_420;
assign u_ca_in_421 = col_in_421;
assign u_ca_in_422 = col_in_422;
assign u_ca_in_423 = col_in_423;
assign u_ca_in_424 = col_in_424;
assign u_ca_in_425 = col_in_425;
assign u_ca_in_426 = col_in_426;
assign u_ca_in_427 = col_in_427;
assign u_ca_in_428 = col_in_428;
assign u_ca_in_429 = col_in_429;
assign u_ca_in_430 = col_in_430;
assign u_ca_in_431 = col_in_431;
assign u_ca_in_432 = col_in_432;
assign u_ca_in_433 = col_in_433;
assign u_ca_in_434 = col_in_434;
assign u_ca_in_435 = col_in_435;
assign u_ca_in_436 = col_in_436;
assign u_ca_in_437 = col_in_437;
assign u_ca_in_438 = col_in_438;
assign u_ca_in_439 = col_in_439;
assign u_ca_in_440 = col_in_440;
assign u_ca_in_441 = col_in_441;
assign u_ca_in_442 = col_in_442;
assign u_ca_in_443 = col_in_443;
assign u_ca_in_444 = col_in_444;
assign u_ca_in_445 = col_in_445;
assign u_ca_in_446 = col_in_446;
assign u_ca_in_447 = col_in_447;
assign u_ca_in_448 = col_in_448;
assign u_ca_in_449 = col_in_449;
assign u_ca_in_450 = col_in_450;
assign u_ca_in_451 = col_in_451;
assign u_ca_in_452 = col_in_452;
assign u_ca_in_453 = col_in_453;
assign u_ca_in_454 = col_in_454;
assign u_ca_in_455 = col_in_455;
assign u_ca_in_456 = col_in_456;
assign u_ca_in_457 = col_in_457;
assign u_ca_in_458 = col_in_458;
assign u_ca_in_459 = col_in_459;
assign u_ca_in_460 = col_in_460;
assign u_ca_in_461 = col_in_461;
assign u_ca_in_462 = col_in_462;
assign u_ca_in_463 = col_in_463;
assign u_ca_in_464 = col_in_464;
assign u_ca_in_465 = col_in_465;
assign u_ca_in_466 = col_in_466;
assign u_ca_in_467 = col_in_467;
assign u_ca_in_468 = col_in_468;
assign u_ca_in_469 = col_in_469;
assign u_ca_in_470 = col_in_470;
assign u_ca_in_471 = col_in_471;
assign u_ca_in_472 = col_in_472;
assign u_ca_in_473 = col_in_473;
assign u_ca_in_474 = col_in_474;
assign u_ca_in_475 = col_in_475;
assign u_ca_in_476 = col_in_476;
assign u_ca_in_477 = col_in_477;
assign u_ca_in_478 = col_in_478;
assign u_ca_in_479 = col_in_479;
assign u_ca_in_480 = col_in_480;
assign u_ca_in_481 = col_in_481;
assign u_ca_in_482 = col_in_482;
assign u_ca_in_483 = col_in_483;
assign u_ca_in_484 = col_in_484;
assign u_ca_in_485 = col_in_485;
assign u_ca_in_486 = col_in_486;
assign u_ca_in_487 = col_in_487;
assign u_ca_in_488 = col_in_488;
assign u_ca_in_489 = col_in_489;
assign u_ca_in_490 = col_in_490;
assign u_ca_in_491 = col_in_491;
assign u_ca_in_492 = col_in_492;
assign u_ca_in_493 = col_in_493;
assign u_ca_in_494 = col_in_494;
assign u_ca_in_495 = col_in_495;
assign u_ca_in_496 = col_in_496;
assign u_ca_in_497 = col_in_497;
assign u_ca_in_498 = col_in_498;
assign u_ca_in_499 = col_in_499;
assign u_ca_in_500 = col_in_500;
assign u_ca_in_501 = col_in_501;
assign u_ca_in_502 = col_in_502;
assign u_ca_in_503 = col_in_503;
assign u_ca_in_504 = col_in_504;
assign u_ca_in_505 = col_in_505;
assign u_ca_in_506 = col_in_506;
assign u_ca_in_507 = col_in_507;
assign u_ca_in_508 = col_in_508;
assign u_ca_in_509 = col_in_509;
assign u_ca_in_510 = col_in_510;
assign u_ca_in_511 = col_in_511;
assign u_ca_in_512 = col_in_512;
assign u_ca_in_513 = col_in_513;
assign u_ca_in_514 = col_in_514;
assign u_ca_in_515 = col_in_515;
assign u_ca_in_516 = col_in_516;
assign u_ca_in_517 = col_in_517;
assign u_ca_in_518 = col_in_518;
assign u_ca_in_519 = col_in_519;
assign u_ca_in_520 = col_in_520;
assign u_ca_in_521 = col_in_521;
assign u_ca_in_522 = col_in_522;
assign u_ca_in_523 = col_in_523;
assign u_ca_in_524 = col_in_524;
assign u_ca_in_525 = col_in_525;
assign u_ca_in_526 = col_in_526;
assign u_ca_in_527 = col_in_527;
assign u_ca_in_528 = col_in_528;
assign u_ca_in_529 = col_in_529;
assign u_ca_in_530 = col_in_530;
assign u_ca_in_531 = col_in_531;
assign u_ca_in_532 = col_in_532;
assign u_ca_in_533 = col_in_533;
assign u_ca_in_534 = col_in_534;
assign u_ca_in_535 = col_in_535;
assign u_ca_in_536 = col_in_536;
assign u_ca_in_537 = col_in_537;
assign u_ca_in_538 = col_in_538;
assign u_ca_in_539 = col_in_539;
assign u_ca_in_540 = col_in_540;
assign u_ca_in_541 = col_in_541;
assign u_ca_in_542 = col_in_542;
assign u_ca_in_543 = col_in_543;
assign u_ca_in_544 = col_in_544;
assign u_ca_in_545 = col_in_545;
assign u_ca_in_546 = col_in_546;
assign u_ca_in_547 = col_in_547;
assign u_ca_in_548 = col_in_548;
assign u_ca_in_549 = col_in_549;
assign u_ca_in_550 = col_in_550;
assign u_ca_in_551 = col_in_551;
assign u_ca_in_552 = col_in_552;
assign u_ca_in_553 = col_in_553;
assign u_ca_in_554 = col_in_554;
assign u_ca_in_555 = col_in_555;
assign u_ca_in_556 = col_in_556;
assign u_ca_in_557 = col_in_557;
assign u_ca_in_558 = col_in_558;
assign u_ca_in_559 = col_in_559;
assign u_ca_in_560 = col_in_560;
assign u_ca_in_561 = col_in_561;
assign u_ca_in_562 = col_in_562;
assign u_ca_in_563 = col_in_563;
assign u_ca_in_564 = col_in_564;
assign u_ca_in_565 = col_in_565;
assign u_ca_in_566 = col_in_566;
assign u_ca_in_567 = col_in_567;
assign u_ca_in_568 = col_in_568;
assign u_ca_in_569 = col_in_569;
assign u_ca_in_570 = col_in_570;
assign u_ca_in_571 = col_in_571;
assign u_ca_in_572 = col_in_572;
assign u_ca_in_573 = col_in_573;
assign u_ca_in_574 = col_in_574;
assign u_ca_in_575 = col_in_575;
assign u_ca_in_576 = col_in_576;
assign u_ca_in_577 = col_in_577;
assign u_ca_in_578 = col_in_578;
assign u_ca_in_579 = col_in_579;
assign u_ca_in_580 = col_in_580;
assign u_ca_in_581 = col_in_581;
assign u_ca_in_582 = col_in_582;
assign u_ca_in_583 = col_in_583;
assign u_ca_in_584 = col_in_584;
assign u_ca_in_585 = col_in_585;
assign u_ca_in_586 = col_in_586;
assign u_ca_in_587 = col_in_587;
assign u_ca_in_588 = col_in_588;
assign u_ca_in_589 = col_in_589;
assign u_ca_in_590 = col_in_590;
assign u_ca_in_591 = col_in_591;
assign u_ca_in_592 = col_in_592;
assign u_ca_in_593 = col_in_593;
assign u_ca_in_594 = col_in_594;
assign u_ca_in_595 = col_in_595;
assign u_ca_in_596 = col_in_596;
assign u_ca_in_597 = col_in_597;
assign u_ca_in_598 = col_in_598;
assign u_ca_in_599 = col_in_599;
assign u_ca_in_600 = col_in_600;
assign u_ca_in_601 = col_in_601;
assign u_ca_in_602 = col_in_602;
assign u_ca_in_603 = col_in_603;
assign u_ca_in_604 = col_in_604;
assign u_ca_in_605 = col_in_605;
assign u_ca_in_606 = col_in_606;
assign u_ca_in_607 = col_in_607;
assign u_ca_in_608 = col_in_608;
assign u_ca_in_609 = col_in_609;
assign u_ca_in_610 = col_in_610;
assign u_ca_in_611 = col_in_611;
assign u_ca_in_612 = col_in_612;
assign u_ca_in_613 = col_in_613;
assign u_ca_in_614 = col_in_614;
assign u_ca_in_615 = col_in_615;
assign u_ca_in_616 = col_in_616;
assign u_ca_in_617 = col_in_617;
assign u_ca_in_618 = col_in_618;
assign u_ca_in_619 = col_in_619;
assign u_ca_in_620 = col_in_620;
assign u_ca_in_621 = col_in_621;
assign u_ca_in_622 = col_in_622;
assign u_ca_in_623 = col_in_623;
assign u_ca_in_624 = col_in_624;
assign u_ca_in_625 = col_in_625;
assign u_ca_in_626 = col_in_626;
assign u_ca_in_627 = col_in_627;
assign u_ca_in_628 = col_in_628;
assign u_ca_in_629 = col_in_629;
assign u_ca_in_630 = col_in_630;
assign u_ca_in_631 = col_in_631;
assign u_ca_in_632 = col_in_632;
assign u_ca_in_633 = col_in_633;
assign u_ca_in_634 = col_in_634;
assign u_ca_in_635 = col_in_635;
assign u_ca_in_636 = col_in_636;
assign u_ca_in_637 = col_in_637;
assign u_ca_in_638 = col_in_638;
assign u_ca_in_639 = col_in_639;
assign u_ca_in_640 = col_in_640;
assign u_ca_in_641 = col_in_641;
assign u_ca_in_642 = col_in_642;
assign u_ca_in_643 = col_in_643;
assign u_ca_in_644 = col_in_644;
assign u_ca_in_645 = col_in_645;
assign u_ca_in_646 = col_in_646;
assign u_ca_in_647 = col_in_647;
assign u_ca_in_648 = col_in_648;
assign u_ca_in_649 = col_in_649;
assign u_ca_in_650 = col_in_650;
assign u_ca_in_651 = col_in_651;
assign u_ca_in_652 = col_in_652;
assign u_ca_in_653 = col_in_653;
assign u_ca_in_654 = col_in_654;
assign u_ca_in_655 = col_in_655;
assign u_ca_in_656 = col_in_656;
assign u_ca_in_657 = col_in_657;
assign u_ca_in_658 = col_in_658;
assign u_ca_in_659 = col_in_659;
assign u_ca_in_660 = col_in_660;
assign u_ca_in_661 = col_in_661;
assign u_ca_in_662 = col_in_662;
assign u_ca_in_663 = col_in_663;
assign u_ca_in_664 = col_in_664;
assign u_ca_in_665 = col_in_665;
assign u_ca_in_666 = col_in_666;
assign u_ca_in_667 = col_in_667;
assign u_ca_in_668 = col_in_668;
assign u_ca_in_669 = col_in_669;
assign u_ca_in_670 = col_in_670;
assign u_ca_in_671 = col_in_671;
assign u_ca_in_672 = col_in_672;
assign u_ca_in_673 = col_in_673;
assign u_ca_in_674 = col_in_674;
assign u_ca_in_675 = col_in_675;
assign u_ca_in_676 = col_in_676;
assign u_ca_in_677 = col_in_677;
assign u_ca_in_678 = col_in_678;
assign u_ca_in_679 = col_in_679;
assign u_ca_in_680 = col_in_680;
assign u_ca_in_681 = col_in_681;
assign u_ca_in_682 = col_in_682;
assign u_ca_in_683 = col_in_683;
assign u_ca_in_684 = col_in_684;
assign u_ca_in_685 = col_in_685;
assign u_ca_in_686 = col_in_686;
assign u_ca_in_687 = col_in_687;
assign u_ca_in_688 = col_in_688;
assign u_ca_in_689 = col_in_689;
assign u_ca_in_690 = col_in_690;
assign u_ca_in_691 = col_in_691;
assign u_ca_in_692 = col_in_692;
assign u_ca_in_693 = col_in_693;
assign u_ca_in_694 = col_in_694;
assign u_ca_in_695 = col_in_695;
assign u_ca_in_696 = col_in_696;
assign u_ca_in_697 = col_in_697;
assign u_ca_in_698 = col_in_698;
assign u_ca_in_699 = col_in_699;
assign u_ca_in_700 = col_in_700;
assign u_ca_in_701 = col_in_701;
assign u_ca_in_702 = col_in_702;
assign u_ca_in_703 = col_in_703;
assign u_ca_in_704 = col_in_704;
assign u_ca_in_705 = col_in_705;
assign u_ca_in_706 = col_in_706;
assign u_ca_in_707 = col_in_707;
assign u_ca_in_708 = col_in_708;
assign u_ca_in_709 = col_in_709;
assign u_ca_in_710 = col_in_710;
assign u_ca_in_711 = col_in_711;
assign u_ca_in_712 = col_in_712;
assign u_ca_in_713 = col_in_713;
assign u_ca_in_714 = col_in_714;
assign u_ca_in_715 = col_in_715;
assign u_ca_in_716 = col_in_716;
assign u_ca_in_717 = col_in_717;
assign u_ca_in_718 = col_in_718;
assign u_ca_in_719 = col_in_719;
assign u_ca_in_720 = col_in_720;
assign u_ca_in_721 = col_in_721;
assign u_ca_in_722 = col_in_722;
assign u_ca_in_723 = col_in_723;
assign u_ca_in_724 = col_in_724;
assign u_ca_in_725 = col_in_725;
assign u_ca_in_726 = col_in_726;
assign u_ca_in_727 = col_in_727;
assign u_ca_in_728 = col_in_728;
assign u_ca_in_729 = col_in_729;
assign u_ca_in_730 = col_in_730;
assign u_ca_in_731 = col_in_731;
assign u_ca_in_732 = col_in_732;
assign u_ca_in_733 = col_in_733;
assign u_ca_in_734 = col_in_734;
assign u_ca_in_735 = col_in_735;
assign u_ca_in_736 = col_in_736;
assign u_ca_in_737 = col_in_737;
assign u_ca_in_738 = col_in_738;
assign u_ca_in_739 = col_in_739;
assign u_ca_in_740 = col_in_740;
assign u_ca_in_741 = col_in_741;
assign u_ca_in_742 = col_in_742;
assign u_ca_in_743 = col_in_743;
assign u_ca_in_744 = col_in_744;
assign u_ca_in_745 = col_in_745;
assign u_ca_in_746 = col_in_746;
assign u_ca_in_747 = col_in_747;
assign u_ca_in_748 = col_in_748;
assign u_ca_in_749 = col_in_749;
assign u_ca_in_750 = col_in_750;
assign u_ca_in_751 = col_in_751;
assign u_ca_in_752 = col_in_752;
assign u_ca_in_753 = col_in_753;
assign u_ca_in_754 = col_in_754;
assign u_ca_in_755 = col_in_755;
assign u_ca_in_756 = col_in_756;
assign u_ca_in_757 = col_in_757;
assign u_ca_in_758 = col_in_758;
assign u_ca_in_759 = col_in_759;
assign u_ca_in_760 = col_in_760;
assign u_ca_in_761 = col_in_761;
assign u_ca_in_762 = col_in_762;
assign u_ca_in_763 = col_in_763;
assign u_ca_in_764 = col_in_764;
assign u_ca_in_765 = col_in_765;
assign u_ca_in_766 = col_in_766;
assign u_ca_in_767 = col_in_767;
assign u_ca_in_768 = col_in_768;
assign u_ca_in_769 = col_in_769;
assign u_ca_in_770 = col_in_770;
assign u_ca_in_771 = col_in_771;
assign u_ca_in_772 = col_in_772;
assign u_ca_in_773 = col_in_773;
assign u_ca_in_774 = col_in_774;
assign u_ca_in_775 = col_in_775;
assign u_ca_in_776 = col_in_776;
assign u_ca_in_777 = col_in_777;
assign u_ca_in_778 = col_in_778;
assign u_ca_in_779 = col_in_779;
assign u_ca_in_780 = col_in_780;
assign u_ca_in_781 = col_in_781;
assign u_ca_in_782 = col_in_782;
assign u_ca_in_783 = col_in_783;
assign u_ca_in_784 = col_in_784;
assign u_ca_in_785 = col_in_785;
assign u_ca_in_786 = col_in_786;
assign u_ca_in_787 = col_in_787;
assign u_ca_in_788 = col_in_788;
assign u_ca_in_789 = col_in_789;
assign u_ca_in_790 = col_in_790;
assign u_ca_in_791 = col_in_791;
assign u_ca_in_792 = col_in_792;
assign u_ca_in_793 = col_in_793;
assign u_ca_in_794 = col_in_794;
assign u_ca_in_795 = col_in_795;
assign u_ca_in_796 = col_in_796;
assign u_ca_in_797 = col_in_797;
assign u_ca_in_798 = col_in_798;
assign u_ca_in_799 = col_in_799;
assign u_ca_in_800 = col_in_800;
assign u_ca_in_801 = col_in_801;
assign u_ca_in_802 = col_in_802;
assign u_ca_in_803 = col_in_803;
assign u_ca_in_804 = col_in_804;
assign u_ca_in_805 = col_in_805;
assign u_ca_in_806 = col_in_806;
assign u_ca_in_807 = col_in_807;
assign u_ca_in_808 = col_in_808;
assign u_ca_in_809 = col_in_809;
assign u_ca_in_810 = col_in_810;
assign u_ca_in_811 = col_in_811;
assign u_ca_in_812 = col_in_812;
assign u_ca_in_813 = col_in_813;
assign u_ca_in_814 = col_in_814;
assign u_ca_in_815 = col_in_815;
assign u_ca_in_816 = col_in_816;
assign u_ca_in_817 = col_in_817;
assign u_ca_in_818 = col_in_818;
assign u_ca_in_819 = col_in_819;
assign u_ca_in_820 = col_in_820;
assign u_ca_in_821 = col_in_821;
assign u_ca_in_822 = col_in_822;
assign u_ca_in_823 = col_in_823;
assign u_ca_in_824 = col_in_824;
assign u_ca_in_825 = col_in_825;
assign u_ca_in_826 = col_in_826;
assign u_ca_in_827 = col_in_827;
assign u_ca_in_828 = col_in_828;
assign u_ca_in_829 = col_in_829;
assign u_ca_in_830 = col_in_830;
assign u_ca_in_831 = col_in_831;
assign u_ca_in_832 = col_in_832;
assign u_ca_in_833 = col_in_833;
assign u_ca_in_834 = col_in_834;
assign u_ca_in_835 = col_in_835;
assign u_ca_in_836 = col_in_836;
assign u_ca_in_837 = col_in_837;
assign u_ca_in_838 = col_in_838;
assign u_ca_in_839 = col_in_839;
assign u_ca_in_840 = col_in_840;
assign u_ca_in_841 = col_in_841;
assign u_ca_in_842 = col_in_842;
assign u_ca_in_843 = col_in_843;
assign u_ca_in_844 = col_in_844;
assign u_ca_in_845 = col_in_845;
assign u_ca_in_846 = col_in_846;
assign u_ca_in_847 = col_in_847;
assign u_ca_in_848 = col_in_848;
assign u_ca_in_849 = col_in_849;
assign u_ca_in_850 = col_in_850;
assign u_ca_in_851 = col_in_851;
assign u_ca_in_852 = col_in_852;
assign u_ca_in_853 = col_in_853;
assign u_ca_in_854 = col_in_854;
assign u_ca_in_855 = col_in_855;
assign u_ca_in_856 = col_in_856;
assign u_ca_in_857 = col_in_857;
assign u_ca_in_858 = col_in_858;
assign u_ca_in_859 = col_in_859;
assign u_ca_in_860 = col_in_860;
assign u_ca_in_861 = col_in_861;
assign u_ca_in_862 = col_in_862;
assign u_ca_in_863 = col_in_863;
assign u_ca_in_864 = col_in_864;
assign u_ca_in_865 = col_in_865;
assign u_ca_in_866 = col_in_866;
assign u_ca_in_867 = col_in_867;
assign u_ca_in_868 = col_in_868;
assign u_ca_in_869 = col_in_869;
assign u_ca_in_870 = col_in_870;
assign u_ca_in_871 = col_in_871;
assign u_ca_in_872 = col_in_872;
assign u_ca_in_873 = col_in_873;
assign u_ca_in_874 = col_in_874;
assign u_ca_in_875 = col_in_875;
assign u_ca_in_876 = col_in_876;
assign u_ca_in_877 = col_in_877;
assign u_ca_in_878 = col_in_878;
assign u_ca_in_879 = col_in_879;
assign u_ca_in_880 = col_in_880;
assign u_ca_in_881 = col_in_881;
assign u_ca_in_882 = col_in_882;
assign u_ca_in_883 = col_in_883;
assign u_ca_in_884 = col_in_884;
assign u_ca_in_885 = col_in_885;
assign u_ca_in_886 = col_in_886;
assign u_ca_in_887 = col_in_887;
assign u_ca_in_888 = col_in_888;
assign u_ca_in_889 = col_in_889;
assign u_ca_in_890 = col_in_890;
assign u_ca_in_891 = col_in_891;
assign u_ca_in_892 = col_in_892;
assign u_ca_in_893 = col_in_893;
assign u_ca_in_894 = col_in_894;
assign u_ca_in_895 = col_in_895;
assign u_ca_in_896 = col_in_896;
assign u_ca_in_897 = col_in_897;
assign u_ca_in_898 = col_in_898;
assign u_ca_in_899 = col_in_899;
assign u_ca_in_900 = col_in_900;
assign u_ca_in_901 = col_in_901;
assign u_ca_in_902 = col_in_902;
assign u_ca_in_903 = col_in_903;
assign u_ca_in_904 = col_in_904;
assign u_ca_in_905 = col_in_905;
assign u_ca_in_906 = col_in_906;
assign u_ca_in_907 = col_in_907;
assign u_ca_in_908 = col_in_908;
assign u_ca_in_909 = col_in_909;
assign u_ca_in_910 = col_in_910;
assign u_ca_in_911 = col_in_911;
assign u_ca_in_912 = col_in_912;
assign u_ca_in_913 = col_in_913;
assign u_ca_in_914 = col_in_914;
assign u_ca_in_915 = col_in_915;
assign u_ca_in_916 = col_in_916;
assign u_ca_in_917 = col_in_917;
assign u_ca_in_918 = col_in_918;
assign u_ca_in_919 = col_in_919;
assign u_ca_in_920 = col_in_920;
assign u_ca_in_921 = col_in_921;
assign u_ca_in_922 = col_in_922;
assign u_ca_in_923 = col_in_923;
assign u_ca_in_924 = col_in_924;
assign u_ca_in_925 = col_in_925;
assign u_ca_in_926 = col_in_926;
assign u_ca_in_927 = col_in_927;
assign u_ca_in_928 = col_in_928;
assign u_ca_in_929 = col_in_929;
assign u_ca_in_930 = col_in_930;
assign u_ca_in_931 = col_in_931;
assign u_ca_in_932 = col_in_932;
assign u_ca_in_933 = col_in_933;
assign u_ca_in_934 = col_in_934;
assign u_ca_in_935 = col_in_935;
assign u_ca_in_936 = col_in_936;
assign u_ca_in_937 = col_in_937;
assign u_ca_in_938 = col_in_938;
assign u_ca_in_939 = col_in_939;
assign u_ca_in_940 = col_in_940;
assign u_ca_in_941 = col_in_941;
assign u_ca_in_942 = col_in_942;
assign u_ca_in_943 = col_in_943;
assign u_ca_in_944 = col_in_944;
assign u_ca_in_945 = col_in_945;
assign u_ca_in_946 = col_in_946;
assign u_ca_in_947 = col_in_947;
assign u_ca_in_948 = col_in_948;
assign u_ca_in_949 = col_in_949;
assign u_ca_in_950 = col_in_950;
assign u_ca_in_951 = col_in_951;
assign u_ca_in_952 = col_in_952;
assign u_ca_in_953 = col_in_953;
assign u_ca_in_954 = col_in_954;
assign u_ca_in_955 = col_in_955;
assign u_ca_in_956 = col_in_956;
assign u_ca_in_957 = col_in_957;
assign u_ca_in_958 = col_in_958;
assign u_ca_in_959 = col_in_959;
assign u_ca_in_960 = col_in_960;
assign u_ca_in_961 = col_in_961;
assign u_ca_in_962 = col_in_962;
assign u_ca_in_963 = col_in_963;
assign u_ca_in_964 = col_in_964;
assign u_ca_in_965 = col_in_965;
assign u_ca_in_966 = col_in_966;
assign u_ca_in_967 = col_in_967;
assign u_ca_in_968 = col_in_968;
assign u_ca_in_969 = col_in_969;
assign u_ca_in_970 = col_in_970;
assign u_ca_in_971 = col_in_971;
assign u_ca_in_972 = col_in_972;
assign u_ca_in_973 = col_in_973;
assign u_ca_in_974 = col_in_974;
assign u_ca_in_975 = col_in_975;
assign u_ca_in_976 = col_in_976;
assign u_ca_in_977 = col_in_977;
assign u_ca_in_978 = col_in_978;
assign u_ca_in_979 = col_in_979;
assign u_ca_in_980 = col_in_980;
assign u_ca_in_981 = col_in_981;
assign u_ca_in_982 = col_in_982;
assign u_ca_in_983 = col_in_983;
assign u_ca_in_984 = col_in_984;
assign u_ca_in_985 = col_in_985;
assign u_ca_in_986 = col_in_986;
assign u_ca_in_987 = col_in_987;
assign u_ca_in_988 = col_in_988;
assign u_ca_in_989 = col_in_989;
assign u_ca_in_990 = col_in_990;
assign u_ca_in_991 = col_in_991;
assign u_ca_in_992 = col_in_992;
assign u_ca_in_993 = col_in_993;
assign u_ca_in_994 = col_in_994;
assign u_ca_in_995 = col_in_995;
assign u_ca_in_996 = col_in_996;
assign u_ca_in_997 = col_in_997;
assign u_ca_in_998 = col_in_998;
assign u_ca_in_999 = col_in_999;
assign u_ca_in_1000 = col_in_1000;
assign u_ca_in_1001 = col_in_1001;
assign u_ca_in_1002 = col_in_1002;
assign u_ca_in_1003 = col_in_1003;
assign u_ca_in_1004 = col_in_1004;
assign u_ca_in_1005 = col_in_1005;
assign u_ca_in_1006 = col_in_1006;
assign u_ca_in_1007 = col_in_1007;
assign u_ca_in_1008 = col_in_1008;
assign u_ca_in_1009 = col_in_1009;
assign u_ca_in_1010 = col_in_1010;
assign u_ca_in_1011 = col_in_1011;
assign u_ca_in_1012 = col_in_1012;
assign u_ca_in_1013 = col_in_1013;
assign u_ca_in_1014 = col_in_1014;
assign u_ca_in_1015 = col_in_1015;
assign u_ca_in_1016 = col_in_1016;
assign u_ca_in_1017 = col_in_1017;
assign u_ca_in_1018 = col_in_1018;
assign u_ca_in_1019 = col_in_1019;
assign u_ca_in_1020 = col_in_1020;
assign u_ca_in_1021 = col_in_1021;
assign u_ca_in_1022 = col_in_1022;
assign u_ca_in_1023 = col_in_1023;

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_6_4 u_ca_6_4_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_6_4 u_ca_6_4_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_6_4 u_ca_6_4_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_6_4 u_ca_6_4_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_6_4 u_ca_6_4_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_6_4 u_ca_6_4_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_6_4 u_ca_6_4_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_6_4 u_ca_6_4_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_6_4 u_ca_6_4_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_6_4 u_ca_6_4_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_6_4 u_ca_6_4_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_6_4 u_ca_6_4_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_6_4 u_ca_6_4_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_6_4 u_ca_6_4_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_6_4 u_ca_6_4_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_6_4 u_ca_6_4_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_6_4 u_ca_6_4_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_6_4 u_ca_6_4_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_6_4 u_ca_6_4_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_6_4 u_ca_6_4_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_6_4 u_ca_6_4_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_6_4 u_ca_6_4_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_6_4 u_ca_6_4_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_6_4 u_ca_6_4_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_6_4 u_ca_6_4_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_6_4 u_ca_6_4_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_6_4 u_ca_6_4_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_6_4 u_ca_6_4_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_6_4 u_ca_6_4_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_6_4 u_ca_6_4_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_6_4 u_ca_6_4_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_6_4 u_ca_6_4_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_6_4 u_ca_6_4_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_6_4 u_ca_6_4_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_6_4 u_ca_6_4_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_6_4 u_ca_6_4_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_6_4 u_ca_6_4_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_6_4 u_ca_6_4_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_6_4 u_ca_6_4_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_6_4 u_ca_6_4_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_6_4 u_ca_6_4_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_6_4 u_ca_6_4_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_6_4 u_ca_6_4_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_6_4 u_ca_6_4_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_6_4 u_ca_6_4_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_6_4 u_ca_6_4_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_6_4 u_ca_6_4_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_6_4 u_ca_6_4_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_6_4 u_ca_6_4_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_6_4 u_ca_6_4_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_6_4 u_ca_6_4_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_6_4 u_ca_6_4_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_6_4 u_ca_6_4_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_6_4 u_ca_6_4_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_6_4 u_ca_6_4_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_6_4 u_ca_6_4_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_6_4 u_ca_6_4_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_6_4 u_ca_6_4_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_6_4 u_ca_6_4_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_6_4 u_ca_6_4_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_6_4 u_ca_6_4_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_6_4 u_ca_6_4_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_6_4 u_ca_6_4_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_6_4 u_ca_6_4_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_6_4 u_ca_6_4_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_6_4 u_ca_6_4_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_6_4 u_ca_6_4_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_6_4 u_ca_6_4_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_6_4 u_ca_6_4_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_6_4 u_ca_6_4_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_6_4 u_ca_6_4_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_6_4 u_ca_6_4_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_6_4 u_ca_6_4_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_6_4 u_ca_6_4_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_6_4 u_ca_6_4_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_6_4 u_ca_6_4_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_6_4 u_ca_6_4_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_6_4 u_ca_6_4_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_6_4 u_ca_6_4_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_6_4 u_ca_6_4_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_6_4 u_ca_6_4_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_6_4 u_ca_6_4_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_6_4 u_ca_6_4_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_6_4 u_ca_6_4_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_6_4 u_ca_6_4_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_6_4 u_ca_6_4_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_6_4 u_ca_6_4_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_6_4 u_ca_6_4_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_6_4 u_ca_6_4_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_6_4 u_ca_6_4_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_6_4 u_ca_6_4_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_6_4 u_ca_6_4_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_6_4 u_ca_6_4_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_6_4 u_ca_6_4_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_6_4 u_ca_6_4_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_6_4 u_ca_6_4_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_6_4 u_ca_6_4_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_6_4 u_ca_6_4_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_6_4 u_ca_6_4_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_6_4 u_ca_6_4_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_6_4 u_ca_6_4_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_6_4 u_ca_6_4_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_6_4 u_ca_6_4_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_6_4 u_ca_6_4_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_6_4 u_ca_6_4_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_6_4 u_ca_6_4_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_6_4 u_ca_6_4_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_6_4 u_ca_6_4_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_6_4 u_ca_6_4_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_6_4 u_ca_6_4_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_6_4 u_ca_6_4_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_6_4 u_ca_6_4_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_6_4 u_ca_6_4_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_6_4 u_ca_6_4_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_6_4 u_ca_6_4_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_6_4 u_ca_6_4_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_6_4 u_ca_6_4_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_6_4 u_ca_6_4_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_6_4 u_ca_6_4_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_6_4 u_ca_6_4_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_6_4 u_ca_6_4_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_6_4 u_ca_6_4_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_6_4 u_ca_6_4_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_6_4 u_ca_6_4_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_6_4 u_ca_6_4_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_6_4 u_ca_6_4_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_6_4 u_ca_6_4_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_6_4 u_ca_6_4_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_6_4 u_ca_6_4_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_6_4 u_ca_6_4_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_6_4 u_ca_6_4_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_6_4 u_ca_6_4_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_6_4 u_ca_6_4_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_6_4 u_ca_6_4_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_6_4 u_ca_6_4_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_6_4 u_ca_6_4_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_6_4 u_ca_6_4_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_6_4 u_ca_6_4_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_6_4 u_ca_6_4_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_6_4 u_ca_6_4_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_6_4 u_ca_6_4_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_6_4 u_ca_6_4_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_6_4 u_ca_6_4_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_6_4 u_ca_6_4_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_6_4 u_ca_6_4_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_6_4 u_ca_6_4_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_6_4 u_ca_6_4_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_6_4 u_ca_6_4_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_6_4 u_ca_6_4_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_6_4 u_ca_6_4_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_6_4 u_ca_6_4_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_6_4 u_ca_6_4_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_6_4 u_ca_6_4_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_6_4 u_ca_6_4_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_6_4 u_ca_6_4_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_6_4 u_ca_6_4_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_6_4 u_ca_6_4_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_6_4 u_ca_6_4_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_6_4 u_ca_6_4_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_6_4 u_ca_6_4_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_6_4 u_ca_6_4_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_6_4 u_ca_6_4_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_6_4 u_ca_6_4_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_6_4 u_ca_6_4_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_6_4 u_ca_6_4_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_6_4 u_ca_6_4_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_6_4 u_ca_6_4_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_6_4 u_ca_6_4_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_6_4 u_ca_6_4_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_6_4 u_ca_6_4_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_6_4 u_ca_6_4_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_6_4 u_ca_6_4_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_6_4 u_ca_6_4_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_6_4 u_ca_6_4_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_6_4 u_ca_6_4_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_6_4 u_ca_6_4_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_6_4 u_ca_6_4_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_6_4 u_ca_6_4_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_6_4 u_ca_6_4_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_6_4 u_ca_6_4_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_6_4 u_ca_6_4_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_6_4 u_ca_6_4_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_6_4 u_ca_6_4_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_6_4 u_ca_6_4_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_6_4 u_ca_6_4_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_6_4 u_ca_6_4_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_6_4 u_ca_6_4_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_6_4 u_ca_6_4_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_6_4 u_ca_6_4_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_6_4 u_ca_6_4_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_6_4 u_ca_6_4_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_6_4 u_ca_6_4_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_6_4 u_ca_6_4_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_6_4 u_ca_6_4_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_6_4 u_ca_6_4_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_6_4 u_ca_6_4_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_6_4 u_ca_6_4_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_6_4 u_ca_6_4_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_6_4 u_ca_6_4_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_6_4 u_ca_6_4_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_6_4 u_ca_6_4_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_6_4 u_ca_6_4_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_6_4 u_ca_6_4_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_6_4 u_ca_6_4_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_6_4 u_ca_6_4_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_6_4 u_ca_6_4_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_6_4 u_ca_6_4_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_6_4 u_ca_6_4_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_6_4 u_ca_6_4_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_6_4 u_ca_6_4_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_6_4 u_ca_6_4_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_6_4 u_ca_6_4_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_6_4 u_ca_6_4_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_6_4 u_ca_6_4_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_6_4 u_ca_6_4_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_6_4 u_ca_6_4_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_6_4 u_ca_6_4_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_6_4 u_ca_6_4_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_6_4 u_ca_6_4_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_6_4 u_ca_6_4_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_6_4 u_ca_6_4_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_6_4 u_ca_6_4_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_6_4 u_ca_6_4_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_6_4 u_ca_6_4_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_6_4 u_ca_6_4_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_6_4 u_ca_6_4_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_6_4 u_ca_6_4_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_6_4 u_ca_6_4_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_6_4 u_ca_6_4_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_6_4 u_ca_6_4_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_6_4 u_ca_6_4_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_6_4 u_ca_6_4_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_6_4 u_ca_6_4_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_6_4 u_ca_6_4_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_6_4 u_ca_6_4_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_6_4 u_ca_6_4_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_6_4 u_ca_6_4_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_6_4 u_ca_6_4_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_6_4 u_ca_6_4_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_6_4 u_ca_6_4_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_6_4 u_ca_6_4_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_6_4 u_ca_6_4_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_6_4 u_ca_6_4_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_6_4 u_ca_6_4_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_6_4 u_ca_6_4_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_6_4 u_ca_6_4_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_6_4 u_ca_6_4_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_6_4 u_ca_6_4_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_6_4 u_ca_6_4_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_6_4 u_ca_6_4_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_6_4 u_ca_6_4_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_6_4 u_ca_6_4_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_6_4 u_ca_6_4_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_6_4 u_ca_6_4_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_6_4 u_ca_6_4_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_6_4 u_ca_6_4_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_6_4 u_ca_6_4_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_6_4 u_ca_6_4_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_6_4 u_ca_6_4_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_6_4 u_ca_6_4_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_6_4 u_ca_6_4_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_6_4 u_ca_6_4_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_6_4 u_ca_6_4_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_6_4 u_ca_6_4_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_6_4 u_ca_6_4_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_6_4 u_ca_6_4_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_6_4 u_ca_6_4_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_6_4 u_ca_6_4_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_6_4 u_ca_6_4_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_6_4 u_ca_6_4_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_6_4 u_ca_6_4_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_6_4 u_ca_6_4_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_6_4 u_ca_6_4_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_6_4 u_ca_6_4_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_6_4 u_ca_6_4_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_6_4 u_ca_6_4_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_6_4 u_ca_6_4_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_6_4 u_ca_6_4_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_6_4 u_ca_6_4_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_6_4 u_ca_6_4_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_6_4 u_ca_6_4_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_6_4 u_ca_6_4_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_6_4 u_ca_6_4_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_6_4 u_ca_6_4_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_6_4 u_ca_6_4_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_6_4 u_ca_6_4_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_6_4 u_ca_6_4_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_6_4 u_ca_6_4_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_6_4 u_ca_6_4_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_6_4 u_ca_6_4_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_6_4 u_ca_6_4_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_6_4 u_ca_6_4_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_6_4 u_ca_6_4_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_6_4 u_ca_6_4_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_6_4 u_ca_6_4_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_6_4 u_ca_6_4_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_6_4 u_ca_6_4_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_6_4 u_ca_6_4_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_6_4 u_ca_6_4_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_6_4 u_ca_6_4_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_6_4 u_ca_6_4_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_6_4 u_ca_6_4_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_6_4 u_ca_6_4_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_6_4 u_ca_6_4_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_6_4 u_ca_6_4_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_6_4 u_ca_6_4_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_6_4 u_ca_6_4_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_6_4 u_ca_6_4_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_6_4 u_ca_6_4_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_6_4 u_ca_6_4_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_6_4 u_ca_6_4_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_6_4 u_ca_6_4_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_6_4 u_ca_6_4_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_6_4 u_ca_6_4_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_6_4 u_ca_6_4_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_6_4 u_ca_6_4_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_6_4 u_ca_6_4_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_6_4 u_ca_6_4_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_6_4 u_ca_6_4_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_6_4 u_ca_6_4_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_6_4 u_ca_6_4_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_6_4 u_ca_6_4_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_6_4 u_ca_6_4_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_6_4 u_ca_6_4_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_6_4 u_ca_6_4_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_6_4 u_ca_6_4_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_6_4 u_ca_6_4_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_6_4 u_ca_6_4_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_6_4 u_ca_6_4_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_6_4 u_ca_6_4_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_6_4 u_ca_6_4_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_6_4 u_ca_6_4_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_6_4 u_ca_6_4_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_6_4 u_ca_6_4_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_6_4 u_ca_6_4_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_6_4 u_ca_6_4_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_6_4 u_ca_6_4_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_6_4 u_ca_6_4_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_6_4 u_ca_6_4_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_6_4 u_ca_6_4_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_6_4 u_ca_6_4_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_6_4 u_ca_6_4_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_6_4 u_ca_6_4_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_6_4 u_ca_6_4_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_6_4 u_ca_6_4_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_6_4 u_ca_6_4_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_6_4 u_ca_6_4_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_6_4 u_ca_6_4_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_6_4 u_ca_6_4_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_6_4 u_ca_6_4_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_6_4 u_ca_6_4_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_6_4 u_ca_6_4_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_6_4 u_ca_6_4_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_6_4 u_ca_6_4_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_6_4 u_ca_6_4_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_6_4 u_ca_6_4_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_6_4 u_ca_6_4_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_6_4 u_ca_6_4_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_6_4 u_ca_6_4_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_6_4 u_ca_6_4_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_6_4 u_ca_6_4_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_6_4 u_ca_6_4_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_6_4 u_ca_6_4_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_6_4 u_ca_6_4_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_6_4 u_ca_6_4_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_6_4 u_ca_6_4_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_6_4 u_ca_6_4_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_6_4 u_ca_6_4_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_6_4 u_ca_6_4_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_6_4 u_ca_6_4_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_6_4 u_ca_6_4_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_6_4 u_ca_6_4_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_6_4 u_ca_6_4_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_6_4 u_ca_6_4_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_6_4 u_ca_6_4_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_6_4 u_ca_6_4_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_6_4 u_ca_6_4_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_6_4 u_ca_6_4_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_6_4 u_ca_6_4_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_6_4 u_ca_6_4_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_6_4 u_ca_6_4_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_6_4 u_ca_6_4_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_6_4 u_ca_6_4_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_6_4 u_ca_6_4_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_6_4 u_ca_6_4_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_6_4 u_ca_6_4_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_6_4 u_ca_6_4_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_6_4 u_ca_6_4_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_6_4 u_ca_6_4_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_6_4 u_ca_6_4_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_6_4 u_ca_6_4_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_6_4 u_ca_6_4_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_6_4 u_ca_6_4_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_6_4 u_ca_6_4_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_6_4 u_ca_6_4_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_6_4 u_ca_6_4_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_6_4 u_ca_6_4_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_6_4 u_ca_6_4_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_6_4 u_ca_6_4_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_6_4 u_ca_6_4_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_6_4 u_ca_6_4_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_6_4 u_ca_6_4_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_6_4 u_ca_6_4_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_6_4 u_ca_6_4_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_6_4 u_ca_6_4_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_6_4 u_ca_6_4_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_6_4 u_ca_6_4_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_6_4 u_ca_6_4_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_6_4 u_ca_6_4_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_6_4 u_ca_6_4_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_6_4 u_ca_6_4_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_6_4 u_ca_6_4_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_6_4 u_ca_6_4_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_6_4 u_ca_6_4_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_6_4 u_ca_6_4_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_6_4 u_ca_6_4_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_6_4 u_ca_6_4_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_6_4 u_ca_6_4_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_6_4 u_ca_6_4_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_6_4 u_ca_6_4_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_6_4 u_ca_6_4_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_6_4 u_ca_6_4_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_6_4 u_ca_6_4_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_6_4 u_ca_6_4_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_6_4 u_ca_6_4_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_6_4 u_ca_6_4_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_6_4 u_ca_6_4_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_6_4 u_ca_6_4_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_6_4 u_ca_6_4_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_6_4 u_ca_6_4_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_6_4 u_ca_6_4_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_6_4 u_ca_6_4_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_6_4 u_ca_6_4_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_6_4 u_ca_6_4_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_6_4 u_ca_6_4_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_6_4 u_ca_6_4_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_6_4 u_ca_6_4_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_6_4 u_ca_6_4_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_6_4 u_ca_6_4_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_6_4 u_ca_6_4_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_6_4 u_ca_6_4_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_6_4 u_ca_6_4_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_6_4 u_ca_6_4_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_6_4 u_ca_6_4_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_6_4 u_ca_6_4_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_6_4 u_ca_6_4_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_6_4 u_ca_6_4_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_6_4 u_ca_6_4_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_6_4 u_ca_6_4_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_6_4 u_ca_6_4_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_6_4 u_ca_6_4_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_6_4 u_ca_6_4_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_6_4 u_ca_6_4_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_6_4 u_ca_6_4_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_6_4 u_ca_6_4_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_6_4 u_ca_6_4_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_6_4 u_ca_6_4_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_6_4 u_ca_6_4_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_6_4 u_ca_6_4_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_6_4 u_ca_6_4_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_6_4 u_ca_6_4_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_6_4 u_ca_6_4_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_6_4 u_ca_6_4_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_6_4 u_ca_6_4_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_6_4 u_ca_6_4_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_6_4 u_ca_6_4_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_6_4 u_ca_6_4_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_6_4 u_ca_6_4_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_6_4 u_ca_6_4_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_6_4 u_ca_6_4_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_6_4 u_ca_6_4_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_6_4 u_ca_6_4_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_6_4 u_ca_6_4_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_6_4 u_ca_6_4_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_6_4 u_ca_6_4_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_6_4 u_ca_6_4_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_6_4 u_ca_6_4_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_6_4 u_ca_6_4_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_6_4 u_ca_6_4_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_6_4 u_ca_6_4_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_6_4 u_ca_6_4_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_6_4 u_ca_6_4_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_6_4 u_ca_6_4_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_6_4 u_ca_6_4_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_6_4 u_ca_6_4_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_6_4 u_ca_6_4_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_6_4 u_ca_6_4_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_6_4 u_ca_6_4_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_6_4 u_ca_6_4_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_6_4 u_ca_6_4_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_6_4 u_ca_6_4_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_6_4 u_ca_6_4_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_6_4 u_ca_6_4_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_6_4 u_ca_6_4_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_6_4 u_ca_6_4_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_6_4 u_ca_6_4_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_6_4 u_ca_6_4_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_6_4 u_ca_6_4_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_6_4 u_ca_6_4_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_6_4 u_ca_6_4_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_6_4 u_ca_6_4_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_6_4 u_ca_6_4_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_6_4 u_ca_6_4_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_6_4 u_ca_6_4_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_6_4 u_ca_6_4_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_6_4 u_ca_6_4_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_6_4 u_ca_6_4_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_6_4 u_ca_6_4_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_6_4 u_ca_6_4_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_6_4 u_ca_6_4_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_6_4 u_ca_6_4_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_6_4 u_ca_6_4_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_6_4 u_ca_6_4_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_6_4 u_ca_6_4_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_6_4 u_ca_6_4_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_6_4 u_ca_6_4_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_6_4 u_ca_6_4_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_6_4 u_ca_6_4_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_6_4 u_ca_6_4_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_6_4 u_ca_6_4_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_6_4 u_ca_6_4_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_6_4 u_ca_6_4_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_6_4 u_ca_6_4_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_6_4 u_ca_6_4_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_6_4 u_ca_6_4_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_6_4 u_ca_6_4_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_6_4 u_ca_6_4_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_6_4 u_ca_6_4_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_6_4 u_ca_6_4_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_6_4 u_ca_6_4_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_6_4 u_ca_6_4_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_6_4 u_ca_6_4_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_6_4 u_ca_6_4_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_6_4 u_ca_6_4_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_6_4 u_ca_6_4_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_6_4 u_ca_6_4_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_6_4 u_ca_6_4_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_6_4 u_ca_6_4_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_6_4 u_ca_6_4_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_6_4 u_ca_6_4_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_6_4 u_ca_6_4_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_6_4 u_ca_6_4_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_6_4 u_ca_6_4_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_6_4 u_ca_6_4_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_6_4 u_ca_6_4_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_6_4 u_ca_6_4_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_6_4 u_ca_6_4_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_6_4 u_ca_6_4_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_6_4 u_ca_6_4_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_6_4 u_ca_6_4_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_6_4 u_ca_6_4_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_6_4 u_ca_6_4_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_6_4 u_ca_6_4_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_6_4 u_ca_6_4_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_6_4 u_ca_6_4_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_6_4 u_ca_6_4_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_6_4 u_ca_6_4_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_6_4 u_ca_6_4_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_6_4 u_ca_6_4_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_6_4 u_ca_6_4_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_6_4 u_ca_6_4_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_6_4 u_ca_6_4_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_6_4 u_ca_6_4_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_6_4 u_ca_6_4_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_6_4 u_ca_6_4_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_6_4 u_ca_6_4_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_6_4 u_ca_6_4_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_6_4 u_ca_6_4_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_6_4 u_ca_6_4_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_6_4 u_ca_6_4_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_6_4 u_ca_6_4_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_6_4 u_ca_6_4_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_6_4 u_ca_6_4_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_6_4 u_ca_6_4_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_6_4 u_ca_6_4_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_6_4 u_ca_6_4_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_6_4 u_ca_6_4_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_6_4 u_ca_6_4_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_6_4 u_ca_6_4_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_6_4 u_ca_6_4_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_6_4 u_ca_6_4_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_6_4 u_ca_6_4_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_6_4 u_ca_6_4_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_6_4 u_ca_6_4_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_6_4 u_ca_6_4_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_6_4 u_ca_6_4_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_6_4 u_ca_6_4_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_6_4 u_ca_6_4_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_6_4 u_ca_6_4_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_6_4 u_ca_6_4_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_6_4 u_ca_6_4_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_6_4 u_ca_6_4_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_6_4 u_ca_6_4_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_6_4 u_ca_6_4_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_6_4 u_ca_6_4_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_6_4 u_ca_6_4_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_6_4 u_ca_6_4_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_6_4 u_ca_6_4_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_6_4 u_ca_6_4_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_6_4 u_ca_6_4_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_6_4 u_ca_6_4_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_6_4 u_ca_6_4_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_6_4 u_ca_6_4_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_6_4 u_ca_6_4_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_6_4 u_ca_6_4_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_6_4 u_ca_6_4_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_6_4 u_ca_6_4_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_6_4 u_ca_6_4_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_6_4 u_ca_6_4_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_6_4 u_ca_6_4_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_6_4 u_ca_6_4_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_6_4 u_ca_6_4_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_6_4 u_ca_6_4_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_6_4 u_ca_6_4_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_6_4 u_ca_6_4_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_6_4 u_ca_6_4_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_6_4 u_ca_6_4_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_6_4 u_ca_6_4_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_6_4 u_ca_6_4_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_6_4 u_ca_6_4_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_6_4 u_ca_6_4_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_6_4 u_ca_6_4_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_6_4 u_ca_6_4_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_6_4 u_ca_6_4_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_6_4 u_ca_6_4_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_6_4 u_ca_6_4_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_6_4 u_ca_6_4_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_6_4 u_ca_6_4_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_6_4 u_ca_6_4_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_6_4 u_ca_6_4_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_6_4 u_ca_6_4_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_6_4 u_ca_6_4_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_6_4 u_ca_6_4_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_6_4 u_ca_6_4_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_6_4 u_ca_6_4_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_6_4 u_ca_6_4_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_6_4 u_ca_6_4_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_6_4 u_ca_6_4_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_6_4 u_ca_6_4_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_6_4 u_ca_6_4_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_6_4 u_ca_6_4_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_6_4 u_ca_6_4_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_6_4 u_ca_6_4_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_6_4 u_ca_6_4_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_6_4 u_ca_6_4_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_6_4 u_ca_6_4_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_6_4 u_ca_6_4_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_6_4 u_ca_6_4_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_6_4 u_ca_6_4_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_6_4 u_ca_6_4_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_6_4 u_ca_6_4_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_6_4 u_ca_6_4_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_6_4 u_ca_6_4_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_6_4 u_ca_6_4_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_6_4 u_ca_6_4_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_6_4 u_ca_6_4_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_6_4 u_ca_6_4_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_6_4 u_ca_6_4_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_6_4 u_ca_6_4_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_6_4 u_ca_6_4_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_6_4 u_ca_6_4_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_6_4 u_ca_6_4_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_6_4 u_ca_6_4_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_6_4 u_ca_6_4_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_6_4 u_ca_6_4_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_6_4 u_ca_6_4_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_6_4 u_ca_6_4_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_6_4 u_ca_6_4_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_6_4 u_ca_6_4_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_6_4 u_ca_6_4_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_6_4 u_ca_6_4_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_6_4 u_ca_6_4_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_6_4 u_ca_6_4_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_6_4 u_ca_6_4_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_6_4 u_ca_6_4_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_6_4 u_ca_6_4_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_6_4 u_ca_6_4_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_6_4 u_ca_6_4_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_6_4 u_ca_6_4_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_6_4 u_ca_6_4_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_6_4 u_ca_6_4_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_6_4 u_ca_6_4_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_6_4 u_ca_6_4_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_6_4 u_ca_6_4_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_6_4 u_ca_6_4_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_6_4 u_ca_6_4_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_6_4 u_ca_6_4_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_6_4 u_ca_6_4_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_6_4 u_ca_6_4_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_6_4 u_ca_6_4_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_6_4 u_ca_6_4_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_6_4 u_ca_6_4_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_6_4 u_ca_6_4_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_6_4 u_ca_6_4_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_6_4 u_ca_6_4_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_6_4 u_ca_6_4_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_6_4 u_ca_6_4_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_6_4 u_ca_6_4_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_6_4 u_ca_6_4_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_6_4 u_ca_6_4_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_6_4 u_ca_6_4_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_6_4 u_ca_6_4_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_6_4 u_ca_6_4_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_6_4 u_ca_6_4_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_6_4 u_ca_6_4_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_6_4 u_ca_6_4_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_6_4 u_ca_6_4_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_6_4 u_ca_6_4_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_6_4 u_ca_6_4_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_6_4 u_ca_6_4_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_6_4 u_ca_6_4_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_6_4 u_ca_6_4_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_6_4 u_ca_6_4_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_6_4 u_ca_6_4_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_6_4 u_ca_6_4_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_6_4 u_ca_6_4_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_6_4 u_ca_6_4_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_6_4 u_ca_6_4_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_6_4 u_ca_6_4_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_6_4 u_ca_6_4_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_6_4 u_ca_6_4_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_6_4 u_ca_6_4_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_6_4 u_ca_6_4_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_6_4 u_ca_6_4_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_6_4 u_ca_6_4_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_6_4 u_ca_6_4_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_6_4 u_ca_6_4_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_6_4 u_ca_6_4_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_6_4 u_ca_6_4_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_6_4 u_ca_6_4_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_6_4 u_ca_6_4_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_6_4 u_ca_6_4_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_6_4 u_ca_6_4_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_6_4 u_ca_6_4_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_6_4 u_ca_6_4_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_6_4 u_ca_6_4_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_6_4 u_ca_6_4_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_6_4 u_ca_6_4_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_6_4 u_ca_6_4_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_6_4 u_ca_6_4_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_6_4 u_ca_6_4_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_6_4 u_ca_6_4_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_6_4 u_ca_6_4_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_6_4 u_ca_6_4_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_6_4 u_ca_6_4_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_6_4 u_ca_6_4_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_6_4 u_ca_6_4_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_6_4 u_ca_6_4_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_6_4 u_ca_6_4_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_6_4 u_ca_6_4_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_6_4 u_ca_6_4_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_6_4 u_ca_6_4_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_6_4 u_ca_6_4_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_6_4 u_ca_6_4_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_6_4 u_ca_6_4_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_6_4 u_ca_6_4_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_6_4 u_ca_6_4_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_6_4 u_ca_6_4_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_6_4 u_ca_6_4_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_6_4 u_ca_6_4_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_6_4 u_ca_6_4_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_6_4 u_ca_6_4_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_6_4 u_ca_6_4_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_6_4 u_ca_6_4_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_6_4 u_ca_6_4_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_6_4 u_ca_6_4_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_6_4 u_ca_6_4_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_6_4 u_ca_6_4_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_6_4 u_ca_6_4_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_6_4 u_ca_6_4_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_6_4 u_ca_6_4_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_6_4 u_ca_6_4_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_6_4 u_ca_6_4_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_6_4 u_ca_6_4_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_6_4 u_ca_6_4_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_6_4 u_ca_6_4_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_6_4 u_ca_6_4_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_6_4 u_ca_6_4_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_6_4 u_ca_6_4_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_6_4 u_ca_6_4_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_6_4 u_ca_6_4_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_6_4 u_ca_6_4_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_6_4 u_ca_6_4_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_6_4 u_ca_6_4_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_6_4 u_ca_6_4_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_6_4 u_ca_6_4_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_6_4 u_ca_6_4_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_6_4 u_ca_6_4_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_6_4 u_ca_6_4_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_6_4 u_ca_6_4_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_6_4 u_ca_6_4_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_6_4 u_ca_6_4_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_6_4 u_ca_6_4_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_6_4 u_ca_6_4_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_6_4 u_ca_6_4_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_6_4 u_ca_6_4_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_6_4 u_ca_6_4_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_6_4 u_ca_6_4_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_6_4 u_ca_6_4_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_6_4 u_ca_6_4_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_6_4 u_ca_6_4_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_6_4 u_ca_6_4_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_6_4 u_ca_6_4_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_6_4 u_ca_6_4_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_6_4 u_ca_6_4_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_6_4 u_ca_6_4_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_6_4 u_ca_6_4_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_6_4 u_ca_6_4_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_6_4 u_ca_6_4_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_6_4 u_ca_6_4_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_6_4 u_ca_6_4_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_6_4 u_ca_6_4_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_6_4 u_ca_6_4_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_6_4 u_ca_6_4_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_6_4 u_ca_6_4_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_6_4 u_ca_6_4_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_6_4 u_ca_6_4_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_6_4 u_ca_6_4_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_6_4 u_ca_6_4_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_6_4 u_ca_6_4_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_6_4 u_ca_6_4_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_6_4 u_ca_6_4_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_6_4 u_ca_6_4_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_6_4 u_ca_6_4_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_6_4 u_ca_6_4_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_6_4 u_ca_6_4_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_6_4 u_ca_6_4_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_6_4 u_ca_6_4_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_6_4 u_ca_6_4_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_6_4 u_ca_6_4_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_6_4 u_ca_6_4_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_6_4 u_ca_6_4_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_6_4 u_ca_6_4_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_6_4 u_ca_6_4_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_6_4 u_ca_6_4_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_6_4 u_ca_6_4_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_6_4 u_ca_6_4_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_6_4 u_ca_6_4_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_6_4 u_ca_6_4_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_6_4 u_ca_6_4_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_6_4 u_ca_6_4_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_6_4 u_ca_6_4_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_6_4 u_ca_6_4_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_6_4 u_ca_6_4_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_6_4 u_ca_6_4_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_6_4 u_ca_6_4_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_6_4 u_ca_6_4_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_6_4 u_ca_6_4_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_6_4 u_ca_6_4_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_6_4 u_ca_6_4_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_6_4 u_ca_6_4_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_6_4 u_ca_6_4_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_6_4 u_ca_6_4_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_6_4 u_ca_6_4_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_6_4 u_ca_6_4_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_6_4 u_ca_6_4_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_6_4 u_ca_6_4_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_6_4 u_ca_6_4_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_6_4 u_ca_6_4_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_6_4 u_ca_6_4_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_6_4 u_ca_6_4_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_6_4 u_ca_6_4_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_6_4 u_ca_6_4_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_6_4 u_ca_6_4_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_6_4 u_ca_6_4_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_6_4 u_ca_6_4_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_6_4 u_ca_6_4_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_6_4 u_ca_6_4_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_6_4 u_ca_6_4_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_6_4 u_ca_6_4_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_6_4 u_ca_6_4_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_6_4 u_ca_6_4_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_6_4 u_ca_6_4_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_6_4 u_ca_6_4_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_6_4 u_ca_6_4_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_6_4 u_ca_6_4_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_6_4 u_ca_6_4_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_6_4 u_ca_6_4_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_6_4 u_ca_6_4_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_6_4 u_ca_6_4_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_6_4 u_ca_6_4_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_6_4 u_ca_6_4_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_6_4 u_ca_6_4_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_6_4 u_ca_6_4_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_6_4 u_ca_6_4_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_6_4 u_ca_6_4_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_6_4 u_ca_6_4_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_6_4 u_ca_6_4_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_6_4 u_ca_6_4_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_6_4 u_ca_6_4_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_6_4 u_ca_6_4_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_6_4 u_ca_6_4_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_6_4 u_ca_6_4_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_6_4 u_ca_6_4_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_6_4 u_ca_6_4_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_6_4 u_ca_6_4_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_6_4 u_ca_6_4_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_6_4 u_ca_6_4_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_6_4 u_ca_6_4_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_6_4 u_ca_6_4_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_6_4 u_ca_6_4_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_6_4 u_ca_6_4_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_6_4 u_ca_6_4_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_6_4 u_ca_6_4_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_6_4 u_ca_6_4_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_6_4 u_ca_6_4_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_6_4 u_ca_6_4_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_6_4 u_ca_6_4_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_6_4 u_ca_6_4_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_6_4 u_ca_6_4_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_6_4 u_ca_6_4_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_6_4 u_ca_6_4_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_6_4 u_ca_6_4_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_6_4 u_ca_6_4_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_6_4 u_ca_6_4_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_6_4 u_ca_6_4_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_6_4 u_ca_6_4_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_6_4 u_ca_6_4_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_6_4 u_ca_6_4_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_6_4 u_ca_6_4_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_6_4 u_ca_6_4_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_6_4 u_ca_6_4_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_6_4 u_ca_6_4_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_6_4 u_ca_6_4_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_6_4 u_ca_6_4_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_6_4 u_ca_6_4_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_6_4 u_ca_6_4_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_6_4 u_ca_6_4_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_6_4 u_ca_6_4_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_6_4 u_ca_6_4_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_6_4 u_ca_6_4_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_6_4 u_ca_6_4_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_6_4 u_ca_6_4_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_6_4 u_ca_6_4_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_6_4 u_ca_6_4_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_6_4 u_ca_6_4_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_6_4 u_ca_6_4_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_6_4 u_ca_6_4_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_6_4 u_ca_6_4_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_6_4 u_ca_6_4_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_6_4 u_ca_6_4_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_6_4 u_ca_6_4_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_6_4 u_ca_6_4_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_6_4 u_ca_6_4_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_6_4 u_ca_6_4_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_6_4 u_ca_6_4_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_6_4 u_ca_6_4_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_6_4 u_ca_6_4_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_6_4 u_ca_6_4_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_6_4 u_ca_6_4_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_6_4 u_ca_6_4_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_6_4 u_ca_6_4_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_6_4 u_ca_6_4_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_6_4 u_ca_6_4_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_6_4 u_ca_6_4_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_6_4 u_ca_6_4_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_6_4 u_ca_6_4_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_6_4 u_ca_6_4_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_6_4 u_ca_6_4_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_6_4 u_ca_6_4_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_6_4 u_ca_6_4_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_6_4 u_ca_6_4_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_6_4 u_ca_6_4_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_6_4 u_ca_6_4_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_6_4 u_ca_6_4_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_6_4 u_ca_6_4_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_6_4 u_ca_6_4_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_6_4 u_ca_6_4_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_6_4 u_ca_6_4_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_6_4 u_ca_6_4_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_6_4 u_ca_6_4_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_6_4 u_ca_6_4_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_6_4 u_ca_6_4_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_6_4 u_ca_6_4_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_6_4 u_ca_6_4_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_6_4 u_ca_6_4_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_6_4 u_ca_6_4_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_6_4 u_ca_6_4_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_6_4 u_ca_6_4_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_6_4 u_ca_6_4_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_6_4 u_ca_6_4_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_6_4 u_ca_6_4_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_6_4 u_ca_6_4_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_6_4 u_ca_6_4_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_6_4 u_ca_6_4_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_6_4 u_ca_6_4_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_6_4 u_ca_6_4_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_6_4 u_ca_6_4_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_6_4 u_ca_6_4_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_6_4 u_ca_6_4_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_6_4 u_ca_6_4_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_6_4 u_ca_6_4_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_6_4 u_ca_6_4_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_6_4 u_ca_6_4_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_6_4 u_ca_6_4_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_6_4 u_ca_6_4_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_6_4 u_ca_6_4_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_6_4 u_ca_6_4_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_6_4 u_ca_6_4_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_6_4 u_ca_6_4_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_6_4 u_ca_6_4_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_6_4 u_ca_6_4_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_6_4 u_ca_6_4_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_6_4 u_ca_6_4_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_6_4 u_ca_6_4_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_6_4 u_ca_6_4_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_6_4 u_ca_6_4_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_6_4 u_ca_6_4_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_6_4 u_ca_6_4_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_6_4 u_ca_6_4_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_6_4 u_ca_6_4_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_6_4 u_ca_6_4_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_6_4 u_ca_6_4_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_6_4 u_ca_6_4_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_6_4 u_ca_6_4_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_6_4 u_ca_6_4_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_6_4 u_ca_6_4_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_6_4 u_ca_6_4_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_6_4 u_ca_6_4_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_6_4 u_ca_6_4_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_6_4 u_ca_6_4_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_6_4 u_ca_6_4_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_6_4 u_ca_6_4_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_6_4 u_ca_6_4_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{2{1'b0}}, u_ca_out_0[1:0]};
assign col_out_1 = {u_ca_out_1[1:0], u_ca_out_0[3:2]};
assign col_out_2 = {u_ca_out_2[1:0], u_ca_out_1[3:2]};
assign col_out_3 = {u_ca_out_3[1:0], u_ca_out_2[3:2]};
assign col_out_4 = {u_ca_out_4[1:0], u_ca_out_3[3:2]};
assign col_out_5 = {u_ca_out_5[1:0], u_ca_out_4[3:2]};
assign col_out_6 = {u_ca_out_6[1:0], u_ca_out_5[3:2]};
assign col_out_7 = {u_ca_out_7[1:0], u_ca_out_6[3:2]};
assign col_out_8 = {u_ca_out_8[1:0], u_ca_out_7[3:2]};
assign col_out_9 = {u_ca_out_9[1:0], u_ca_out_8[3:2]};
assign col_out_10 = {u_ca_out_10[1:0], u_ca_out_9[3:2]};
assign col_out_11 = {u_ca_out_11[1:0], u_ca_out_10[3:2]};
assign col_out_12 = {u_ca_out_12[1:0], u_ca_out_11[3:2]};
assign col_out_13 = {u_ca_out_13[1:0], u_ca_out_12[3:2]};
assign col_out_14 = {u_ca_out_14[1:0], u_ca_out_13[3:2]};
assign col_out_15 = {u_ca_out_15[1:0], u_ca_out_14[3:2]};
assign col_out_16 = {u_ca_out_16[1:0], u_ca_out_15[3:2]};
assign col_out_17 = {u_ca_out_17[1:0], u_ca_out_16[3:2]};
assign col_out_18 = {u_ca_out_18[1:0], u_ca_out_17[3:2]};
assign col_out_19 = {u_ca_out_19[1:0], u_ca_out_18[3:2]};
assign col_out_20 = {u_ca_out_20[1:0], u_ca_out_19[3:2]};
assign col_out_21 = {u_ca_out_21[1:0], u_ca_out_20[3:2]};
assign col_out_22 = {u_ca_out_22[1:0], u_ca_out_21[3:2]};
assign col_out_23 = {u_ca_out_23[1:0], u_ca_out_22[3:2]};
assign col_out_24 = {u_ca_out_24[1:0], u_ca_out_23[3:2]};
assign col_out_25 = {u_ca_out_25[1:0], u_ca_out_24[3:2]};
assign col_out_26 = {u_ca_out_26[1:0], u_ca_out_25[3:2]};
assign col_out_27 = {u_ca_out_27[1:0], u_ca_out_26[3:2]};
assign col_out_28 = {u_ca_out_28[1:0], u_ca_out_27[3:2]};
assign col_out_29 = {u_ca_out_29[1:0], u_ca_out_28[3:2]};
assign col_out_30 = {u_ca_out_30[1:0], u_ca_out_29[3:2]};
assign col_out_31 = {u_ca_out_31[1:0], u_ca_out_30[3:2]};
assign col_out_32 = {u_ca_out_32[1:0], u_ca_out_31[3:2]};
assign col_out_33 = {u_ca_out_33[1:0], u_ca_out_32[3:2]};
assign col_out_34 = {u_ca_out_34[1:0], u_ca_out_33[3:2]};
assign col_out_35 = {u_ca_out_35[1:0], u_ca_out_34[3:2]};
assign col_out_36 = {u_ca_out_36[1:0], u_ca_out_35[3:2]};
assign col_out_37 = {u_ca_out_37[1:0], u_ca_out_36[3:2]};
assign col_out_38 = {u_ca_out_38[1:0], u_ca_out_37[3:2]};
assign col_out_39 = {u_ca_out_39[1:0], u_ca_out_38[3:2]};
assign col_out_40 = {u_ca_out_40[1:0], u_ca_out_39[3:2]};
assign col_out_41 = {u_ca_out_41[1:0], u_ca_out_40[3:2]};
assign col_out_42 = {u_ca_out_42[1:0], u_ca_out_41[3:2]};
assign col_out_43 = {u_ca_out_43[1:0], u_ca_out_42[3:2]};
assign col_out_44 = {u_ca_out_44[1:0], u_ca_out_43[3:2]};
assign col_out_45 = {u_ca_out_45[1:0], u_ca_out_44[3:2]};
assign col_out_46 = {u_ca_out_46[1:0], u_ca_out_45[3:2]};
assign col_out_47 = {u_ca_out_47[1:0], u_ca_out_46[3:2]};
assign col_out_48 = {u_ca_out_48[1:0], u_ca_out_47[3:2]};
assign col_out_49 = {u_ca_out_49[1:0], u_ca_out_48[3:2]};
assign col_out_50 = {u_ca_out_50[1:0], u_ca_out_49[3:2]};
assign col_out_51 = {u_ca_out_51[1:0], u_ca_out_50[3:2]};
assign col_out_52 = {u_ca_out_52[1:0], u_ca_out_51[3:2]};
assign col_out_53 = {u_ca_out_53[1:0], u_ca_out_52[3:2]};
assign col_out_54 = {u_ca_out_54[1:0], u_ca_out_53[3:2]};
assign col_out_55 = {u_ca_out_55[1:0], u_ca_out_54[3:2]};
assign col_out_56 = {u_ca_out_56[1:0], u_ca_out_55[3:2]};
assign col_out_57 = {u_ca_out_57[1:0], u_ca_out_56[3:2]};
assign col_out_58 = {u_ca_out_58[1:0], u_ca_out_57[3:2]};
assign col_out_59 = {u_ca_out_59[1:0], u_ca_out_58[3:2]};
assign col_out_60 = {u_ca_out_60[1:0], u_ca_out_59[3:2]};
assign col_out_61 = {u_ca_out_61[1:0], u_ca_out_60[3:2]};
assign col_out_62 = {u_ca_out_62[1:0], u_ca_out_61[3:2]};
assign col_out_63 = {u_ca_out_63[1:0], u_ca_out_62[3:2]};
assign col_out_64 = {u_ca_out_64[1:0], u_ca_out_63[3:2]};
assign col_out_65 = {u_ca_out_65[1:0], u_ca_out_64[3:2]};
assign col_out_66 = {u_ca_out_66[1:0], u_ca_out_65[3:2]};
assign col_out_67 = {u_ca_out_67[1:0], u_ca_out_66[3:2]};
assign col_out_68 = {u_ca_out_68[1:0], u_ca_out_67[3:2]};
assign col_out_69 = {u_ca_out_69[1:0], u_ca_out_68[3:2]};
assign col_out_70 = {u_ca_out_70[1:0], u_ca_out_69[3:2]};
assign col_out_71 = {u_ca_out_71[1:0], u_ca_out_70[3:2]};
assign col_out_72 = {u_ca_out_72[1:0], u_ca_out_71[3:2]};
assign col_out_73 = {u_ca_out_73[1:0], u_ca_out_72[3:2]};
assign col_out_74 = {u_ca_out_74[1:0], u_ca_out_73[3:2]};
assign col_out_75 = {u_ca_out_75[1:0], u_ca_out_74[3:2]};
assign col_out_76 = {u_ca_out_76[1:0], u_ca_out_75[3:2]};
assign col_out_77 = {u_ca_out_77[1:0], u_ca_out_76[3:2]};
assign col_out_78 = {u_ca_out_78[1:0], u_ca_out_77[3:2]};
assign col_out_79 = {u_ca_out_79[1:0], u_ca_out_78[3:2]};
assign col_out_80 = {u_ca_out_80[1:0], u_ca_out_79[3:2]};
assign col_out_81 = {u_ca_out_81[1:0], u_ca_out_80[3:2]};
assign col_out_82 = {u_ca_out_82[1:0], u_ca_out_81[3:2]};
assign col_out_83 = {u_ca_out_83[1:0], u_ca_out_82[3:2]};
assign col_out_84 = {u_ca_out_84[1:0], u_ca_out_83[3:2]};
assign col_out_85 = {u_ca_out_85[1:0], u_ca_out_84[3:2]};
assign col_out_86 = {u_ca_out_86[1:0], u_ca_out_85[3:2]};
assign col_out_87 = {u_ca_out_87[1:0], u_ca_out_86[3:2]};
assign col_out_88 = {u_ca_out_88[1:0], u_ca_out_87[3:2]};
assign col_out_89 = {u_ca_out_89[1:0], u_ca_out_88[3:2]};
assign col_out_90 = {u_ca_out_90[1:0], u_ca_out_89[3:2]};
assign col_out_91 = {u_ca_out_91[1:0], u_ca_out_90[3:2]};
assign col_out_92 = {u_ca_out_92[1:0], u_ca_out_91[3:2]};
assign col_out_93 = {u_ca_out_93[1:0], u_ca_out_92[3:2]};
assign col_out_94 = {u_ca_out_94[1:0], u_ca_out_93[3:2]};
assign col_out_95 = {u_ca_out_95[1:0], u_ca_out_94[3:2]};
assign col_out_96 = {u_ca_out_96[1:0], u_ca_out_95[3:2]};
assign col_out_97 = {u_ca_out_97[1:0], u_ca_out_96[3:2]};
assign col_out_98 = {u_ca_out_98[1:0], u_ca_out_97[3:2]};
assign col_out_99 = {u_ca_out_99[1:0], u_ca_out_98[3:2]};
assign col_out_100 = {u_ca_out_100[1:0], u_ca_out_99[3:2]};
assign col_out_101 = {u_ca_out_101[1:0], u_ca_out_100[3:2]};
assign col_out_102 = {u_ca_out_102[1:0], u_ca_out_101[3:2]};
assign col_out_103 = {u_ca_out_103[1:0], u_ca_out_102[3:2]};
assign col_out_104 = {u_ca_out_104[1:0], u_ca_out_103[3:2]};
assign col_out_105 = {u_ca_out_105[1:0], u_ca_out_104[3:2]};
assign col_out_106 = {u_ca_out_106[1:0], u_ca_out_105[3:2]};
assign col_out_107 = {u_ca_out_107[1:0], u_ca_out_106[3:2]};
assign col_out_108 = {u_ca_out_108[1:0], u_ca_out_107[3:2]};
assign col_out_109 = {u_ca_out_109[1:0], u_ca_out_108[3:2]};
assign col_out_110 = {u_ca_out_110[1:0], u_ca_out_109[3:2]};
assign col_out_111 = {u_ca_out_111[1:0], u_ca_out_110[3:2]};
assign col_out_112 = {u_ca_out_112[1:0], u_ca_out_111[3:2]};
assign col_out_113 = {u_ca_out_113[1:0], u_ca_out_112[3:2]};
assign col_out_114 = {u_ca_out_114[1:0], u_ca_out_113[3:2]};
assign col_out_115 = {u_ca_out_115[1:0], u_ca_out_114[3:2]};
assign col_out_116 = {u_ca_out_116[1:0], u_ca_out_115[3:2]};
assign col_out_117 = {u_ca_out_117[1:0], u_ca_out_116[3:2]};
assign col_out_118 = {u_ca_out_118[1:0], u_ca_out_117[3:2]};
assign col_out_119 = {u_ca_out_119[1:0], u_ca_out_118[3:2]};
assign col_out_120 = {u_ca_out_120[1:0], u_ca_out_119[3:2]};
assign col_out_121 = {u_ca_out_121[1:0], u_ca_out_120[3:2]};
assign col_out_122 = {u_ca_out_122[1:0], u_ca_out_121[3:2]};
assign col_out_123 = {u_ca_out_123[1:0], u_ca_out_122[3:2]};
assign col_out_124 = {u_ca_out_124[1:0], u_ca_out_123[3:2]};
assign col_out_125 = {u_ca_out_125[1:0], u_ca_out_124[3:2]};
assign col_out_126 = {u_ca_out_126[1:0], u_ca_out_125[3:2]};
assign col_out_127 = {u_ca_out_127[1:0], u_ca_out_126[3:2]};
assign col_out_128 = {u_ca_out_128[1:0], u_ca_out_127[3:2]};
assign col_out_129 = {u_ca_out_129[1:0], u_ca_out_128[3:2]};
assign col_out_130 = {u_ca_out_130[1:0], u_ca_out_129[3:2]};
assign col_out_131 = {u_ca_out_131[1:0], u_ca_out_130[3:2]};
assign col_out_132 = {u_ca_out_132[1:0], u_ca_out_131[3:2]};
assign col_out_133 = {u_ca_out_133[1:0], u_ca_out_132[3:2]};
assign col_out_134 = {u_ca_out_134[1:0], u_ca_out_133[3:2]};
assign col_out_135 = {u_ca_out_135[1:0], u_ca_out_134[3:2]};
assign col_out_136 = {u_ca_out_136[1:0], u_ca_out_135[3:2]};
assign col_out_137 = {u_ca_out_137[1:0], u_ca_out_136[3:2]};
assign col_out_138 = {u_ca_out_138[1:0], u_ca_out_137[3:2]};
assign col_out_139 = {u_ca_out_139[1:0], u_ca_out_138[3:2]};
assign col_out_140 = {u_ca_out_140[1:0], u_ca_out_139[3:2]};
assign col_out_141 = {u_ca_out_141[1:0], u_ca_out_140[3:2]};
assign col_out_142 = {u_ca_out_142[1:0], u_ca_out_141[3:2]};
assign col_out_143 = {u_ca_out_143[1:0], u_ca_out_142[3:2]};
assign col_out_144 = {u_ca_out_144[1:0], u_ca_out_143[3:2]};
assign col_out_145 = {u_ca_out_145[1:0], u_ca_out_144[3:2]};
assign col_out_146 = {u_ca_out_146[1:0], u_ca_out_145[3:2]};
assign col_out_147 = {u_ca_out_147[1:0], u_ca_out_146[3:2]};
assign col_out_148 = {u_ca_out_148[1:0], u_ca_out_147[3:2]};
assign col_out_149 = {u_ca_out_149[1:0], u_ca_out_148[3:2]};
assign col_out_150 = {u_ca_out_150[1:0], u_ca_out_149[3:2]};
assign col_out_151 = {u_ca_out_151[1:0], u_ca_out_150[3:2]};
assign col_out_152 = {u_ca_out_152[1:0], u_ca_out_151[3:2]};
assign col_out_153 = {u_ca_out_153[1:0], u_ca_out_152[3:2]};
assign col_out_154 = {u_ca_out_154[1:0], u_ca_out_153[3:2]};
assign col_out_155 = {u_ca_out_155[1:0], u_ca_out_154[3:2]};
assign col_out_156 = {u_ca_out_156[1:0], u_ca_out_155[3:2]};
assign col_out_157 = {u_ca_out_157[1:0], u_ca_out_156[3:2]};
assign col_out_158 = {u_ca_out_158[1:0], u_ca_out_157[3:2]};
assign col_out_159 = {u_ca_out_159[1:0], u_ca_out_158[3:2]};
assign col_out_160 = {u_ca_out_160[1:0], u_ca_out_159[3:2]};
assign col_out_161 = {u_ca_out_161[1:0], u_ca_out_160[3:2]};
assign col_out_162 = {u_ca_out_162[1:0], u_ca_out_161[3:2]};
assign col_out_163 = {u_ca_out_163[1:0], u_ca_out_162[3:2]};
assign col_out_164 = {u_ca_out_164[1:0], u_ca_out_163[3:2]};
assign col_out_165 = {u_ca_out_165[1:0], u_ca_out_164[3:2]};
assign col_out_166 = {u_ca_out_166[1:0], u_ca_out_165[3:2]};
assign col_out_167 = {u_ca_out_167[1:0], u_ca_out_166[3:2]};
assign col_out_168 = {u_ca_out_168[1:0], u_ca_out_167[3:2]};
assign col_out_169 = {u_ca_out_169[1:0], u_ca_out_168[3:2]};
assign col_out_170 = {u_ca_out_170[1:0], u_ca_out_169[3:2]};
assign col_out_171 = {u_ca_out_171[1:0], u_ca_out_170[3:2]};
assign col_out_172 = {u_ca_out_172[1:0], u_ca_out_171[3:2]};
assign col_out_173 = {u_ca_out_173[1:0], u_ca_out_172[3:2]};
assign col_out_174 = {u_ca_out_174[1:0], u_ca_out_173[3:2]};
assign col_out_175 = {u_ca_out_175[1:0], u_ca_out_174[3:2]};
assign col_out_176 = {u_ca_out_176[1:0], u_ca_out_175[3:2]};
assign col_out_177 = {u_ca_out_177[1:0], u_ca_out_176[3:2]};
assign col_out_178 = {u_ca_out_178[1:0], u_ca_out_177[3:2]};
assign col_out_179 = {u_ca_out_179[1:0], u_ca_out_178[3:2]};
assign col_out_180 = {u_ca_out_180[1:0], u_ca_out_179[3:2]};
assign col_out_181 = {u_ca_out_181[1:0], u_ca_out_180[3:2]};
assign col_out_182 = {u_ca_out_182[1:0], u_ca_out_181[3:2]};
assign col_out_183 = {u_ca_out_183[1:0], u_ca_out_182[3:2]};
assign col_out_184 = {u_ca_out_184[1:0], u_ca_out_183[3:2]};
assign col_out_185 = {u_ca_out_185[1:0], u_ca_out_184[3:2]};
assign col_out_186 = {u_ca_out_186[1:0], u_ca_out_185[3:2]};
assign col_out_187 = {u_ca_out_187[1:0], u_ca_out_186[3:2]};
assign col_out_188 = {u_ca_out_188[1:0], u_ca_out_187[3:2]};
assign col_out_189 = {u_ca_out_189[1:0], u_ca_out_188[3:2]};
assign col_out_190 = {u_ca_out_190[1:0], u_ca_out_189[3:2]};
assign col_out_191 = {u_ca_out_191[1:0], u_ca_out_190[3:2]};
assign col_out_192 = {u_ca_out_192[1:0], u_ca_out_191[3:2]};
assign col_out_193 = {u_ca_out_193[1:0], u_ca_out_192[3:2]};
assign col_out_194 = {u_ca_out_194[1:0], u_ca_out_193[3:2]};
assign col_out_195 = {u_ca_out_195[1:0], u_ca_out_194[3:2]};
assign col_out_196 = {u_ca_out_196[1:0], u_ca_out_195[3:2]};
assign col_out_197 = {u_ca_out_197[1:0], u_ca_out_196[3:2]};
assign col_out_198 = {u_ca_out_198[1:0], u_ca_out_197[3:2]};
assign col_out_199 = {u_ca_out_199[1:0], u_ca_out_198[3:2]};
assign col_out_200 = {u_ca_out_200[1:0], u_ca_out_199[3:2]};
assign col_out_201 = {u_ca_out_201[1:0], u_ca_out_200[3:2]};
assign col_out_202 = {u_ca_out_202[1:0], u_ca_out_201[3:2]};
assign col_out_203 = {u_ca_out_203[1:0], u_ca_out_202[3:2]};
assign col_out_204 = {u_ca_out_204[1:0], u_ca_out_203[3:2]};
assign col_out_205 = {u_ca_out_205[1:0], u_ca_out_204[3:2]};
assign col_out_206 = {u_ca_out_206[1:0], u_ca_out_205[3:2]};
assign col_out_207 = {u_ca_out_207[1:0], u_ca_out_206[3:2]};
assign col_out_208 = {u_ca_out_208[1:0], u_ca_out_207[3:2]};
assign col_out_209 = {u_ca_out_209[1:0], u_ca_out_208[3:2]};
assign col_out_210 = {u_ca_out_210[1:0], u_ca_out_209[3:2]};
assign col_out_211 = {u_ca_out_211[1:0], u_ca_out_210[3:2]};
assign col_out_212 = {u_ca_out_212[1:0], u_ca_out_211[3:2]};
assign col_out_213 = {u_ca_out_213[1:0], u_ca_out_212[3:2]};
assign col_out_214 = {u_ca_out_214[1:0], u_ca_out_213[3:2]};
assign col_out_215 = {u_ca_out_215[1:0], u_ca_out_214[3:2]};
assign col_out_216 = {u_ca_out_216[1:0], u_ca_out_215[3:2]};
assign col_out_217 = {u_ca_out_217[1:0], u_ca_out_216[3:2]};
assign col_out_218 = {u_ca_out_218[1:0], u_ca_out_217[3:2]};
assign col_out_219 = {u_ca_out_219[1:0], u_ca_out_218[3:2]};
assign col_out_220 = {u_ca_out_220[1:0], u_ca_out_219[3:2]};
assign col_out_221 = {u_ca_out_221[1:0], u_ca_out_220[3:2]};
assign col_out_222 = {u_ca_out_222[1:0], u_ca_out_221[3:2]};
assign col_out_223 = {u_ca_out_223[1:0], u_ca_out_222[3:2]};
assign col_out_224 = {u_ca_out_224[1:0], u_ca_out_223[3:2]};
assign col_out_225 = {u_ca_out_225[1:0], u_ca_out_224[3:2]};
assign col_out_226 = {u_ca_out_226[1:0], u_ca_out_225[3:2]};
assign col_out_227 = {u_ca_out_227[1:0], u_ca_out_226[3:2]};
assign col_out_228 = {u_ca_out_228[1:0], u_ca_out_227[3:2]};
assign col_out_229 = {u_ca_out_229[1:0], u_ca_out_228[3:2]};
assign col_out_230 = {u_ca_out_230[1:0], u_ca_out_229[3:2]};
assign col_out_231 = {u_ca_out_231[1:0], u_ca_out_230[3:2]};
assign col_out_232 = {u_ca_out_232[1:0], u_ca_out_231[3:2]};
assign col_out_233 = {u_ca_out_233[1:0], u_ca_out_232[3:2]};
assign col_out_234 = {u_ca_out_234[1:0], u_ca_out_233[3:2]};
assign col_out_235 = {u_ca_out_235[1:0], u_ca_out_234[3:2]};
assign col_out_236 = {u_ca_out_236[1:0], u_ca_out_235[3:2]};
assign col_out_237 = {u_ca_out_237[1:0], u_ca_out_236[3:2]};
assign col_out_238 = {u_ca_out_238[1:0], u_ca_out_237[3:2]};
assign col_out_239 = {u_ca_out_239[1:0], u_ca_out_238[3:2]};
assign col_out_240 = {u_ca_out_240[1:0], u_ca_out_239[3:2]};
assign col_out_241 = {u_ca_out_241[1:0], u_ca_out_240[3:2]};
assign col_out_242 = {u_ca_out_242[1:0], u_ca_out_241[3:2]};
assign col_out_243 = {u_ca_out_243[1:0], u_ca_out_242[3:2]};
assign col_out_244 = {u_ca_out_244[1:0], u_ca_out_243[3:2]};
assign col_out_245 = {u_ca_out_245[1:0], u_ca_out_244[3:2]};
assign col_out_246 = {u_ca_out_246[1:0], u_ca_out_245[3:2]};
assign col_out_247 = {u_ca_out_247[1:0], u_ca_out_246[3:2]};
assign col_out_248 = {u_ca_out_248[1:0], u_ca_out_247[3:2]};
assign col_out_249 = {u_ca_out_249[1:0], u_ca_out_248[3:2]};
assign col_out_250 = {u_ca_out_250[1:0], u_ca_out_249[3:2]};
assign col_out_251 = {u_ca_out_251[1:0], u_ca_out_250[3:2]};
assign col_out_252 = {u_ca_out_252[1:0], u_ca_out_251[3:2]};
assign col_out_253 = {u_ca_out_253[1:0], u_ca_out_252[3:2]};
assign col_out_254 = {u_ca_out_254[1:0], u_ca_out_253[3:2]};
assign col_out_255 = {u_ca_out_255[1:0], u_ca_out_254[3:2]};
assign col_out_256 = {u_ca_out_256[1:0], u_ca_out_255[3:2]};
assign col_out_257 = {u_ca_out_257[1:0], u_ca_out_256[3:2]};
assign col_out_258 = {u_ca_out_258[1:0], u_ca_out_257[3:2]};
assign col_out_259 = {u_ca_out_259[1:0], u_ca_out_258[3:2]};
assign col_out_260 = {u_ca_out_260[1:0], u_ca_out_259[3:2]};
assign col_out_261 = {u_ca_out_261[1:0], u_ca_out_260[3:2]};
assign col_out_262 = {u_ca_out_262[1:0], u_ca_out_261[3:2]};
assign col_out_263 = {u_ca_out_263[1:0], u_ca_out_262[3:2]};
assign col_out_264 = {u_ca_out_264[1:0], u_ca_out_263[3:2]};
assign col_out_265 = {u_ca_out_265[1:0], u_ca_out_264[3:2]};
assign col_out_266 = {u_ca_out_266[1:0], u_ca_out_265[3:2]};
assign col_out_267 = {u_ca_out_267[1:0], u_ca_out_266[3:2]};
assign col_out_268 = {u_ca_out_268[1:0], u_ca_out_267[3:2]};
assign col_out_269 = {u_ca_out_269[1:0], u_ca_out_268[3:2]};
assign col_out_270 = {u_ca_out_270[1:0], u_ca_out_269[3:2]};
assign col_out_271 = {u_ca_out_271[1:0], u_ca_out_270[3:2]};
assign col_out_272 = {u_ca_out_272[1:0], u_ca_out_271[3:2]};
assign col_out_273 = {u_ca_out_273[1:0], u_ca_out_272[3:2]};
assign col_out_274 = {u_ca_out_274[1:0], u_ca_out_273[3:2]};
assign col_out_275 = {u_ca_out_275[1:0], u_ca_out_274[3:2]};
assign col_out_276 = {u_ca_out_276[1:0], u_ca_out_275[3:2]};
assign col_out_277 = {u_ca_out_277[1:0], u_ca_out_276[3:2]};
assign col_out_278 = {u_ca_out_278[1:0], u_ca_out_277[3:2]};
assign col_out_279 = {u_ca_out_279[1:0], u_ca_out_278[3:2]};
assign col_out_280 = {u_ca_out_280[1:0], u_ca_out_279[3:2]};
assign col_out_281 = {u_ca_out_281[1:0], u_ca_out_280[3:2]};
assign col_out_282 = {u_ca_out_282[1:0], u_ca_out_281[3:2]};
assign col_out_283 = {u_ca_out_283[1:0], u_ca_out_282[3:2]};
assign col_out_284 = {u_ca_out_284[1:0], u_ca_out_283[3:2]};
assign col_out_285 = {u_ca_out_285[1:0], u_ca_out_284[3:2]};
assign col_out_286 = {u_ca_out_286[1:0], u_ca_out_285[3:2]};
assign col_out_287 = {u_ca_out_287[1:0], u_ca_out_286[3:2]};
assign col_out_288 = {u_ca_out_288[1:0], u_ca_out_287[3:2]};
assign col_out_289 = {u_ca_out_289[1:0], u_ca_out_288[3:2]};
assign col_out_290 = {u_ca_out_290[1:0], u_ca_out_289[3:2]};
assign col_out_291 = {u_ca_out_291[1:0], u_ca_out_290[3:2]};
assign col_out_292 = {u_ca_out_292[1:0], u_ca_out_291[3:2]};
assign col_out_293 = {u_ca_out_293[1:0], u_ca_out_292[3:2]};
assign col_out_294 = {u_ca_out_294[1:0], u_ca_out_293[3:2]};
assign col_out_295 = {u_ca_out_295[1:0], u_ca_out_294[3:2]};
assign col_out_296 = {u_ca_out_296[1:0], u_ca_out_295[3:2]};
assign col_out_297 = {u_ca_out_297[1:0], u_ca_out_296[3:2]};
assign col_out_298 = {u_ca_out_298[1:0], u_ca_out_297[3:2]};
assign col_out_299 = {u_ca_out_299[1:0], u_ca_out_298[3:2]};
assign col_out_300 = {u_ca_out_300[1:0], u_ca_out_299[3:2]};
assign col_out_301 = {u_ca_out_301[1:0], u_ca_out_300[3:2]};
assign col_out_302 = {u_ca_out_302[1:0], u_ca_out_301[3:2]};
assign col_out_303 = {u_ca_out_303[1:0], u_ca_out_302[3:2]};
assign col_out_304 = {u_ca_out_304[1:0], u_ca_out_303[3:2]};
assign col_out_305 = {u_ca_out_305[1:0], u_ca_out_304[3:2]};
assign col_out_306 = {u_ca_out_306[1:0], u_ca_out_305[3:2]};
assign col_out_307 = {u_ca_out_307[1:0], u_ca_out_306[3:2]};
assign col_out_308 = {u_ca_out_308[1:0], u_ca_out_307[3:2]};
assign col_out_309 = {u_ca_out_309[1:0], u_ca_out_308[3:2]};
assign col_out_310 = {u_ca_out_310[1:0], u_ca_out_309[3:2]};
assign col_out_311 = {u_ca_out_311[1:0], u_ca_out_310[3:2]};
assign col_out_312 = {u_ca_out_312[1:0], u_ca_out_311[3:2]};
assign col_out_313 = {u_ca_out_313[1:0], u_ca_out_312[3:2]};
assign col_out_314 = {u_ca_out_314[1:0], u_ca_out_313[3:2]};
assign col_out_315 = {u_ca_out_315[1:0], u_ca_out_314[3:2]};
assign col_out_316 = {u_ca_out_316[1:0], u_ca_out_315[3:2]};
assign col_out_317 = {u_ca_out_317[1:0], u_ca_out_316[3:2]};
assign col_out_318 = {u_ca_out_318[1:0], u_ca_out_317[3:2]};
assign col_out_319 = {u_ca_out_319[1:0], u_ca_out_318[3:2]};
assign col_out_320 = {u_ca_out_320[1:0], u_ca_out_319[3:2]};
assign col_out_321 = {u_ca_out_321[1:0], u_ca_out_320[3:2]};
assign col_out_322 = {u_ca_out_322[1:0], u_ca_out_321[3:2]};
assign col_out_323 = {u_ca_out_323[1:0], u_ca_out_322[3:2]};
assign col_out_324 = {u_ca_out_324[1:0], u_ca_out_323[3:2]};
assign col_out_325 = {u_ca_out_325[1:0], u_ca_out_324[3:2]};
assign col_out_326 = {u_ca_out_326[1:0], u_ca_out_325[3:2]};
assign col_out_327 = {u_ca_out_327[1:0], u_ca_out_326[3:2]};
assign col_out_328 = {u_ca_out_328[1:0], u_ca_out_327[3:2]};
assign col_out_329 = {u_ca_out_329[1:0], u_ca_out_328[3:2]};
assign col_out_330 = {u_ca_out_330[1:0], u_ca_out_329[3:2]};
assign col_out_331 = {u_ca_out_331[1:0], u_ca_out_330[3:2]};
assign col_out_332 = {u_ca_out_332[1:0], u_ca_out_331[3:2]};
assign col_out_333 = {u_ca_out_333[1:0], u_ca_out_332[3:2]};
assign col_out_334 = {u_ca_out_334[1:0], u_ca_out_333[3:2]};
assign col_out_335 = {u_ca_out_335[1:0], u_ca_out_334[3:2]};
assign col_out_336 = {u_ca_out_336[1:0], u_ca_out_335[3:2]};
assign col_out_337 = {u_ca_out_337[1:0], u_ca_out_336[3:2]};
assign col_out_338 = {u_ca_out_338[1:0], u_ca_out_337[3:2]};
assign col_out_339 = {u_ca_out_339[1:0], u_ca_out_338[3:2]};
assign col_out_340 = {u_ca_out_340[1:0], u_ca_out_339[3:2]};
assign col_out_341 = {u_ca_out_341[1:0], u_ca_out_340[3:2]};
assign col_out_342 = {u_ca_out_342[1:0], u_ca_out_341[3:2]};
assign col_out_343 = {u_ca_out_343[1:0], u_ca_out_342[3:2]};
assign col_out_344 = {u_ca_out_344[1:0], u_ca_out_343[3:2]};
assign col_out_345 = {u_ca_out_345[1:0], u_ca_out_344[3:2]};
assign col_out_346 = {u_ca_out_346[1:0], u_ca_out_345[3:2]};
assign col_out_347 = {u_ca_out_347[1:0], u_ca_out_346[3:2]};
assign col_out_348 = {u_ca_out_348[1:0], u_ca_out_347[3:2]};
assign col_out_349 = {u_ca_out_349[1:0], u_ca_out_348[3:2]};
assign col_out_350 = {u_ca_out_350[1:0], u_ca_out_349[3:2]};
assign col_out_351 = {u_ca_out_351[1:0], u_ca_out_350[3:2]};
assign col_out_352 = {u_ca_out_352[1:0], u_ca_out_351[3:2]};
assign col_out_353 = {u_ca_out_353[1:0], u_ca_out_352[3:2]};
assign col_out_354 = {u_ca_out_354[1:0], u_ca_out_353[3:2]};
assign col_out_355 = {u_ca_out_355[1:0], u_ca_out_354[3:2]};
assign col_out_356 = {u_ca_out_356[1:0], u_ca_out_355[3:2]};
assign col_out_357 = {u_ca_out_357[1:0], u_ca_out_356[3:2]};
assign col_out_358 = {u_ca_out_358[1:0], u_ca_out_357[3:2]};
assign col_out_359 = {u_ca_out_359[1:0], u_ca_out_358[3:2]};
assign col_out_360 = {u_ca_out_360[1:0], u_ca_out_359[3:2]};
assign col_out_361 = {u_ca_out_361[1:0], u_ca_out_360[3:2]};
assign col_out_362 = {u_ca_out_362[1:0], u_ca_out_361[3:2]};
assign col_out_363 = {u_ca_out_363[1:0], u_ca_out_362[3:2]};
assign col_out_364 = {u_ca_out_364[1:0], u_ca_out_363[3:2]};
assign col_out_365 = {u_ca_out_365[1:0], u_ca_out_364[3:2]};
assign col_out_366 = {u_ca_out_366[1:0], u_ca_out_365[3:2]};
assign col_out_367 = {u_ca_out_367[1:0], u_ca_out_366[3:2]};
assign col_out_368 = {u_ca_out_368[1:0], u_ca_out_367[3:2]};
assign col_out_369 = {u_ca_out_369[1:0], u_ca_out_368[3:2]};
assign col_out_370 = {u_ca_out_370[1:0], u_ca_out_369[3:2]};
assign col_out_371 = {u_ca_out_371[1:0], u_ca_out_370[3:2]};
assign col_out_372 = {u_ca_out_372[1:0], u_ca_out_371[3:2]};
assign col_out_373 = {u_ca_out_373[1:0], u_ca_out_372[3:2]};
assign col_out_374 = {u_ca_out_374[1:0], u_ca_out_373[3:2]};
assign col_out_375 = {u_ca_out_375[1:0], u_ca_out_374[3:2]};
assign col_out_376 = {u_ca_out_376[1:0], u_ca_out_375[3:2]};
assign col_out_377 = {u_ca_out_377[1:0], u_ca_out_376[3:2]};
assign col_out_378 = {u_ca_out_378[1:0], u_ca_out_377[3:2]};
assign col_out_379 = {u_ca_out_379[1:0], u_ca_out_378[3:2]};
assign col_out_380 = {u_ca_out_380[1:0], u_ca_out_379[3:2]};
assign col_out_381 = {u_ca_out_381[1:0], u_ca_out_380[3:2]};
assign col_out_382 = {u_ca_out_382[1:0], u_ca_out_381[3:2]};
assign col_out_383 = {u_ca_out_383[1:0], u_ca_out_382[3:2]};
assign col_out_384 = {u_ca_out_384[1:0], u_ca_out_383[3:2]};
assign col_out_385 = {u_ca_out_385[1:0], u_ca_out_384[3:2]};
assign col_out_386 = {u_ca_out_386[1:0], u_ca_out_385[3:2]};
assign col_out_387 = {u_ca_out_387[1:0], u_ca_out_386[3:2]};
assign col_out_388 = {u_ca_out_388[1:0], u_ca_out_387[3:2]};
assign col_out_389 = {u_ca_out_389[1:0], u_ca_out_388[3:2]};
assign col_out_390 = {u_ca_out_390[1:0], u_ca_out_389[3:2]};
assign col_out_391 = {u_ca_out_391[1:0], u_ca_out_390[3:2]};
assign col_out_392 = {u_ca_out_392[1:0], u_ca_out_391[3:2]};
assign col_out_393 = {u_ca_out_393[1:0], u_ca_out_392[3:2]};
assign col_out_394 = {u_ca_out_394[1:0], u_ca_out_393[3:2]};
assign col_out_395 = {u_ca_out_395[1:0], u_ca_out_394[3:2]};
assign col_out_396 = {u_ca_out_396[1:0], u_ca_out_395[3:2]};
assign col_out_397 = {u_ca_out_397[1:0], u_ca_out_396[3:2]};
assign col_out_398 = {u_ca_out_398[1:0], u_ca_out_397[3:2]};
assign col_out_399 = {u_ca_out_399[1:0], u_ca_out_398[3:2]};
assign col_out_400 = {u_ca_out_400[1:0], u_ca_out_399[3:2]};
assign col_out_401 = {u_ca_out_401[1:0], u_ca_out_400[3:2]};
assign col_out_402 = {u_ca_out_402[1:0], u_ca_out_401[3:2]};
assign col_out_403 = {u_ca_out_403[1:0], u_ca_out_402[3:2]};
assign col_out_404 = {u_ca_out_404[1:0], u_ca_out_403[3:2]};
assign col_out_405 = {u_ca_out_405[1:0], u_ca_out_404[3:2]};
assign col_out_406 = {u_ca_out_406[1:0], u_ca_out_405[3:2]};
assign col_out_407 = {u_ca_out_407[1:0], u_ca_out_406[3:2]};
assign col_out_408 = {u_ca_out_408[1:0], u_ca_out_407[3:2]};
assign col_out_409 = {u_ca_out_409[1:0], u_ca_out_408[3:2]};
assign col_out_410 = {u_ca_out_410[1:0], u_ca_out_409[3:2]};
assign col_out_411 = {u_ca_out_411[1:0], u_ca_out_410[3:2]};
assign col_out_412 = {u_ca_out_412[1:0], u_ca_out_411[3:2]};
assign col_out_413 = {u_ca_out_413[1:0], u_ca_out_412[3:2]};
assign col_out_414 = {u_ca_out_414[1:0], u_ca_out_413[3:2]};
assign col_out_415 = {u_ca_out_415[1:0], u_ca_out_414[3:2]};
assign col_out_416 = {u_ca_out_416[1:0], u_ca_out_415[3:2]};
assign col_out_417 = {u_ca_out_417[1:0], u_ca_out_416[3:2]};
assign col_out_418 = {u_ca_out_418[1:0], u_ca_out_417[3:2]};
assign col_out_419 = {u_ca_out_419[1:0], u_ca_out_418[3:2]};
assign col_out_420 = {u_ca_out_420[1:0], u_ca_out_419[3:2]};
assign col_out_421 = {u_ca_out_421[1:0], u_ca_out_420[3:2]};
assign col_out_422 = {u_ca_out_422[1:0], u_ca_out_421[3:2]};
assign col_out_423 = {u_ca_out_423[1:0], u_ca_out_422[3:2]};
assign col_out_424 = {u_ca_out_424[1:0], u_ca_out_423[3:2]};
assign col_out_425 = {u_ca_out_425[1:0], u_ca_out_424[3:2]};
assign col_out_426 = {u_ca_out_426[1:0], u_ca_out_425[3:2]};
assign col_out_427 = {u_ca_out_427[1:0], u_ca_out_426[3:2]};
assign col_out_428 = {u_ca_out_428[1:0], u_ca_out_427[3:2]};
assign col_out_429 = {u_ca_out_429[1:0], u_ca_out_428[3:2]};
assign col_out_430 = {u_ca_out_430[1:0], u_ca_out_429[3:2]};
assign col_out_431 = {u_ca_out_431[1:0], u_ca_out_430[3:2]};
assign col_out_432 = {u_ca_out_432[1:0], u_ca_out_431[3:2]};
assign col_out_433 = {u_ca_out_433[1:0], u_ca_out_432[3:2]};
assign col_out_434 = {u_ca_out_434[1:0], u_ca_out_433[3:2]};
assign col_out_435 = {u_ca_out_435[1:0], u_ca_out_434[3:2]};
assign col_out_436 = {u_ca_out_436[1:0], u_ca_out_435[3:2]};
assign col_out_437 = {u_ca_out_437[1:0], u_ca_out_436[3:2]};
assign col_out_438 = {u_ca_out_438[1:0], u_ca_out_437[3:2]};
assign col_out_439 = {u_ca_out_439[1:0], u_ca_out_438[3:2]};
assign col_out_440 = {u_ca_out_440[1:0], u_ca_out_439[3:2]};
assign col_out_441 = {u_ca_out_441[1:0], u_ca_out_440[3:2]};
assign col_out_442 = {u_ca_out_442[1:0], u_ca_out_441[3:2]};
assign col_out_443 = {u_ca_out_443[1:0], u_ca_out_442[3:2]};
assign col_out_444 = {u_ca_out_444[1:0], u_ca_out_443[3:2]};
assign col_out_445 = {u_ca_out_445[1:0], u_ca_out_444[3:2]};
assign col_out_446 = {u_ca_out_446[1:0], u_ca_out_445[3:2]};
assign col_out_447 = {u_ca_out_447[1:0], u_ca_out_446[3:2]};
assign col_out_448 = {u_ca_out_448[1:0], u_ca_out_447[3:2]};
assign col_out_449 = {u_ca_out_449[1:0], u_ca_out_448[3:2]};
assign col_out_450 = {u_ca_out_450[1:0], u_ca_out_449[3:2]};
assign col_out_451 = {u_ca_out_451[1:0], u_ca_out_450[3:2]};
assign col_out_452 = {u_ca_out_452[1:0], u_ca_out_451[3:2]};
assign col_out_453 = {u_ca_out_453[1:0], u_ca_out_452[3:2]};
assign col_out_454 = {u_ca_out_454[1:0], u_ca_out_453[3:2]};
assign col_out_455 = {u_ca_out_455[1:0], u_ca_out_454[3:2]};
assign col_out_456 = {u_ca_out_456[1:0], u_ca_out_455[3:2]};
assign col_out_457 = {u_ca_out_457[1:0], u_ca_out_456[3:2]};
assign col_out_458 = {u_ca_out_458[1:0], u_ca_out_457[3:2]};
assign col_out_459 = {u_ca_out_459[1:0], u_ca_out_458[3:2]};
assign col_out_460 = {u_ca_out_460[1:0], u_ca_out_459[3:2]};
assign col_out_461 = {u_ca_out_461[1:0], u_ca_out_460[3:2]};
assign col_out_462 = {u_ca_out_462[1:0], u_ca_out_461[3:2]};
assign col_out_463 = {u_ca_out_463[1:0], u_ca_out_462[3:2]};
assign col_out_464 = {u_ca_out_464[1:0], u_ca_out_463[3:2]};
assign col_out_465 = {u_ca_out_465[1:0], u_ca_out_464[3:2]};
assign col_out_466 = {u_ca_out_466[1:0], u_ca_out_465[3:2]};
assign col_out_467 = {u_ca_out_467[1:0], u_ca_out_466[3:2]};
assign col_out_468 = {u_ca_out_468[1:0], u_ca_out_467[3:2]};
assign col_out_469 = {u_ca_out_469[1:0], u_ca_out_468[3:2]};
assign col_out_470 = {u_ca_out_470[1:0], u_ca_out_469[3:2]};
assign col_out_471 = {u_ca_out_471[1:0], u_ca_out_470[3:2]};
assign col_out_472 = {u_ca_out_472[1:0], u_ca_out_471[3:2]};
assign col_out_473 = {u_ca_out_473[1:0], u_ca_out_472[3:2]};
assign col_out_474 = {u_ca_out_474[1:0], u_ca_out_473[3:2]};
assign col_out_475 = {u_ca_out_475[1:0], u_ca_out_474[3:2]};
assign col_out_476 = {u_ca_out_476[1:0], u_ca_out_475[3:2]};
assign col_out_477 = {u_ca_out_477[1:0], u_ca_out_476[3:2]};
assign col_out_478 = {u_ca_out_478[1:0], u_ca_out_477[3:2]};
assign col_out_479 = {u_ca_out_479[1:0], u_ca_out_478[3:2]};
assign col_out_480 = {u_ca_out_480[1:0], u_ca_out_479[3:2]};
assign col_out_481 = {u_ca_out_481[1:0], u_ca_out_480[3:2]};
assign col_out_482 = {u_ca_out_482[1:0], u_ca_out_481[3:2]};
assign col_out_483 = {u_ca_out_483[1:0], u_ca_out_482[3:2]};
assign col_out_484 = {u_ca_out_484[1:0], u_ca_out_483[3:2]};
assign col_out_485 = {u_ca_out_485[1:0], u_ca_out_484[3:2]};
assign col_out_486 = {u_ca_out_486[1:0], u_ca_out_485[3:2]};
assign col_out_487 = {u_ca_out_487[1:0], u_ca_out_486[3:2]};
assign col_out_488 = {u_ca_out_488[1:0], u_ca_out_487[3:2]};
assign col_out_489 = {u_ca_out_489[1:0], u_ca_out_488[3:2]};
assign col_out_490 = {u_ca_out_490[1:0], u_ca_out_489[3:2]};
assign col_out_491 = {u_ca_out_491[1:0], u_ca_out_490[3:2]};
assign col_out_492 = {u_ca_out_492[1:0], u_ca_out_491[3:2]};
assign col_out_493 = {u_ca_out_493[1:0], u_ca_out_492[3:2]};
assign col_out_494 = {u_ca_out_494[1:0], u_ca_out_493[3:2]};
assign col_out_495 = {u_ca_out_495[1:0], u_ca_out_494[3:2]};
assign col_out_496 = {u_ca_out_496[1:0], u_ca_out_495[3:2]};
assign col_out_497 = {u_ca_out_497[1:0], u_ca_out_496[3:2]};
assign col_out_498 = {u_ca_out_498[1:0], u_ca_out_497[3:2]};
assign col_out_499 = {u_ca_out_499[1:0], u_ca_out_498[3:2]};
assign col_out_500 = {u_ca_out_500[1:0], u_ca_out_499[3:2]};
assign col_out_501 = {u_ca_out_501[1:0], u_ca_out_500[3:2]};
assign col_out_502 = {u_ca_out_502[1:0], u_ca_out_501[3:2]};
assign col_out_503 = {u_ca_out_503[1:0], u_ca_out_502[3:2]};
assign col_out_504 = {u_ca_out_504[1:0], u_ca_out_503[3:2]};
assign col_out_505 = {u_ca_out_505[1:0], u_ca_out_504[3:2]};
assign col_out_506 = {u_ca_out_506[1:0], u_ca_out_505[3:2]};
assign col_out_507 = {u_ca_out_507[1:0], u_ca_out_506[3:2]};
assign col_out_508 = {u_ca_out_508[1:0], u_ca_out_507[3:2]};
assign col_out_509 = {u_ca_out_509[1:0], u_ca_out_508[3:2]};
assign col_out_510 = {u_ca_out_510[1:0], u_ca_out_509[3:2]};
assign col_out_511 = {u_ca_out_511[1:0], u_ca_out_510[3:2]};
assign col_out_512 = {u_ca_out_512[1:0], u_ca_out_511[3:2]};
assign col_out_513 = {u_ca_out_513[1:0], u_ca_out_512[3:2]};
assign col_out_514 = {u_ca_out_514[1:0], u_ca_out_513[3:2]};
assign col_out_515 = {u_ca_out_515[1:0], u_ca_out_514[3:2]};
assign col_out_516 = {u_ca_out_516[1:0], u_ca_out_515[3:2]};
assign col_out_517 = {u_ca_out_517[1:0], u_ca_out_516[3:2]};
assign col_out_518 = {u_ca_out_518[1:0], u_ca_out_517[3:2]};
assign col_out_519 = {u_ca_out_519[1:0], u_ca_out_518[3:2]};
assign col_out_520 = {u_ca_out_520[1:0], u_ca_out_519[3:2]};
assign col_out_521 = {u_ca_out_521[1:0], u_ca_out_520[3:2]};
assign col_out_522 = {u_ca_out_522[1:0], u_ca_out_521[3:2]};
assign col_out_523 = {u_ca_out_523[1:0], u_ca_out_522[3:2]};
assign col_out_524 = {u_ca_out_524[1:0], u_ca_out_523[3:2]};
assign col_out_525 = {u_ca_out_525[1:0], u_ca_out_524[3:2]};
assign col_out_526 = {u_ca_out_526[1:0], u_ca_out_525[3:2]};
assign col_out_527 = {u_ca_out_527[1:0], u_ca_out_526[3:2]};
assign col_out_528 = {u_ca_out_528[1:0], u_ca_out_527[3:2]};
assign col_out_529 = {u_ca_out_529[1:0], u_ca_out_528[3:2]};
assign col_out_530 = {u_ca_out_530[1:0], u_ca_out_529[3:2]};
assign col_out_531 = {u_ca_out_531[1:0], u_ca_out_530[3:2]};
assign col_out_532 = {u_ca_out_532[1:0], u_ca_out_531[3:2]};
assign col_out_533 = {u_ca_out_533[1:0], u_ca_out_532[3:2]};
assign col_out_534 = {u_ca_out_534[1:0], u_ca_out_533[3:2]};
assign col_out_535 = {u_ca_out_535[1:0], u_ca_out_534[3:2]};
assign col_out_536 = {u_ca_out_536[1:0], u_ca_out_535[3:2]};
assign col_out_537 = {u_ca_out_537[1:0], u_ca_out_536[3:2]};
assign col_out_538 = {u_ca_out_538[1:0], u_ca_out_537[3:2]};
assign col_out_539 = {u_ca_out_539[1:0], u_ca_out_538[3:2]};
assign col_out_540 = {u_ca_out_540[1:0], u_ca_out_539[3:2]};
assign col_out_541 = {u_ca_out_541[1:0], u_ca_out_540[3:2]};
assign col_out_542 = {u_ca_out_542[1:0], u_ca_out_541[3:2]};
assign col_out_543 = {u_ca_out_543[1:0], u_ca_out_542[3:2]};
assign col_out_544 = {u_ca_out_544[1:0], u_ca_out_543[3:2]};
assign col_out_545 = {u_ca_out_545[1:0], u_ca_out_544[3:2]};
assign col_out_546 = {u_ca_out_546[1:0], u_ca_out_545[3:2]};
assign col_out_547 = {u_ca_out_547[1:0], u_ca_out_546[3:2]};
assign col_out_548 = {u_ca_out_548[1:0], u_ca_out_547[3:2]};
assign col_out_549 = {u_ca_out_549[1:0], u_ca_out_548[3:2]};
assign col_out_550 = {u_ca_out_550[1:0], u_ca_out_549[3:2]};
assign col_out_551 = {u_ca_out_551[1:0], u_ca_out_550[3:2]};
assign col_out_552 = {u_ca_out_552[1:0], u_ca_out_551[3:2]};
assign col_out_553 = {u_ca_out_553[1:0], u_ca_out_552[3:2]};
assign col_out_554 = {u_ca_out_554[1:0], u_ca_out_553[3:2]};
assign col_out_555 = {u_ca_out_555[1:0], u_ca_out_554[3:2]};
assign col_out_556 = {u_ca_out_556[1:0], u_ca_out_555[3:2]};
assign col_out_557 = {u_ca_out_557[1:0], u_ca_out_556[3:2]};
assign col_out_558 = {u_ca_out_558[1:0], u_ca_out_557[3:2]};
assign col_out_559 = {u_ca_out_559[1:0], u_ca_out_558[3:2]};
assign col_out_560 = {u_ca_out_560[1:0], u_ca_out_559[3:2]};
assign col_out_561 = {u_ca_out_561[1:0], u_ca_out_560[3:2]};
assign col_out_562 = {u_ca_out_562[1:0], u_ca_out_561[3:2]};
assign col_out_563 = {u_ca_out_563[1:0], u_ca_out_562[3:2]};
assign col_out_564 = {u_ca_out_564[1:0], u_ca_out_563[3:2]};
assign col_out_565 = {u_ca_out_565[1:0], u_ca_out_564[3:2]};
assign col_out_566 = {u_ca_out_566[1:0], u_ca_out_565[3:2]};
assign col_out_567 = {u_ca_out_567[1:0], u_ca_out_566[3:2]};
assign col_out_568 = {u_ca_out_568[1:0], u_ca_out_567[3:2]};
assign col_out_569 = {u_ca_out_569[1:0], u_ca_out_568[3:2]};
assign col_out_570 = {u_ca_out_570[1:0], u_ca_out_569[3:2]};
assign col_out_571 = {u_ca_out_571[1:0], u_ca_out_570[3:2]};
assign col_out_572 = {u_ca_out_572[1:0], u_ca_out_571[3:2]};
assign col_out_573 = {u_ca_out_573[1:0], u_ca_out_572[3:2]};
assign col_out_574 = {u_ca_out_574[1:0], u_ca_out_573[3:2]};
assign col_out_575 = {u_ca_out_575[1:0], u_ca_out_574[3:2]};
assign col_out_576 = {u_ca_out_576[1:0], u_ca_out_575[3:2]};
assign col_out_577 = {u_ca_out_577[1:0], u_ca_out_576[3:2]};
assign col_out_578 = {u_ca_out_578[1:0], u_ca_out_577[3:2]};
assign col_out_579 = {u_ca_out_579[1:0], u_ca_out_578[3:2]};
assign col_out_580 = {u_ca_out_580[1:0], u_ca_out_579[3:2]};
assign col_out_581 = {u_ca_out_581[1:0], u_ca_out_580[3:2]};
assign col_out_582 = {u_ca_out_582[1:0], u_ca_out_581[3:2]};
assign col_out_583 = {u_ca_out_583[1:0], u_ca_out_582[3:2]};
assign col_out_584 = {u_ca_out_584[1:0], u_ca_out_583[3:2]};
assign col_out_585 = {u_ca_out_585[1:0], u_ca_out_584[3:2]};
assign col_out_586 = {u_ca_out_586[1:0], u_ca_out_585[3:2]};
assign col_out_587 = {u_ca_out_587[1:0], u_ca_out_586[3:2]};
assign col_out_588 = {u_ca_out_588[1:0], u_ca_out_587[3:2]};
assign col_out_589 = {u_ca_out_589[1:0], u_ca_out_588[3:2]};
assign col_out_590 = {u_ca_out_590[1:0], u_ca_out_589[3:2]};
assign col_out_591 = {u_ca_out_591[1:0], u_ca_out_590[3:2]};
assign col_out_592 = {u_ca_out_592[1:0], u_ca_out_591[3:2]};
assign col_out_593 = {u_ca_out_593[1:0], u_ca_out_592[3:2]};
assign col_out_594 = {u_ca_out_594[1:0], u_ca_out_593[3:2]};
assign col_out_595 = {u_ca_out_595[1:0], u_ca_out_594[3:2]};
assign col_out_596 = {u_ca_out_596[1:0], u_ca_out_595[3:2]};
assign col_out_597 = {u_ca_out_597[1:0], u_ca_out_596[3:2]};
assign col_out_598 = {u_ca_out_598[1:0], u_ca_out_597[3:2]};
assign col_out_599 = {u_ca_out_599[1:0], u_ca_out_598[3:2]};
assign col_out_600 = {u_ca_out_600[1:0], u_ca_out_599[3:2]};
assign col_out_601 = {u_ca_out_601[1:0], u_ca_out_600[3:2]};
assign col_out_602 = {u_ca_out_602[1:0], u_ca_out_601[3:2]};
assign col_out_603 = {u_ca_out_603[1:0], u_ca_out_602[3:2]};
assign col_out_604 = {u_ca_out_604[1:0], u_ca_out_603[3:2]};
assign col_out_605 = {u_ca_out_605[1:0], u_ca_out_604[3:2]};
assign col_out_606 = {u_ca_out_606[1:0], u_ca_out_605[3:2]};
assign col_out_607 = {u_ca_out_607[1:0], u_ca_out_606[3:2]};
assign col_out_608 = {u_ca_out_608[1:0], u_ca_out_607[3:2]};
assign col_out_609 = {u_ca_out_609[1:0], u_ca_out_608[3:2]};
assign col_out_610 = {u_ca_out_610[1:0], u_ca_out_609[3:2]};
assign col_out_611 = {u_ca_out_611[1:0], u_ca_out_610[3:2]};
assign col_out_612 = {u_ca_out_612[1:0], u_ca_out_611[3:2]};
assign col_out_613 = {u_ca_out_613[1:0], u_ca_out_612[3:2]};
assign col_out_614 = {u_ca_out_614[1:0], u_ca_out_613[3:2]};
assign col_out_615 = {u_ca_out_615[1:0], u_ca_out_614[3:2]};
assign col_out_616 = {u_ca_out_616[1:0], u_ca_out_615[3:2]};
assign col_out_617 = {u_ca_out_617[1:0], u_ca_out_616[3:2]};
assign col_out_618 = {u_ca_out_618[1:0], u_ca_out_617[3:2]};
assign col_out_619 = {u_ca_out_619[1:0], u_ca_out_618[3:2]};
assign col_out_620 = {u_ca_out_620[1:0], u_ca_out_619[3:2]};
assign col_out_621 = {u_ca_out_621[1:0], u_ca_out_620[3:2]};
assign col_out_622 = {u_ca_out_622[1:0], u_ca_out_621[3:2]};
assign col_out_623 = {u_ca_out_623[1:0], u_ca_out_622[3:2]};
assign col_out_624 = {u_ca_out_624[1:0], u_ca_out_623[3:2]};
assign col_out_625 = {u_ca_out_625[1:0], u_ca_out_624[3:2]};
assign col_out_626 = {u_ca_out_626[1:0], u_ca_out_625[3:2]};
assign col_out_627 = {u_ca_out_627[1:0], u_ca_out_626[3:2]};
assign col_out_628 = {u_ca_out_628[1:0], u_ca_out_627[3:2]};
assign col_out_629 = {u_ca_out_629[1:0], u_ca_out_628[3:2]};
assign col_out_630 = {u_ca_out_630[1:0], u_ca_out_629[3:2]};
assign col_out_631 = {u_ca_out_631[1:0], u_ca_out_630[3:2]};
assign col_out_632 = {u_ca_out_632[1:0], u_ca_out_631[3:2]};
assign col_out_633 = {u_ca_out_633[1:0], u_ca_out_632[3:2]};
assign col_out_634 = {u_ca_out_634[1:0], u_ca_out_633[3:2]};
assign col_out_635 = {u_ca_out_635[1:0], u_ca_out_634[3:2]};
assign col_out_636 = {u_ca_out_636[1:0], u_ca_out_635[3:2]};
assign col_out_637 = {u_ca_out_637[1:0], u_ca_out_636[3:2]};
assign col_out_638 = {u_ca_out_638[1:0], u_ca_out_637[3:2]};
assign col_out_639 = {u_ca_out_639[1:0], u_ca_out_638[3:2]};
assign col_out_640 = {u_ca_out_640[1:0], u_ca_out_639[3:2]};
assign col_out_641 = {u_ca_out_641[1:0], u_ca_out_640[3:2]};
assign col_out_642 = {u_ca_out_642[1:0], u_ca_out_641[3:2]};
assign col_out_643 = {u_ca_out_643[1:0], u_ca_out_642[3:2]};
assign col_out_644 = {u_ca_out_644[1:0], u_ca_out_643[3:2]};
assign col_out_645 = {u_ca_out_645[1:0], u_ca_out_644[3:2]};
assign col_out_646 = {u_ca_out_646[1:0], u_ca_out_645[3:2]};
assign col_out_647 = {u_ca_out_647[1:0], u_ca_out_646[3:2]};
assign col_out_648 = {u_ca_out_648[1:0], u_ca_out_647[3:2]};
assign col_out_649 = {u_ca_out_649[1:0], u_ca_out_648[3:2]};
assign col_out_650 = {u_ca_out_650[1:0], u_ca_out_649[3:2]};
assign col_out_651 = {u_ca_out_651[1:0], u_ca_out_650[3:2]};
assign col_out_652 = {u_ca_out_652[1:0], u_ca_out_651[3:2]};
assign col_out_653 = {u_ca_out_653[1:0], u_ca_out_652[3:2]};
assign col_out_654 = {u_ca_out_654[1:0], u_ca_out_653[3:2]};
assign col_out_655 = {u_ca_out_655[1:0], u_ca_out_654[3:2]};
assign col_out_656 = {u_ca_out_656[1:0], u_ca_out_655[3:2]};
assign col_out_657 = {u_ca_out_657[1:0], u_ca_out_656[3:2]};
assign col_out_658 = {u_ca_out_658[1:0], u_ca_out_657[3:2]};
assign col_out_659 = {u_ca_out_659[1:0], u_ca_out_658[3:2]};
assign col_out_660 = {u_ca_out_660[1:0], u_ca_out_659[3:2]};
assign col_out_661 = {u_ca_out_661[1:0], u_ca_out_660[3:2]};
assign col_out_662 = {u_ca_out_662[1:0], u_ca_out_661[3:2]};
assign col_out_663 = {u_ca_out_663[1:0], u_ca_out_662[3:2]};
assign col_out_664 = {u_ca_out_664[1:0], u_ca_out_663[3:2]};
assign col_out_665 = {u_ca_out_665[1:0], u_ca_out_664[3:2]};
assign col_out_666 = {u_ca_out_666[1:0], u_ca_out_665[3:2]};
assign col_out_667 = {u_ca_out_667[1:0], u_ca_out_666[3:2]};
assign col_out_668 = {u_ca_out_668[1:0], u_ca_out_667[3:2]};
assign col_out_669 = {u_ca_out_669[1:0], u_ca_out_668[3:2]};
assign col_out_670 = {u_ca_out_670[1:0], u_ca_out_669[3:2]};
assign col_out_671 = {u_ca_out_671[1:0], u_ca_out_670[3:2]};
assign col_out_672 = {u_ca_out_672[1:0], u_ca_out_671[3:2]};
assign col_out_673 = {u_ca_out_673[1:0], u_ca_out_672[3:2]};
assign col_out_674 = {u_ca_out_674[1:0], u_ca_out_673[3:2]};
assign col_out_675 = {u_ca_out_675[1:0], u_ca_out_674[3:2]};
assign col_out_676 = {u_ca_out_676[1:0], u_ca_out_675[3:2]};
assign col_out_677 = {u_ca_out_677[1:0], u_ca_out_676[3:2]};
assign col_out_678 = {u_ca_out_678[1:0], u_ca_out_677[3:2]};
assign col_out_679 = {u_ca_out_679[1:0], u_ca_out_678[3:2]};
assign col_out_680 = {u_ca_out_680[1:0], u_ca_out_679[3:2]};
assign col_out_681 = {u_ca_out_681[1:0], u_ca_out_680[3:2]};
assign col_out_682 = {u_ca_out_682[1:0], u_ca_out_681[3:2]};
assign col_out_683 = {u_ca_out_683[1:0], u_ca_out_682[3:2]};
assign col_out_684 = {u_ca_out_684[1:0], u_ca_out_683[3:2]};
assign col_out_685 = {u_ca_out_685[1:0], u_ca_out_684[3:2]};
assign col_out_686 = {u_ca_out_686[1:0], u_ca_out_685[3:2]};
assign col_out_687 = {u_ca_out_687[1:0], u_ca_out_686[3:2]};
assign col_out_688 = {u_ca_out_688[1:0], u_ca_out_687[3:2]};
assign col_out_689 = {u_ca_out_689[1:0], u_ca_out_688[3:2]};
assign col_out_690 = {u_ca_out_690[1:0], u_ca_out_689[3:2]};
assign col_out_691 = {u_ca_out_691[1:0], u_ca_out_690[3:2]};
assign col_out_692 = {u_ca_out_692[1:0], u_ca_out_691[3:2]};
assign col_out_693 = {u_ca_out_693[1:0], u_ca_out_692[3:2]};
assign col_out_694 = {u_ca_out_694[1:0], u_ca_out_693[3:2]};
assign col_out_695 = {u_ca_out_695[1:0], u_ca_out_694[3:2]};
assign col_out_696 = {u_ca_out_696[1:0], u_ca_out_695[3:2]};
assign col_out_697 = {u_ca_out_697[1:0], u_ca_out_696[3:2]};
assign col_out_698 = {u_ca_out_698[1:0], u_ca_out_697[3:2]};
assign col_out_699 = {u_ca_out_699[1:0], u_ca_out_698[3:2]};
assign col_out_700 = {u_ca_out_700[1:0], u_ca_out_699[3:2]};
assign col_out_701 = {u_ca_out_701[1:0], u_ca_out_700[3:2]};
assign col_out_702 = {u_ca_out_702[1:0], u_ca_out_701[3:2]};
assign col_out_703 = {u_ca_out_703[1:0], u_ca_out_702[3:2]};
assign col_out_704 = {u_ca_out_704[1:0], u_ca_out_703[3:2]};
assign col_out_705 = {u_ca_out_705[1:0], u_ca_out_704[3:2]};
assign col_out_706 = {u_ca_out_706[1:0], u_ca_out_705[3:2]};
assign col_out_707 = {u_ca_out_707[1:0], u_ca_out_706[3:2]};
assign col_out_708 = {u_ca_out_708[1:0], u_ca_out_707[3:2]};
assign col_out_709 = {u_ca_out_709[1:0], u_ca_out_708[3:2]};
assign col_out_710 = {u_ca_out_710[1:0], u_ca_out_709[3:2]};
assign col_out_711 = {u_ca_out_711[1:0], u_ca_out_710[3:2]};
assign col_out_712 = {u_ca_out_712[1:0], u_ca_out_711[3:2]};
assign col_out_713 = {u_ca_out_713[1:0], u_ca_out_712[3:2]};
assign col_out_714 = {u_ca_out_714[1:0], u_ca_out_713[3:2]};
assign col_out_715 = {u_ca_out_715[1:0], u_ca_out_714[3:2]};
assign col_out_716 = {u_ca_out_716[1:0], u_ca_out_715[3:2]};
assign col_out_717 = {u_ca_out_717[1:0], u_ca_out_716[3:2]};
assign col_out_718 = {u_ca_out_718[1:0], u_ca_out_717[3:2]};
assign col_out_719 = {u_ca_out_719[1:0], u_ca_out_718[3:2]};
assign col_out_720 = {u_ca_out_720[1:0], u_ca_out_719[3:2]};
assign col_out_721 = {u_ca_out_721[1:0], u_ca_out_720[3:2]};
assign col_out_722 = {u_ca_out_722[1:0], u_ca_out_721[3:2]};
assign col_out_723 = {u_ca_out_723[1:0], u_ca_out_722[3:2]};
assign col_out_724 = {u_ca_out_724[1:0], u_ca_out_723[3:2]};
assign col_out_725 = {u_ca_out_725[1:0], u_ca_out_724[3:2]};
assign col_out_726 = {u_ca_out_726[1:0], u_ca_out_725[3:2]};
assign col_out_727 = {u_ca_out_727[1:0], u_ca_out_726[3:2]};
assign col_out_728 = {u_ca_out_728[1:0], u_ca_out_727[3:2]};
assign col_out_729 = {u_ca_out_729[1:0], u_ca_out_728[3:2]};
assign col_out_730 = {u_ca_out_730[1:0], u_ca_out_729[3:2]};
assign col_out_731 = {u_ca_out_731[1:0], u_ca_out_730[3:2]};
assign col_out_732 = {u_ca_out_732[1:0], u_ca_out_731[3:2]};
assign col_out_733 = {u_ca_out_733[1:0], u_ca_out_732[3:2]};
assign col_out_734 = {u_ca_out_734[1:0], u_ca_out_733[3:2]};
assign col_out_735 = {u_ca_out_735[1:0], u_ca_out_734[3:2]};
assign col_out_736 = {u_ca_out_736[1:0], u_ca_out_735[3:2]};
assign col_out_737 = {u_ca_out_737[1:0], u_ca_out_736[3:2]};
assign col_out_738 = {u_ca_out_738[1:0], u_ca_out_737[3:2]};
assign col_out_739 = {u_ca_out_739[1:0], u_ca_out_738[3:2]};
assign col_out_740 = {u_ca_out_740[1:0], u_ca_out_739[3:2]};
assign col_out_741 = {u_ca_out_741[1:0], u_ca_out_740[3:2]};
assign col_out_742 = {u_ca_out_742[1:0], u_ca_out_741[3:2]};
assign col_out_743 = {u_ca_out_743[1:0], u_ca_out_742[3:2]};
assign col_out_744 = {u_ca_out_744[1:0], u_ca_out_743[3:2]};
assign col_out_745 = {u_ca_out_745[1:0], u_ca_out_744[3:2]};
assign col_out_746 = {u_ca_out_746[1:0], u_ca_out_745[3:2]};
assign col_out_747 = {u_ca_out_747[1:0], u_ca_out_746[3:2]};
assign col_out_748 = {u_ca_out_748[1:0], u_ca_out_747[3:2]};
assign col_out_749 = {u_ca_out_749[1:0], u_ca_out_748[3:2]};
assign col_out_750 = {u_ca_out_750[1:0], u_ca_out_749[3:2]};
assign col_out_751 = {u_ca_out_751[1:0], u_ca_out_750[3:2]};
assign col_out_752 = {u_ca_out_752[1:0], u_ca_out_751[3:2]};
assign col_out_753 = {u_ca_out_753[1:0], u_ca_out_752[3:2]};
assign col_out_754 = {u_ca_out_754[1:0], u_ca_out_753[3:2]};
assign col_out_755 = {u_ca_out_755[1:0], u_ca_out_754[3:2]};
assign col_out_756 = {u_ca_out_756[1:0], u_ca_out_755[3:2]};
assign col_out_757 = {u_ca_out_757[1:0], u_ca_out_756[3:2]};
assign col_out_758 = {u_ca_out_758[1:0], u_ca_out_757[3:2]};
assign col_out_759 = {u_ca_out_759[1:0], u_ca_out_758[3:2]};
assign col_out_760 = {u_ca_out_760[1:0], u_ca_out_759[3:2]};
assign col_out_761 = {u_ca_out_761[1:0], u_ca_out_760[3:2]};
assign col_out_762 = {u_ca_out_762[1:0], u_ca_out_761[3:2]};
assign col_out_763 = {u_ca_out_763[1:0], u_ca_out_762[3:2]};
assign col_out_764 = {u_ca_out_764[1:0], u_ca_out_763[3:2]};
assign col_out_765 = {u_ca_out_765[1:0], u_ca_out_764[3:2]};
assign col_out_766 = {u_ca_out_766[1:0], u_ca_out_765[3:2]};
assign col_out_767 = {u_ca_out_767[1:0], u_ca_out_766[3:2]};
assign col_out_768 = {u_ca_out_768[1:0], u_ca_out_767[3:2]};
assign col_out_769 = {u_ca_out_769[1:0], u_ca_out_768[3:2]};
assign col_out_770 = {u_ca_out_770[1:0], u_ca_out_769[3:2]};
assign col_out_771 = {u_ca_out_771[1:0], u_ca_out_770[3:2]};
assign col_out_772 = {u_ca_out_772[1:0], u_ca_out_771[3:2]};
assign col_out_773 = {u_ca_out_773[1:0], u_ca_out_772[3:2]};
assign col_out_774 = {u_ca_out_774[1:0], u_ca_out_773[3:2]};
assign col_out_775 = {u_ca_out_775[1:0], u_ca_out_774[3:2]};
assign col_out_776 = {u_ca_out_776[1:0], u_ca_out_775[3:2]};
assign col_out_777 = {u_ca_out_777[1:0], u_ca_out_776[3:2]};
assign col_out_778 = {u_ca_out_778[1:0], u_ca_out_777[3:2]};
assign col_out_779 = {u_ca_out_779[1:0], u_ca_out_778[3:2]};
assign col_out_780 = {u_ca_out_780[1:0], u_ca_out_779[3:2]};
assign col_out_781 = {u_ca_out_781[1:0], u_ca_out_780[3:2]};
assign col_out_782 = {u_ca_out_782[1:0], u_ca_out_781[3:2]};
assign col_out_783 = {u_ca_out_783[1:0], u_ca_out_782[3:2]};
assign col_out_784 = {u_ca_out_784[1:0], u_ca_out_783[3:2]};
assign col_out_785 = {u_ca_out_785[1:0], u_ca_out_784[3:2]};
assign col_out_786 = {u_ca_out_786[1:0], u_ca_out_785[3:2]};
assign col_out_787 = {u_ca_out_787[1:0], u_ca_out_786[3:2]};
assign col_out_788 = {u_ca_out_788[1:0], u_ca_out_787[3:2]};
assign col_out_789 = {u_ca_out_789[1:0], u_ca_out_788[3:2]};
assign col_out_790 = {u_ca_out_790[1:0], u_ca_out_789[3:2]};
assign col_out_791 = {u_ca_out_791[1:0], u_ca_out_790[3:2]};
assign col_out_792 = {u_ca_out_792[1:0], u_ca_out_791[3:2]};
assign col_out_793 = {u_ca_out_793[1:0], u_ca_out_792[3:2]};
assign col_out_794 = {u_ca_out_794[1:0], u_ca_out_793[3:2]};
assign col_out_795 = {u_ca_out_795[1:0], u_ca_out_794[3:2]};
assign col_out_796 = {u_ca_out_796[1:0], u_ca_out_795[3:2]};
assign col_out_797 = {u_ca_out_797[1:0], u_ca_out_796[3:2]};
assign col_out_798 = {u_ca_out_798[1:0], u_ca_out_797[3:2]};
assign col_out_799 = {u_ca_out_799[1:0], u_ca_out_798[3:2]};
assign col_out_800 = {u_ca_out_800[1:0], u_ca_out_799[3:2]};
assign col_out_801 = {u_ca_out_801[1:0], u_ca_out_800[3:2]};
assign col_out_802 = {u_ca_out_802[1:0], u_ca_out_801[3:2]};
assign col_out_803 = {u_ca_out_803[1:0], u_ca_out_802[3:2]};
assign col_out_804 = {u_ca_out_804[1:0], u_ca_out_803[3:2]};
assign col_out_805 = {u_ca_out_805[1:0], u_ca_out_804[3:2]};
assign col_out_806 = {u_ca_out_806[1:0], u_ca_out_805[3:2]};
assign col_out_807 = {u_ca_out_807[1:0], u_ca_out_806[3:2]};
assign col_out_808 = {u_ca_out_808[1:0], u_ca_out_807[3:2]};
assign col_out_809 = {u_ca_out_809[1:0], u_ca_out_808[3:2]};
assign col_out_810 = {u_ca_out_810[1:0], u_ca_out_809[3:2]};
assign col_out_811 = {u_ca_out_811[1:0], u_ca_out_810[3:2]};
assign col_out_812 = {u_ca_out_812[1:0], u_ca_out_811[3:2]};
assign col_out_813 = {u_ca_out_813[1:0], u_ca_out_812[3:2]};
assign col_out_814 = {u_ca_out_814[1:0], u_ca_out_813[3:2]};
assign col_out_815 = {u_ca_out_815[1:0], u_ca_out_814[3:2]};
assign col_out_816 = {u_ca_out_816[1:0], u_ca_out_815[3:2]};
assign col_out_817 = {u_ca_out_817[1:0], u_ca_out_816[3:2]};
assign col_out_818 = {u_ca_out_818[1:0], u_ca_out_817[3:2]};
assign col_out_819 = {u_ca_out_819[1:0], u_ca_out_818[3:2]};
assign col_out_820 = {u_ca_out_820[1:0], u_ca_out_819[3:2]};
assign col_out_821 = {u_ca_out_821[1:0], u_ca_out_820[3:2]};
assign col_out_822 = {u_ca_out_822[1:0], u_ca_out_821[3:2]};
assign col_out_823 = {u_ca_out_823[1:0], u_ca_out_822[3:2]};
assign col_out_824 = {u_ca_out_824[1:0], u_ca_out_823[3:2]};
assign col_out_825 = {u_ca_out_825[1:0], u_ca_out_824[3:2]};
assign col_out_826 = {u_ca_out_826[1:0], u_ca_out_825[3:2]};
assign col_out_827 = {u_ca_out_827[1:0], u_ca_out_826[3:2]};
assign col_out_828 = {u_ca_out_828[1:0], u_ca_out_827[3:2]};
assign col_out_829 = {u_ca_out_829[1:0], u_ca_out_828[3:2]};
assign col_out_830 = {u_ca_out_830[1:0], u_ca_out_829[3:2]};
assign col_out_831 = {u_ca_out_831[1:0], u_ca_out_830[3:2]};
assign col_out_832 = {u_ca_out_832[1:0], u_ca_out_831[3:2]};
assign col_out_833 = {u_ca_out_833[1:0], u_ca_out_832[3:2]};
assign col_out_834 = {u_ca_out_834[1:0], u_ca_out_833[3:2]};
assign col_out_835 = {u_ca_out_835[1:0], u_ca_out_834[3:2]};
assign col_out_836 = {u_ca_out_836[1:0], u_ca_out_835[3:2]};
assign col_out_837 = {u_ca_out_837[1:0], u_ca_out_836[3:2]};
assign col_out_838 = {u_ca_out_838[1:0], u_ca_out_837[3:2]};
assign col_out_839 = {u_ca_out_839[1:0], u_ca_out_838[3:2]};
assign col_out_840 = {u_ca_out_840[1:0], u_ca_out_839[3:2]};
assign col_out_841 = {u_ca_out_841[1:0], u_ca_out_840[3:2]};
assign col_out_842 = {u_ca_out_842[1:0], u_ca_out_841[3:2]};
assign col_out_843 = {u_ca_out_843[1:0], u_ca_out_842[3:2]};
assign col_out_844 = {u_ca_out_844[1:0], u_ca_out_843[3:2]};
assign col_out_845 = {u_ca_out_845[1:0], u_ca_out_844[3:2]};
assign col_out_846 = {u_ca_out_846[1:0], u_ca_out_845[3:2]};
assign col_out_847 = {u_ca_out_847[1:0], u_ca_out_846[3:2]};
assign col_out_848 = {u_ca_out_848[1:0], u_ca_out_847[3:2]};
assign col_out_849 = {u_ca_out_849[1:0], u_ca_out_848[3:2]};
assign col_out_850 = {u_ca_out_850[1:0], u_ca_out_849[3:2]};
assign col_out_851 = {u_ca_out_851[1:0], u_ca_out_850[3:2]};
assign col_out_852 = {u_ca_out_852[1:0], u_ca_out_851[3:2]};
assign col_out_853 = {u_ca_out_853[1:0], u_ca_out_852[3:2]};
assign col_out_854 = {u_ca_out_854[1:0], u_ca_out_853[3:2]};
assign col_out_855 = {u_ca_out_855[1:0], u_ca_out_854[3:2]};
assign col_out_856 = {u_ca_out_856[1:0], u_ca_out_855[3:2]};
assign col_out_857 = {u_ca_out_857[1:0], u_ca_out_856[3:2]};
assign col_out_858 = {u_ca_out_858[1:0], u_ca_out_857[3:2]};
assign col_out_859 = {u_ca_out_859[1:0], u_ca_out_858[3:2]};
assign col_out_860 = {u_ca_out_860[1:0], u_ca_out_859[3:2]};
assign col_out_861 = {u_ca_out_861[1:0], u_ca_out_860[3:2]};
assign col_out_862 = {u_ca_out_862[1:0], u_ca_out_861[3:2]};
assign col_out_863 = {u_ca_out_863[1:0], u_ca_out_862[3:2]};
assign col_out_864 = {u_ca_out_864[1:0], u_ca_out_863[3:2]};
assign col_out_865 = {u_ca_out_865[1:0], u_ca_out_864[3:2]};
assign col_out_866 = {u_ca_out_866[1:0], u_ca_out_865[3:2]};
assign col_out_867 = {u_ca_out_867[1:0], u_ca_out_866[3:2]};
assign col_out_868 = {u_ca_out_868[1:0], u_ca_out_867[3:2]};
assign col_out_869 = {u_ca_out_869[1:0], u_ca_out_868[3:2]};
assign col_out_870 = {u_ca_out_870[1:0], u_ca_out_869[3:2]};
assign col_out_871 = {u_ca_out_871[1:0], u_ca_out_870[3:2]};
assign col_out_872 = {u_ca_out_872[1:0], u_ca_out_871[3:2]};
assign col_out_873 = {u_ca_out_873[1:0], u_ca_out_872[3:2]};
assign col_out_874 = {u_ca_out_874[1:0], u_ca_out_873[3:2]};
assign col_out_875 = {u_ca_out_875[1:0], u_ca_out_874[3:2]};
assign col_out_876 = {u_ca_out_876[1:0], u_ca_out_875[3:2]};
assign col_out_877 = {u_ca_out_877[1:0], u_ca_out_876[3:2]};
assign col_out_878 = {u_ca_out_878[1:0], u_ca_out_877[3:2]};
assign col_out_879 = {u_ca_out_879[1:0], u_ca_out_878[3:2]};
assign col_out_880 = {u_ca_out_880[1:0], u_ca_out_879[3:2]};
assign col_out_881 = {u_ca_out_881[1:0], u_ca_out_880[3:2]};
assign col_out_882 = {u_ca_out_882[1:0], u_ca_out_881[3:2]};
assign col_out_883 = {u_ca_out_883[1:0], u_ca_out_882[3:2]};
assign col_out_884 = {u_ca_out_884[1:0], u_ca_out_883[3:2]};
assign col_out_885 = {u_ca_out_885[1:0], u_ca_out_884[3:2]};
assign col_out_886 = {u_ca_out_886[1:0], u_ca_out_885[3:2]};
assign col_out_887 = {u_ca_out_887[1:0], u_ca_out_886[3:2]};
assign col_out_888 = {u_ca_out_888[1:0], u_ca_out_887[3:2]};
assign col_out_889 = {u_ca_out_889[1:0], u_ca_out_888[3:2]};
assign col_out_890 = {u_ca_out_890[1:0], u_ca_out_889[3:2]};
assign col_out_891 = {u_ca_out_891[1:0], u_ca_out_890[3:2]};
assign col_out_892 = {u_ca_out_892[1:0], u_ca_out_891[3:2]};
assign col_out_893 = {u_ca_out_893[1:0], u_ca_out_892[3:2]};
assign col_out_894 = {u_ca_out_894[1:0], u_ca_out_893[3:2]};
assign col_out_895 = {u_ca_out_895[1:0], u_ca_out_894[3:2]};
assign col_out_896 = {u_ca_out_896[1:0], u_ca_out_895[3:2]};
assign col_out_897 = {u_ca_out_897[1:0], u_ca_out_896[3:2]};
assign col_out_898 = {u_ca_out_898[1:0], u_ca_out_897[3:2]};
assign col_out_899 = {u_ca_out_899[1:0], u_ca_out_898[3:2]};
assign col_out_900 = {u_ca_out_900[1:0], u_ca_out_899[3:2]};
assign col_out_901 = {u_ca_out_901[1:0], u_ca_out_900[3:2]};
assign col_out_902 = {u_ca_out_902[1:0], u_ca_out_901[3:2]};
assign col_out_903 = {u_ca_out_903[1:0], u_ca_out_902[3:2]};
assign col_out_904 = {u_ca_out_904[1:0], u_ca_out_903[3:2]};
assign col_out_905 = {u_ca_out_905[1:0], u_ca_out_904[3:2]};
assign col_out_906 = {u_ca_out_906[1:0], u_ca_out_905[3:2]};
assign col_out_907 = {u_ca_out_907[1:0], u_ca_out_906[3:2]};
assign col_out_908 = {u_ca_out_908[1:0], u_ca_out_907[3:2]};
assign col_out_909 = {u_ca_out_909[1:0], u_ca_out_908[3:2]};
assign col_out_910 = {u_ca_out_910[1:0], u_ca_out_909[3:2]};
assign col_out_911 = {u_ca_out_911[1:0], u_ca_out_910[3:2]};
assign col_out_912 = {u_ca_out_912[1:0], u_ca_out_911[3:2]};
assign col_out_913 = {u_ca_out_913[1:0], u_ca_out_912[3:2]};
assign col_out_914 = {u_ca_out_914[1:0], u_ca_out_913[3:2]};
assign col_out_915 = {u_ca_out_915[1:0], u_ca_out_914[3:2]};
assign col_out_916 = {u_ca_out_916[1:0], u_ca_out_915[3:2]};
assign col_out_917 = {u_ca_out_917[1:0], u_ca_out_916[3:2]};
assign col_out_918 = {u_ca_out_918[1:0], u_ca_out_917[3:2]};
assign col_out_919 = {u_ca_out_919[1:0], u_ca_out_918[3:2]};
assign col_out_920 = {u_ca_out_920[1:0], u_ca_out_919[3:2]};
assign col_out_921 = {u_ca_out_921[1:0], u_ca_out_920[3:2]};
assign col_out_922 = {u_ca_out_922[1:0], u_ca_out_921[3:2]};
assign col_out_923 = {u_ca_out_923[1:0], u_ca_out_922[3:2]};
assign col_out_924 = {u_ca_out_924[1:0], u_ca_out_923[3:2]};
assign col_out_925 = {u_ca_out_925[1:0], u_ca_out_924[3:2]};
assign col_out_926 = {u_ca_out_926[1:0], u_ca_out_925[3:2]};
assign col_out_927 = {u_ca_out_927[1:0], u_ca_out_926[3:2]};
assign col_out_928 = {u_ca_out_928[1:0], u_ca_out_927[3:2]};
assign col_out_929 = {u_ca_out_929[1:0], u_ca_out_928[3:2]};
assign col_out_930 = {u_ca_out_930[1:0], u_ca_out_929[3:2]};
assign col_out_931 = {u_ca_out_931[1:0], u_ca_out_930[3:2]};
assign col_out_932 = {u_ca_out_932[1:0], u_ca_out_931[3:2]};
assign col_out_933 = {u_ca_out_933[1:0], u_ca_out_932[3:2]};
assign col_out_934 = {u_ca_out_934[1:0], u_ca_out_933[3:2]};
assign col_out_935 = {u_ca_out_935[1:0], u_ca_out_934[3:2]};
assign col_out_936 = {u_ca_out_936[1:0], u_ca_out_935[3:2]};
assign col_out_937 = {u_ca_out_937[1:0], u_ca_out_936[3:2]};
assign col_out_938 = {u_ca_out_938[1:0], u_ca_out_937[3:2]};
assign col_out_939 = {u_ca_out_939[1:0], u_ca_out_938[3:2]};
assign col_out_940 = {u_ca_out_940[1:0], u_ca_out_939[3:2]};
assign col_out_941 = {u_ca_out_941[1:0], u_ca_out_940[3:2]};
assign col_out_942 = {u_ca_out_942[1:0], u_ca_out_941[3:2]};
assign col_out_943 = {u_ca_out_943[1:0], u_ca_out_942[3:2]};
assign col_out_944 = {u_ca_out_944[1:0], u_ca_out_943[3:2]};
assign col_out_945 = {u_ca_out_945[1:0], u_ca_out_944[3:2]};
assign col_out_946 = {u_ca_out_946[1:0], u_ca_out_945[3:2]};
assign col_out_947 = {u_ca_out_947[1:0], u_ca_out_946[3:2]};
assign col_out_948 = {u_ca_out_948[1:0], u_ca_out_947[3:2]};
assign col_out_949 = {u_ca_out_949[1:0], u_ca_out_948[3:2]};
assign col_out_950 = {u_ca_out_950[1:0], u_ca_out_949[3:2]};
assign col_out_951 = {u_ca_out_951[1:0], u_ca_out_950[3:2]};
assign col_out_952 = {u_ca_out_952[1:0], u_ca_out_951[3:2]};
assign col_out_953 = {u_ca_out_953[1:0], u_ca_out_952[3:2]};
assign col_out_954 = {u_ca_out_954[1:0], u_ca_out_953[3:2]};
assign col_out_955 = {u_ca_out_955[1:0], u_ca_out_954[3:2]};
assign col_out_956 = {u_ca_out_956[1:0], u_ca_out_955[3:2]};
assign col_out_957 = {u_ca_out_957[1:0], u_ca_out_956[3:2]};
assign col_out_958 = {u_ca_out_958[1:0], u_ca_out_957[3:2]};
assign col_out_959 = {u_ca_out_959[1:0], u_ca_out_958[3:2]};
assign col_out_960 = {u_ca_out_960[1:0], u_ca_out_959[3:2]};
assign col_out_961 = {u_ca_out_961[1:0], u_ca_out_960[3:2]};
assign col_out_962 = {u_ca_out_962[1:0], u_ca_out_961[3:2]};
assign col_out_963 = {u_ca_out_963[1:0], u_ca_out_962[3:2]};
assign col_out_964 = {u_ca_out_964[1:0], u_ca_out_963[3:2]};
assign col_out_965 = {u_ca_out_965[1:0], u_ca_out_964[3:2]};
assign col_out_966 = {u_ca_out_966[1:0], u_ca_out_965[3:2]};
assign col_out_967 = {u_ca_out_967[1:0], u_ca_out_966[3:2]};
assign col_out_968 = {u_ca_out_968[1:0], u_ca_out_967[3:2]};
assign col_out_969 = {u_ca_out_969[1:0], u_ca_out_968[3:2]};
assign col_out_970 = {u_ca_out_970[1:0], u_ca_out_969[3:2]};
assign col_out_971 = {u_ca_out_971[1:0], u_ca_out_970[3:2]};
assign col_out_972 = {u_ca_out_972[1:0], u_ca_out_971[3:2]};
assign col_out_973 = {u_ca_out_973[1:0], u_ca_out_972[3:2]};
assign col_out_974 = {u_ca_out_974[1:0], u_ca_out_973[3:2]};
assign col_out_975 = {u_ca_out_975[1:0], u_ca_out_974[3:2]};
assign col_out_976 = {u_ca_out_976[1:0], u_ca_out_975[3:2]};
assign col_out_977 = {u_ca_out_977[1:0], u_ca_out_976[3:2]};
assign col_out_978 = {u_ca_out_978[1:0], u_ca_out_977[3:2]};
assign col_out_979 = {u_ca_out_979[1:0], u_ca_out_978[3:2]};
assign col_out_980 = {u_ca_out_980[1:0], u_ca_out_979[3:2]};
assign col_out_981 = {u_ca_out_981[1:0], u_ca_out_980[3:2]};
assign col_out_982 = {u_ca_out_982[1:0], u_ca_out_981[3:2]};
assign col_out_983 = {u_ca_out_983[1:0], u_ca_out_982[3:2]};
assign col_out_984 = {u_ca_out_984[1:0], u_ca_out_983[3:2]};
assign col_out_985 = {u_ca_out_985[1:0], u_ca_out_984[3:2]};
assign col_out_986 = {u_ca_out_986[1:0], u_ca_out_985[3:2]};
assign col_out_987 = {u_ca_out_987[1:0], u_ca_out_986[3:2]};
assign col_out_988 = {u_ca_out_988[1:0], u_ca_out_987[3:2]};
assign col_out_989 = {u_ca_out_989[1:0], u_ca_out_988[3:2]};
assign col_out_990 = {u_ca_out_990[1:0], u_ca_out_989[3:2]};
assign col_out_991 = {u_ca_out_991[1:0], u_ca_out_990[3:2]};
assign col_out_992 = {u_ca_out_992[1:0], u_ca_out_991[3:2]};
assign col_out_993 = {u_ca_out_993[1:0], u_ca_out_992[3:2]};
assign col_out_994 = {u_ca_out_994[1:0], u_ca_out_993[3:2]};
assign col_out_995 = {u_ca_out_995[1:0], u_ca_out_994[3:2]};
assign col_out_996 = {u_ca_out_996[1:0], u_ca_out_995[3:2]};
assign col_out_997 = {u_ca_out_997[1:0], u_ca_out_996[3:2]};
assign col_out_998 = {u_ca_out_998[1:0], u_ca_out_997[3:2]};
assign col_out_999 = {u_ca_out_999[1:0], u_ca_out_998[3:2]};
assign col_out_1000 = {u_ca_out_1000[1:0], u_ca_out_999[3:2]};
assign col_out_1001 = {u_ca_out_1001[1:0], u_ca_out_1000[3:2]};
assign col_out_1002 = {u_ca_out_1002[1:0], u_ca_out_1001[3:2]};
assign col_out_1003 = {u_ca_out_1003[1:0], u_ca_out_1002[3:2]};
assign col_out_1004 = {u_ca_out_1004[1:0], u_ca_out_1003[3:2]};
assign col_out_1005 = {u_ca_out_1005[1:0], u_ca_out_1004[3:2]};
assign col_out_1006 = {u_ca_out_1006[1:0], u_ca_out_1005[3:2]};
assign col_out_1007 = {u_ca_out_1007[1:0], u_ca_out_1006[3:2]};
assign col_out_1008 = {u_ca_out_1008[1:0], u_ca_out_1007[3:2]};
assign col_out_1009 = {u_ca_out_1009[1:0], u_ca_out_1008[3:2]};
assign col_out_1010 = {u_ca_out_1010[1:0], u_ca_out_1009[3:2]};
assign col_out_1011 = {u_ca_out_1011[1:0], u_ca_out_1010[3:2]};
assign col_out_1012 = {u_ca_out_1012[1:0], u_ca_out_1011[3:2]};
assign col_out_1013 = {u_ca_out_1013[1:0], u_ca_out_1012[3:2]};
assign col_out_1014 = {u_ca_out_1014[1:0], u_ca_out_1013[3:2]};
assign col_out_1015 = {u_ca_out_1015[1:0], u_ca_out_1014[3:2]};
assign col_out_1016 = {u_ca_out_1016[1:0], u_ca_out_1015[3:2]};
assign col_out_1017 = {u_ca_out_1017[1:0], u_ca_out_1016[3:2]};
assign col_out_1018 = {u_ca_out_1018[1:0], u_ca_out_1017[3:2]};
assign col_out_1019 = {u_ca_out_1019[1:0], u_ca_out_1018[3:2]};
assign col_out_1020 = {u_ca_out_1020[1:0], u_ca_out_1019[3:2]};
assign col_out_1021 = {u_ca_out_1021[1:0], u_ca_out_1020[3:2]};
assign col_out_1022 = {u_ca_out_1022[1:0], u_ca_out_1021[3:2]};
assign col_out_1023 = {u_ca_out_1023[1:0], u_ca_out_1022[3:2]};
assign col_out_1024 = {{2{1'b0}}, u_ca_out_1023[3:2]};

//---------------------------------------------------------


endmodule
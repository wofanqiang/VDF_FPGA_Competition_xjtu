module xpb_5_110
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5d2e3ffa4315d9f8b41f139c00ff726eab8c34bf110a4ea775fdaf29b43f6b1a8b2efe18df518f983fd29a09a70aedff48adc372d500b06ee31cda6e2a1683d670b92a4b913d101826f344101aa8f3cfb34fd36ce0a5f6775cac9bc73d0319ce0e96b574229c5d3bb64591d44ae8f0d37e7a5825e8f1616c7c6ae56716b9e355;
    5'b00010 : xpb = 1024'h9af3a9ec43d7f289d38af60f1a49d8be5a2664d4c9cfcd76e1ea4fdb57c292d13157eb8f47ca0a1e046f4cc6ab7cb342d415eff874e9092159a757e195a92fb6d231fe872e922eb3b4c857d9c76236e729aad4134c5bfde03cca593bfdb9109ee25d8be946fc1e9e5cb3cc99e01bb7dae1ad169819765a8b2664fc9a491603f;
    5'b00011 : xpb = 1024'h66dd7a99075359215157c2fcf2a40ffa912e9b0c5da74b7ee41c542769bb94479e447cd1d3ce303a20198ed611c2b93375ef22725c4f4100f8b74fec437116d1dddc4a3404263303623fc98db71f173e25ea80ae156bb6556079415afcdeaad7fcbc8e32b70c1f259c10ce9de8eaac512c95298f6a88c7152ed13530bb4b4394;
    5'b00100 : xpb = 1024'h135e753d887afe513a715ec1e3493b17cb44cc9a9939f9aedc3d49fb6af8525a262afd71e8f94143c08de998d56f96685a82bdff0e9d21242b34eafc32b525f6da463fd0e5d245d676990afb38ec46dce5355a82698b7fbc07994b277fb72213dc4bb17d28df83d3cb9679933c0376fb5c35a2d3032ecb5164cc9f934922c07e;
    5'b00101 : xpb = 1024'h708cb537cb90d849ee90725de448ad8676d10159aa444856523af9251f37bd74b159fb8ac84ad0dc006083a27c7a8467a3308171e39dd1930e51c56a5ccba9cd4aff6a1c770f55ee9d8c4f0b53953aac98852def4a3176336445e6eebcba3be1eae266f14b7be10f81dc0b6786ec67cedaaffaf8ec202cbde13784fa5fdca3d3;
    5'b00110 : xpb = 1024'h1d0dafdc4cb87d79d7aa0e22d4edd8a3b0e732e7e5d6f6864a5beef920747b8739407c2add75e1e5a0d4de654027619c87c41cfe95ebb1b640cf607a4c0fb8f247695fb958bb68c1b1e59078d5626a4b57d007c39e513f9a0b65f0bb3f92b31dca718a3bbd4f45bdb161b65cda0532790a50743c84c630fa1732ef5cedb420bd;
    5'b00111 : xpb = 1024'h7a3befd68fce57728bc921bed5ed4b125c7367a6f6e1452dc0599e22d4b3e6a1c46f7a43bcc7717de0a7786ee7324f9bd071e0716aec622523ec3ae876263cc8b8228a04e9f878d9d8d8d488f00b5e1b0b1fdb307ef7361168128c827c95ccebd9083fafdfeba2f967a7483124ee234c88cacc626db79266939dd4c4046e0412;
    5'b01000 : xpb = 1024'h26bcea7b10f5fca274e2bd83c692762f968999353273f35db87a93f6d5f0a4b44c55fae3d1f28287811bd331aadf2cd0b5057bfe1d3a42485669d5f8656a4bedb48c7fa1cba48baced3215f671d88db9ca6ab504d316ff780f32964eff6e4427b89762fa51bf07a7972cf3267806edf6b86b45a6065d96a2c9993f26924580fc;
    5'b01001 : xpb = 1024'h83eb2a75540bd69b2901d11fc791e89e4215cdf4437e42052e7843208a300fced784f8fcb144121fc0ee6d3b51ea1acffdb33f70f23af2b73986b0668f80cfc42545a9ed5ce19bc514255a068c8181897dba8871b3bcf5ef6bdf32163c715df5c72e186e745b64e34d7284fac2efdeca36e59dcbef4ef80f4604248da8ff6451;
    5'b01010 : xpb = 1024'h306c2519d5337bcb121b6ce4b83713bb7c2bff827f10f035269938f48b6ccde15f6b799cc66f23296162c7fe1596f804e246dafda488d2da6c044b767ec4dee921af9f8a3e8dae98287e9b740e4eb1283d05624607dcbf5612ff3be2bf49d531a6bd3bb8e62ec9917cf82ff01608a9746686170f87f4fc4b7bff8ef036d6e13b;
    5'b01011 : xpb = 1024'h8d9a6514184955c3c63a8080b936862a27b83441901b3edc9c96e81e3fac38fbea9a77b5a5c0b2c1a1356207bca1e6042af49e70798983494f2125e4a8db62bf9268c9d5cfcabeb04f71df8428f7a4f7f05535b2e882b5cd6fabd7a9fc4ceeffb553f12d08cb26cd333dc1c460f19a47e5006f3570e65db7f86a74574d90c490;
    5'b01100 : xpb = 1024'h3a1b5fb89970faf3af541c45a9dbb14761ce65cfcbaded0c94b7ddf240e8f70e7280f855baebc3cb41a9bcca804ec3390f8839fd2bd7636c819ec0f4981f71e48ed2bf72b176d18363cb20f1aac4d496afa00f873ca27f3416cbe1767f25663b94e314777a9e8b7b62c36cb9b40a64f214a0e879098c61f42e65deb9db68417a;
    5'b01101 : xpb = 1024'h97499fb2dc86d4ec63732fe1aadb23b60d5a9a8edcb83bb40ab58d1bf5286228fdaff66e9a3d5363817c56d42759b1385835fd7000d813db64bb9b62c235f5baff8be9be42b3e19b8abe6501c56dc86662efe2f41d4875ab73787d3dbc288009a379c9eb9d3ae8b71908fe8dfef355c5931b409ef27dc360aad0c420f22224cf;
    5'b01110 : xpb = 1024'h43ca9a575dae7a1c4c8ccba69b804ed34770cc1d184ae9e402d682eff665203b8596770eaf68646d21f0b196eb068e6d3cc998fcb325f3fe97393672b17a04dffbf5df5b245ff46e9f17a66f473af805223abcc871683f121a98870a3f00f7458308ed360f0e4d65488ea983520c206fc2bbb9e28b23c79ce0cc2e837ff9a1b9;
    5'b01111 : xpb = 1024'ha0f8da51a0c4541500abdf429c7fc141f2fd00dc2955388b78d43219aaa48b5610c575278eb9f40561c34ba092117c6c85775c6f8826a46d7a5610e0db9088b66caf09a6b59d0486c60aea7f61e3ebd4d58a9035520e3589774522d17c041113919fa2aa31aaaaa0fed43b579cf5114341361208741529095d3713ea96b3850e;
    5'b10000 : xpb = 1024'h4d79d4f621ebf944e9c57b078d24ec5f2d13326a64e7e6bb70f527edabe1496898abf5c7a3e5050f0237a66355be59a16a0af7fc3a748490acd3abf0cad497db6918ff4397491759da642bece3b11b7394d56a09a62dfef01e652c9dfedc884f712ec5f4a37e0f4f2e59e64cf00ddbed70d68b4c0cbb2d4593327e4d248b01f8;
    5'b10001 : xpb = 1024'haaa814f06501d33d9de48ea38e245ecdd89f672975f23562e6f2d7176020b48323daf3e0833694a7420a406cfcc947a0b2b8bb6f0f7534ff8ff0865ef4eb1bb1d9d2298f2886277201576ffcfe5a0f4348253d7686d3f5677b11c8653bdfa21d7fc57b68c61a6c8ae49f78213af6ccc0ef50e371f5ac8eb20f9d63b43b44e54d;
    5'b10010 : xpb = 1024'h57290f94e629786d86fe2a687ec989eb12b598b7b184e392df13cceb615d7295abc174809861a5b0e27e9b2fc07624d5974c56fbc1c31522c26e216ee42f2ad6d63c1f2c0a323a4515b0b16a80273ee20770174adaf3bece2231d231beb819595f549eb337edd139142523168e0f976b1ef15cb58e5292ee4598ce16c91c6237;
    5'b10011 : xpb = 1024'h3aa0a3967511d9d7017c62d6f6eb5084ccbca45ed1791c2d734c2bf629a30a833a7f520ad8cb6ba82f2f5f28423020a7bdff2887410f545f4ebbc7ed37339fbd2a614c8ebde4d182a09f2d801f46e80c6baf11f2f138834c951dbfe419090953ee3c1fda9c135e743aace0be12862154e91d5f926f8972a7b94387956f3df21;
    5'b10100 : xpb = 1024'h60d84a33aa66f7962436d9c9706e2776f857ff04fe21e06a4d3271e916d99bc2bed6f3398cde4652c2c58ffc2b2df009c48db5fb4911a5b4d80896ecfd89bdd2435f3f147d1b5d3050fd36e81c9d62507a0ac48c0fb97eac25fe77c57e93aa634d7a7771cc5d9322f9f05fe02c1152e8cd0c2e1f0fe9f896f7ff1de06dadc276;
    5'b10101 : xpb = 1024'hd5944d82b8e9cc60d50758e61135294326e309339b48e9a455367bd181659d546bd73d9a209575c6339eabeeedacd3ea9215187fb5f85d80a8631fceccdccf73fc934b15ec77003655678559e6a91ef39559e6063d94812cd1e8192016c219f2d099abc3e30f7d129760ad57f2a1d92fcaca762a88ffcd32dfa8842fb853f60;
    5'b10110 : xpb = 1024'h6a8784d26ea476bec16f892a6212c502ddfa65524abedd41bb5116e6cc55c4efd1ec71f2815ae6f4a30c84c895e5bb3df1cf14fad0603646eda30c6b16e450cdb0825efcf004801b8c49bc65b91385beeca571cd447f3e8a29cb1d593e6f3b6d3ba0503060cd550cdfbb9ca9ca130e667b26ff8891815e3faa656daa123f22b5;
    5'b10111 : xpb = 1024'h17087f76efcc1beeaa8924ef52b7f020181096e086518b71b3720cbacd92830259d2f2929685f7fe4380df8b59929872d662b08782ae166a2020a77b06285ff2acec5499d1b092eea0a2fdd33ae0b55dabf04ba1989f07f0d0eb2725c147b2a91b2f737ad2a0b9bb0f41479f1d2bd910aac778cc2a27627be060d80ca0169f9f;
    5'b11000 : xpb = 1024'h7436bf7132e1f5e75ea8388b53b7628ec39ccb9f975bda19296fbbe481d1ee1ce501f0ab75d7879683537995009d86721f1073fa57aec6d9033d81e9303ee3c91da57ee562eda306c79641e35589a92d5f401f0e7944fe682d97c2ecfe4acc7729c628eef53d16f6c586d9736814c9e42941d0f21318c3e85ccbbd73b6d082f4;
    5'b11001 : xpb = 1024'h20b7ba15b4099b1747c1d450445c8dabfdb2fd2dd2ee88492190b1b8830eac2f6ce8714b8b0298a023c7d457c44a63a703a40f8709fca6fc35bb1cf91f82f2ee1a0f74824499b5d9dbef8350d756d8cc1e8af8e2cd64c7ced4b7ccb9812343b309554c3967107ba4f50c8468bb2d948e58e24a35abbec82492c727d644a7ffde;
    5'b11010 : xpb = 1024'h7de5fa0ff71f750ffbe0e7ec455c001aa93f31ece3f8d6f0978e60e2374e1749f8176f646a542838639a6e616b5551a64c51d2f9defd576b18d7f767499976c48ac89ecdd5d6c5f202e2c760f1ffcc9bd1dacc4fae0abe4631646880be265d8117ec01ad89acd8e0ab52163d06168561d75ca25b94b029910f320d3d5b61e333;
    5'b11011 : xpb = 1024'h2a66f4b478471a3fe4fa83b136012b37e355637b1f8b85208faf56b6388ad55c7ffdf0047f7f3942040ec9242f022edb30e56e86914b378e4b55927738dd85e98732946ab782d8c5173c08ce73ccfc3a9125a624022a87acd884724d40fed4bcf77b24f7fb803d8edad7c132592f500c06fd1b9f2d562dcd452d779fe939601d;
    5'b11100 : xpb = 1024'h879534aebb5cf4389919974d37009da68ee1983a3095d3c805ad05dfecca40770b2cee1d5ed0c8da43e1632dd60d1cda799331f9664be7fd2e726ce562f409bff7ebbeb648bfe8dd3e2f4cde8e75f00a44757990e2d07e2435310e147e01ee8b0611da6c1e1c9aca911d5306a41840df857773c516478f39c1985d06fff34372;
    5'b11101 : xpb = 1024'h34162f533c8499688233331227a5c8c3c8f7c9c86c2881f7fdcdfbb3ee06fe8993136ebd73fbd9e3e455bdf099b9fa0f5e26cd861899c82060f007f5523818e4f455b4532a6bfbb052888e4c10431fa903c0536536f0478adc5117e100da65c6e5a0fdb68fefff78c0a2fdfbf7310b89b517ed08aeed9375f793c7698dcac05c;
    5'b11110 : xpb = 1024'h91446f4d7f9a7361365246ae28a53b327483fe877d32d09f73cbaadda24669a41e426cd6534d697c242857fa40c4e80ea6d490f8ed9a788f440ce2637c4e9cbb650ede9ebba90bc8797bd25c2aec1378b71026d217963e0238fdb3a83ddd7f94f437b32ab28c5cb476e88fd04219fc5d3392452e97def4e273feacd0a484a3b1;
    5'b11111 : xpb = 1024'h3dc569f200c218911f6be273194a664fae9a3015b8c57ecf6beca0b1a38327b6a628ed7668787a85c49cb2bd0471c5438b682c859fe858b2768a7d736b92abe06178d43b9d551e9b8dd513c9acb94317765b00a66bb60768e01dbd74c0b5f6d0d3c6d675245fc162a66e3ac59532c7076332be723084f91ea9fa1733325c209b;
    endcase
end

endmodule

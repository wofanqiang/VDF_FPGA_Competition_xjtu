module xpb_5_960
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h724dba974c4ea5a204f914483b7d57a206fe7f72b452eba7add72ccb0b9817d5d9d76d486fa7468c84ca0fae60919ffcce7572e42565141c345812739f550e06149c4df373764d0b6f126774eebe706f7bea7597e46942b2587a1f5bde45c86dc8862fb7d45849333c6a98f40767f453a50b6cbcd5e4ac2bdb9ef2884a47934a;
    5'b00010 : xpb = 1024'h33ee2fd8d6af167b3eecb0b966a067f29c86fbb4932e36d7ddd1a040642d82a3b0665d1815280e8a6a35e015ddc52f2f38d0bde2281757ecb810e58903d7a75ab4e96738375b9cd1cb8acc4744a11cae03cff1973c4c5853fb67acbd0260ee496204cd45f7e799d8f2154b0916ffc27dfb3cfa975b7dfb2770ce6a0c0bacc029;
    5'b00011 : xpb = 1024'ha63bea7022fdbc1d43e5c501a21dbf94a3857b274781227f8ba8cd0b6fc59a798a3dca6084cf5516eeffefc43e56cf2c074630c64d7c6c08ec68f7fca32cb560c985b52baad1e9dd3a9d33bc335f8d1d7fba672f20b59b0653e1cc18e0a6b6b72a8afcfdcc3fe30c2e7fe3fd1e67b6d1a04867543162a7534c6d5c9455f45373;
    5'b00100 : xpb = 1024'h67dc5fb1ad5e2cf67dd96172cd40cfe5390df769265c6dafbba34080c85b054760ccba302a501d14d46bc02bbb8a5e5e71a17bc4502eafd97021cb1207af4eb569d2ce706eb739a39715988e8942395c079fe32e7898b0a7f6cf597a04c1dc92c4099a8befcf33b1e42a96122dff84fbf679f52eb6fbf64ee19cd41817598052;
    5'b00101 : xpb = 1024'h297cd4f337be9dcfb7ccfde3f863e035ce9673ab0537b8dfeb9db3f620f07015375ba9ffcfd0e512b9d7909338bded90dbfcc6c252e0f3a9f3da9e276c31e80a0a1fe7b5329c8969f38dfd60df24e59a8f855f2dd07bc64999bce6db28dd026e5d88381a135e845799d548273d9753264cab83093c95454a76cc4b9bd8bead31;
    5'b00110 : xpb = 1024'h9bca8f8a840d4371bcc6122c33e137d7d594f31db98aa4879974e0c12c8887eb113317483f782b9f3ea1a041994f8d8daa7239a6784607c62832b09b0b86f6101ebc35a8a612d67562a064d5cde3560a0b6fd4c5b4e508fbf23706370722cadc260e67d1e7b6cd8ad63fe11b44ff4779f1b6efc61279f176526b3e242306407b;
    5'b00111 : xpb = 1024'h5d6b04cc0e6db44af6b9ae9d5f0448286b1d6f5f9865efb7c96f5436851df2b8e7c20717e4f8f39d240d70a916831cc014cd84a47af84b96abeb83b070098f64bf094eed69f8263bbf18c9a823c60248935550c50cc81e9d952493982b3df0b7bf8d05600b461e308bea9330549715a447e87da098134071e79ab5a7e46b6d5a;
    5'b01000 : xpb = 1024'h1f0b7a0d98ce252430ad4b0e8a27587900a5eba177413ae7f969c7abddb35d86be50f6e78a79bb9b0979411093b6abf27f28cfa27daa8f672fa456c5d48c28b95f5668322ddd76021b912e7a79a8ae871b3accc464ab343f381220f94f591693590ba2ee2ed56ed641954545642ee3ce9e1a0b7b1dac8f6d7cca2d2ba5d09a39;
    5'b01001 : xpb = 1024'h915934a4e51ccac635a65f56c5a4b01b07a46b142b94268fa740f476e94b755c9828642ffa2102278e4350bef4484bef4d9e4286a30fa38363fc693973e136bf73f2b625a153c30d8aa395ef68671ef69725425c491476f1908c40552d9edf012191d2a6032db8097dffde396b96d82243257837f3913b9958691fb3f0182d83;
    5'b01010 : xpb = 1024'h52f9a9e66f7d3b9f6f99fbc7f0c7c06b9d2ce7560a6f71bfd73b67ec41e0e02a6eb753ff9fa1ca2573af2126717bdb21b7f98d84a5c1e753e7b53c4ed863d014143fcf6a653912d3e71bfac1be49cb351f0abe5ba0f78c933379cdb651ba04dcbb10703426bd08af33aa904e7b2ea64c99570612792a8a94ed989737b17d5a62;
    5'b01011 : xpb = 1024'h149a1f27f9ddac78a98d98391bead0bc32b56397e94abcf00735db619a764af8454643cf45229223591af18deeaf6a542254d882a8742b246b6e0f643ce66968b48ce8af291e629a43945f94142c7773a6f03a5af8daa234d6675b1775d52ab8548f0dc24a4c5954e95542638ac67476ef8893ecfec3d99082c80ebb72e28741;
    5'b01100 : xpb = 1024'h86e7d9bf462c521aae86ac815768285e39b3e30a9d9da897b50d082ca60e62ce1f1db117b4c9d8afdde5013c4f410a50f0ca4b66cdd93f409fc621d7dc3b776ec92936a29c94afa5b2a6c70902eae7e322daaff2dd43e4e72ee17a73541af3261d153d7a1ea4a28825bfdb57922e68ca949400a9d4a885bc5e670143bd2a1a8b;
    5'b01101 : xpb = 1024'h48884f00d08cc2f3e87a48f2828b38aecf3c5f4c7c78f3c7e5077ba1fea3cd9bf5aca0e75a4aa0adc350d1a3cc7499835b259664d08b8311237ef4ed40be10c369764fe76079ff6c0f1f2bdb58cd9421aac02bf23526fa88d1cf07d478361901b693db084233f32ddb6a8d6ca1c636f4eac58e845a41d4b7f39678c77e8f476a;
    5'b01110 : xpb = 1024'ha28c4425aed33cd226de563adae48ff64c4db8e5b543ef81501ef1757393869cc3b90b6ffcb68aba8bca20b49a828b5c580e162d33dc6e1a737c802a540aa1809c3692c245f4f326b9790adaeb0406032a5a7f18d0a102a74bc95359c513edd5012789665c343d391153f81b15e051f40f71c5edfdb23b388c5f04b3ff47449;
    5'b01111 : xpb = 1024'h7c767ed9a73bd96f2766f9abe92ba0a16bc35b010fa72a9fc2d91be262d1503fa612fdff6f72af382d86b1b9aa39c8b293f65446f8a2dafddb8fda764495b81e1e5fb71f97d59c3ddaa9f8229d6eb0cfae901d89717352dccd36b4917a97074b1898a84e3a1b8d06cd7fd875b8c5f972e602891bb5bfcfdf6464e2d38a3c0793;
    5'b10000 : xpb = 1024'h3e16f41b319c4a48615a961d144eb0f2014bd742ee8275cff2d38f57bb66bb0d7ca1edcf14f3773612f28221276d57e4fe519f44fb551ece5f48ad8ba9185172beacd0645bbaec0437225cf4f3515d0e36759988c956687e702441f29eb22d26b21745dc5daaddac832a8a8ac85dc79d3c3416f63b591edaf9945a574ba13472;
    5'b10001 : xpb = 1024'hb064aeb27deaefea6653aa654fcc0894084a56b5a2d56177a0aabc22c6fed2e356795b17849abdc297bc91cf87fef7e1ccc7122920ba32ea93a0bfff486d5f78d3491e57cf31390fa634c469e20fcd7db2600f20adbfab30c89e614e7cf7f5947a9d7594320326dfbf95237ecfc5bbf0e13f83b3113dcb06d5334cdf95e8c7bc;
    5'b10010 : xpb = 1024'h720523f4084b60c3a04746d67aef18e49dd2d2f781b0aca7d0a52f981f943db12d084ae72a1b85c07d2862370532871437225d27236c76bb17599314aceff8cd7396379c931688d602ad293c37f279bc3a458b2005a2c0d26b8beeafa1131b70141c132255927785753fd593df5d8a1b3771118d96d71a026a62c463574df49b;
    5'b10011 : xpb = 1024'h33a5993592abd19cda3ae347a6122935335b4f39608bf7d8009fa30d7829a87f03973ab6cf9c4dbe6294329e82661646a17da825261eba8b9b12662a1172922213e350e156fbd89c5f258e0e8dd525fac22b071f5d85d6740e797c10c52e414bad9ab0b07921c82b2aea87a8eef558458da29f681c7068fdff923be718b3217a;
    5'b10100 : xpb = 1024'ha5f353ccdefa773edf33f78fe18f80d73a59ceac14dee37fae76cfd883c1c054dd6ea7ff3f43944ae75e424ce2f7b6436ff31b094b83cea7cf6a789db0c7a028287f9ed4ca7225a7ce37f5837c93966a3e157cb741ef192666f39b6ca37409b97620e0684d7a115e6755209cf65d4c9932ae0c24f2551529db312e6f62fab4c4;
    5'b10101 : xpb = 1024'h6793c90e695ae818192794010cb29127cfe24aedf3ba2eafde71434ddc572b22b3fd97cee4c45c48ccca12b4602b4575da4e66074e36127853234bb3154a397cc8ccb8198e57756e2ab05a55d27642a8c5faf8b699d22ec809e128cdc78f2f950f9f7df6710962041cffd2b205f51ac388df99ff77ee64257060a5f3245fe1a3;
    5'b10110 : xpb = 1024'h29343e4ff3bb58f1531b307237d5a178656ac72fd29579e00e6bb6c334ec95f08a8c879e8a452446b235e31bdd5ed4a844a9b10550e85648d6dc1ec879ccd2d16919d15e523cc5348728bf282858eee74de074b5f1b54469acceb62eebaa5570a91e1b849498b2a9d2aa84c7158ce8eddf1127d9fd87b32105901d76e5c50e82;
    5'b10111 : xpb = 1024'h9b81f8e74009fe93581444ba7352f91a6c6946a286e86587bc42e38e4084adc66463f4e6f9ec6ad336fff2ca3df074a5131f23e9764d6a650b34313c1921e0d77db61f51c5b3123ff63b269d17175f56c9caea4dd61e871c0548d58ac9f01dde71a44b3c68f0fbdd0f151dbb1cf4dd41841c9496d36c5f4ce12f0fff300ca1cc;
    5'b11000 : xpb = 1024'h5d226e28ca6a6f6c9207e12b9e76096b01f1c2e465c3b0b7ec3d5703991a18943af2e4b69f6d32d11c6bc331bb2403d77d7a6ee778ffae358eed04517da47a2c1e0338968998620652b38b6f6cfa0b9551b0664d2e019cbda83662ebee0b43ba0b22e8ca8c804c82c4bfcfd02c8cab6bda4e22715905ae48765e8782f171ceab;
    5'b11001 : xpb = 1024'h1ec2e36a54cae045cbfb7d9cc99919bb977a3f26449efbe81c37ca78f1af83621181d48644edfacf01d7939938579309e7d5b9e57bb1f20612a5d766e2271380be5051db4d7db1ccaf2bf041c2dcb7d3d995e24c85e4b25f4b23f04d12266995a4a18658b00f9d287a6a81e53c247996307fb04bde9efd440b8dff06b2d6fb8a;
    5'b11010 : xpb = 1024'h91109e01a11985e7d0f491e50516715d9e78be98f8f1e78fca0ef743fd479b37eb5941ceb495415b86a1a34798e93306b64b2cc9a117062246fde9da817c2186d2ec9fcec0f3fed81e3e57b6b19b2843558057e46a4df511a39e0fa8f06c32036d27b6108467e65bb6d51ad9438c6de9d58b1d08b483a96fe72cf18efd1e8ed4;
    5'b11011 : xpb = 1024'h52b113432b79f6c10ae82e56303981ae34013adad7cd32bffa096ab955dd0605c1e8319e5a1609596c0d73af161cc23920a677c7a3c949f2cab6bcefe5febadb7339b91384d94e9e7ab6bc89077dd481dd65d3e3c2310ab3468b9d0a148757df06a6539ea7f737016c7fccee53243c142bbcaae33a1cf86b7c5c6912be83bbb3;
    5'b11100 : xpb = 1024'h14518884b5da679a44dbcac75b5c91fec989b71cb6a87df02a03de2eae7270d39877216dff96d157517944169350516b8b01c2c5a67b8dc34e6f90054a8154301386d25848be9e64d72f215b5d6080c0654b4fe31a142054e9792a6b38a27dbaa024f12ccb8687a7222a7f0362bc0a3e81ee38bdbfb64767118be0967fe8e892;
    5'b11101 : xpb = 1024'h869f431c02290d3c49d4df0f96d9e9a0d088368f6afb6997d7db0af9ba0a88a9724e8eb66f3e17e3d64353c4f3e1f168597735a9cbe0a1df82c7a278e9d662362823204bbc34eb70464188d04c1ef12fe135c57afe7d630741f349c716e8462868ab20e49fded0da5e9517f76a23fe9226f9a57a959af392ed2ad31eca307bdc;
    5'b11110 : xpb = 1024'h483fb85d8c897e1583c87b80c1fcf9f16610b2d149d6b4c807d57e6f129ff37748dd7e8614bedfe1bbaf242c7115809ac3d280a7ce92e5b00680758e4e58fb8ac8703990801a3b36a2b9eda2a2019d6e691b417a566078a8e4e0d7283b036c040229be72c36e2180143fca0c79bbccbc7d2b33551b34428e825a4aa28b95a8bb;
    5'b11111 : xpb = 1024'h9e02d9f16e9eeeebdbc17f1ed200a41fb992f1328b1fff837cff1e46b355e451f6c6e55ba3fa7dfa11af493ee490fcd2e2dcba5d14529808a3948a3b2db94df68bd52d543ff8afcff325274f7e449acf100bd79ae438e4a87ce64895f1e91df9ba85c00e6fd7225c9ea7c2189539ae6d35cc12fa0cd918a1789c2264cfad59a;
    endcase
end

endmodule

module xpb_5_440
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1e55b72e7d399d1ecee6be4701d18ca1d93df595d78ba7c263a5a7050d4944b9038838d1f085d2b7303b5714e31f6c49719e23e7f36dd17c52db940f79a7435415aed90e2d18578ad482af94dce14350e97dbeb6ed07bb4e2bb902b702ce36a7a1edb629891714f7b6272e7866922b32b738edad835c86040fe2bf4b5ae0dab7;
    5'b00010 : xpb = 1024'h3cab6e5cfa733a3d9dcd7c8e03a31943b27beb2baf174f84c74b4e0a1a928972071071a3e10ba56e6076ae29c63ed892e33c47cfe6dba2f8a5b7281ef34e86a82b5db21c5a30af15a9055f29b9c286a1d2fb7d6dda0f769c5772056e059c6d4f43db6c53122e29ef6c4e5cf0cd2456656e71db5b06b90c081fc57e96b5c1b56e;
    5'b00011 : xpb = 1024'h5b01258b77acd75c6cb43ad50574a5e58bb9e0c186a2f7472af0f50f27dbce2b0a98aa75d191782590b2053ea95e44dc54da6bb7da497474f892bc2e6cf5c9fc410c8b2a874906a07d880ebe96a3c9f2bc793c24c71731ea832b0825086aa3f6e5c9227c9b453ee722758b6933b6819825aac9088a15920c2fa83de210a29025;
    5'b00100 : xpb = 1024'h7956dcb9f4e6747b3b9af91c0746328764f7d6575e2e9f098e969c14352512e40e20e347c2174adcc0ed5c538c7db125c6788f9fcdb745f14b6e503de69d0d5056bb6438b4615e2b520abe5373850d43a5f6fadbb41eed38aee40adc0b38da9e87b6d8a6245c53ded89cb9e19a48accadce3b6b60d7218103f8afd2d6b836adc;
    5'b00101 : xpb = 1024'h97ac93e87220119a0a81b7630917bf293e35cbed35ba46cbf23c4319426e579d11a91c19b29d1d93f128b3686f9d1d6f3816b387c125176d9e49e44d604450a46c6a3d46e179b5b6268d6de8506650948f74b992a126a886da9d0d930e07114629a48ecfad7368d68ec3e85a00dad7fd941ca46390ce9e144f6dbc78c6644593;
    5'b00110 : xpb = 1024'h55505c12d6b79f00e62fdd2fa8f0479a5fdbe5237ce4e16d80530c89cb4ef4e11e8d772d8fc71bc8205cb366f5e78ee459aaf8991e0189e408638fe9f191f470dc9e1a65f010ffbe8761ada946bcfb484ed7eb101a836c450c97e4f56aaa55b9c8ab2cf85c18540be2b2ff36f9cdd06fc7bb32ec3dfc6e818e100bf9862b9df;
    5'b00111 : xpb = 1024'h23aabcefaaa5170edd49bc19fc60911b7f3bb3e80f59f5d93baad7cda9fe340715711044c9824473b241224b527de537b738d371854dea1a9361cd0e18c0629b2378bab48c196786bcf8ca6f714d13056e6b3d67eeaff2127c8281065978dc033e7868f90ed89a3874525e6bd62f0839b3b4a0dc473c4cec28c3c00af3439496;
    5'b01000 : xpb = 1024'h4200741e27deb42dac307a60fe321dbd5879a97de6e59d9b9f507ed2b74778c018f94916ba08172ae27c7960359d518128d6f75978bbbb96e63d611d9267a5ef392793c2b931bf11917b7a044e2e565657e8fc1edbb7ad60a83b83bd5c4712aae0661f2297efaf302a798ce43cc1336c6aed8e89ca98d2f038a67f564e246f4d;
    5'b01001 : xpb = 1024'h60562b4ca518514c7b1738a80003aa5f31b79f13be71455e02f625d7c490bd791c8181e8aa8de9e212b7d07518bcbdca9a751b416c298d133918f52d0c0ee9434ed66cd0e64a169c65fe29992b0f99a74166bad5c8bf68aed3f486745f1549528253d54c2106c427e0a0bb5ca3535e9f22267c374df558f448893ea1a9054a04;
    5'b01010 : xpb = 1024'h7eabe27b2251ee6b49fdf6ef01d537010af594a995fced20669bccdcd1da02322009baba9b13bc9942f32789fbdc2a140c133f295f975e8f8bf4893c85b62c97648545df13626e273a80d92e07f0dcf82ae4798cb5c723fcffad892b61e37ffa24418b75aa1dd91f96c7e9d509e589d1d95f69e4d151def8586bfded03e624bb;
    5'b01011 : xpb = 1024'h9d0199a99f8b8b8a18e4b53603a6c3a2e4338a3f6d8894e2ca4173e1df2346eb2391f38c8b998f50732e7e9edefb965d7db163115305300bded01d4bff5d6feb7a341eed407ac5b20f0388c2e4d2204914623843a2cedf4b2b668be264b1b6a1c62f419f3334ee174cef184d7077b5049098579254ae64fc684ebd385ec6ff72;
    5'b01100 : xpb = 1024'haaa0b825ad6f3e01cc5fba5f51e08f34bfb7ca46f9c9c2db00a61913969de9c23d1aee5b1f8e379040b966cdebcf1dc8b355f1323c0313c810c71fd3e323e8e1b93c34cbe021ff7d0ec35b528d79f6909dafd6203506d88a192fc9ead554ab73915659f0b830a817c565fe6df39ba0df8f7665d87bf8dd031c2017f30c573be;
    5'b01101 : xpb = 1024'h28ffc2b0d81090feebacb9ecf6ef95952539723a472843f013b0089646b323552759e7b7a27eb6303446ed81c1dc5e25fcd382fb172e02b8d3e8060cb7d981e231429c5aeb1a7782a56ee54a05b8e2b9f358bc18f05828d6cd4bff55b023815edb031bc8949a1f79327d8e5f45cbe540b030540b0b1c13d441a4c0ca8ba64e75;
    5'b01110 : xpb = 1024'h475579df554a2e1dba937833f8c12236fe7767d01eb3ebb27755af9b53fc680e2ae22089930488e764824496a4fbca6f6e71a6e30a9bd43526c39a1c3180c53646f175691832cf0d79f194dee29a260adcd67acfdd5fe424f905020cb2f1b8067cf0d1f21db13470e8a4bcd7ac5e1073676941b88e7899d851878015e687292c;
    5'b01111 : xpb = 1024'h65ab310dd283cb3c897a367afa92aed8d7b55d65f63f9374dafb56a06145acc72e6a595b838a5b9e94bd9bab881b36b8e00fcacafe09a5b1799f2e2bab28088a5ca04e77454b26984e744473bf7b695bc6543986ca679f7324be04c3b5bfeeae1ede881ba6c849689ecbeb5012f03ba61ea22f6611d51fdc616a3f61416803e3;
    5'b10000 : xpb = 1024'h8400e83c4fbd685b5860f4c1fc643b7ab0f352fbcdcb3b373ea0fda56e8ef18031f2922d74102e55c4f8f2c06b3aa30251adeeb2f177772dcc7ac23b24cf4bde724f278572637e2322f6f4089c5cacacafd1f83db76f5ac15077077ab88e2555c0cc3e452fdf5e6054f319c8798266d8d5db1d139531a5e0714cfeac9c48de9a;
    5'b10001 : xpb = 1024'ha2569f6accf7057a2747b308fe35c81c8a314891a556e2f9a246a4aa7bd83639357acaff6496010cf53449d54e5a0f4bc34c129ae4e548aa1f56564a9e768f3287fe00939f7bd5adf779a39d793deffd994fb6f4a477160f7c300a31bb5c5bfd62b9f46eb8f673580b1a4840e014920b8d140ac1188e2be4812fbdf7f729b951;
    5'b10010 : xpb = 1024'hfff114388426dd02b28f978efad0d6cf1f93af6a76aea44880f9259d61ecdea35ba86588af55535861161a34e1b6acad0d00e9cb5a049dac192aafbdd4b5dd5295da4f31d032ff3b962508fbd436f1d8ec87c1304f8a44cf25c7aee03fff012d5a0186e91448fc23a818fda4ed69714f573198c4b9f54b84aa3023ec9282d9d;
    5'b10011 : xpb = 1024'h2e54c872057c0aeefa0fb7bff17e9a0ecb37308c7ef69206ebb5395ee36812a33942bf2a7b7b27ecb64cb8b8313ad714426e3284a90e1b57146e3f0b56f2a1293f0c7e014a1b877e8de500249a24b26e78463ac9f2005f9b1e157da506ce26ba778dce981a5ba4b9f0a8be52b568c247acac0739cefbdabc5a85c18a24090854;
    5'b10100 : xpb = 1024'h4caa7fa082b5a80dc8f67606f35026b0a4752622568239c94f5ae063f0b1575c3ccaf7fc6c00faa3e6880fcd145a435db40c566c9c7becd36749d31ad099e47d54bb570f7733df096267afb97705f5bf61c3f980df081ae949ce805c099c5d62197b84c1a372b9b1a6cfeccb1bfaed7a63e4f4e7525860c06a6880d57ee9e30b;
    5'b10101 : xpb = 1024'h6b0036ceffef452c97dd344df521b3527db31bb82e0de18bb3008768fdfa9c15405330ce5c86cd5b16c366e1f779afa725aa7a548fe9be4fba25672a4a4127d16a6a301da44c369436ea5f4e53e739104b41b837cc0fd637758783130c6a9409bb693aeb2c89cea95cf71b43828d18ad1b1de294d5b4e6c47a4b4020d9cabdc2;
    5'b10110 : xpb = 1024'h8955edfd7d28e24b66c3f294f6f33ff456f1114e0599894e16a62e6e0b43e0ce43db69a04d0ca01246febdf6da991bf097489e3c83578fcc0d00fb39c3e86b258019092bd1648e1f0b6d0ee330c87c6134bf76eeb9179185a14085ca0f38cab15d56f114b5a0e3a1131e49bbe91f43dfd256d04259116cc88a2dff6c34ab9879;
    5'b10111 : xpb = 1024'ha7aba52bfa627f6a35aab0dbf8c4cc96302f06e3dd2531107a4bd573188d25874763a2723d9272c9773a150bbdb8883a08e6c22476c561485fdc8f493d8fae7995c7e239fe7ce5a9dfefbe780da9bfb21e3d35a5a61f4cd3ccf9888112070158ff44a73e3eb7f898c94578344fb16f12898fbdefdc6df2cc9a10beb78f8c7330;
    5'b11000 : xpb = 1024'h15541704b5ade7c0398bf74bea3c11e697f6f948df39385b6014c32272d3bd3847a35dcb63f1c6f208172cd9bd79e3b9166abe26478062790218e3fa7c647d1c372786997c043fefa1d86b6a51af3ed213b5fac406a0db114325f93d5aaa956e722acb3e17061502f8acbfcdbe73741bf1eeccbb0f7f1ba0638402fe618ae77c;
    5'b11001 : xpb = 1024'h33a9ce3332e784df0872b592ec0d9e887134eedeb6c4e01dc3ba6a27801d01f14b2b969d547799a9385283eea09950028808e20e3aee33f554f47809f60bc0704cd65fa7a91c977a765b1aff2e908222fd33b97af3a8965f6edefbf45d78cc1614188167a01d29faaed3ee4625059f4ea927ba6892dba1a47366c249bc6bc233;
    5'b11010 : xpb = 1024'h51ff8561b02121fdd75973d9eddf2b2a4a72e4748e5087e02760112c8d6646aa4eb3cf6f44fd6c60688ddb0383b8bc4bf9a705f62e5c0571a7d00c196fb303c4628538b5d634ef054addca940b71c573e6b17831e0b051ad9a97feab604702bdb606379129343ef264fb1cbe8b97ca816060a816163827a883498195174c9cea;
    5'b11011 : xpb = 1024'h70553c902d5abf1ca6403220efb0b7cc23b0da0a65dc2fa28b05b8319aaf8b63523c084135833f1798c9321866d828956b4529de21c9d6edfaaba028e95a4718783411c4034d46901f607a28e85308c4d02f36e8cdb80cfbc65101626315396557f3edbab24b53ea1b224b36f229f5b4179995c39994adac932c40e0722d77a1;
    5'b11100 : xpb = 1024'h8eaaf3beaa945c3b7526f067f182446dfceecfa03d67d764eeab5f36a7f8d01c55c44113260911cec904892d49f794dedce34dc61537a86a4d87343863018a6c8de2ead230659e1af3e329bdc5344c15b9acf59fbabfc849f20a041965e3700cf9e1a3e43b6268e1d14979af58bc20e6ced283711cf133b0a30f002bcd0e5258;
    5'b11101 : xpb = 1024'had00aaed27cdf95a440daeaef353d10fd62cc53614f37f275251063bb54214d5594c79e5168ee485f93fe0422d1701284e8171ae08a579e6a062c847dca8cdc0a391c3e05d7df5a5c865d952a2158f66a32ab456a7c783981dc306d068b1a6b49bcf5a0dc4797dd98770a827bf4e4c19860b711ea04db9b4b2f1bf7727ef2d0f;
    5'b11110 : xpb = 1024'h1aa91cc5e31961b047eef51ee4cb16603df4b79b170786723819f3eb0f88ac86598c353e3cee38ae8a1cf8102cd85ca75c056dafd9607b17429f1cf91b7d9c6344f1683fdb054feb8a4e8644e61b0e8698a37975084911d593ef778cb1553aca0eb57e0d9cc79a43b6d7efc12e105122ee6a7fe9d35ee2887c6503bdf9eda15b;
    5'b11111 : xpb = 1024'h38fed3f46052fecf16d5b365e69ca3021732ad30ee932e349bbf9af01cd1f13f5d146e102d740b65ba584f250ff7c8f0cda39197ccce4c93957ab1089524dfb75aa0414e081da7765ed135d9c2fc51d78221382bf550cd23bfa87a43b4237171b0a3343725deaf3b6cff1e3994a27c55a5a36d9756bb688c8c47c30954ce7c12;
    endcase
end

endmodule

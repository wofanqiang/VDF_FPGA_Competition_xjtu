module xpb_5_340
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9811fdd24de17adbd3b805de8716fb1f5cd03829fcd35963651b8213194c24981c8060bf473f97d0656695b1adebec717132e6f63da42b90dde9208bba625d0bd13aea29cf3b235311b7a8d02d2b69450922bda425e1b9519fa8f4c8f332c982161101553a2b4717c7aadc7d58a52ea10b84a656217aab31f4b3c83e06216dea;
    5'b00010 : xpb = 1024'h7f76b64ed9d4c0eedc6a93e5fdd3aeed482a6d23242f124f4c5a4ad07f959c2835b84405c458b1122b6eec1c7879c8187e4ba606589586d60b3301b939f245662e269fa4eee5496110d54efdc17b0e591e4081afbf3d459289c557972c3af071fd1a7080c38d95a20895d21bb97a3718c82f6dc9f2a9f933a2f8157783607569;
    5'b00011 : xpb = 1024'h66db6ecb65c80701e51d21ed749062bb3384a21c4b8acb3b3399138de5df13b84ef0274c4171ca53f17742874307a3bf8b6465167386e21b387ce2e6b9822dc08b1255200e8f6f6f0ff2f52b55cab36d335e45bb5898d1d373e1ba6565431761e423dfac4cefe42c4980c7ba1a4f3f9084da353dc3d94735513c62b1009f7ce8;
    5'b00100 : xpb = 1024'h4e402747f1bb4d14edcfaff4eb4d16891eded71572e684271ad7dc4b4c288b4868280a92be8ae395b77f98f20d957f66987d24268e783d6065c6c4143912161ae7fe0a9b2e39957d0f109b58ea1a5881487c09c6f1f45e145dfe1d339e4b3e51cb2d4ed7d65232b68a6bbd587b2448084184fcb195089536ff80afea7dde8467;
    5'b00101 : xpb = 1024'h35a4dfc47dae9327f6823dfc6209ca570a390c0e9a423d130216a508b27202d8815fedd93ba3fcd77d87ef5cd8235b0da595e336a96998a59310a541b8a1fe7544e9c0164de3bb8b0e2e41867e69fd955d99cdd28b4fea55481a8001d7536541b236be035fb48140cb56b2f6dbf9507ffe2fc4256637e338adc4fd23fb1d8be6;
    5'b00110 : xpb = 1024'h1d09984109a1d93aff34cc03d8c67e24f5934107c19df5fee9556dc618bb7a689a97d11fb8bd1619439045c7a2b136b4b2aea246c45af3eac05a866f3831e6cfa1d575916d8de1990d4be7b412b9a2a972b791de24ab76963236e2d0105b8c3199402d2ee916cfcb0c41a8953cce58f7bada8b993767313a5c094a5d785c9365;
    5'b00111 : xpb = 1024'h46e50bd95951f4e07e75a0b4f8331f2e0ed7600e8f9aeead09436837f04f1f8b3cfb46635d62f5b09989c326d3f125bbfc76156df4c4f2feda4679cb7c1cf29fec12b0c8d3807a70c698de1a70947bd87d555e9be0702d71c53459e4963b32180499c5a72791e554d2c9e339da3616f7785530d08967f3c0a4d9796f59b9ae4;
    5'b01000 : xpb = 1024'h9c804e8fe3769a29db9f5fe9d69a2d123dbdae2ae5cd084e35afb89698511690d05015257d15c72b6eff31e41b2afecd30fa484d1cf07ac0cb8d882872242c35cffc15365c732afa1e2136b1d434b10290f8138de3e8bc28bbfc3a673c967ca3965a9dafaca4656d14d77ab0f64890108309f9632a112a6dff015fd4fbbd08ce;
    5'b01001 : xpb = 1024'h83e5070c6f69e03ce451edf14d56e0e02917e3240d28c13a1cee8153fe9a8e20e987f86bfa2ee06d3507884ee5b8da743e13075d37e1d605f8d76955f1b414902ce7cab17c1d51081d3edcdf68845616a615d7997d444869a6189d35759ea3937d640cdb3606b3f755c2704f571d98883fb4c0d6fb40786fad45ad0e78fc104d;
    5'b01010 : xpb = 1024'h6b49bf88fb5d264fed047bf8c41394ae1472181d34847a26042d4a1164e405b102bfdbb27747f9aefb0fdeb9b046b61b4b2bc66d52d3314b26214a837143fcea89d3802c9bc777161c5c830cfcd3fb2abb339ba5169fd4aa90350003aea6ca83646d7c06bf69028196ad65edb7f2a0fffc5f884acc6fc6715b89fa47f63b17cc;
    5'b01011 : xpb = 1024'h52ae780587506c62f5b70a003ad0487bffcc4d165be03311eb6c12cecb2d7d411bf7bef8f46112f0c11835247ad491c25844857d6dc48c90536b2bb0f0d3e544e6bf35a7bb719d241b7a293a9123a03ed0515fb0affb60eb7a5162d1e7aef1734b76eb3248cb510bd7985b8c18c7a977b90a4fbe9d9f147309ce4781737a1f4b;
    5'b01100 : xpb = 1024'h3a1330821343b275fe699807b18cfc49eb26820f833bebfdd2aadb8c3176f4d1352fa23f717a2c3287208b8f45626d69655d448d88b5e7d580b50cde7063cd9f43aaeb22db1bc3321a97cf6825734552e56f23bc4956ed2c646dc5a020b7186332805a5dd22d9f961883512a799cb1ef75b517326ece6274b81294baf0b926ca;
    5'b01101 : xpb = 1024'h2177e8fe9f36f889071c260f2849b017d680b708aa97a4e9b9e9a44997c06c614e678585ee9345744d28e1fa0ff049107276039da3a7431aadfeee0beff3b5f9a096a09dfac5e94019b57595b9c2ea66fa8ce7c7e2b2796d4e8a286e59bf3f531989c9895b8fee20596e46c8da71ba67325fdea63ffdb0766656e1f46df82e49;
    5'b01110 : xpb = 1024'h8dca17b2b2a3e9c0fceb4169f0663e5c1daec01d1f35dd5a1286d06fe09e3f1679f68cc6bac5eb613313864da7e24b77f8ec2adbe989e5fdb48cf396f839e53fd8256191a700f4e18d31bc34e128f7b0faaabd37c0e05ae38a68b3c92c76643009338b4e4f23caa9a593c673b46c2deef0aa61a112cfe78149b2f2deb3735c8;
    5'b01111 : xpb = 1024'ha0ee9f4d790bb977e386b9f5261d5f051eab242bcec6b7390643ef1a17560889841fc98bb2ebf6867897ce16886a1128f0c1a9a3fc3cc9f0b931efc529e5fb5fcebd4042e9ab32a12a8ac4937b3df8c018cd6977a1efbeffd84f800585fa2fc516a43a0a1f1d83c2620418e493ebf17ffa8f4c7032a7a9aa094ef76bf158a3b2;
    5'b10000 : xpb = 1024'h885357ca04feff8aec3947fc9cda12d30a055924f6227024ed82b7d77d9f80199d57acd230050fc83ea0248152f7eccffdda68b4172e2535e67bd0f2a975e3ba2ba8f5be095558af29a86ac10f8d9dd42deb2d833b4b4b40c26be2d3bf0256b4fdada935a87fd24ca2ef0e82f4c0f9f7b73a13e403d6f7abb79344a56e97ab31;
    5'b10001 : xpb = 1024'h6fb8104690f2459df4ebd6041396c6a0f55f8e1e1d7e2910d4c18094e3e8f7a9b68f9018ad1e290a04a87aec1d85c8770af327c4321f807b13c5b2202905cc148894ab3928ff7ebd28c610eea3dd42e84308f18ed4a6d781ac8845a1f80a7da4e4b7186131e220d6e3da04215596026f73e4db57d50645ad65d791deebd6b2b0;
    5'b10010 : xpb = 1024'h571cc8c31ce58bb0fd9e640b8a537a6ee0b9c31744d9e1fcbc0049524a326f39cfc7735f2a37424bcab0d156e813a41e180be6d44d10dbc0410f934da895b46ee58060b448a9a4cb27e3b71c382ce7fc5826b59a6e0263c296a4a8703112a494cbc0878cbb446f6124c4f9bfb66b0ae7308fa2cba63593af141bdf186915ba2f;
    5'b10011 : xpb = 1024'h3e81813fa8d8d1c40650f21301102e3ccc13f8106c359ae8a33f120fb07be6c9e8ff56a5a7505b8d90b927c1b2a17fc52524a5e4680237056e59747b28259cc9426c162f6853cad927015d49cc7c8d106d4479a6075df00380c10b3e6a1acb84b2c9f6b844a6bdeb65afef5e1740135eed3a6a3f7764e1b0c2602c51e654c1ae;
    5'b10100 : xpb = 1024'h25e639bc34cc17d70f03801a77cce20ab76e2d09939153d48a7ddacd16c55e5a023739ec246974cf56c17e2c7d2f5b6c323d64f482f3924a9ba355a8a7b585239f57cbaa87fdf0e7261f037760cc322482623db1a0b97c446add6e0ca322f27499d365e3ce090c75a69ae4fc78151bd6a9e531b348942fb270a4798b6393c92d;
    5'b10101 : xpb = 1024'hd4af238c0bf5dea17b60e21ee8995d8a2c86202baed0cc071bca38a7d0ed5ea1b6f1d32a1828e111cc9d49747bd37133f5624049de4ed8fc8ed36d627456d7dfc438125a7a816f5253ca9a4f51bd738978001bd3a15088554f9d0dadc2b196480dcd50f576b5affe785da9ad8ea244e668ff92719c37db41ee8c6c4e0d2d0ac;
    5'b10110 : xpb = 1024'ha55cf00b0ea0d8c5eb6e140075a090f7ff989a2cb7c06623d6d8259d965afa8237ef7df1e8c225e182306a48f5a92384b0890afadb891920a6d65761e1a7ca89cd7e6b4f76e33a4836f452752247407da0a2bf615ff6c1d6f4a2c5a3cf5de2e696edd6649196a217af30b718318f52ef72149f7d3b3e28e6139c8f02e6f43e96;
    5'b10111 : xpb = 1024'h8cc1a8879a941ed8f420a207ec5d44c5eaf2cf25df1c1f0fbe16ee5afca472125127613865db3f234838c0b3c036ff2bbda1ca0af67a7465d420388f6137b2e42a6a20ca968d60563611f8a2b696e591b5c0836cf9524e17debf2872086609d67df745901af8f0a1f01bacb692645b672ebf66f10c6d76e7c1e0dc3c64334615;
    5'b11000 : xpb = 1024'h74266104268764ebfcd3300f6319f893d64d041f0677d7fba555b71862ede9a26a5f447ee2f458650e41171e8ac4dad2caba891b116bcfab016a19bce0c79b3e8755d645b6378664352f9ed04ae68aa5cade477892adda58c8db8b40416e30c66500b4bba45b3f2c3106a254f33963deeb6a2e64dd9cc4e970252975e1724d94;
    5'b11001 : xpb = 1024'h5b8b1980b27aaaff0585be16d9d6ac61c1a739182dd390e78c947fd5c9376132839727c5600d71a6d4496d895552b679d7d3482b2c5d2af02eb3faea60578398e4418bc0d5e1ac72344d44fddf362fb9dffc0b842c096699b2f7ee0e7a7657b64c0a23e72dbd8db671f197f3540e6c56a814f5d8aecc12eb1e6976af5eb15513;
    5'b11010 : xpb = 1024'h42efd1fd3e6df1120e384c1e5093602fad016e11552f49d373d348932f80d8c29ccf0b0bdd268ae89a51c3f41fe09220e4ec073b474e86355bfddc17dfe76bf3412d413bf58bd280336aeb2b7385d4cdf519cf8fc564f2da9d1450dcb37e7ea633139312b71fdc40b2dc8d91b4e374ce64bfbd4c7ffb60ecccadc3e8dbf05c92;
    5'b11011 : xpb = 1024'h2a548a79ca61372516eada25c75013fd985ba30a7c8b02bf5b12115095ca5052b606ee525a3fa42a605a1a5eea6e6dc7f204c64b623fe17a8947bd455f77544d9e18f6b71535f88e3288915907d579e20a37939b5ec07f1b8730b3aaec86a5961a1d023e40822acaf3c7833015b87d46216a84c0512aaeee7af21122592f6411;
    5'b11100 : xpb = 1024'h11b942f656547d381f9d682d3e0cc7cb83b5d803a3e6bbab4250da0dfc13c7e2cf3ed198d758bd6c266270c9b4fc496eff1d855b7d313cbfb6919e72df073ca7fb04ac3234e01e9c31a637869c251ef61f5557a6f81c0b5c714d1679258ecc8601267169c9e4795534b278ce768d85bdde154c342259fcf029365e5bd66e6b90;
    5'b11101 : xpb = 1024'ha9cb40c8a435f813f3556e0bc523c2eae086102da0ba150ea76c5c21155fec7aebbf32581e98553c8bc9067b62e835e070506c51bad56850947abefe996999b3cc3f965c041b41ef435de056c950883b2878154b1dfdc4ae10f60b4218c19608173772bf040fc06cfc5d554bcf32b45ee999f28a43d4a8221dea2699dc8fd97a;
    5'b11110 : xpb = 1024'h912ff94530293e26fc07fc133be076b8cbe04526c815cdfa8eab24de7ba9640b04f7159e9bb16e7e51d15ce62d7611877d692b61d5c6c395c1c4a02c18f9820e292b4bd723c567fd427b86845da02d4f3d95d956b75950eefb126e1051c9bcf7fe40e1ea8d720ef73d484aea3007bcd6a644b9fe1503f623cc2e73d359cee0f9;
    5'b11111 : xpb = 1024'h7894b1c1bc1c843a04ba8a1ab29d2a86b73a7a1fef7186e675e9ed9be1f2db9b1e2ef8e518ca87c017d9b350f803ed2e8a81ea71f0b81edaef0e815998896a6886170152436f8e0b41992cb1f1efd26352b39d6250b4dd2fe52ed0de8ad1e3e7e54a511616d45d817e33408890dcc54e62ef8171e63344257a72c10cd70de878;
    endcase
end

endmodule

module xpb_5_965
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7c2de83663389490c2b52c3a289d61e40297ae85dd04eb9fe5a71eaf76cd761af943db9e29e6ee6c25e504424edaafc9fca33e89f6aa3d9cbe915b175230a2e57d59a0c8b775d8086e44b9e9e6a2ba1c6ceb331192acd0fce04883e53d645a4d642e8bb8bb55bb590655151590bb8f3a78682dec76b23db5f328b4ae974268e4;
    5'b00010 : xpb = 1024'h47ae8b170482f458ba64e09d40e07c7693b959dae49236c84d7184093a983f2def3f39c389a75e49ac6bc93dba574ec9952c552dcaa1aaedcc8376d0698ed11986640ce2bf5ab2cbc9ef71313469b007e5d16c8a98d374e90b0475cfc09e120899558547c5e27e2485ea434c29a6f84ba1f67cf69d191e3b9fe1ee58a5a26b5d;
    5'b00011 : xpb = 1024'h132f2df7a5cd5420b21495005923970924db052fec1f81f0b53be962fe630840e53a97e8e967ce2732f28e3925d3edc92db56bd19e99183eda75928980ecff4d8f6e78fcc73f8d8f259a28788230a5f35eb7a6039efa18d535c067ba43d7c9c3ce7c7ed6d06f40f0057f7182c292615ccb84cc00c37ffec14c9b2802b4026dd6;
    5'b00100 : xpb = 1024'h8f5d162e0905e8b174c9c13a81c0f8ed2772b3b5c9246d909ae3081275307e5bde7e7387134ebc9358d7927b74ae9d932a58aa5b954355db9906eda0d31da2330cc819c57eb5659793dee26268d3600fcba2d91531a6e9d21608eb9f813c241132ab0a8f8bc4fc490bd48698534df09743ecf9ed3a323c773fc3dcb14b44d6ba;
    5'b00101 : xpb = 1024'h5addb90eaa5048796c79759d9a04137fb8945f0ad0b1b8b902ad6d6c38fb476ed479d1ac730f2c70df5e5776e02b3c92c2e1c0ff693ac32ca6f90959ea7bd06715d285df869a405aef8999a9b69a55fb4489128e37cd8dbe40c4dd8a0475dbcc67d2041e9651bf148b69b4ceec3959a86d7b48f760991cfcec7d165b59a4d933;
    5'b00110 : xpb = 1024'h265e5bef4b9aa84164292a00b2472e1249b60a5fd83f03e16a77d2c5fcc61081ca752fd1d2cf9c4e65e51c724ba7db925b6ad7a33d32307db4eb251301d9fe9b1edcf1f98e7f1b1e4b3450f104614be6bd6f4c073df431aa6b80cf7487af93879cf8fdada0de81e00afee3058524c2b99709980186fffd82993650056804dbac;
    5'b00111 : xpb = 1024'ha28c4425aed33cd226de563adae48ff64c4db8e5b543ef81501ef1757393869cc3b90b6ffcb68aba8bca20b49a828b5c580e162d33dc6e1a737c802a540aa1809c3692c245f4f326b9790adaeb0406032a5a7f18d0a102a74bc95359c513edd5012789665c343d391153f81b15e051f40f71c5edfdb23b388c5f04b3ff474490;
    5'b01000 : xpb = 1024'h6e0ce706501d9c9a1e8e0a9df327aa88dd6f643abcd13aa9b7e956cf375e4fafb9b469955c76fa981250e5b005ff2a5bf0972cd107d3db6b816e9be36b68cfb4a540fedc4dd9cdea1523c22238cafbeea340b891d6c7a69376854544484da590364e82f566c1000490e92651aecbbb05390014f824191bbe39183e5e0da74709;
    5'b01001 : xpb = 1024'h398d89e6f167fc62163dbf010b6ac51b6e910f8fc45e85d21fb3bc28fb2918c2afafc7babc376a7598d7aaab717bc95b89204374dbcb48bc8f60b79c82c6fde8ae4b6af655bea8ad70ce79698691f1da1c26f20adcee4a7fa141372ecb875d4b6b757c84714dc2d0107e548847b72416628e64024a7ffc43e5d178081c074982;
    5'b01010 : xpb = 1024'h50e2cc792b25c2a0ded736423addfadffb2bae4cbebd0fa877e2182bef3e1d5a5ab25e01bf7da531f5e6fa6dcf8685b21a95a18afc2b60d9d52d3559a252c1cb755d7105da38370cc7930b0d458e7c5950d2b83e314ee6bcbfd29194ec11506a09c76137bda859b901382bee0a28d278c1cb30c70e6dcc9928ab1b22a674bfb;
    5'b01011 : xpb = 1024'h813c14fdf5eaf0bad0a29f9e4c4b4192024a696aa8f0bc9a6d25403235c157f09eef017e45dec8bf454373e92bd318251e4c98a2a66cf3aa5be42e6cec55cf0234af77d915195b793abdea9abafba1e201f85e9575c1bf68ac45acfe8c256f5404cb01cc373040f4966897d4715e1c620484e0f8e7991a7f85b36660c1a9b4df;
    5'b01100 : xpb = 1024'h4cbcb7de97355082c8525401648e5c24936c14bfb07e07c2d4efa58bf98c210394ea5fa3a59f389ccbca38e4974fb724b6d5af467a6460fb69d64a2603b3fd363db9e3f31cfe363c9668a1e208c297cd7ade980e7be86354d7019ee90f5f270f39f1fb5b41bd03c015fdc60b0a4985732e1330030dfffb05326ca00ad009b758;
    5'b01101 : xpb = 1024'h183d5abf387fb04ac00208647cd176b7248dc014b80b52eb3cba0ae5bd56ea168ae5bdc9055fa87a5250fde002cc56244f5ec5ea4e5bce4c77c865df1b122b6a46c4500d24e310fff213592956898db8f3c4d187820f074101bd90d39298deca6f18f4ea4c49c68b9592f441a334ee8457a17f0d3466db8adf25d9b4de69b9d1;
    5'b01110 : xpb = 1024'h946b42f59bb844db82b7349ea56ed89b27256e9a95103e8b2261299534246031842999672f4696e67836022251a705ee4c02047445060be93659c0f66d42ce4fc41df0d5dc58e908605813133d2c47d560b0049914bbd83de20614b8cffd3917d34780a3079f81e49be8095733f07dbed009acf9ab191940d24e8e6375ac22b5;
    5'b01111 : xpb = 1024'h5febe5d63d02a4a37a66e901bdb1f32db84719ef9c9d89b38a2b8eeef7ef29447a24f78c8f0706c3febcc71dbd23a4ede48b1b1818fd793a444bdcaf84a0fc83cd285cefe43dc3cbbc02ca5a8af33dc0d9963e121ae27c2a0cc206a35336f0d3086e7a32122c44b01b7d378dccdbe6cff997fc03d17ff9c67f07c80d840c252e;
    5'b10000 : xpb = 1024'h2b6c88b6de4d046b72169d64d5f50dc04968c544a42ad4dbf1f5f448bbb9f257702055b1eec776a185438c1928a043ed7d1431bbecf4e68b523df8689bff2ab7d632c909ec229e8f17ad81a1d8ba33ac527c778b21092016377df88dd670a88e3d9573c11cb9077b9b1265c465c74fe123264b0df7e6da4c2bc101b7926c27a7;
    5'b10001 : xpb = 1024'ha79a70ed418598fc34cbc99efe926fa44c0073ca812fc07bd79d12f8328768726964315018ae650dab28905b777af3b779b77045e39f242810cf537fee2fcd9d538c69d2a398769785f23b8bbf5cedc8bf67aa9cb3b5f11317c67c7313d502dba1c3ff79d80ec2d4a1677ad9f682df1b9b8e78fa6e9918021ee9b66629ae908b;
    5'b10010 : xpb = 1024'h731b13cde2cff8c42c7b7e0216d58a36dd221f1f88bd0ba43f677851f65231855f5f8f75786ed4eb31af5556e2f792b7124086e9b79691791ec16f39058dfbd15c96d5ecab7d515ae19cf2d30d23e3b4384de415b9dc94ff42826e5d970eba96d6eaf908e29b85a020fca9108f6e482cc51cc80494fff887cba2f010380e9304;
    5'b10011 : xpb = 1024'h3e9bb6ae841a588c242b32652f18a4c96e43ca74904a56cca731ddabba1cfa98555aed9ad82f44c8b8361a524e7431b6aac99d8d8b8dfeca2cb38af21cec2a0565a14206b3622c1e3d47aa1a5aead99fb1341d8ec00338eb6d3e60481a4872520c11f297ed28486ba091d7472859b13deeab170ebb66d90d785c29ba466e957d;
    5'b10100 : xpb = 1024'ha1c598f2564b8541bdae6c8475bbf5bff6575c997d7a1f50efc43057de7c3ab4b564bc037efb4a63ebcdf4db9f0d0b64352b4315f856c1b3aa5a6ab344a58396eabae20bb4706e198f26161a8b1cf8b2a1a5707c629dcd797fa52329d822a0d4138ec26f7b50b372027057dc1451a4f18396618e1cdb9932515636454ce97f6;
    5'b10101 : xpb = 1024'h864a41c5889d4ce4de9013026ff9214001fd244f74dc8d94f4a361b4f4b539c6449a275e61d6a31264a1e39008cb80803ff5f2bb562fa9b7f93701c2867afb1eec054ee972bcdeea07371b4b8f5489a797058a1958d6add47842d617dae6845aa56777dfb30ac690267c1a935200a98990a19405587ff749183e1812ec1100da;
    5'b10110 : xpb = 1024'h51cae4a629e7acacd63fc765883c3bd2931ecfa47c69d8bd5c6dc70eb88002d93a958583c19712efeb28a88b74481f7fd87f095f2a27170907291d7b9dd92952f50fbb037aa1b9ad62e1d292dd1b7f930febc3925efd51c0a2fec8025e203c15da8e716ebd97895ba61148c9eaec129aba2fe30f7ee6d7cec4f751bcfa710353;
    5'b10111 : xpb = 1024'h1d4b8786cb320c74cdef7bc8a07f566524407af983f723e5c4382c687c4acbec3090e3a9215782cd71af6d86dfc4be7f71082002fe1e845a151b3934b5375786fe1a271d82869470be8c89da2ae2757e88d1fd0b6523f5accdbab9ece159f3d10fb56afdc8244c2725a6770083d77babe3be3219a54db85471b08b6708d105cc;
    5'b11000 : xpb = 1024'h99796fbd2e6aa10590a4a802c91cb84926d8297f60fc0f85a9df4b17f318420729d4bf474b3e7139979471c92e9f6e496dab5e8cf4c8c1f6d3ac944c0767fa6c7b73c7e639fc6c792cd143c411852f9af5bd301cf7d0c6a9ae033dd21ebe4e1e73e3f6b6837a07802bfb8c1614930ae65c2660061bfff60a64d94015a0136eb0;
    5'b11001 : xpb = 1024'h64fa129dcfb500cd88545c65e15fd2dbb7f9d4d468895aae11a9b071b6e30b1a1fd01d6caafee1171e1b36c49a1c0d4906347530c8c02f47e19eb0051ec628a0847e340041e1473c887bfb0b5f4c25866ea36995fdf76a95d8bf2fbca1f805d9a90af0458e06ca4bab90ba4cad7e73f785b4af104266d690119279bfae737129;
    5'b11010 : xpb = 1024'h307ab57e70ff6095800410c8f9a2ed6e491b80297016a5d6797415cb7aadd42d15cb7b920abf50f4a4a1fbc00598ac489ebd8bd49cb79c98ef90cbbe362456d48d88a01a49c621ffe426b252ad131b71e789a30f041e0e82037b21a72531bd94de31e9d498938d172b25e8834669dd08af42fe1a68cdb715be4bb369bcd373a2;
    5'b11011 : xpb = 1024'haca89db4d437f52642b93d0322404f524bb32eaf4d1b91765f1b347af17b4a480f0f573034a63f60ca87000254735c129b60ca5e9361da35ae2226d58854f9ba0ae240e3013bfa08526b6c3c93b5d58e5474d62096cadf7ee3c3a58c629617e24260758d53e94870317afd98d7256c4327ab2c06df7ff4cbb17468185415dc86;
    5'b11100 : xpb = 1024'h78294095758254ee3a68f1663a8369e4dcd4da0454a8dc9ec6e599d4b546135b050ab5559466af3e510dc4fdbfeffb1233e9e10267594786bc14428e9fb327ee13ecacfd0920d4cbae162383e17ccb79cd5b0f999cf1836b0e7f9776e5cfcf9d77876f1c5e760b3bb1102bcf7010d55451397b1105e6d5515e2da1c26275deff;
    5'b11101 : xpb = 1024'h43a9e37616ccb4b63218a5c952c684776df685595c3627c72eafff2e7910dc6dfb06137af4271f1bd79489f92b6c9a11cc72f7a63b50b4d7ca065e47b71156221cf719171105af8f09c0dacb2f43c16546414912a3182757393b896169098758acae68ab6902ce0730a55a0608fc3e657ac7ca1b2c4db5d70ae6db6c70d5e178;
    5'b11110 : xpb = 1024'hf2a8656b817147e29c85a2c6b099f09ff1830ae63c372ef967a64883cdba580f10171a053e78ef95e1b4ef496e9391164fc0e4a0f482228d7f87a00ce6f84562601853118ea8a52656b92127d0ab750bf27828ba93ecb4363f77b4bec433f13e1d5623a738f90d2b03a883ca1e7a776a456192552b4965cb7a015167f35e3f1;
    5'b11111 : xpb = 1024'h8b586e8d1b4fa90eec7d866693a700ee01afdf3440c85e8f7c218337b3a91b9bea454d3e7dce7d6584005336e5c3e8db619f4cd405f25fc59689d51820a0273ba35b25f9d060625ad3b04bfc63ad716d2c12b59d3beb9c40443fff3129a799614603edf32ee54c2bb68f9d5232a336b11cbe4711c966d412aac8c9c516784cd5;
    endcase
end

endmodule

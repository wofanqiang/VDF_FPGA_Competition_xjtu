module xpb_5_320
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1774601716f27865b61a6470e028868c6c680a90337f47ed867e7f37cbbb76e5743a15b92ab101edc03ee1309e5ae80d1f024c7a646f5d0f6908e7e0004b8b3633139f5ff5cef6450941fd6048a4228d9ebf48252754f3d2651105dd265aa76560e0ac8d432e779abd328efcac117a553b82eec619626d540af2dcb1da005f8f;
    5'b00010 : xpb = 1024'h2ee8c02e2de4f0cb6c34c8e1c0510d18d8d0152066fe8fdb0cfcfe6f9776edcae8742b72556203db807dc2613cb5d01a3e0498f4c8deba1ed211cfc00097166c66273ebfeb9dec8a1283fac09148451b3d7e904a4ea9e7a4ca220bba4cb54ecac1c1591a865cef357a651df95822f4aa7705dd8c32c4daa815e5b963b400bf1e;
    5'b00011 : xpb = 1024'h465d204544d76931224f2d52a07993a545381fb09a7dd7c8937b7da7633264b05cae412b801305c940bca391db10b8275d06e56f2d4e172e3b1ab7a000e2a1a2993ade1fe16ce2cf1bc5f820d9ec67a8dc3dd86f75fedb772f331197730ff63022a205a7c98b66d03797acf604346effb288cc524c2747fc20d896158e011ead;
    5'b00100 : xpb = 1024'h5dd1805c5bc9e196d86991c380a21a31b1a02a40cdfd1fb619f9fcdf2eeddb95d0e856e4aac407b700fb84c2796ba0347c0931e991bd743da4239f80012e2cd8cc4e7d7fd73bd9142507f58122908a367afd20949d53cf4994441774996a9d958382b2350cb9de6af4ca3bf2b045e954ee0bbb186589b5502bcb72c768017e3c;
    5'b00101 : xpb = 1024'h7545e07372bc59fc8e83f63460caa0be1e0834d1017c67a3a0787c16faa9527b45226c9dd57509a4c13a65f317c688419b0b7e63f62cd14d0d2c87600179b80eff621cdfcd0acf592e49f2e16b34acc419bc68b9c4a8c31bf9551d51bfc544fae4635ec24fe85605b1fccaef5c5763aa298ea9de7eec22a436be4f794201ddcb;
    5'b00110 : xpb = 1024'h8cba408a89aed262449e5aa540f3274a8a703f6134fbaf9126f6fb4ec664c960b95c825700260b9281794723b621704eba0dcade5a9c2e5c76356f4001c543453275bc3fc2d9c59e378bf041b3d8cf51b87bb0deebfdb6ee5e66232ee61fec6045440b4f9316cda06f2f59ec0868ddff651198a4984e8ff841b12c2b1c023d5a;
    5'b00111 : xpb = 1024'ha42ea0a1a0a14ac7fab8bf16211badd6f6d849f1687af77ead757a86922040462d9698102ad70d8041b82854547c585bd9101758bf0b8b6bdf3e57200210ce7b65895b9fb8a8bbe340cdeda1fc7cf1df573af9041352aac0c377290c0c7a93c5a624b7dcd645453b2c61e8e8b47a5854a094876ab1b0fd4c4ca408dcf6029ce9;
    5'b01000 : xpb = 1024'haf5bb62f5a58e64e5cdabaff0e9ed11f1ca5150c6829ef4b6174068aad90a239e8830508b6190df6298ca3e0f792f9e93f83bed00c8182f97a7ffa1c789e500244dc650fee6b4e33775e85fac45503c01f54790ae21718272fb9cee78aa9898d7fdd24068aac44862d4910668bbac808d3d974e7ac80d7011276a8a4720960d;
    5'b01001 : xpb = 1024'h226a1b7a0c9806ca9be81020d112739e5e325be0fa01e6e23c95bfa07694810912c24609b61292cd22d7ab6eadd417abb2fa88676537753f00b0e781c7d57036576165b0f4b5ab2840b7e5bff4e972c9a0b48fb5d5766554d80ca2cb9f053ffe38de7ecdabd93be32007200314cd26d5c8c08614942a7ac41c1a473c2120f59c;
    5'b01010 : xpb = 1024'h39de7b91238a7f3052027491b13afa2aca9a66712d812ecfc3143ed8424ff7ee86fc5bc2e0c394bae3168c9f4c2effb8d1fcd4e1c9a6d24e69b9cf61c820fb6c8a750510ea84a16d49f9e3203d8d95573f73d7dafccb59273d1da8a8c55fe76399bf2b5aef07b37ddd39aeffc0dea12b044374daad8ce818270d23edfb21552b;
    5'b01011 : xpb = 1024'h5152dba83a7cf796081cd902916380b737027101610076bd4992be100e0b6ed3fb36717c0b7496a8a3556dcfea89e7c5f0ff215c2e162f5dd2c2b741c86c86a2bd88a470e05397b2533be0808631b7e4de33200024204cf9a22eae85ebba8ec8fa9fd7e832362b189a6c3dfc6cf01b803fc663a0c6ef556c3200009fd521b4ba;
    5'b01100 : xpb = 1024'h68c73bbf516f6ffbbe373d73718c0743a36a7b91947fbeaad0113d47d9c6e5b96f7087353625989663944f0088e4cfd310016dd692858c6d3bcb9f21c8b811d8f09c43d0d6228df75c7ddde0ced5da727cf268254b7540cc073fb4631215362e5b8084757564a2b3579eccf9190195d57b495266e051c2c03cf2dd51af221449;
    5'b01101 : xpb = 1024'h803b9bd66861e8617451a1e451b48dd00fd28621c7ff0698568fbc7fa5825c9ee3aa9cee60d69a8423d33031273fb7e02f03ba50f6f4e97ca4d48701c9039d0f23afe330cbf1843c65bfdb411779fd001bb1b04a72ca349e6c50ba40386fdd93bc613102b8931a4e14d15bf5c513102ab6cc412cf9b4301447e5ba03892273d8;
    5'b01110 : xpb = 1024'h97affbed7f5460c72a6c065531dd145c7c3a90b1fb7e4e85dd0e3bb7713dd38457e4b2a78b879c71e4121161c59a9fed4e0606cb5b64468c0ddd6ee1c94f284556c38290c1c07a816f01d8a1601e1f8dba70f86f9a1f2870d161c01d5eca84f91d41dd8ffbc191e8d203eaf271248a7ff24f2ff313169d6852d896b56322d367;
    5'b01111 : xpb = 1024'haf245c049646d92ce0866ac612059ae8e8a29b422efd9673638cbaef3cf94a69cc1ec860b6389e5fa450f29263f587fa6d085345bfd3a39b76e656c1c99ab37b89d721f0b78f70c67843d601a8c2421b59304094c1741c433672c5fa85252c5e7e228a1d3ef009838f3679ef1d3604d52dd21eb92c790abc5dcb73673d2332f6;
    5'b10000 : xpb = 1024'h15eb76c5eb4b1cc9cb9b575fe1d3da23e394a2a18d053de96c2e80d155b214473d1060a116c321bec531947c1ef25f3d27f077da0190305f2f4fff438f13ca00489b8ca1fdcd69c66eebd0bf588aa07803ea8f215c42e304e5f739dcf1553131affba480d1558890c5a9220cd17759011a7b2e9cf5901ae0224ed5148e412c1a;
    5'b10001 : xpb = 1024'h2d5fd6dd023d952f81b5bbd0c1fc60b04ffcad31c08485d6f2ad0009216d8b2cb14a765a417423ac857075acbd4d474a46f2c45465ff8d6e9858e7238f5f55367baf2c01f39c600b782dce1fa12ec305a2a9d7468397d6d74b083fba17afd89710dc510e1484002b82dbb1097d88d35655fe1d630ef288342d41b1c668418ba9;
    5'b10010 : xpb = 1024'h44d436f419300d9537d02041a224e73cbc64b7c1f403cdc4792b7f40ed29021225848c136c25259a45af56dd5ba82f5765f510ceca6eea7e0161cf038faae06caec2cb61e96b5650816fcb7fe9d2e59341691f6baaeccaa9b01945973e0a7ffc71bcfd9b57b277c6400e4006299a4dab91810c292854f58838348e784241eb38;
    5'b10011 : xpb = 1024'h5c48970b302285faedea84b2824d6dc928ccc252278315b1ffa9fe78b8e478f799bea1cc96d6278805ee380dfa03176484f75d492ede478d6a6ab6e38ff66ba2e1d66ac1df3a4c958ab1c8e032770820e0286790d241be7c152a4b7464652761d29daa289ae0ef60fd40cf02d5abc800cd03faef41b762dc43276b2a1c424ac7;
    5'b10100 : xpb = 1024'h73bcf7224714fe60a404e9236275f4559534cce25b025d9f86287db0849fefdd0df8b785c1872975c62d193e985dff71a3f9a9c3934da49cd3739ec39041f6d914ea0a21d50942da93f3c6407b1b2aae7ee7afb5f996b24e7a3b51518abfcec7337e56b5de0f66fbba735dff81bd42560886e9b55b19d0304e1a47dbf642aa56;
    5'b10101 : xpb = 1024'h8b3157395e0776c65a1f4d94429e7ae2019cd7728e81a58d0ca6fce8505b66c28232cd3eec382b63866bfa6f36b8e77ec2fbf63df7bd01ac3c7c86a3908d820f47fda981cad8391f9d35c3a0c3bf4d3c1da6f7db20eba620df4c572eb11a762c945f0343213dde9677a5ecfc2dcebcab4409d87b747c3d84590d248dd04309e5;
    5'b10110 : xpb = 1024'ha2a5b75074f9ef2c1039b20522c7016e6e04e202c200ed7a93257c201c16dda7f66ce2f816e92d5146aadb9fd513cf8be1fe42b85c2c5ebba5856e8390d90d457b1148e1c0a72f64a677c1010c636fc9bc664000484099f3445d5d0bd7751d91f53fafd0646c563134d87bf8d9e037007f8cc7418ddeaad86400013faa436974;
    5'b10111 : xpb = 1024'h96cd211c9fe32c8fb4e9e9ef29540a968f6e962200894f09bc7420234cfa785675e7b387773b0b0678b7d899010a6ce9ce6674c9de8eb7f5def1705565223ca39d5b39306e528649d1fbbbebc2bce2667208e8ce30f60b4f3e1d0ee43a522652718ca33f6d1d53e6b4b24168e218b2c6c35d72556f5bafc288362ecfb616298;
    5'b11000 : xpb = 1024'h20e13228e0f0ab2eb169030fd2bdc735d55ef3f25387dcde2245c13a008b1e6adb9890f1a224b29e27ca5eba2e6b8edbbbe8b3c70258488ec6f7fee5569daf006ce952f2fcb41ea9a661b91f04cff0b405dfd6b20a64548758f2d6cb69ffc9ca87f976c13a004cd9287db3133a330581a7b8c5eb7058285033763f9ed561c227;
    5'b11001 : xpb = 1024'h3855923ff7e3239467836780b2e64dc241c6fe82870724cba8c44071cc4695504fd2a6aaccd5b48be8093feaccc676e8daeb004166c7a59e3000e6c556e93a369ffcf252f28314eeafa3b67f4d741341a49f1ed731b94859be03dca8905a712fe8da234e7d2ec473e5b0420fe6447fd6e33bb4b189ba95a43e691c50af6221b6;
    5'b11010 : xpb = 1024'h4fc9f2570ed59bfa1d9dcbf1930ed44eae2f0912ba866cb92f42bfa998020c35c40cbc63f786b679a848211b6b215ef5f9ed4cbbcb3702ad9909cea55734c56cd31091b2e8520b33b8e5b3df961835cf435e66fc590e3c2c2314e285b6b5189549bacfdbc05d3c0ea2e2d10c9255fa2c1ebea377a31d02f8495bf90289628145;
    5'b11011 : xpb = 1024'h673e526e25c8145fd3b8306273375adb1a9713a2ee05b4a6b5c13ee163bd831b3846d21d2237b8676887024c097c470318ef99362fa65fbd0212b685578050a306243112de210178c227b13fdebc585ce21daf2180632ffe8825e862dd0fbffaaa9b7c69038bb3a9601560093e6774815a41923dbc7f704c544ed5b46362e0d4;
    5'b11100 : xpb = 1024'h7eb2b2853cba8cc589d294d3535fe16786ff1e332184fc943c3fbe192f78fa00ac80e7d64ce8ba5528c5e37ca7d72f1037f1e5b09415bccc6b1b9e6557cbdbd93937d072d3eff7bdcb69aea027607aea80dcf746a7b823d0ed36ee40036a67600b7c28f646ba2b441d47ef05ea78eed695c48103d5e1dda05f41b2663d634063;
    5'b11101 : xpb = 1024'h9627129c53ad052b3fecf944338867f3f36728c355044481c2be3d50fb3470e620bafd8f7799bc42e904c4ad4632171d56f4322af88519dbd42486455817670f6c4b6fd2c9beee02d4abac0070049d781f9c3f6bcf0d17a35247f41d29c50ec56c5cd58389e8a2deda7a7e02968a692bd1476fc9ef444af46a348f1817639ff2;
    5'b11110 : xpb = 1024'had9b72b36a9f7d90f6075db513b0ee805fcf335388838c6f493cbc88c6efe7cb94f51348a24abe30a943a5dde48cff2a75f67ea55cf476eb3d2d6e255862f2459f5f0f32bf8de447ddeda960b8a8c005be5b8790f6620b75b758f9fa501fb62acd3d8210cd171a7997ad0cff429be3810cca5e9008a6b84875276bc9f163ff81;
    5'b11111 : xpb = 1024'h14628d74bfa3c12de11c4a4ee37f2dbb5ac13ab2e68b33e551de826adfa8b1a905e6ab8902d5418fca2447c79f89d66d30dea3399eb103aef59716a71ddc08ca5e2379e405cbdd47d495a41e68711e626915d61d9130d23766dd6ddcbc4fbafdff169c745f7c9986ce1fb51cf6dd37acf9736e73d1bdc86c39aacd774281f8a5;
    endcase
end

endmodule

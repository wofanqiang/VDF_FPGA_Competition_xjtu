module xpb_5_310
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9de4b0cc66cf564884d6a96e8814b55ba93d4d5c86cb8474c1189a3b21a792faa24c14a31cec91d66c5786c2e3d1e43adc3a1fba021a6376e5ec8e196b0fa0a85e3a8b3aef5e420d09a16e5a22288897617321d918daba01a2d29fb241232f6df8de3c05e4085fb65cd7462f7b1a4277fe840ea46ac5b02037f2d9e379c6cd1c;
    5'b00010 : xpb = 1024'h8b1c1c430bb077c83ea7db05ffcf2365e1049788381f687204547b20904c78ed414fabcd6fb2a51e3950ce3ee445b7ab545a178de181f6a21b39dcd49b4ccc9f4825e1c72f2b86d500a8da11ab754cfdcee14a19a52f46f29018ad69c81bbc49c2b4e5e21747c6df32eea57ffe645ec6ae2e3e6685400310297638c26aab33cd;
    5'b00011 : xpb = 1024'h785387b9b0919947f8790c9d7789917018cbe1b3e9734c6f47905c05fef15edfe05342f7c278b866064a15bae4b98b1bcc7a0f61c0e989cd50872b8fcb89f896321138536ef8cb9cf7b045c934c211643c4f725a3183d3e37d5ebb214f1449258c8b8fbe4a872e08090604d081ae7b155dd86e289fba56001af997a15b8f9a7e;
    5'b00100 : xpb = 1024'h658af3305572bac7b24a3e34ef43ff7a50932bdf9ac7306c8acc3ceb6d9644d27f56da22153ecbadd3435d36e52d5e8c449a0735a0511cf885d47a4afbc7248d1bfc8edfaec61064eeb7b180be0ed5caa9bd9a9abdd860d46aa4c8d8d60cd6015662399a7dc69530df1d642104f897640d829deaba34a8f00c7cf6804c74012f;
    5'b00101 : xpb = 1024'h52c25ea6fa53dc476c1b6fcc66fe6d84885a760b4c1b1469ce081dd0dc3b2ac51e5a714c6804def5a03ca4b2e5a131fcbcb9ff097fb8b023bb21c9062c04508405e7e56bee93552ce5bf1d38475b9a31172bc2db4a2cedc557ead6905d0562dd2038e376b105fc59b534c3718842b3b2bd2ccdacd4aefbdffe00555f3d5867e0;
    5'b00110 : xpb = 1024'h3ff9ca1d9f34fdc725eca163deb8db8ec021c036fd6ef8671143feb64ae010b7bd5e0876bacaf23d6d35ec2ee615056d34d9f6dd5f20434ef06f17c15c417c7aefd33bf82e6099f4dcc688efd0a85e978499eb1bd6817ab64530e447e3fdefb8ea0f8d52e44563828b4c22c20b8cd0016cd6fd6eef294ecfef83b43e2e3cce91;
    5'b00111 : xpb = 1024'h2d31359444161f46dfbdd2fb56734998f7e90a62aec2dc64547fdf9bb984f6aa5c619fa10d9105853a2f33aae688d8ddacf9eeb13e87d67a25bc667c8c7ea871d9be92846e2ddebcd3cdf4a759f522fdf208135c62d607a73276f1ff6af67c94b3e6372f1784caab616382128ed6ec501c812d3109a3a1bfe107131d1f213542;
    5'b01000 : xpb = 1024'h1a68a10ae8f740c6998f0492ce2db7a32fb0548e6016c06197bbc0812829dc9cfb6536cb605718cd07287b26e6fcac4e2519e6851def69a55b09b537bcbbd468c3a9e910adfb2384cad5605ee341e7645f763b9cef2a94981fbcffb6f1ef09707dbce10b4ac431d4377ae1631221089ecc2b5cf3241df4afd28a71fc10059bf3;
    5'b01001 : xpb = 1024'h7a00c818dd862465360362a45e825ad67779eba116aa45edaf7a16696cec28f9a68cdf5b31d2c14d421c2a2e7707fbe9d39de58fd56fcd0905703f2ecf9005fad953f9cedc8684cc1dccc166c8eabcacce463dd7b7f21890d030d6e78e7964c47938ae77e0398fd0d9240b3956b24ed7bd58cb53e98479fc40dd0db00ea02a4;
    5'b01010 : xpb = 1024'ha584bd4df4a7b88ed836df98cdfcdb0910b4ec16983628d39c103ba1b876558a3cb4e298d009bdeb40794965cb4263f97973fe12ff7160477643920c5808a1080bcfcad7dd26aa59cb7e3a708eb734622e5785b69459db8aafd5ad20ba0ac5ba4071c6ed620bf8b36a6986e3108567657a599b59a95df7bffc00aabe7ab0cfc0;
    5'b01011 : xpb = 1024'h92bc28c49988da0e9208113045b74913487c3642498a0cd0df4c1c87271b3b7cdbb879c322cfd1330d7290e1cbb63769f193f5e6ded8f372ab90e0c78845ccfef5bb21641cf3ef21c285a6281803f8c89bc5adf720ae687b9d1bbad8410352960a4870c9954b5fdc4080e63393cf83b42a03cb1bc3d84aafed84099d6b953671;
    5'b01100 : xpb = 1024'h7ff3943b3e69fb8e4bd942c7bd71b71d8043806dfaddf0ce2287fd6c95c0216f7abc10ed7595e47ada6bd85dcc2a0ada69b3edbabe40869de0de2f82b882f8f5dfa677f05cc133e9b98d11dfa150bd2f0933d637ad02f56c8a61c88fc7fbdf71d41f1aa5c88ac705169845841719a002d9adfaddde529d9fdf07687c5c799d22;
    5'b01101 : xpb = 1024'h6d2affb1e34b1d0e05aa745f352c2527b80aca99ac31d4cb65c3de520465076219bfa817c85bf7c2a7651fd9cc9dde4ae1d3e58e9da819c9162b7e3de8c024ecc991ce7c9c8e78b1b0947d972a9d819576a1fe783957825d77a7d6474ef46c4d9df5c481fbca2e2decafa4d49a63bc5189582a9ff8ccf08fd08ac75b4d5e03d3;
    5'b01110 : xpb = 1024'h5a626b28882c3e8dbf7ba5f6ace69331efd214c55d85b8c8a8ffbf377309ed54b8c33f421b220b0a745e6755cd11b1bb59f3dd627d0facf44b78ccf918fd50e3b37d2508dc5bbd79a79be94eb3ea45fbe41026b8c5ac0f4e64ede3fed5ecf92967cc6e5e2f099556c2c704251dadd8a039025a621347437fc20e263a3e426a84;
    5'b01111 : xpb = 1024'h4799d69f2d0d600d794cd78e24a1013c27995ef10ed99cc5ec3ba01ce1aed34757c6d66c6de81e524157aed1cd85852bd213d5365c77401f80c61bb4493a7cda9d687b951c2902419ea355063d370a62517e4ef952009c3f5233f1b65ce5860531a3183a6248fc7f98de6375a0f7f4eee8ac8a242dc1966fb39185192f26d135;
    5'b10000 : xpb = 1024'h34d14215d1ee818d331e09259c5b6f465f60a91cc02d80c32f7781025053b939f6ca6d96c0ae319a0e50f64dcdf9589c4a33cd0a3bded34ab6136a6f7977a8d18753d2215bf6470995aac0bdc683cec8beec7739de5529303f79ff6de3de12e0fb79c216958863a86ef5c2c62442113d9856b9e6483be95fa514e3f8200b37e6;
    5'b10001 : xpb = 1024'h2208ad8c76cfa30cecef3abd1415dd509727f348718164c072b361e7bef89f2c95ce04c1137444e1db4a3dc9ce6d2c0cc253c4de1b466675eb60b92aa9b4d4c8713f28ad9bc38bd18cb22c754fd0932f2c5a9f7a6aa9b6212cc00d256ad69fbcc5506bf2c8c7cad1450d2216a78c2d8c4800e9a862b63c4f969842d710ef9e97;
    5'b10010 : xpb = 1024'hf4019031bb0c48ca6c06c548bd04b5aceef3d7422d548bdb5ef42cd2d9d851f34d19beb663a5829a8438545cee0ff7d3a73bcb1faadf9a120ae07e5d9f200bf5b2a7f39db90d09983b9982cd91d579599c8c7baf6fe43121a061adcf1cf2c988f2715cefc0731fa1b2481672ad649daf7ab196a7d308f3f881ba1b601d40548;
    5'b10011 : xpb = 1024'had24c9cf82801ad52b9715c313e500b6782c8ad0a9a0cd327707dd084f451819d71db08e8326ea00149b0c08b2b2e3b816addc6bfcc85d18069a95ff4501a167b9650a74caef12a68d5b0686fb45e02cfb3be9940fd8fd13bcd8ba8f32f25c06880551d4e00f91b077fbc796a5f08c52f62f280ee7f63f5fc00e7b997b9ad264;
    5'b10100 : xpb = 1024'h9a5c354627613c54e568475a8b9f6ec0aff3d4fc5af4b12fba43bdedbde9fe0c762147b8d5ecfd47e1945384b326b7288ecdd43fdc2ff0433be7e4ba753ecd5ea35061010abc576e8462723e8492a49368aa11d49c2d8a04aa1ec846b9eae8e251dbfbb1134ef8d94e1326e7293aa8a1a5d957d10270924fb191da786c7f3915;
    5'b10101 : xpb = 1024'h8793a0bccc425dd49f3978f20359dccae7bb1f280c48952cfd7f9ed32c8ee3ff1524dee328b3108fae8d9b00b39a8a9906edcc13bb97836e71353375a57bf9558d3bb78d4a899c367b69ddf60ddf68f9d6183a15288216f59764d5fe40e375be1bb2a58d468e6002242a8637ac84c4f0558387931ceae53fa31539575d639fc6;
    5'b10110 : xpb = 1024'h74cb0c3371237f54590aaa897b144ad51f826953bd9c792a40bb7fb89b33c9f1b428760d7b7923d77b86e27cb40e5e097f0dc3e79aff1699a6828230d5b9254c77270e198a56e0fe727149ad972c2d6043866255b4d6a3e684aae3b5c7dc0299e5894f6979cdc72afa41e5882fcee13f052db7553765382f949898364e480677;
    5'b10111 : xpb = 1024'h620277aa1604a0d412dbdc20f2ceb8df5749b37f6ef05d2783f7609e09d8afe4532c0d37ce3f371f488029f8b4823179f72dbbbb7a66a9c4dbcfd0ec05f65143611264a5ca2425c66978b5652078f1c6b0f48a96412b30d771f0f16d4ed48f75af5ff945ad0d2e53d05944d8b318fd8db4d7e71751df8b1f861bf7153f2c6d28;
    5'b11000 : xpb = 1024'h4f39e320bae5c253ccad0db86a8926e98f10fdab20444124c7334183787d95d6f22fa46221054a6715797174b4f604ea6f4db38f59ce3cf0111d1fa736337d3a4afdbb3209f16a8e6080211ca9c5b62d1e62b2d6cd7fbdc85f36ff24d5cd1c517936a321e04c957ca670a429366319dc648216d96c59de0f779f55f43010d3d9;
    5'b11001 : xpb = 1024'h3c714e975fc6e3d3867e3f4fe24394f3c6d847d6d19825220a6f2268e7227bc991333b8c73cb5daee272b8f0b569d85ae76dab633935d01b466a6e626670a93134e911be49beaf5657878cd433127a938bd0db1759d44ab94c7d0cdc5cc5a92d430d4cfe138bfca57c880379b9ad362b142c469b86d430ff6922b4d320f53a8a;
    5'b11010 : xpb = 1024'h29a8ba0e04a80553404f70e759fe02fdfe9f920282ec091f4dab034e55c761bc3036d2b6c69170f6af6c006cb5ddabcb5f8da337189d63467bb7bd1d96add5281ed4684a898bf41e4e8ef88bbc5f3ef9f93f0357e628d7aa39c31a93e3be36090ce3f6da46cb63ce529f62ca3cf75279c3d6765da14e83ef5aa613b211d9a13b;
    5'b11011 : xpb = 1024'h16e02584a98926d2fa20a27ed1b871083666dc2e343fed1c90e6e433c46c47aecf3a69e11957843e7c6547e8b6517f3bd7ad9b0af804f671b1050bd8c6eb011f08bfbed6c95938e64596644345ac036066ad2b98727d649b2709284b6ab6c2e4d6baa0b67a0acaf728b6c21ac0416ec87380a61fbbc8d6df4c29729102be07ec;
    5'b11100 : xpb = 1024'h41790fb4e6a4852b3f1d4164972df126e2e2659e593d119d422c51933112da16e3e010b6c1d9786495e8f64b6c552ac4fcd92ded76c899ce6525a93f7282d15f2ab156309267dae3c9dcffacef8c7c6d41b53d8fed1f18c144f3602f1af4fc0a0914a92ad4a321ffece216b438b8b17232ad5e1d64329cf3dacd16ff3a26e9d;
    5'b11101 : xpb = 1024'ha1fc41c7b5399e9b38c87d84d187946e176b73b66c5f558e953b5f5454b8c09c108a15ae890a295cb5b616279a9736e72c07b298d986ed13cc3ee8ad6237cdbe50e5a09df884bfbb463f3e54f121505e358e75b217acab8db721d5b532d27f2e996f8698915291d65ba5679abea5cd8f21aee4864108d9ef759fab536d693bb9;
    5'b11110 : xpb = 1024'h8f33ad3e5a1ac01af299af1c494202784f32bde21db3398bd8774039c35da68eaf8dacd8dbd03ca482af5da39b0b0a57a427aa6cb8ee803f018c37689274f9b53ad0f72a385204833d46aa0c7a6e14c4a2fc9df2a401387ea467e36cb9cb0c0a63463074c491f8ff31bcc6eb41efe9ddd15914485b832cdf67230a325e4da26a;
    5'b11111 : xpb = 1024'h7c6b18b4fefbe19aac6ae0b3c0fc708286fa080dcf071d891bb3211f32028c814e9144032e964fec4fa8a51f9b7eddc81c47a2409856136a36d98623c2b225ac24bc4db6781f494b344e15c403bad92b106ac6333055c56f91adf12440c398e62d1cda50f7d1602807d4263bc53a062c8103440a75fd7fcf58a669114f32091b;
    endcase
end

endmodule

module xpb_5_345
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5ff96a3e480fca4d0d6d18222959de54a294af1916cd3fd25d28b659483c532b3766dc2b95e3a101dde209bbc291c8d5979aa9820ba97a201c586287181952c2e302b6cd6319b41940b6d2df863f777767d1616dea106970cf4b33acc3da0ad7cc53c041a036ac0bbf1e3626f1b1cdc61f9a48e5b762922728b70e46544ceff7;
    5'b00010 : xpb = 1024'hf458f26ce315fd14fd4b86d42597557d3b35b015822df2d3c74b35cdd75f94e6b853ade61a0c3751c65d430a1c580e0cb1b2b1df4a023f4881185aff56030d451b638ec16a26aed6ed3a31c73a32abddb9dc943479aa5d0e909d55ecd89731d699fee598fa45f89f77c856eeb937562f05ab2e91e79c71e0afea1881fb77983;
    5'b00011 : xpb = 1024'h6f3ef96516412a1e5d41d08f6bb353ac76480a1a6ef01eff999d69b625b24c79a2ec1709f7846476fa47ddec645749b662b5d4a000499e14a469e8370d79839734b8efb979bc1f06af8a75fbf9e2a235436f2ab131ab0f41b855090b91637df535f3ae9b2fdb0b95b69abb95dd4543290ff4fbced5dc594533b5afce7404697a;
    5'b00100 : xpb = 1024'h1e8b1e4d9c62bfa29fa970da84b2eaafa766b602b045be5a78e966b9baebf29cd70a75bcc34186ea38cba861438b01c19636563be94047e910230b5feac061a8a36c71d82d44d5dadda74638e746557bb73b92868f354ba1d213aabd9b12e63ad33fdcb31f48bf13eef90addd726eac5e0b565d23cf38e3c15fd43103f6ef306;
    5'b00101 : xpb = 1024'h7e84888be47289efad1688fcae0cc90449fb651bc712fe2cd6121d13032845c80e7151e8592527ec16adb21d061cca972dd0ffbdf4e9c2092c7b6de702d9b46b866f28a5905e89f41e5e19186d85ccf31f0cf3f47945b512a15ede6a5eecf1129f939cf4bf7f6b1fae174104c8d8b88c004faeb7f45620633eb4515693bbe2fd;
    5'b00110 : xpb = 1024'h2dd0ad746a941f73ef7e2947c70c60077b1a110408689d87b55e1a169861ebeb428fb09b24e24a5f55317c91e55082a261518159dde06bdd9834910fe020927cf522aac443e740c84c7ae9555ae9803992d95bc9d6cff172bb1d801c689c59583cdfcb0caeed1e9de675904cc2ba6028d11018bb5b6d555a20fbe4985f266c89;
    5'b00111 : xpb = 1024'h8dca17b2b2a3e9c0fceb4169f0663e5c1daec01d1f35dd5a1286d06fe09e3f1679f68cc6bac5eb613313864da7e24b77f8ec2adbe989e5fdb48cf396f839e53fd8256191a700f4e18d31bc34e128f7b0faaabd37c0e05ae38a68b3c92c76643009338b4e4f23caa9a593c673b46c2deef0aa61a112cfe78149b2f2deb3735c80;
    5'b01000 : xpb = 1024'h3d163c9b38c57f453f52e1b50965d55f4ecd6c05608b7cb4f1d2cd7375d7e539ae14eb7986830dd4719750c2871603832c6cac77d2808fd2204616bfd580c35146d8e3b05a89abb5bb4e8c71ce8caaf76e77250d1e6a9743a427557b3625cc75a67fb9663e917e27ddf215bbae4dd58bc16acba479e71c782bfa86207edde60c;
    5'b01001 : xpb = 1024'h9d0fa6d980d549924cbff9d732bfb3b3f1621b1e7758bc874efb83ccbe143864e57bc7a51c66aed64f795a7e49a7cc58c40755f9de2a09f23c9e7946ed9a161429db9a7dbda35fcefc055f5154cc226ed648867b087b00b473728927f9ffd74d72d379a7dec82a339d104be29fffa351e105148a3149ae9f54b19466d32ad603;
    5'b01010 : xpb = 1024'h4c5bcbc206f6df168f279a224bbf4ab72280c706b8ae5be22e4780d0534dde88199a2657e823d1498dfd24f328db8463f787d795c720b3c6a8579c6fcae0f425988f1c9c712c16a32a222f8e422fd5b54a14ee5066053d148d312ada03af3f93101fa7bfce35ddb1d56e9b2a99e14aeeb1c57e8d9860e39636f927a89e955f8f;
    5'b01011 : xpb = 1024'hac5536004f06a9639c94b2447519290bc515761fcf7b9bb48b7037299b8a31b3510102837e07724b6bdf2eaeeb6d4d398f228117d2ca2de6c4affef6e2fa46e87b91d369d445cabc6ad9026dc86f4d2cb1e64fbe5015a6855c7c5e86c7894a6adc7368016e6c89bd948cd1518b9318b4d15fc7734fc375bd5fb035eef2e24f86;
    5'b01100 : xpb = 1024'h5ba15ae8d5283ee7defc528f8e18c00ef634220810d13b0f6abc342d30c3d7d6851f613649c494beaa62f923caa10544c2a302b3bbc0d7bb3069221fc04124f9ea45558887ce819098f5d2aab5d3007325b2b793ad9fe2e5763b0038d138b2b079bf96195dda3d3bcceb20998574c051a2203176b6daaab441f7c930be4cd912;
    5'b01101 : xpb = 1024'haed7fd15b49d46c2163f2daa71857122752cdf05226da6a4a083130c5fd7df9b93dbfe91581b731e8e6c398a9d4bd4ff623844fa4b7818f9c2245489d88030b58f8d7a73b573864c712a2e7a336b3b9997f1f690b2a1f458ff9a1eadae81af6170bc4314d47f0ba05496fe17f5667ee72e09b7a1df1dfab243f5c7289b7629e;
    5'b01110 : xpb = 1024'h6ae6ea0fa3599eb92ed10afcd0723566c9e77d0968f41a3ca730e78a0e39d124f0a49c14ab655833c6c8cd546c6686258dbe2dd1b060fbafb87aa7cfb5a155ce3bfb8e749e70ec7e07c975c729762b31015080d6f53a88b65f44d5979ec225cde35f8472ed7e9cc5c467a608710835b4927ae45fd55471d24cf66ab8de045295;
    5'b01111 : xpb = 1024'h1a330ef8297b343d7138ab47e971cc69fb0628f1aa49b997867ce48da373774824c2fac777227aa7054c97c94b9a3e30c13eaf6d9957a5842433caf892e833dfaaaf109351f9a35235e6460416d9de77751ce8ac52c4c51679037749a8718e1380abb28adcec5043fcc5f5506ae9dd51633b4e633c6ba6c92f3dfdfaa96edc21;
    5'b10000 : xpb = 1024'h7a2c7936718afe8a7ea5c36a12cbaabe9d9ad80ac116f969e3a59ae6ebafca735c29d6f30d061ba8e32ea1850e2c070658d958efa5011fa4408c2d7fab0186a28db1c760b513576b769d18e39d1955eedcee4a1a3cd52e87484eaaf66c4b98eb4cff72cc7d22fc4fbbe42b775c9bab1782d59748f3ce38f057f50c40fdbbcc18;
    5'b10001 : xpb = 1024'h29789e1ef7ac940ec10d63b52bcb41c1ceb983f3026c98c4c2f197ea80e97096904835a5d8c33e1c21b26bf9ed5fbf118c59da8b8df7c978ac4550a8884864b3fc65497f689c0e3fa4b9e9208a7d093550bab1ef9a5f6ae7620d4ca875fb0130ea4ba0e46c90afcdf4427abf567d52b45396014c5ae56de73a3c9f82c92655a4;
    5'b10010 : xpb = 1024'h8972085d3fbc5e5bce7a7bd755252016714e330c1939d897201a4e43c925c3c1c7af11d16ea6df1dff9475b5aff187e723f4840d99a14398c89db32fa061b776df68004ccbb5c258e570bc0010bc80acb88c135d846fd4583158805539d50c08b69f61260cc75bd9b360b0e6482f207a73304a321248000e62f3adc91d73459b;
    5'b10011 : xpb = 1024'h38be2d45c5ddf3e010e21c226e24b719a26cdef45a8f77f1ff664b475e5f69e4fbcd70843a6401913e18402a8f253ff2577505a98297ed6d3456d6587da895884e1b826b7f3e792d138d8c3cfe2033f32c587b32e1fa10b84b1722074384744e53eb8f3dfc350f57ebbf002e4210c81743f0b435795f3505453b410ae8ddcf27;
    5'b10100 : xpb = 1024'h98b797840dedbe2d1e4f3444977e956e45018e0d715cb7c45c8f01a0a69bbd1033344cafd047a2931bfa49e651b708c7ef0faf2b8e41678d50af38df95c1e84b311e3938e2582d4654445f1c845fab6a9429dca0cc0a7a291a6255b4075e7f26203f4f7f9c6bbb63aadd365533c295dd638afd1b30c1c72c6df24f513d2abf1e;
    5'b10101 : xpb = 1024'h4803bc6c940f53b160b6d48fb07e2c71762039f5b2b2571f3bdafea43bd563336752ab629c04c5065a7e145b30eac0d3229030c777381161bc685c087308c65c9fd1bb5795e0e41a82612f5971c35eb107f644762994b6893420f766110de76bbd8b7d978bd96ee1e33b859d2da43d7a344b671e97d8fc235039e293089548aa;
    5'b10110 : xpb = 1024'ha7fd26aadc1f1dfe6e23ecb1d9d80ac618b4e90ec97f96f19903b4fd8411b65e9eb9878e31e8660838601e16f37c89a8ba2ada4982e18b81d8c0be8f8b22191f82d47224f8fa9833c3180238f802d6286fc7a5e413a51ffa036c2b12d4e7f24389df3dd92c101aeda259bbc41f560b4053e5b0044f3b8e4a78f0f0d95ce238a1;
    5'b10111 : xpb = 1024'h57494b936240b382b08b8cfcf2d7a1c949d394f70ad5364c784fb201194b5c81d2d7e640fda5887b76e3e88bd2b041b3edab5be56bd835564479e1b86868f730f187f443ac834f07f134d275e566896ee3940db9712f5c5a1d2accc4de975a89272b6bf11b7dce6bdab80b0c1937b2dd24a61a07b652c3415b38841b284cc22d;
    5'b11000 : xpb = 1024'h695707be8624906f2f32d480bd738cc7af240df4c2ad5a7579baf04ae8502a506f644f3c962aaeeb567b300b1e3f9bf212bdd8154cedf2ab03304e145afd542603b7662600c05dc1f51a2b2d2ca3cb55760758eceb998ba36e96e76e846c2cec4779a090aeb81ea13165a5413195a79f566840b1d69f8383d80175cf3b74bb9;
    5'b11001 : xpb = 1024'h668edaba307213540060456a353117211d86eff862f81579b4c4655df6c155d03e5d211f5f464bf09349bcbc7475c294b8c687036078594acc8b67685dc92805433e2d2fc325b9f5600875925909b42cbf31d6fcb8ca022b0634a223ac20cda690cb5a4aab222df5d234907b04cb28401500ccf0d4cc8a5f663725a348043bb0;
    5'b11010 : xpb = 1024'h15daffa2b693a8d842c7e5b54e30ae244ea59be0a44db4d4941062618bfafbf3727b7fd22b036e63d1cd873153a97a9fec47089f496f031f38448a913b100616b1f1af4e76ae70c98e2545cf466d677332fe3ed216543e8b1ff343d5b5d035ec2e1788629a8fe1740a92dfc2feaccfdce5c136f43be3bf56487eb8e5136ec53c;
    5'b11011 : xpb = 1024'h75d469e0fea373255034fdd7778a8c78f13a4af9bb1af4a6f13918bad4374f1ea9e25bfdc0e70f65afaf90ed163b437583e1b22155187d3f549ced18532958d994f4661bd9c824e2cedc18aeccacdeea9acfa0400064a7fbef3e778279aa40c3fa6b48a43ac68d7fc9b115e9f05e9da3055b7fd9f346517d7135c72b67bbb533;
    5'b11100 : xpb = 1024'h25208ec984c508a9929c9e22908a237c2258f6e1fc709401d08515be6970f541de00bab08ca431d8ee335b61f56efb80b76233bd3e0f2713c0561041307036eb03a7e83a8d50dbb6fcf8e8ebba1092310e9c08155deee45c08fd19348359a90997b776bc2a3440fe020f6531ea40453fd61be9dd5a5d8674537d5a6d33263ebf;
    5'b11101 : xpb = 1024'h8519f907ccd4d2f6a009b644b9e401d0c4eda5fb133dd3d42dadcc17b1ad486d156796dc2287d2dacc15651db800c4564efcdd3f49b8a133dcae72c8488989ade6aa9f07f06a8fd03dafbbcb405009a8766d698347ff4dccd8484ce14733b3e1640b36fdca6aed09c12d9b58dbf21305f5b632c311c0189b7c3468b387732eb6;
    5'b11110 : xpb = 1024'h34661df052f6687ae271568fd2e398d3f60c51e35493732f0cf9c91b46e6ee904985f58eee44f54e0a992f9297347c61827d5edb32af4b08486795f125d067bf555e2126a3f346a46bcc8c082db3bceeea39d158a5898a2cf206ee9350e31c2701576515b9d8a087f98beaa0d5d3baa2c6769cc678d74d925e7bfbf552ddb842;
    5'b11111 : xpb = 1024'h945f882e9b0632c7efde6eb1fc3d772898a100fc6b60b3016a227f748f2341bb80ecd1ba8428964fe87b394e59c645371a18085d3e58c52864bff8783de9ba823860d7f4070cfabdac835ee7b3f33466520b32c68f99f39dc152224014bd26fecdab25575a0f4c93b8aa20c7c7858868e610e5ac3039dfb987330a3ba72aa839;
    endcase
end

endmodule

module xpb_5_715
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h902dfdbceeb0a218bd444deb1b9fbdc3362636d0093a597d052770f41a688a3c9c19dc07e5cb3e92b7d79303cec47e2dbfde50cddbc32868dc65204b5e18bfb75360ee070046cdda7838e9b0e180d61feadabbc49577b48062935b445b86ef74b8a4e516f9292b1f817cb518c49db346e77d30087db0c6681a696f303dee5632;
    5'b00010 : xpb = 1024'h6faeb6241b730f68af8323ff26e53434fad66a6f3cfd12828c72289281ce677134eb3a97016ffe96d050e6c0ba2aeb911ba279b594d38086082b0138815f0abd3272a75f50fc9e6fddd7d0bf2a25e80ee1b07df09e693bf00f9a248dfce33c574242380441895db17c398352916b40648020812eab162f9fee63635bf2fa45f9;
    5'b00011 : xpb = 1024'h4f2f6e8b48357cb8a1c1fa13322aaaa6bf869e0e70bfcb8813bce030e93444a5cdbc99261d14be9ae8ca3a7da59158f47766a29d4de3d8a333f0e225a4a555c3118460b7a1b26f054376b7cd72caf9fdd886401ca75ac35fbca0edd79e3f8939cbdf8af189e9904376f6518c5e38cd8218c3d254d87b98d7c25d5787a80635c0;
    5'b00100 : xpb = 1024'h2eb026f274f7ea089400d0273d7021188436d1ada482848d9b0797cf509a21da668df7b538b97e9f01438e3a90f7c657d32acb8506f430c05fb6c312c7eba0c8f0961a0ff2683f9aa9159edbbb700beccf5c0248b04c4acf69a7b7213f9bd61c557cddded249c2d571b31fc62b065a9fb167237b05e1020f96574bb35d122587;
    5'b00101 : xpb = 1024'he30df59a1ba5758863fa63b48b5978a48e7054cd8453d9322524f6db7ffff0eff5f5644545e3ea319bce1f77c5e33bb2eeef46cc00488dd8b7ca3ffeb31ebcecfa7d368431e10300eb485ea04151ddbc631c474b93dd23f16ae806ae0f822fedf1a30cc1aa9f5676c6fedfff7d3e7bd4a0a74a133466b476a513fdf121e154e;
    5'b00110 : xpb = 1024'h9e5edd16906af9714383f4266455554d7f0d3c1ce17f97102779c061d268894b9b79324c3a297d35d19474fb4b22b1e8eecd453a9bc7b14667e1c44b494aab862308c16f4364de0a86ed6f9ae595f3fbb10c80394eb586bf7941dbaf3c7f127397bf15e313d32086edeca318bc719b043187a4a9b0f731af84baaf0f500c6b80;
    5'b00111 : xpb = 1024'h7ddf957dbd2d66c135c2ca3a6f9acbbf43bd6fbc15425015aec4780039ce6680344a90db55ce3d39ea0dc8b836891f4c4a916e2254d8096393a7a5386c90f68c021a7ac7941aae9fec8c56a92e3b05eaa7e2426557a70e2f2648a4f8dddb5f56215c68d05c335318e8a97152893f2821ca2af5cfde5c9ae758b4a33b05185b47;
    5'b01000 : xpb = 1024'h5d604de4e9efd4112801a04e7ae04231086da35b4905091b360f2f9ea13443b4cd1bef6a7172fd3e02871c7521ef8cafa655970a0de86180bf6d86258fd74191e12c341fe4d07f35522b3db776e017d99eb804916098959ed34f6e427f37ac38aaf9bbbda49385aae3663f8c560cb53f62ce46f60bc2041f2cae9766ba244b0e;
    5'b01001 : xpb = 1024'h3ce1064c16b241611a4076628625b8a2cd1dd6fa7cc7c220bd59e73d089a20e965ed4df98d17bd421b0070320d55fa130219bff1c6f8b99deb336712b31d8c97c03ded7835864fcab7ca24c5bf8529c8958dc6bd698a1d0e8056378c2093f91b34970eaaecf3b83cde230dc622da425cfb71981c39276d5700a88b926f303ad5;
    5'b01010 : xpb = 1024'h1c61beb34374aeb10c7f4c76916b2f1491ce0a99b08a7b2644a49edb6ffffe1dfebeac88a8bc7d463379c3eef8bc67765ddde8d9800911bb16f947ffd663d79d9f4fa6d0863c20601d690bd4082a3bb78c6388e9727ba47e2d5d00d5c1f045fdbe3461983553eaced8dfdbffefa7cf7a9414e942668cd68ed4a27fbe243c2a9c;
    5'b01011 : xpb = 1024'hac8fbc70322550c9c9c39a61ad0aecd7c7f44169b9c4d4a349cc0fcf8a68885a9ad888908e87bbd8eb5156f2c780e5a41dbc39a75bcc3a23f35e684b347c9754f2b094d78682ee3a95a1f584e9ab11d7773e44ae07f358fe8ff05c1a1d77357276d946af2e7d15ee5a5c9118b44582c17b92194ae43d9cf6ef0beeee622a80ce;
    5'b01100 : xpb = 1024'h8c1074d75ee7be19bc027075b85063498ca47508ed878da8d116c76df1ce658f33a9e71faa2c7bdd03caaaafb2e753077980628f14dc92411f24493857c2e25ad1c24e2fd738becffb40dc93325023c66e1406da10e4e06e3cf72563bed382550076999c76dd488055195f5281130fdf14356a7111a3062ec305e31a17367095;
    5'b01101 : xpb = 1024'h6b912d3e8baa2b69ae414689c395d9bb5154a8a8214a46ae58617f0c593442c3cc7b45aec5d13be11c43fe6c9e4dc06ad5448b76cdecea5e4aea2a257b092d60b0d4078827ee8f6560dfc3a17af535b564e9c90619d667dde9fdeead602fcf378a13ec89bf3d7b124fd62d8c4de09cfcacd8bb973f086f6696ffd745cc42605c;
    5'b01110 : xpb = 1024'h4b11e5a5b86c98b9a0801c9dcedb502d1604dc47550cffb3dfac36aac09a1ff8654ca43de175fbe534bd522989b42dce3108b45e86fd427b76b00b129e4f78668fe5c0e078a45ffac67eaaafc39a47a45bbf8b3222c7ef4d9704b7f7018c1c1a13b13f77079dada44a92fbc61aae2a1a457c0cbd6c6dd89e6af9cb71814e5023;
    5'b01111 : xpb = 1024'h2a929e0ce52f060992bef2b1da20c69edab50fe688cfb8b966f6ee4927fffd2cfe1e02ccfd1abbe94d36a5e6751a9b318cccdd46400d9a98a275ebffc195c36c6ef77a38c95a30902c1d91be0c3f599352954d5e2bb976bd440b8140a2e868fc9d4e92644ffde036454fc9ffe77bb737de1f5de399d341d63ef3bf9d365a3fea;
    5'b10000 : xpb = 1024'ha13567411f1735984fdc8c5e5663d109f654385bc9271beee41a5e78f65da6196ef615c18bf7bed65aff9a360810894e891062df91df2b5ce3bccece4dc0e724e0933911a10012591bc78cc54e46b82496b0f8a34aafe2cf1124a8a4444b5df26ebe551985e12c8400c9839b449445576c2af09c738ab0e12edb3c8eb662fb1;
    5'b10001 : xpb = 1024'h9a41543100a21572424216b10105fad3d58b7a55c5cccb3bf36916dba9ce649e33093d63fe8aba801d878ca72f4586c2a86f56fbd4e11b1eaaa0ed3842f4ce29a16a21981a56cf0009f5627d366541a23445cb4eca22b2ad53a5a5ce9fcba553df90ca6891873de7c1894d5278e6f79c5e3fdf1244e971762d5722f9295485e3;
    5'b10010 : xpb = 1024'h79c20c982d6482c23480ecc50c4b71459a3badf4f98f84417ab3ce7a113441d2cbda9bf31a2f7a843600e0641aabf42604337fe38df1733bd666ce25663b192f807bdaf06b0c9f956f94498b7f0a53912b1b8d7ad3143a1d00ac6f184127f236692e1d55d9e77079bc461b8c45b484b9f6e33038724edaae01511724de6075aa;
    5'b10011 : xpb = 1024'h5942c4ff5a26f01226bfc2d91790e7b75eebe1942d523d4701fe8618789a1f0764abfa8235d43a884e7a3421061261895ff7a8cb4701cb59022caf12898164355f8d9448bbc2702ad5333099c7af658021f14fa6dc05c18cadb33861e2843f18f2cb70432247a30bb702e9c6128211d78f86815e9fb443e5d54b0b50936c6571;
    5'b10100 : xpb = 1024'h38c37d6686e95d6218fe98ed22d65e29239c15336114f64c89493db6dffffc3bfd7d59115178fa8c66f387ddf178ceecbbbbd1b3001223762df28fffacc7af3b3e9f4da10c7840c03ad217a81054776f18c711d2e4f748fc5aba01ab83e08bfb7c68c3306aa7d59db1bfb7ffdf4f9ef52829d284cd19ad1da944ff7c48785538;
    5'b10101 : xpb = 1024'h184435cdb3abcab20b3d6f012e1bd49ae84c48d294d7af521093f5554765d970964eb7a06d1dba907f6cdb9adcdf3c50177ffa9ab9227b9359b870ecd00dfa411db106f95d2e1155a070feb658f9895e0f9cd3feede8d06c07c0caf5253cd8de0606161db308082fac7c8639ac1d2c12c0cd23aafa7f16557d3ef3a7fd8444ff;
    5'b10110 : xpb = 1024'ha872338aa25c6ccac881bcec49bb925e1e727fa29e1208cf15bb664961ce63ad326893a852e8f92337446e9eaba3ba7dd75e4b6894e5a3fc361d91382e26b9f87111f5005d74df3018a9e8673a7a5f7dfa778fc3836084ec6a54263980c3c852beaafb34ac31334f2df93b5270badf59a84a53b3782fdcbd97a862d83b729b31;
    5'b10111 : xpb = 1024'h87f2ebf1cf1eda1abac09300550108cfe322b341d1d4c1d49d061de7c93440e1cb39f2376e8db9274fbdc25b970a27e1332274504df5fc1961e37225516d04fe5023ae58ae2aafc57e48cf75831f716cf14d51ef8c520c5c175aef832220153548484e21f49165e128b6098c3d886c7740eda4d9a59545f56ba25703f07e8af8;
    5'b11000 : xpb = 1024'h6773a458fbe1476aacff691460467f41a7d2e6e105977ada2450d586309a1e16640b50c68a32792b68371618827095448ee69d38070654368da9531274b350042f3567b0fee0805ae3e7b683cbc4835be823141b954393cbc461b8ccc37c6217d1e5a10f3cf198732372d7c60a55f994d990f5ffd2faaf2d3f9c4b2fa58a7abf;
    5'b11001 : xpb = 1024'h46f45cc028a3b4ba9f3e3f286b8bf5b36c831a80395a33dfab9b8d2497fffb4afcdcaf55a5d7392f80b069d56dd702a7eaaac61fc016ac53b96f33ff97f99b0a0e4721094f9650f049869d921469954adef8d6479e351b3b7168821664d8aefa5b82f3fc8551cb051e2fa5ffd72386b2723447260060186513963f5b5a966a86;
    5'b11010 : xpb = 1024'h267515275566220a917d153c76d16c2531334e1f6d1cece532e644c2ff65d87f95ae0de4c17bf9339929bd92593d700b466eef0779270470e53514ecbb3fe60fed58da61a04c2185af2584a05d0ea739d5ce9873a726a2ab1e6f4b600634fbdce52046e9cdb1fd9718ec7439a3f113d00ad7984c2dc5819ce79033870fa25a4d;
    5'b11011 : xpb = 1024'h5f5cd8e82288f5a83bbeb508216e296f5e381bea0dfa5eaba30fc6166cbb5b42e7f6c73dd20b937b1a3114f44a3dd6ea23317ef32375c8e10faf5d9de863115cc6a93b9f101f21b14c46baea5b3b928cca45a9fb0182a1acb7614a9a79148bf6ebd99d71612302913a9427370bea0eda37ae9725b2aead4bb8a27b2c4ae4a14;
    5'b11100 : xpb = 1024'h9623cb4b70d931734100393b9db6a05a2c09b88eaa19ff67bf586d5581343ff0ca99487bc2ebf7ca697aa45313685b9c621168bd0dfa84f6ed6016253c9ef0cd1fcb81c0f148bff58cfd555f87348f48b77f1664458fde9b2e096fee0318383427627eee0f3b5b489525f78c355c54348af8197ad8dbb13cd5f396e3029ca046;
    5'b11101 : xpb = 1024'h75a483b29d9b9ec3333f0f4fa8fc16cbf0b9ec2ddddcb86d46a324f3e89a1d25636aa70ade90b7ce81f3f80ffecec8ffbdd591a4c70add141925f7125fe53bd2fedd3b1941fe908af29c3c6dcfd9a137ae54d8904e81660adb103937a4748516b0ffd1db579b8dda8fe2c5c60229e152239b6aa106411a74a9ed8b0eb7a8900d;
    5'b11110 : xpb = 1024'h55253c19ca5e0c13257de563b4418d3db56a1fcd119f7172cdeddc924ffffa59fc3c0599fa3577d29a6d4bccea3536631999ba8c801b353144ebd7ff832b86d8ddeef47192b46120583b237c187eb326a52a9abc5772ed7a8817028145d0d1f93a9d24c89ffbc06c8a9f93ffcef76e6fbc3ebbc733a683ac7de77f3a6cb47fd4;
    5'b11111 : xpb = 1024'h34a5f480f720796317bcbb77bf8703af7a1a536c45622a7855389430b765d78e950d642915da37d6b2e69f89d59ba3c6755de374392b8d4e70b1b8eca671d1debd00adc9e36a31b5bdda0a8a6123c5159c005ce8606474ea351dcbcae72d1edbc43a77b5e85bf2fe855c62399bc4fb8d54e20ced610bece451e1736621c06f9b;
    endcase
end

endmodule

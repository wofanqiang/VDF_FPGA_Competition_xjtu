module xpb_5_585
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4ac7e7a6618a0df520c2360931ffcffeb4aa7fcc35b2f6cb7170ee02ee1017f11318f1e8f1940f2ba17482554d2cf63dd124ef12f1a99ed54e89b048fd5ec1454c7903b2d9752300d429c1271ffe3f8d6be4635264e2f734da7bd9a7e2a04a8ebf69b81f45077d3a7fbb667203db9e1b1a0993cc88c75ec54fb3f5c2198a37c1;
    5'b00010 : xpb = 1024'h958fcf4cc3141bea41846c1263ff9ffd6954ff986b65ed96e2e1dc05dc202fe22631e3d1e3281e5742e904aa9a59ec7ba249de25e3533daa9d136091fabd828a98f20765b2ea4601a853824e3ffc7f1ad7c8c6a4c9c5ee69b4f7b34fc540951d7ed3703e8a0efa74ff76cce407b73c3634132799118ebd8a9f67eb8433146f82;
    5'b00011 : xpb = 1024'h2faa719d62aff51697412a4485a528aaac897c33cba143ead67610b3172d9acb360258420a95aef444ff47b90428d1ef0f54a552b24a0c343afdd17cbd49cf1e711bd669dcce6bbd69e340d2c71efa774fa8305ea222b88dd9e6fafcedb63d1a0f3596341e4d7f21f8724c7713c2b427ff42dc834a0abf1fa8ac6641c3bc40d8;
    5'b00100 : xpb = 1024'h7a725943c43a030bb803604db7a4f8a96133fc0001543ab647e6feb6053db2bc491b4a2afc29be1fe673ca0e5155c82ce0799465a3f3ab09898781c5baa89063bd94da1cb6438ebe3e0d01f9e71d3a04bb8c93b10705afc2b462d4a4d05687a8ce9f4e536354fc5c782db2e9179e5243194c704fd2d21de4f8605c03dd467899;
    5'b00101 : xpb = 1024'h148cfb9463d5dc380dc01e7fd94a8156a468789b618f910a3b7b3363404b1da558ebbe9b23974ebce88a0d1cbb24ada04d845b9272ea79932771f2b07d34dcf795bea920e027b479ff9cc07e6e3fb561336bfd6adf6279e6d9521c51f8cc2fa55f017448f79381097129327c23a9ca34e47c253a0b4e1f7a01a4d6c16dee49ef;
    5'b00110 : xpb = 1024'h5f54e33ac55fea2d2e8254890b4a51555912f867974287d5acec21662e5b35966c04b084152b5de889fe8f720851a3de1ea94aa56494186875fba2f97a939e3ce237acd3b99cd77ad3c681a58e3df4ee9f5060bd4445711bb3cdf5f9db6c7a341e6b2c683c9afe43f0e498ee2785684ffe85b90694157e3f5158cc83877881b0;
    5'b00111 : xpb = 1024'haa1ccae126e9f8224f448a923d4a21540dbd7833ccf57ea11e5d0f691c6b4d877f1da26d06bf6d142b7311c7557e9a1befce39b8563db73dc485534277f25f822eb0b0869311fa7ba7f042ccae3c347c0b34c40fa92868508e49cfa1be0cc4c2ddd4e48781a27b7e709fff602b61066b188f4cd31cdcdd04a10cc245a102b971;
    5'b01000 : xpb = 1024'h44376d31c685d14ea50148c45eefaa0150f1f4cf2d30d4f511f144165778b8708eee16dd2e2cfdb12d8954d5bf4d7f8f5cd900e5253485c7626fc42d3a7eac1606da7f8abcf6203769800151355eafd883142dc981853274b339174ee6826cbf6e370a7d15e1002b699b7ef3376c7e5ce3bf01bd5558de99aa513d0331aa8ac7;
    5'b01001 : xpb = 1024'h8eff54d8280fdf43c5c37ecd90ef7a00059c749b62e3cbc0836232194588d061a20708c61fc10cdccefdd72b0c7a75cd2dfdeff816de249cb0f9747637dd6d5b5353833d966b43383da9c278555cef65eef8911be66829a98db4f0f6c922b74e2da0c29c5ae87d65e956e5653b481c77fdc89589de203d5efa0532c54b34c288;
    5'b01010 : xpb = 1024'h2919f728c7abb8701b803cffb29502ad48d0f136c31f221476f666c680963b4ab1d77d36472e9d79d1141a3976495b409b08b724e5d4f3264ee3e560fa69b9ef2b7d5241c04f68f3ff3980fcdc7f6ac266d7fad5bec4f3cdb2a438a3f1985f4abe02e891ef270212e25264f847539469c8f84a74169c3ef40349ad82dbdc93de;
    5'b01011 : xpb = 1024'h73e1decf2935c6653c427308e494d2abfd7b7102f8d218dfe86754c96ea6533bc4f06f1f38c2aca572889c8ec376517e6c2da637d77e91fb9d6d95a9f7c87b3477f655f499c48bf4d3634223fc7daa4fd2bc5e2823a7eb028d20124bd438a9d97d6ca0b1342e7f4d620dcb6a4b2f3284e301de409f639db952fda344f566cb9f;
    5'b01100 : xpb = 1024'hdfc811fc8d19f9191ff313b063a5b5940afed9e590d6f33dbfb8976a9b3be24d4c0e38f60303d42749edf9d2d4536f1d9386d64a67560853b580694ba54c7c8502024f8c3a8b1b094f300a883a025ac4a9bc7e1fc04b526b20f59f8fcae51d60dcec6a6c86d03fa5b094afd573aaa76ae31932ad7df9f4e5c421e02860e9cf5;
    5'b01101 : xpb = 1024'h58c468c62a5bad86b2c16744383a2b57f55a6d6a8ec065ff4d6c777997c3d615e7d9d57851c44c6e161361f27a722d2faa5d5c77981eff5a89e1b6ddb7b3890d9c9928ab9d1dd4b1691cc1cfa39e6539b6802b3460e7ac5b8c8b33a0df4e9c64cd387ec60d748134dac4b16f5b164891c83b26f760a6fe13abf613c49f98d4b6;
    5'b01110 : xpb = 1024'ha38c506c8be5bb7bd3839d4d6a39fb56aa04ed36c4735ccabedd657c85d3ee06faf2c76143585b99b787e447c79f236d7b824b8a89c89e2fd86b6726b5124a52e9122c5e7692f7b23d4682f6c39ca4c722648e86c5caa39067070d48c1eee6f38ca236e5527bfe6f5a8017e15ef1e6ace244bac3e96e5cd8fbaa0986b9230c77;
    5'b01111 : xpb = 1024'h3da6f2bd2b8194a829405b7f8bdf8403ed3969d224aeb31eb2719a29c0e158f00ac33bd16ac5ec36b99e2756316e08e0e88d12b758bf6cb97655d811779e96e6c13bfb62a0771d6dfed6417b4abf20239a43f8409e276db48bf654f5ea648ef01d045cdae6ba831c537b97746afd5e9ead746fae21ea5e6e04ee844449caddcd;
    5'b10000 : xpb = 1024'h886eda638d0ba29d4a029188bddf5402a1e3e99e5a61a9ea23e2882caef170e11ddc2dba5c59fb625b12a9ab7e9aff1eb9b201ca4a690b8ec4df885a74fd582c0db4ff1579ec406ed30002a26abd5fb106285b93030a64e966722e9dcd04d97edc6e14fa2bc20056d336fde66ed8fcb9c77e037aaab1bd3354a27a066355158e;
    5'b10001 : xpb = 1024'h22897cb42ca77bc99fbf4fbadf84dcafe5186639ba9d003e1776bcd9e9fedbca2daca22a83c78bff5d28ecb9e869e49226bcc8f7195fda1862c9f9453789a4bfe5dece19a3d0662a948fc126f1dfdb0d7e07c54cdb672f0d8b61764af57a817b6cd03aefc0008503cc327d797ae474ab92adb864e32dbec85de6f4c3f3fce6e4;
    5'b10010 : xpb = 1024'h6d51645a8e3189bec08185c41184acae99c2e605f04ff70988e7aadcd80ef3bb40c59413755b9b2afe9d6f0f3596dacff7e1b80a0b0978edb153a98e34e866053257d1cc7d45892b68b9824e11de1a9ae9ec289f404a264265dd4ff2d81acc0a2c39f30f0508023e4bede3eb7ec012c6acb74c316bf51d8dad9aea860d871ea5;
    5'b10011 : xpb = 1024'h76c06ab2dcd62eb163e43f6332a355bdcf762a1508b4d5d7c7bdf8a131c5ea4509608839cc92bc800b3b21d9f65c04364ec7f36da0047774f3e1a78f774b2990a81a0d0a729aee72a4940d2990095f761cb925918a6f0668acc97a000907406bc9c1904994686eb44e9637e8acb8ab877e7011ba4711f22b6df65439e2eeffb;
    5'b10100 : xpb = 1024'h5233ee518f5770e0370079ff652a055a91a1e26d863e4428edeccd8d012c769563aefa6c8e5d3af3a2283472ec92b68136116e49cba9e64c9dc7cac1f4d373de56faa483809ed1e7fe7301f9b8fed584cdaff5ab7d89e79b65487147e330be957c05d123de4e0425c4a4c9f08ea728d391f094e82d387de806935b05b7b927bc;
    5'b10101 : xpb = 1024'h9cfbd5f7f0e17ed557c2b0089729d559464c6239bbf13af45f5dbb8fef3c8e8676c7ec557ff14a1f439cb6c839bfacbf07365d5cbd538521ec517b0af2323523a373a8365a13f4e8d29cc320d8fd1512399458fde26cded03fc44aefc5d109243b6f894323558160446030629282c6eeabfa28b4b5ffdcad564750c7d1435f7d;
    5'b10110 : xpb = 1024'h37167848907d5801ad7f6e3ab8cf5e068980ded51c2c914852f1f03d2a49f96f869860c5a75edabc45b2f9d6a38e9232744124898c4a53ab8a3bebf5b4be81b77b9d773a83f81aa4942c81a5601f906eb173c2b7bac9a8f464b3929cee46b120cbd1af38b794060d3d5baff59e8e3ee07729dd9eee7bde425f8bcb8561eb30d3;
    5'b10111 : xpb = 1024'h81de5feef20765f6ce41a443eacf2e053e2b5ea151df8813c462de40185a116099b152ae98f2e9e7e7277c2bf0bb88704566139c7df3f280d8c59c3eb21d42fcc8167aed5d6d3da5685642cc801dcffc1d58260a1faca0293f2f6c44d0e6fbaf8b3b6757fc9b8347bd171667a269dcfb9133716b77433d07af3fc1477b756894;
    5'b11000 : xpb = 1024'h1bf9023f91a33f2323fe62760c74b6b2815fdb3cb21ade67b7f712ed53677c49a981c71ec0607a84e93dbf3a5a8a6de3b270dac94ceac10a76b00d2974a98f90a04049f18751636129e6015107404b5895378fc3f8096a4d641eb3f1f95ca3ac1b9d8d4d90da07f4b61295faae7554ed5c632655afbf3e9cb8843c050c1d39ea;
    5'b11001 : xpb = 1024'h66c0e9e5f32d4d1844c0987f3e7486b1360a5b08e7cdd533296800f04177943abc9ab907b1f489b08ab2418fa7b764218395c9dc3e945fdfc539bd72720850d5ecb94da460c68661fe0fc278273e8ae6011bf3165cec61823e9a8d99dbfcee3adb07456cd5e1852f35cdfc6cb250f308766cba2238869d62083831c725a771ab;
    5'b11010 : xpb = 1024'hdb8c3692c926449a7d56b1601a0f5e793ed7a448092b871cfc359d7c84ff23cc6b2d77d9621a4d8cc8849e11864994f0a091090d8b2e6963242e5d34949d69c4e31ca88aaaac1dbf9f80fcae61064278fb5cd035492ba66389d547047296376b696b626a2009dc2ec97bffbe5c6afa419c6f0c71029ef7117cac84b64f4301;
    5'b11011 : xpb = 1024'h4ba373dcf4533439bb3f8cba9219df5d2de957707dbc22528e6d23a06a951714df841f60caf629792e3d06f35eb33fd2c1c5801bff34cd3eb1addea631f35eaf115c205b641fcf1e93c94223ce5f45cfe4dfc0229a2c22db3e05aeeee712e0c62ad32381af278716ae84e271c23809155ba602d8f9c9fdbc6130a246cfd97ac2;
    5'b11100 : xpb = 1024'h966b5b8355dd422edc01c2c3c419af5be293d73cb36f191dffde11a358a52f05f29d1149bc8a38a4cfb18948abe0361092ea6f2ef0de6c1400378eef2f521ff45dd5240e3d94f21f67f3034aee5d855d50c42374ff0f1a1018818896c9b32b54ea3cdba0f42f04512e4048e3c613a73075af96a582915c81b0e49808e963b283;
    5'b11101 : xpb = 1024'h3085fdd3f5791b5b31be80f5e5bf380925c853d813aa6f71f372465093b299ef026d85b9e3f7c941d1c7cc5715af1b83fff5365bbfd53a9d9e21ffd9f1de6c8835fef312677917db2982c1cf758000b9c8a38d2ed76be4343d70d043f228d3517a9f0196886d88fe273bc876d21f1f2240df4b8fbb0d5e16ba2912c67a0b83d9;
    5'b11110 : xpb = 1024'h7b4de57a570329505280b6ff17bf0807da72d3a4495d663d64e3345381c2b1e0158677a2d58bd86d733c4eac62dc11c1d11a256eb17ed972ecabb022ef3d2dcd8277f6c540ee3adbfdac82f6957e40473487f0813c4edb6917eca9ebd4c91de03a08b9b5cd750638a6f72ee8d5fabd3d5ae8df5c43d4bcdc09dd08889395bb9a;
    5'b11111 : xpb = 1024'h156887caf69f027ca83d7531396490b51da7503fa998bc9158776900bcd01cc92556ec12fcf9690a755291baccaaf7353e24ec9b8075a7fc8a96210db1c97a615aa1c5c96ad26097bf3c417b1ca0bba3ac675a3b14aba58d3cdbf198fd3ec5dcca6adfab61b38ae59ff2ae7be206352f261894467c50be7113218346243d8cf0;
    endcase
end

endmodule

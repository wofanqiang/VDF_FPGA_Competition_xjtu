module xpb_5_330
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha620cc228543c0f559af9117027e95becaee920d6b0a17169a9722fd877256972d1cb9f829baf9caf0d16417850559c13f66df35712865b9ffa5155029314f37f8b8b7b8a66384b838be1d63f4a5c0aa4e80f52b390d85c486f679613e21da6cb5b421107fe35852bb09331b9725352576d68f0d31f72bb6a6a8e803d21a3993;
    5'b00010 : xpb = 1024'h9b9452ef48994d21e859aa56f4a2e42c246720ea009c8db5b7518ca55be2002656f0f677894f7507424488e826aca2b81ab39684bf9dfb284eaaeb42179029be7d223ac29d360c2b5ee23825506fbd23a8fcf0bde594de78586060c7c21912473c60aff74efdb817ef527f58367a44219ed33f3813a2fa3d06e255031b520cbb;
    5'b00011 : xpb = 1024'h9107d9bc0beed94e7703c396e6c732997ddfafc6962f0454d40bf64d3051a9b580c532f6e8e3f04393b7adb8c853ebaef6004dd40e1390969db0c13405ef0445018bbdcc9408939e850652e6ac39b99d0378ec50921c372c29ca482e46104a21c30d3ede1e1817dd239bcb94d5cf531dc6cfef62f54ec8c3671bc2026489dfe3;
    5'b00100 : xpb = 1024'h867b6088cf44657b05addcd6d8eb8106d7583ea32bc17af3f0c65ff504c15344aa996f7648786b7fe52ad28969fb34a5d14d05235c892604ecb69725f44ddecb85f540d68adb1b11ab2a6da80803b6165df4e7e33ea38fdffb342f94ca0781fc49b9cdc4ed3277a257e517d175246219eecc9f8dd6fa9749c7552f01adc1b30b;
    5'b00101 : xpb = 1024'h7beee7559299f1a79457f616cb0fcf7430d0cd7fc153f1930d80c99cd930fcd3d46dabf5a80ce6bc369df75a0ba27d9cac99bc72aafebb733bbc6d17e2acb9520a5ec3e081ada284d14e886963cdb28fb870e375eb2ae893cc9e16fb4dfeb9d6d0665cabbc4cd7678c2e640e1479711616c94fb8b8a665d0278e9c00f6f98633;
    5'b00110 : xpb = 1024'h71626e2255ef7dd423020f56bd341de18a495c5c56e668322a3b3344ada0a662fe41e87507a161f888111c2aad49c69387e673c1f97450e18ac24309d10b93d88ec846ea788029f7f772a32abf97af0912ecdf0897b241479e07fe61d1f5f1b15712eb928b67372cc077b04ab3ce80123ec5ffe39a52345687c809004031595b;
    5'b00111 : xpb = 1024'h66d5f4ef19450a00b1ac2896af586c4ee3c1eb38ec78ded146f59cec82104ff2281624f46735dd34d98440fb4ef10f8a63332b1147e9e64fd9c818fbbf6a6e5f1331c9f46f52b16b1d96bdec1b61ab826d68da9b443999fb6f71e5c855ed298bddbf7a795a8196f1f4c0fc8753238f0e66c2b00e7bfe02dce80175ff89692c83;
    5'b01000 : xpb = 1024'h5c497bbbdc9a962d405641d6a17cbabc3d3a7a15820b557063b00694567ff98151ea6173c6ca58712af765cbf09858813e7fe260965f7bbe28cdeeedadc948e5979b4cfe662538de43bad8ad772ba7fbc7e4d62df0c0f2af40dbcd2ed9e46166646c0960299bf6b7290a48c3f2789e0a8ebf60395da9d163483ae2fed2a0ffab;
    5'b01001 : xpb = 1024'h51bd02889ff02259cf005b1693a1092996b308f2179dcc0f806a703c2aefa3107bbe9df3265ed3ad7c6a8a9c923fa17819cc99afe4d5112c77d3c4df9c28236c1c04d0085cf7c05169def36ed2f5a4752260d1c09d484b631245b4955ddb9940eb189846f8b6567c5d53950091cdad06b6bc10643f559fe9a8744ffe1bd8d2d3;
    5'b01010 : xpb = 1024'h473089556345ae865daa745685c55796f02b97cead3042ae9d24d9e3ff5f4c9fa592da7285f34ee9cdddaf6d33e6ea6ef51950ff334aa69ac6d99ad18a86fdf2a06e531253ca47c490030e302ebfa0ee7cdccd5349cfa416e3af9bfbe1d2d11b71c5272dc7d0b641919ce13d3122bc02deb8c08f21016e7008adbcfd6510a5fb;
    5'b01011 : xpb = 1024'h3ca41022269b3ab2ec548d9677e9a60449a426ab42c2b94db9df438bd3cef62ecf6716f1e587ca261f50d43dd58e3365d066084e81c03c0915df70c378e5d87924d7d61c4a9ccf37b62728f18a899d67d758c8e5f656fccab519836265ca08f5f871b61496eb1606c5e62d79d077caff06b570ba02ad3cf668e729fcae487923;
    5'b01100 : xpb = 1024'h321796eee9f0c6df7afea6d66a0df471a31cb587d8552fecd699ad33a83e9fbdf93b5371451c456270c3f90e77357c5cabb2bf9dd035d17764e546b56744b2ffa9415926416f56aadc4b43b2e65399e131d4c478a2de557e86836ac8e9c140d07f1e44fb660575cbfa2f79b66fccd9fb2eb220e4e4590b7cc92096fbf7804c4b;
    5'b01101 : xpb = 1024'h278b1dbbad46530c09a8c0165c3242defc9544646de7a68bf35416db7cae494d230f8ff0a4b0c09ec2371ddf18dcc55386ff76ed1eab66e5b3eb1ca755a38d862daadc303841de1e026f5e74421d965a8c50c00b4f65ae3257ed522f6db878ab05cad3e2351fd5912e78c5f30f21e8f756aed10fc604da03295a03fb40b81f73;
    5'b01110 : xpb = 1024'h1cfea488709bdf389852d9564e56914c560dd341037a1d2b100e8083511df2dc4ce3cc7004453bdb13aa42afba840e4a624c2e3c6d20fc5402f0f2994402680cb2145f3a2f146591289379359de792d3e6ccbb9dfbed06e629573995f1afb0858c7762c9043a355662c2122fae76f7f37eab813aa7b0a889899370fa89eff29b;
    5'b01111 : xpb = 1024'h12722b5533f16b6526fcf296407adfb9af86621d990c93ca2cc8ea2b258d9c6b76b808ef63d9b717651d67805c2b57413d98e58bbb9691c251f6c88b32614293367de24425e6ed044eb793f6f9b18f4d4148b730a8745f99fac120fc75a6e8601323f1afd354951b970b5e6c4dcc06efa6a83165895c770fe9ccddf9d327c5c3;
    5'b10000 : xpb = 1024'h7e5b221f746f791b5a70bd6329f2e2708fef0fa2e9f0a69498353d2f9fd45faa08c456ec36e3253b6908c50fdd2a03818e59cdb0a0c2730a0fc9e7d20c01d19bae7654e1cb9747774dbaeb8557b8bc69bc4b2c354fbb84dcc2b0862f99e203a99d08096a26ef4e0cb54aaa8ed2115ebcea4e1906b0845964a064af91c5f98eb;
    5'b10001 : xpb = 1024'hae067e447c8ab8870f569ced351dc3e5d3ed830799a9217fe41a76d0816f9c91cda8ff66ed292c1ea761f06882d7f9f9584c7c107b348ceaa0a1b3cd49f16c51b3a01d06c31cf92fad99cc1c4a214c70ea45a7ee8e093e12532181c437bffaa74f84a1a722524d33865dddc484464b11457b709d9cff714cf0af32fcee79d27e;
    5'b10010 : xpb = 1024'ha37a05113fe044b39e00b62d274212532d6611e42f3b981f00d4e07855df4620f77d3be64cbda75af8d51539247f42f03399335fc9aa2258efa789bf385046d83809a010b9ef80a2d3bde6dda5eb48ea44c1a3813a9096c6248b692abbb73281d631308df16cacf8baa72a01239b5a0d6d7820c87eab3fd350e89ffc37b1a5a6;
    5'b10011 : xpb = 1024'h98ed8bde0335d0e02caacf6d196660c086dea0c0c4ce0ebe1d8f4a202a4eefb021517865ac5222974a483a09c6268be70ee5eaaf181fb7c73ead5fb126af215ebc73231ab0c20815f9e2019f01b545639f3d9f13e717ef79f5f550913fae6a5c5cddbf74c0870cbdeef0763dc2f069099574d0f360570e59b1220cfb80e978ce;
    5'b10100 : xpb = 1024'h8e6112aac68b5d0cbb54e8ad0b8aaf2de0572f9d5a60855d3a49b3c7febe993f4b25b4e50be69dd39bbb5eda67cdd4ddea32a1fe66954d358db335a3150dfbe540dca624a7948f8920061c605d7f41dcf9b99aa6939f482dc75f37f7c3a5a236e38a4e5b8fa16c832339c27a62457805bd71811e4202dce0115b79faca214bf6;
    5'b10101 : xpb = 1024'h83d4997789e0e93949ff01ecfdaefd9b39cfbe79eff2fbfc57041d6fd32e42ce74f9f1646b7b190fed2e83ab09751dd4c57f594db50ae2a3dcb90b95036cd66bc546292e9e6716fc462a3721b9493e56543596394026a0e198c91f5e479cda116a36dd425ebbcc4857830eb7019a8701e56e314923aeab667194e6fa13591f1e;
    5'b10110 : xpb = 1024'h794820444d367565d8a91b2cefd34c0893484d568585729b73be8717a79dec5d9ece2de3cb0f944c3ea1a87bab1c66cba0cc109d038078122bbee186f1cbb0f249afac3895399e6f6c4e51e315133acfaeb191cbecadf9956a3306c4cb9411ebf0e36c292dd62c0d8bcc5af3a0ef95fe0d6ae174055a79ecd1ce53f95c90f246;
    5'b10111 : xpb = 1024'h6ebba711108c01926753346ce1f79a75ecc0dc331b17e93a9078f0bf7c0d95ecc8a26a632aa40f889014cd4c4cc3afc27c18c7ec51f60d807ac4b778e02a8b78ce192f428c0c25e292726ca470dd3749092d8d5e993552493b9cee2b4f8b49c6778ffb0ffcf08bd2c015a7304044a4fa3567919ee70648733207c0f8a5c8c56e;
    5'b11000 : xpb = 1024'h642f2dddd3e18dbef5fd4dacd41be8e346396b0fb0aa5fd9ad335a67507d3f7bf276a6e28a388ac4e187f21cee6af8b957657f3ba06ba2eec9ca8d6ace8965ff5282b24c82dead55b8968765cca733c263a988f145bcaafd0d06d591d38281a0fe3c89f6cc0aeb97f45ef36cdf99b3f65d6441c9c8b216f992412df7ef009896;
    5'b11001 : xpb = 1024'h59a2b4aa973719eb84a766ecc64037509fb1f9ec463cd678c9edc40f24ece90b1c4ae361e9cd060132fb16ed901241b032b2368aeee1385d18d0635cbce84085d6ec355679b134c8debaa2272871303bbe258483f24403b0de70bcf85779b97b84e918dd9b254b5d28a83fa97eeec2f28560f1f4aa5de57ff27a9af738386bbe;
    5'b11010 : xpb = 1024'h4f163b775a8ca6181351802cb86485bdf92a88c8dbcf4d17e6a82db6f95c929a461f1fe14961813d846e3bbe31b98aa70dfeedda3d56cdcb67d6394eab471b0c5b55b8607083bc3c04debce8843b2cb518a180169ecb5c64afdaa45edb70f1560b95a7c46a3fab225cf18be61e43d1eead5da21f8c09b40652b407f681703ee6;
    5'b11011 : xpb = 1024'h4489c2441de23244a1fb996caa88d42b52a317a57161c3b70362975ecdcc3c296ff35c60a8f5fc79d5e1608ed360d39de94ba5298bcc6339b6dc0f4099a5f592dfbf3b6a675643af2b02d7a9e005292e731d7ba94b52b51881448bc55f682930924236ab395a0ae7913ad822bd98e0ead55a524a6db5828cb2ed74f5caa8120e;
    5'b11100 : xpb = 1024'h39fd4910e137be7130a5b2ac9cad2298ac1ba68206f43a56201d0106a23be5b899c798e0088a77b62754855f75081c94c4985c78da41f8a805e1e5328804d0196428be745e28cb225126f26b3bcf25a7cd99773bf7da0dcc52ae732be35f610b18eec59208746aacc584245f5cedefe6fd5702754f6151131326e1f513dfe536;
    5'b11101 : xpb = 1024'h2f70cfdda48d4a9dbf4fcbec8ed171060594355e9c86b0f53cd76aae76ab8f47c39bd55f681ef2f278c7aa3016af658b9fe513c828b78e1654e7bb247663aa9fe892417e54fb5295774b0d2c97992221281572cea461668024185a92675698e59f9b5478d78eca71f9cd709bfc42fee32553b2a0310d1f9973604ef45d17b85e;
    5'b11110 : xpb = 1024'h24e456aa67e2d6ca4df9e52c80f5bf735f0cc43b321927945991d4564b1b38d6ed7011dec7b36e2eca3acf00b856ae827b31cb17772d2384a3ed911664c285266cfbc4884bcdda089d6f27edf3631e9a82916e6150e8bf33f58241f8eb4dd0c02647e35fa6a92a372e16bcd89b980ddf4d5062cb12b8ee1fd399bbf3a64f8b86;
    5'b11111 : xpb = 1024'h1a57dd772b3862f6dca3fe6c731a0de0b8855317c7ab9e33764c3dfe1f8ae26617444e5e2747e96b1badf3d159fdf779567e8266c5a2b8f2f2f3670853215facf165479242a0617bc39342af4f2d1b13dd0d69f3fd7017e7c6ec295f6f45089aacf4724675c389fc626009153aed1cdb754d12f5f464bca633d328f2ef875eae;
    endcase
end

endmodule

module xpb_5_495
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6cf1ecd3d6723fc74f4bd09f15edf490a7cfd9b208032a50e3c52d149f9da032bc142f8c3214631df6b26053e7fbf84547dd82ce43d2bfd8a8241db1e520530062e658635d72b7b72790fa61976da63da759a4ded9555b1794737acbed88d90c3286e75c783c922027e2419b1b52ce36df44f8ea874da095807bf1f0badf6d70;
    5'b00010 : xpb = 1024'h29369451eaf64ac5d39229671b81a1cfde29b0333a8eb42a49ada0d38c38935d74dfe19f9a0247ad4e068160ec99dfc02ba0ddb664f2af659fa8fc058f6e314f517d7c180b5472293c87f22095ff884a5aae50252624891e735a639d20e70f8636063c8f3fb02bb2c9049c573ed576446fb012f2be4fe3faba8868dcecdc7475;
    5'b00011 : xpb = 1024'h96288125c1688a8d22ddfa06316f966085f989e54291de7b2d72cde82bd6339030f4112bcc16aacb44b8e1b4d495d805737e6084a8c56f3e47cd19b7748e844fb463d47b68c729e06418ec822d6d2e880207f503ff79e43607cdde690e6fe892688d23ebb7ecbdd2f0e6ddf25a28447b4ef50bdd459d84903b045acda7bbe1e5;
    5'b00100 : xpb = 1024'h526d28a3d5ec958ba72452ce3703439fbc536066751d6854935b41a7187126bae9bfc33f34048f5a9c0d02c1d933bf805741bb6cc9e55ecb3f51f80b1edc629ea2faf83016a8e452790fe4412bff1094b55ca04a4c49123ce6b4c73a41ce1f0c6c0c791e7f605765920938ae7daaec88df6025e57c9fc7f57510d1b9d9b8e8ea;
    5'b00101 : xpb = 1024'heb1d021ea70a08a2b6aab963c96f0def2ad36e7a7a8f22df943b566050c19e5a28b75529bf273e9f36123ceddd1a6fb3b051654eb054e5836d6d65ec92a40ed91921be4c48a9ec48e06dc002a90f2a168b14b9099184043c59bb00b752c55866f8bce5146d3f0f8332b936aa12d94966fcb3fedb3a20b5aaf1d48a60bb5efef;
    5'b00110 : xpb = 1024'h7ba3bcf5c0e2e0517ab67c355284e56f9a7d1099afac1c7edd08e27aa4a9ba185e9fa4dece06d707ea138422c5cd9f4082e299232ed80e30defaf410ae4a93edf478744821fd567bb597d661c1fe98df100af06f726d9b5b5a0f2ad762b52e92a212b5adbf1083185b0dd505bc8062cd4f1038d83aefabf02f993a96c6955d5f;
    5'b00111 : xpb = 1024'h37e86473d566eb4ffefcd4fd581892aed0d6e71ae237a65842f156399144ad43176b56f235f4bb974167a52fca6b86bb66a5f40b4ff7fdbdd67fd2645898723ce30f97fccfdf10edca8ece20c0907aebc35f9bb5bf3cc96238f613a89613650ca5920ae086841caafc302fc1e0030adadf7b52e071f1ef5569a5b182f8926464;
    5'b01000 : xpb = 1024'ha4da5147abd92b174e48a59c6e06873f78a6c0ccea3ad0a926b6834e30e24d75d37f867e68091eb5381a0583b2677f00ae8376d993cabd967ea3f0163db8c53d45f5f0602d51c8a4f21fc88257fe21296ab9409498922479cd698e74839c3e18d818f23cfec0aecb2412715cfb55d911bec04bcaf93f8feaea21a373b371d1d4;
    5'b01001 : xpb = 1024'h611ef8c5c05d3615d28efe64739a347eaf00974e1cc65a828c9ef70d1d7d40a08c4b3891cff703448f6e2690b705667b9246d1c1b4eaad237628ce69e806a38c348d1414db3383170716c041569003361e0debdae5615280ac507745b6fa7492db98476fc634485dc534cc191ed8811f4f2b65d33041d350242e1a5fe56ed8d9;
    5'b01010 : xpb = 1024'h1d63a043d4e1411456d5572c792de1bde55a6dcf4f51e45bf2876acc0a1833cb4516eaa537e4e7d3e6c2479dbba34df6760a2ca9d60a9cb06dadacbd925481db232437c989153d891c0db8005521e542d1629721323080878b376016ea58ab0cdf179ca28da7e1f0665726d5425b292cdf967fdb674416b55e3a914c176bdfde;
    5'b01011 : xpb = 1024'h8a558d17ab5380dba62127cb8f1bd64e8d2a478157550eacd64c97e0a9b5d3fe012b1a3169f94af1dd74a7f1a39f463bbde7af7819dd5c8915d1ca6f7774d4db860a902ce687f540439eb261ec8f8b8078bc3c000b85db9f1faadae2d7e18419119e83ff05e474108e3968705dadf763bedb78c5ee91b74adeb6833cd24b4d4e;
    5'b01100 : xpb = 1024'h469a3495bfd78bda2a67809394af838dc3841e0289e098863c350b9f9650c728b9f6cc44d1e72f8134c8c8fea83d2db6a1ab0a603afd4c160d56a8c321c2b32a74a1b3e19469afb25895aa20eb216d8d2c10e746585509a5fe91c3b40b3fba93151dd931cd580da32f5bc32c81309f714f4692ce2593fab018c2fa2904485453;
    5'b01101 : xpb = 1024'h2dedc13d45b96d8aeadd95b9a4330ccf9ddf483bc6c225fa21d7f5e82ebba5372c27e5839d514108c1cea0bacdb1531856e65485c1d3ba304db8716cc1091796338d796424b6a246d8ca1dfe9b34f99df65928ca52437acdd78ac853e9df10d189d2e6494cba735d07e1de8a4b3477edfb1acd65c963e1552cf711536455b58;
    5'b01110 : xpb = 1024'h6fd0c8e7aacdd69ffdf9a9fab031255da1adce35c46f4cb085e2ac7322895a862ed6ade46be9772e82cf4a5f94d70d76cd4be8169feffb7bacffa4c8b130e479c61f2ff99fbe21db951d9c418120f5d786bf376b7e7992c471ec27512c26ca194b2415c10d083955f8605f83c00615b5bef6a5c0e3e3deaad34b6305f124c8c8;
    5'b01111 : xpb = 1024'h2c157065bf51e19e824002c2b5c4d29cd807a4b6f6fad689ebcb20320f244db0e7a25ff7d3d75bbdda236b6c9974f4f1b10f42fec10feb08a484831c5b7ec2c8b4b653ae4d9fdc4daa1494007fb2d7e43a13e2b1cb48c0cb50d310225f8500934ea36af3d47bd2e89982ba3fe388bdc34f61bfc91ae622100d57d9f22321cfcd;
    5'b10000 : xpb = 1024'h99075d3995c42165d18bd361cbb2c72d7fd77e68fefe00dacf904d46aec1ede3a3b68f8405ebbedbd0d5cbc08170ed36f8ecc5cd04e2aae14ca8a0ce409f15c9179cac11ab129404d1a58e6217207e21e16d8790a49e1be2e5468aee4d0dd99f812a52504cb86508c164fbdafedb8bfa2ea6b8b3a233c2a58dd3cbe2de013d3d;
    5'b10001 : xpb = 1024'h554c04b7aa482c6455d22c29d146746cb63154ea31898ab43578c1059b5ce10e5c8241976dd9a36b2829eccd860ed4b1dcb020b526029a6e442d7f21eaecf4180633cfc658f44e76e69c862115b2602e94c232d6f16d49e9c42d73bf806c101984a9a783142bfe9b62875697225e3407bf11d2bbd936060ac7e042cf0ffe4442;
    5'b10010 : xpb = 1024'h1190ac35becc3762da1884f1d6da21abec8b2b6b6415148d9b6134c487f7d439154df3aad5c787fa7f7e0dda8aacbc2cc0737b9d472289fb3bb25d75953ad266f4caf37b06d608e8fb937de01444423b4816de1d3e3c77f0a3145c90b3ca46938828fcb5db9f982e03a9b15345e0dc154f7cecc41038497001ecb9bb41fb4b47;
    5'b10011 : xpb = 1024'h7e829909953e772a29645590ecc8163c945b051d6c183ede7f2661d92795746bd162233707dbeb1876306e2e72a8b4720850fe6b8af549d3e3d67b277a5b256757b14bde6448c0a023247841abb1e878ef7082fc1791d3083787d75ca1531f9fbaafe41253dc2a4e2b8bf2ee6133aa4c2ec1e5ae9785ea058268ababfcdab8b7;
    5'b10100 : xpb = 1024'h3ac74087a9c28228adaaae58f25bc37bcab4db9e9ea3c8b7e50ed598143067968a2dd54a6fc9cfa7cd848f3b77469becec145953ac153960db5b597b24a903b646486f93122a7b12381b7000aa43ca85a2c52e426461010f166ec02dd4b15619be2f39451b4fc3e0ccae4daa84b65259bf2cffb6ce882d6abc7522982ed7bfbc;
    5'b10101 : xpb = 1024'ha7b92d5b8034c1effcf67ef80849b80c7284b550a6a6f308c8d402acb3ce07c9464204d6a1de32c5c436ef8f5f42943233f1dc21efe7f939837f772d09c956b6a92ec7f66f9d32c95fac6a6241b170c34a1ed3213db65c26aae23af9c23a2f25f0b620a1938c5600f4908f45a00920909e71f8a155d5ce003cf11488e9b72d2c;
    5'b10110 : xpb = 1024'h63fdd4d994b8ccee813cd7c00ddd654ba8de8bd1d9327ce22ebc766ba068faf3ff0db6ea09cc17551b8b109c63e07bad17b5370a1107e8c67b045580b417350597c5ebab1d7eed3b74a36221404352cffd737e678a858a2d89c923caf598659ff43575d45affef9395b2ea01c38bc89e2edd12a98cd8116576fd8b751bb43431;
    5'b10111 : xpb = 1024'h20427c57a93cd7ed058330881371128adf3862530bbe06bb94a4ea2a8d03ee1eb7d968fd71b9fbe472df31a9687e6327fb7891f23227d853728933d45e651354865d0f5fcb60a7ad899a59e03ed534dcb0c829add754b83468b00c9c28f69c19f7b4cb072273892636d544bde70e70abbf482cb1c3da54cab10a02614db13b36;
    5'b11000 : xpb = 1024'h8d34692b7faf17b454cf0127295f071b87083c0513c1310c786a173f2ca18e5173ed9889a3ce5f02699191fd507a5b6d435614c075fa982c1aad518643856654e94367c328d35f64b12b5441d642db1a5821ce8cb0aa134bfd238768167f75262a3bb2639ab01b465eb7865902613ee29e8d259c4b27f5603185f4520890a8a6;
    5'b11001 : xpb = 1024'h497910a9943322b2d91559ef2ef2b45abd621286464cbae5de528afe193c817c2cb94a9d0bbc4391c0e5b30a551842e827196fa8971a87b912322fd9edd344a3d7da8b77d6b519d6c6224c00d4d4bd270b7679d2fd794152dc0a703949ddaba02dbb07966223b4d8ffd9e11525e3e6f02ef83fa4822a38c56b926b3e3a8dafab;
    5'b11010 : xpb = 1024'h5bdb827a8b72db15d5bb2b734866199f3bbe90778d844bf443afebd05d774a6e584fcb073aa28211839d41759b62a630adcca90b83a774609b70e2d982122f2c671af2c8496d448db1943bfd3669f33becb25194a486f59baf1590a7d3be21a313a5cc929974e6ba0fc3bd149668efdbf6359acb92c7c2aa59ee22a6c8ab6b0;
    5'b11011 : xpb = 1024'h72afa4fb7f296d78aca783564a74562a9b8bc2b980db6f1028002bd1a57514d9a1992c3ca5be8b3f0eec346b41b222a852ba4d5efc0d371eb1db2bdf7d4175f32958078fe2098c0002aa3e216ad445716624c9f8239dca714f64d3d66ac4bb2663c14425a1d3e08bc8de7d6c64b95d349ea85297407a1cc0261ad41b276a2420;
    5'b11100 : xpb = 1024'h2ef44c7993ad787730eddc1e50080369d1e5993ab366f8e98de89f90921008045a64de500dac6fce6640557846500a23367da8471d2d26aba9600a33278f544217ef2b448feb467217a135e06966277e1979753e706cf8782e4bbca79e22f1a06740995869477a1e6a00d828883c05422f136c9f777c602560274b0759672b25;
    5'b11101 : xpb = 1024'h9be6394d6a1fb83e8039acbd65f5f7fa79b572ecbb6a233a71adcca531ada83716790ddc3fc0d2ec5cf2b5cc2e4c02687e5b2b1560ffe684518427e50cafa7427ad583a7ed5dfe293f32304200d3cdbbc0d31a1d49c2538fc2bf37738babcaac99c780b4e1840c3e91e319c3a38ed3790e586589feca00bae0a33cf814469895;
    5'b11110 : xpb = 1024'h582ae0cb7ea3c33d048005856b89a539b00f496dedf5ad13d79640641e489b61cf44bfefa7aeb77bb446d6d932e9e9e3621e85fd821fd61149090638b6fd8591696ca75c9b3fb89b54292800ff65afc87427c56396918196a1a62044bf0a01269d46d5e7a8f7a5d13305747fc7117b869ec37f9235cc44201aafb3e446439f9a;
    5'b11111 : xpb = 1024'h146f88499327ce3b88c65e4d711d5278e6691fef208136ed3d7eb4230ae38e8c881072030f9c9c0b0b9af7e63787d15e45e1e0e5a33fc59e408de48c614b63e05803cb114921730d69201fbffdf791d5277c70a9e360af9d808d0915f26837a0a0c62b1a706b3f63d427cf3bea9423942f2e999a6cce878554bc2ad07840a69f;
    endcase
end

endmodule

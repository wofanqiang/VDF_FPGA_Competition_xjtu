module xpb_5_460
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2cda3ef69c54ec927df3a3977efb458b1cb825d713fd78462e089e6b2ae94569a0683aef9893fa0ad23797c2c20ca716fe17c8cb3932f4d5707c2866c1498b3b5ddea50ff185678088e967d821048907cada0795ef7b38237ad4f14288cde4eeb2dafbcc6c3bf449acee4854f45bae44f0fa849c7094ebcd5d811ef0f2a9029;
    5'b00010 : xpb = 1024'h59b47ded38a9d924fbe7472efdf68b1639704bae27faf08c5c113cd655d28ad340d075df3127f415a46f2f8584194e2dfc2f91967265e9aae0f850cd82931676bbbd4a1fe30acf0111d2cfb04209120f95b40f2bdef67046f5a9e285119bc9dd65b5f798d877e89359dc90a9e8b75c89e1f50938e129d79abb023de1e552052;
    5'b00011 : xpb = 1024'h868ebce3d4fec5b779daeac67cf1d0a1562871853bf868d28a19db4180bbd03ce138b0cec9bbee2076a6c7484625f544fa475a61ab98de805174793443dca1b2199bef2fd49036819abc3788630d9b17608e16c1ce71a86a707ed3c79a69aecc1890f36544b3dcdd06cad8fedd130aced2ef8dd551bec36818835cd2d7fb07b;
    5'b00100 : xpb = 1024'hb368fbda7153b249f7ce8e5dfbed162c72e0975c4ff5e118b82279acaba515a681a0ebbe624fe82b48de5f0b08329c5bf85f232ce4cbd355c1f0a19b05262ced777a943fc6159e0223a59f608412241f2b681e57bdece08deb53c50a233793bacb6bef31b0efd126b3b92153d16eb913c3ea1271c253af3576047bc3caa40a4;
    5'b00101 : xpb = 1024'he0433ad10da89edc75c231f57ae85bb78f98bd3363f3595ee62b1817d68e5b10220926adfae3e2361b15f6cdca3f4372f676ebf81dfec82b326cca01c66fb828d559394fb79b0582ac8f0738a516ad26f64225edad6818b16628b64cac0578a97e46eafe1d2bc57060a769a8c5ca6758b4e4970e32e89b02d3859ab4bd4d0cd;
    5'b00110 : xpb = 1024'h10d1d79c7a9fd8b6ef3b5d58cf9e3a142ac50e30a77f0d1a51433b6830177a079c271619d9377dc40ed4d8e908c4bea89f48eb4c35731bd00a2e8f26887b943643337de5fa9206d0335786f10c61b362ec11c2d839ce350d4e0fda78f34d35d983121e6ca8967b9ba0d95b1fdba26159da5df1baaa37d86d03106b9a5aff60f6;
    5'b00111 : xpb = 1024'h139f7b8be4652780171a9792478dee6cdc90908e18bee49eb423c54ee2c60e5e362d99c8d2c0bd64bbf8526534e5891a0f2a67d8e9064b1d613651acf4902ce9f9116836f9aa5d483be61d6e8e71fbf368bf635198c5e88f85bd298d1bda14286e3fce296f5a3ae03ba83fa52ae81c3e296d9a0471412729d8e87d896a29f11f;
    5'b01000 : xpb = 1024'h166d1f7b4e2a76493ef9d1cbbf7da2c58e5c12eb89febc2317044f359574a2b4d0341d77cc49fd05691bcbe16106538b7f0be4659c997a6ab83e143360a4c59daeef5287f8c2b3c04474b3ec10824483e56d03caf7bd9c11bd6a78a14466f277596d7de6361dfa24d677242a7a2dd722787d424e384a75e6aec08f7879548148;
    5'b01001 : xpb = 1024'h193ac36ab7efc51266d90c05376d571e40279548fb3e93a779e4d91c4823370b6a3aa126c5d33ca6163f455d8d271dfceeed60f2502ca9b80f45d6b9ccb95e5164cd3cd8f7db0a384d034a6992928d14621aa44456b54f93f517c7b56cf3d0c6449b2da2fce1b969714608afc9739206c78cea97ff53c4a38498a167887f1171;
    5'b01010 : xpb = 1024'h1c08675a21b513db8eb8463eaf5d0b76f1f317a66c7e6b2bdcc56302fad1cb62044124d5bf5c7c46c362bed9b947e86e5ecedd7f03bfd905664d994038cdf7051aab2729f6f360b05591e0e714a2d5a4dec844bdb5ad03162cc516c99580af152fc8dd5fc3a578ae0c14ed3518b94ceb169c92e1c65d13605a70b35697a9a19a;
    5'b01011 : xpb = 1024'h1ed60b498b7a62a4b6978078274cbfcfa3be9a03ddbe42b03fa5ece9ad805fb89e47a884b8e5bbe770863855e568b2dfceb05a0bb7530852bd555bc6a4e28fb8d089117af60bb7285e20776496b31e355b75e53714a4b698647265ddbe0d8d641af68d1c8a6937f2a6e3d1ba67ff07cf65ac3b2b8d66621d3048c545a6d431c3;
    5'b01100 : xpb = 1024'h21a3af38f53fb16dde76bab19f3c7428558a1c614efe1a34a28676d0602ef40f384e2c33b26efb881da9b1d211897d513e91d6986ae637a0145d1e4d10f7286c8666fbcbf5240da066af0de218c366c5d82385b0739c6a1a9c1fb4f1e69a6bb306243cd9512cf73741b2b63fb744c2b3b4bbe375546fb0da0620d734b5fec1ec;
    5'b01101 : xpb = 1024'h247153285f0500370655f4eb172c288107559ebec03df1b9056700b712dd8865d254afe2abf83b28cacd2b4e3daa47c2ae7353251e7966ed6b64e0d37d0bc1203c44e61cf43c64186f3da45f9ad3af5654d12629d2941d9cd3cd04060f274a01f151ec9617f0b67bdc819ac5068a7d9803cb8bbf1b78ff96dbf8e923c5295215;
    5'b01110 : xpb = 1024'h273ef717c8ca4f002e352f248f1bdcd9b921211c317dc93d68478a9dc58c1cbc6c5b3391a5817ac977f0a4ca69cb12341e54cfb1d20c963ac26ca359e92059d3f222d06df354ba9077cc3add1ce3f7e6d17ec6a3318bd11f0b7a531a37b42850dc7f9c52deb475c077507f4a55d0387c52db3408e2824e53b1d0fb12d453e23e;
    5'b01111 : xpb = 1024'h2a0c9b07328f9dc95614695e070b91326aeca379a2bda0c1cb281484783ab1130661b7409f0aba6a25141e4695ebdca58e364c3e859fc588197465e05534f287a800babef26d1108805ad15a9ef440774e2c671c908384a14327a22e6041069fc7ad4c0fa5783505121f63cfa515f360a1eadc52a98b9d1087a90d01e37e7267;
    5'b10000 : xpb = 1024'h2cda3ef69c54ec927df3a3977efb458b1cb825d713fd78462e089e6b2ae94569a0683aef9893fa0ad23797c2c20ca716fe17c8cb3932f4d5707c2866c1498b3b5ddea50ff185678088e967d821048907cada0795ef7b38237ad4f14288cde4eeb2dafbcc6c3bf449acee4854f45bae44f0fa849c7094ebcd5d811ef0f2a90290;
    5'b10001 : xpb = 1024'h2fa7e2e6061a3b5ba5d2ddd0f6eaf9e3ce83a834853d4fca90e92851dd97d9c03a6ebe9e921d39ab7f5b113eee2d71886df94557ecc62422c783eaed2d5e23ef13bc8f60f09dbdf89177fe55a314d1984787a80f4e72eba5b2824056b15ac33d9e08ab8932ffb38e47bd2cda43a16929400a2ce6379e3a8a335930e001d392b9;
    5'b10010 : xpb = 1024'h327586d56fdf8a24cdb2180a6edaae3c804f2a91f67d274ef3c9b23890466e16d475424d8ba6794c2c7e8abb1a4e3bf9dddac1e4a05953701e8bad739972bca2c99a79b1efb614709a0694d325251a28c4354888ad6a9f27ea2f8f6ad9e7a18c89365b45f9c372d2e28c115f92e7240d8f19d52ffea78947093142cf10fe22e2;
    5'b10011 : xpb = 1024'h35432ac4d9a4d8edf5915243e6ca6295321aacef67bcfed356aa3c1f42f5026d6e7bc5fc852fb8ecd9a20437466f066b4dbc3e7153ec82bd75936ffa058755567f786402eece6ae8a2952b50a73562b940e2e9020c6252aa21dcde7f02747fdb74640b02c08732177d5af5e4e22cdef1de297d79c5b0d803df0954be2028b30b;
    5'b10100 : xpb = 1024'h3810ceb4436a27b71d708c7d5eba16ede3e62f4cd8fcd657b98ac605f5a396c4088249ab7eb8f88d86c57db3728fd0dcbd9dbafe077fb20acc9b3280719bee0a35564e53ede6c160ab23c1ce2945ab49bd90897b6b5a062c598a2d932b015e2a5f91babf874af15c1829da6a317299d62d3925c38cba26c0b4e166ad2f534334;
    5'b10101 : xpb = 1024'h3ade72a3ad2f7680454fc6b6d6a9cb4695b1b1aa4a3caddc1c6b4feca8522b1aa288cd5a7842382e33e8f72f9eb09b4e2d7f378abb12e15823a2f506ddb086bdeb3438a4ecff17d8b3b2584bab55f3da3a3e29f4ca51b9ae91377ca7538e3c794abf6a7c4e0eb0a0b2f8beef80b854ba7c48ce0d53c3757d8ab9789c3e7dd35d;
    5'b10110 : xpb = 1024'h3dac169316f4c5496d2f00f04e997f9f477d3407bb7c85607f4bd9d35b00bf713c8f510971cb77cee10c70abcad165bf9d60b4176ea610a57aaab78d49c51f71a11222f5ec176e50bc40eec92d663c6ab6ebca6e29496d30c8e4cbbb7c1b1ac835ed1a3914d26fe54dc7a374cffe0f9ecb5876571accc43a60918a8b4da86386;
    5'b10111 : xpb = 1024'h4079ba8280ba1412950e3b29c68933f7f948b6652cbc5ce4e22c63ba0daf53c7d695d4b86b54b76f8e2fea27f6f230310d4230a422393ff2d1b27a13b5d9b82556f00d46eb2fc4c8c4cf8546af7684fb33996ae7884120b300921acfa4a7f917211ac9f5db962f29e89687fa1f43ca831a681ea0e1d612f736699c7a5cd2f3af;
    5'b11000 : xpb = 1024'h43475e71ea7f62dbbced75633e78e850ab1438c29dfc3469450ceda0c05de81e709c586764ddf7103b5363a42312faa27d23ad30d5cc6f4028ba3c9a21ee50d90ccdf797ea481b40cd5e1bc43186cd8bb0470b60e738d435383f69e3cd34d7660c4879b2a259ee6e83656c7f6e8985676977c6eaa8df61b40c41ae696bfd83d8;
    5'b11001 : xpb = 1024'h461502615444b1a4e4ccaf9cb6689ca95cdfbb200f3c0beda7ed7787730c7c750aa2dc165e6736b0e876dd204f33c513ed0529bd895f9e8d7fc1ff208e02e98cc2abe1e8e96071b8d5ecb241b397161c2cf4abda463087b76fecb8f7f5c1b5b4f776296f691dadb31e345104bdcf404bb8876f346fe8b070e219c0587b281401;
    5'b11010 : xpb = 1024'h48e2a650be0a006e0cabe9d62e5851020eab3d7d807be3720ace016e25bb10cba4a95fc557f07651959a569c7b548f855ce6a64a3cf2cddad6c9c1a6fa1782407889cc39e878c830de7b48bf35a75eaca9a24c53a5283b39a79a080c1e4e9403e2a3d92c2fe16cf7b903358a0d14fb300797177e36f1ff2db7f1d2478a52a42a;
    5'b11011 : xpb = 1024'h4bb04a4027cf4f37348b240fa648055ac076bfdaf1bbbaf66dae8b54d869a5223eafe3745179b5f242bdd018a77559f6ccc822d6f085fd282dd1842d662c1af42e67b68ae7911ea8e709df3cb7b7a73d264feccd041feebbdf47572046db7252cdd188e8f6a52c3c53d21a0f5c5ab61456a6bfc7fdfb4dea8dc9e436997d3453;
    5'b11100 : xpb = 1024'h4e7dee2f91949e005c6a5e491e37b9b37242423862fb927ad08f153b8b183978d8b667234b02f592efe14994d39624683ca99f63a4192c7584d946b3d240b3a7e445a0dbe6a97520ef9875ba39c7efcda2fd8d466317a23e16f4a6346f6850a1b8ff38a5bd68eb80eea0fe94aba070f8a5b66811c5049ca763a1f625a8a7c47c;
    5'b11101 : xpb = 1024'h514b921efb59ecc98449988296276e0c240dc495d43b69ff336f9f223dc6cdcf72bcead2448c35339d04c310ffb6eed9ac8b1bf057ac5bc2dbe1093a3e554c5b9a238b2ce5c1cb98f8270c37bbd8385e1fab2dbfc20f55c04ea1f54897f52ef0a42ce862842caac5896fe319fae62bdcf4c6105b8c0deb64397a0814b7d254a5;
    5'b11110 : xpb = 1024'h5419360e651f3b92ac28d2bc0e172264d5d946f3457b418396502908f07562260cc36e813e1574d44a283c8d2bd7b94b1c6c987d0b3f8b1032e8cbc0aa69e50f5001757de4da221100b5a2b53de880ee9c58ce3921070942864f445cc0820d3f8f5a981f4af06a0a243ec79f4a2be6c143d5b8a553173a210f521a03c6fce4ce;
    5'b11111 : xpb = 1024'h56e6d9fdcee48a5bd4080cf58606d6bd87a4c950b6bb1907f930b2efa323f67ca6c9f230379eb474f74bb60957f883bc8c4e1509bed2ba5d89f08e47167e7dc305df5fcee3f2788909443932bff8c97f19066eb27ffebcc4bdfc9370e90eeb8e7a8847dc11b4294ebf0dac249971a1a592e560ef1a2088dde52a2bf2d62774f7;
    endcase
end

endmodule

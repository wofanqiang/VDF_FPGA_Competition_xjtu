module xpb_1024
(
    input [1023:0] data_in, 

    output [1023:0] data_out_0,
    output [1023:0] data_out_1,
    output [1023:0] data_out_2,
    output [1023:0] data_out_3,
    output [1023:0] data_out_4,
    output [1023:0] data_out_5,
    output [1023:0] data_out_6,
    output [1023:0] data_out_7,
    output [1023:0] data_out_8,
    output [1023:0] data_out_9,
    output [1023:0] data_out_10,
    output [1023:0] data_out_11,
    output [1023:0] data_out_12,
    output [1023:0] data_out_13,
    output [1023:0] data_out_14,
    output [1023:0] data_out_15,
    output [1023:0] data_out_16,
    output [1023:0] data_out_17,
    output [1023:0] data_out_18,
    output [1023:0] data_out_19,
    output [1023:0] data_out_20,
    output [1023:0] data_out_21,
    output [1023:0] data_out_22,
    output [1023:0] data_out_23,
    output [1023:0] data_out_24,
    output [1023:0] data_out_25,
    output [1023:0] data_out_26,
    output [1023:0] data_out_27,
    output [1023:0] data_out_28,
    output [1023:0] data_out_29,
    output [1023:0] data_out_30,
    output [1023:0] data_out_31,
    output [1023:0] data_out_32,
    output [1023:0] data_out_33,
    output [1023:0] data_out_34,
    output [1023:0] data_out_35,
    output [1023:0] data_out_36,
    output [1023:0] data_out_37,
    output [1023:0] data_out_38,
    output [1023:0] data_out_39,
    output [1023:0] data_out_40,
    output [1023:0] data_out_41,
    output [1023:0] data_out_42,
    output [1023:0] data_out_43,
    output [1023:0] data_out_44,
    output [1023:0] data_out_45,
    output [1023:0] data_out_46,
    output [1023:0] data_out_47,
    output [1023:0] data_out_48,
    output [1023:0] data_out_49,
    output [1023:0] data_out_50,
    output [1023:0] data_out_51,
    output [1023:0] data_out_52,
    output [1023:0] data_out_53,
    output [1023:0] data_out_54,
    output [1023:0] data_out_55,
    output [1023:0] data_out_56,
    output [1023:0] data_out_57,
    output [1023:0] data_out_58,
    output [1023:0] data_out_59,
    output [1023:0] data_out_60,
    output [1023:0] data_out_61,
    output [1023:0] data_out_62,
    output [1023:0] data_out_63,
    output [1023:0] data_out_64,
    output [1023:0] data_out_65,
    output [1023:0] data_out_66,
    output [1023:0] data_out_67,
    output [1023:0] data_out_68,
    output [1023:0] data_out_69,
    output [1023:0] data_out_70,
    output [1023:0] data_out_71,
    output [1023:0] data_out_72,
    output [1023:0] data_out_73,
    output [1023:0] data_out_74,
    output [1023:0] data_out_75,
    output [1023:0] data_out_76,
    output [1023:0] data_out_77,
    output [1023:0] data_out_78,
    output [1023:0] data_out_79,
    output [1023:0] data_out_80,
    output [1023:0] data_out_81,
    output [1023:0] data_out_82,
    output [1023:0] data_out_83,
    output [1023:0] data_out_84,
    output [1023:0] data_out_85,
    output [1023:0] data_out_86,
    output [1023:0] data_out_87,
    output [1023:0] data_out_88,
    output [1023:0] data_out_89,
    output [1023:0] data_out_90,
    output [1023:0] data_out_91,
    output [1023:0] data_out_92,
    output [1023:0] data_out_93,
    output [1023:0] data_out_94,
    output [1023:0] data_out_95,
    output [1023:0] data_out_96,
    output [1023:0] data_out_97,
    output [1023:0] data_out_98,
    output [1023:0] data_out_99,
    output [1023:0] data_out_100,
    output [1023:0] data_out_101,
    output [1023:0] data_out_102,
    output [1023:0] data_out_103,
    output [1023:0] data_out_104,
    output [1023:0] data_out_105,
    output [1023:0] data_out_106,
    output [1023:0] data_out_107,
    output [1023:0] data_out_108,
    output [1023:0] data_out_109,
    output [1023:0] data_out_110,
    output [1023:0] data_out_111,
    output [1023:0] data_out_112,
    output [1023:0] data_out_113,
    output [1023:0] data_out_114,
    output [1023:0] data_out_115,
    output [1023:0] data_out_116,
    output [1023:0] data_out_117,
    output [1023:0] data_out_118,
    output [1023:0] data_out_119,
    output [1023:0] data_out_120,
    output [1023:0] data_out_121,
    output [1023:0] data_out_122,
    output [1023:0] data_out_123,
    output [1023:0] data_out_124,
    output [1023:0] data_out_125,
    output [1023:0] data_out_126,
    output [1023:0] data_out_127,
    output [1023:0] data_out_128,
    output [1023:0] data_out_129,
    output [1023:0] data_out_130,
    output [1023:0] data_out_131,
    output [1023:0] data_out_132,
    output [1023:0] data_out_133,
    output [1023:0] data_out_134,
    output [1023:0] data_out_135,
    output [1023:0] data_out_136,
    output [1023:0] data_out_137,
    output [1023:0] data_out_138,
    output [1023:0] data_out_139,
    output [1023:0] data_out_140,
    output [1023:0] data_out_141,
    output [1023:0] data_out_142,
    output [1023:0] data_out_143,
    output [1023:0] data_out_144,
    output [1023:0] data_out_145,
    output [1023:0] data_out_146,
    output [1023:0] data_out_147,
    output [1023:0] data_out_148,
    output [1023:0] data_out_149,
    output [1023:0] data_out_150,
    output [1023:0] data_out_151,
    output [1023:0] data_out_152,
    output [1023:0] data_out_153,
    output [1023:0] data_out_154,
    output [1023:0] data_out_155,
    output [1023:0] data_out_156,
    output [1023:0] data_out_157,
    output [1023:0] data_out_158,
    output [1023:0] data_out_159,
    output [1023:0] data_out_160,
    output [1023:0] data_out_161,
    output [1023:0] data_out_162,
    output [1023:0] data_out_163,
    output [1023:0] data_out_164,
    output [1023:0] data_out_165,
    output [1023:0] data_out_166,
    output [1023:0] data_out_167,
    output [1023:0] data_out_168,
    output [1023:0] data_out_169,
    output [1023:0] data_out_170,
    output [1023:0] data_out_171,
    output [1023:0] data_out_172,
    output [1023:0] data_out_173,
    output [1023:0] data_out_174,
    output [1023:0] data_out_175,
    output [1023:0] data_out_176,
    output [1023:0] data_out_177,
    output [1023:0] data_out_178,
    output [1023:0] data_out_179,
    output [1023:0] data_out_180,
    output [1023:0] data_out_181,
    output [1023:0] data_out_182,
    output [1023:0] data_out_183,
    output [1023:0] data_out_184,
    output [1023:0] data_out_185,
    output [1023:0] data_out_186,
    output [1023:0] data_out_187,
    output [1023:0] data_out_188,
    output [1023:0] data_out_189,
    output [1023:0] data_out_190,
    output [1023:0] data_out_191,
    output [1023:0] data_out_192,
    output [1023:0] data_out_193,
    output [1023:0] data_out_194,
    output [1023:0] data_out_195,
    output [1023:0] data_out_196,
    output [1023:0] data_out_197,
    output [1023:0] data_out_198,
    output [1023:0] data_out_199,
    output [1023:0] data_out_200,
    output [1023:0] data_out_201,
    output [1023:0] data_out_202,
    output [1023:0] data_out_203,
    output [1023:0] data_out_204

);





xpb_5_0  u_xpb_5_0 (
.data_in( data_in[4 : 0]),
.data_out(data_out_0)
);

xpb_5_5  u_xpb_5_5 (
.data_in( data_in[9 : 5]),
.data_out(data_out_1)
);

xpb_5_10  u_xpb_5_10 (
.data_in( data_in[14 : 10]),
.data_out(data_out_2)
);

xpb_5_15  u_xpb_5_15 (
.data_in( data_in[19 : 15]),
.data_out(data_out_3)
);

xpb_5_20  u_xpb_5_20 (
.data_in( data_in[24 : 20]),
.data_out(data_out_4)
);

xpb_5_25  u_xpb_5_25 (
.data_in( data_in[29 : 25]),
.data_out(data_out_5)
);

xpb_5_30  u_xpb_5_30 (
.data_in( data_in[34 : 30]),
.data_out(data_out_6)
);

xpb_5_35  u_xpb_5_35 (
.data_in( data_in[39 : 35]),
.data_out(data_out_7)
);

xpb_5_40  u_xpb_5_40 (
.data_in( data_in[44 : 40]),
.data_out(data_out_8)
);

xpb_5_45  u_xpb_5_45 (
.data_in( data_in[49 : 45]),
.data_out(data_out_9)
);

xpb_5_50  u_xpb_5_50 (
.data_in( data_in[54 : 50]),
.data_out(data_out_10)
);

xpb_5_55  u_xpb_5_55 (
.data_in( data_in[59 : 55]),
.data_out(data_out_11)
);

xpb_5_60  u_xpb_5_60 (
.data_in( data_in[64 : 60]),
.data_out(data_out_12)
);

xpb_5_65  u_xpb_5_65 (
.data_in( data_in[69 : 65]),
.data_out(data_out_13)
);

xpb_5_70  u_xpb_5_70 (
.data_in( data_in[74 : 70]),
.data_out(data_out_14)
);

xpb_5_75  u_xpb_5_75 (
.data_in( data_in[79 : 75]),
.data_out(data_out_15)
);

xpb_5_80  u_xpb_5_80 (
.data_in( data_in[84 : 80]),
.data_out(data_out_16)
);

xpb_5_85  u_xpb_5_85 (
.data_in( data_in[89 : 85]),
.data_out(data_out_17)
);

xpb_5_90  u_xpb_5_90 (
.data_in( data_in[94 : 90]),
.data_out(data_out_18)
);

xpb_5_95  u_xpb_5_95 (
.data_in( data_in[99 : 95]),
.data_out(data_out_19)
);

xpb_5_100  u_xpb_5_100 (
.data_in( data_in[104 : 100]),
.data_out(data_out_20)
);

xpb_5_105  u_xpb_5_105 (
.data_in( data_in[109 : 105]),
.data_out(data_out_21)
);

xpb_5_110  u_xpb_5_110 (
.data_in( data_in[114 : 110]),
.data_out(data_out_22)
);

xpb_5_115  u_xpb_5_115 (
.data_in( data_in[119 : 115]),
.data_out(data_out_23)
);

xpb_5_120  u_xpb_5_120 (
.data_in( data_in[124 : 120]),
.data_out(data_out_24)
);

xpb_5_125  u_xpb_5_125 (
.data_in( data_in[129 : 125]),
.data_out(data_out_25)
);

xpb_5_130  u_xpb_5_130 (
.data_in( data_in[134 : 130]),
.data_out(data_out_26)
);

xpb_5_135  u_xpb_5_135 (
.data_in( data_in[139 : 135]),
.data_out(data_out_27)
);

xpb_5_140  u_xpb_5_140 (
.data_in( data_in[144 : 140]),
.data_out(data_out_28)
);

xpb_5_145  u_xpb_5_145 (
.data_in( data_in[149 : 145]),
.data_out(data_out_29)
);

xpb_5_150  u_xpb_5_150 (
.data_in( data_in[154 : 150]),
.data_out(data_out_30)
);

xpb_5_155  u_xpb_5_155 (
.data_in( data_in[159 : 155]),
.data_out(data_out_31)
);

xpb_5_160  u_xpb_5_160 (
.data_in( data_in[164 : 160]),
.data_out(data_out_32)
);

xpb_5_165  u_xpb_5_165 (
.data_in( data_in[169 : 165]),
.data_out(data_out_33)
);

xpb_5_170  u_xpb_5_170 (
.data_in( data_in[174 : 170]),
.data_out(data_out_34)
);

xpb_5_175  u_xpb_5_175 (
.data_in( data_in[179 : 175]),
.data_out(data_out_35)
);

xpb_5_180  u_xpb_5_180 (
.data_in( data_in[184 : 180]),
.data_out(data_out_36)
);

xpb_5_185  u_xpb_5_185 (
.data_in( data_in[189 : 185]),
.data_out(data_out_37)
);

xpb_5_190  u_xpb_5_190 (
.data_in( data_in[194 : 190]),
.data_out(data_out_38)
);

xpb_5_195  u_xpb_5_195 (
.data_in( data_in[199 : 195]),
.data_out(data_out_39)
);

xpb_5_200  u_xpb_5_200 (
.data_in( data_in[204 : 200]),
.data_out(data_out_40)
);

xpb_5_205  u_xpb_5_205 (
.data_in( data_in[209 : 205]),
.data_out(data_out_41)
);

xpb_5_210  u_xpb_5_210 (
.data_in( data_in[214 : 210]),
.data_out(data_out_42)
);

xpb_5_215  u_xpb_5_215 (
.data_in( data_in[219 : 215]),
.data_out(data_out_43)
);

xpb_5_220  u_xpb_5_220 (
.data_in( data_in[224 : 220]),
.data_out(data_out_44)
);

xpb_5_225  u_xpb_5_225 (
.data_in( data_in[229 : 225]),
.data_out(data_out_45)
);

xpb_5_230  u_xpb_5_230 (
.data_in( data_in[234 : 230]),
.data_out(data_out_46)
);

xpb_5_235  u_xpb_5_235 (
.data_in( data_in[239 : 235]),
.data_out(data_out_47)
);

xpb_5_240  u_xpb_5_240 (
.data_in( data_in[244 : 240]),
.data_out(data_out_48)
);

xpb_5_245  u_xpb_5_245 (
.data_in( data_in[249 : 245]),
.data_out(data_out_49)
);

xpb_5_250  u_xpb_5_250 (
.data_in( data_in[254 : 250]),
.data_out(data_out_50)
);

xpb_5_255  u_xpb_5_255 (
.data_in( data_in[259 : 255]),
.data_out(data_out_51)
);

xpb_5_260  u_xpb_5_260 (
.data_in( data_in[264 : 260]),
.data_out(data_out_52)
);

xpb_5_265  u_xpb_5_265 (
.data_in( data_in[269 : 265]),
.data_out(data_out_53)
);

xpb_5_270  u_xpb_5_270 (
.data_in( data_in[274 : 270]),
.data_out(data_out_54)
);

xpb_5_275  u_xpb_5_275 (
.data_in( data_in[279 : 275]),
.data_out(data_out_55)
);

xpb_5_280  u_xpb_5_280 (
.data_in( data_in[284 : 280]),
.data_out(data_out_56)
);

xpb_5_285  u_xpb_5_285 (
.data_in( data_in[289 : 285]),
.data_out(data_out_57)
);

xpb_5_290  u_xpb_5_290 (
.data_in( data_in[294 : 290]),
.data_out(data_out_58)
);

xpb_5_295  u_xpb_5_295 (
.data_in( data_in[299 : 295]),
.data_out(data_out_59)
);

xpb_5_300  u_xpb_5_300 (
.data_in( data_in[304 : 300]),
.data_out(data_out_60)
);

xpb_5_305  u_xpb_5_305 (
.data_in( data_in[309 : 305]),
.data_out(data_out_61)
);

xpb_5_310  u_xpb_5_310 (
.data_in( data_in[314 : 310]),
.data_out(data_out_62)
);

xpb_5_315  u_xpb_5_315 (
.data_in( data_in[319 : 315]),
.data_out(data_out_63)
);

xpb_5_320  u_xpb_5_320 (
.data_in( data_in[324 : 320]),
.data_out(data_out_64)
);

xpb_5_325  u_xpb_5_325 (
.data_in( data_in[329 : 325]),
.data_out(data_out_65)
);

xpb_5_330  u_xpb_5_330 (
.data_in( data_in[334 : 330]),
.data_out(data_out_66)
);

xpb_5_335  u_xpb_5_335 (
.data_in( data_in[339 : 335]),
.data_out(data_out_67)
);

xpb_5_340  u_xpb_5_340 (
.data_in( data_in[344 : 340]),
.data_out(data_out_68)
);

xpb_5_345  u_xpb_5_345 (
.data_in( data_in[349 : 345]),
.data_out(data_out_69)
);

xpb_5_350  u_xpb_5_350 (
.data_in( data_in[354 : 350]),
.data_out(data_out_70)
);

xpb_5_355  u_xpb_5_355 (
.data_in( data_in[359 : 355]),
.data_out(data_out_71)
);

xpb_5_360  u_xpb_5_360 (
.data_in( data_in[364 : 360]),
.data_out(data_out_72)
);

xpb_5_365  u_xpb_5_365 (
.data_in( data_in[369 : 365]),
.data_out(data_out_73)
);

xpb_5_370  u_xpb_5_370 (
.data_in( data_in[374 : 370]),
.data_out(data_out_74)
);

xpb_5_375  u_xpb_5_375 (
.data_in( data_in[379 : 375]),
.data_out(data_out_75)
);

xpb_5_380  u_xpb_5_380 (
.data_in( data_in[384 : 380]),
.data_out(data_out_76)
);

xpb_5_385  u_xpb_5_385 (
.data_in( data_in[389 : 385]),
.data_out(data_out_77)
);

xpb_5_390  u_xpb_5_390 (
.data_in( data_in[394 : 390]),
.data_out(data_out_78)
);

xpb_5_395  u_xpb_5_395 (
.data_in( data_in[399 : 395]),
.data_out(data_out_79)
);

xpb_5_400  u_xpb_5_400 (
.data_in( data_in[404 : 400]),
.data_out(data_out_80)
);

xpb_5_405  u_xpb_5_405 (
.data_in( data_in[409 : 405]),
.data_out(data_out_81)
);

xpb_5_410  u_xpb_5_410 (
.data_in( data_in[414 : 410]),
.data_out(data_out_82)
);

xpb_5_415  u_xpb_5_415 (
.data_in( data_in[419 : 415]),
.data_out(data_out_83)
);

xpb_5_420  u_xpb_5_420 (
.data_in( data_in[424 : 420]),
.data_out(data_out_84)
);

xpb_5_425  u_xpb_5_425 (
.data_in( data_in[429 : 425]),
.data_out(data_out_85)
);

xpb_5_430  u_xpb_5_430 (
.data_in( data_in[434 : 430]),
.data_out(data_out_86)
);

xpb_5_435  u_xpb_5_435 (
.data_in( data_in[439 : 435]),
.data_out(data_out_87)
);

xpb_5_440  u_xpb_5_440 (
.data_in( data_in[444 : 440]),
.data_out(data_out_88)
);

xpb_5_445  u_xpb_5_445 (
.data_in( data_in[449 : 445]),
.data_out(data_out_89)
);

xpb_5_450  u_xpb_5_450 (
.data_in( data_in[454 : 450]),
.data_out(data_out_90)
);

xpb_5_455  u_xpb_5_455 (
.data_in( data_in[459 : 455]),
.data_out(data_out_91)
);

xpb_5_460  u_xpb_5_460 (
.data_in( data_in[464 : 460]),
.data_out(data_out_92)
);

xpb_5_465  u_xpb_5_465 (
.data_in( data_in[469 : 465]),
.data_out(data_out_93)
);

xpb_5_470  u_xpb_5_470 (
.data_in( data_in[474 : 470]),
.data_out(data_out_94)
);

xpb_5_475  u_xpb_5_475 (
.data_in( data_in[479 : 475]),
.data_out(data_out_95)
);

xpb_5_480  u_xpb_5_480 (
.data_in( data_in[484 : 480]),
.data_out(data_out_96)
);

xpb_5_485  u_xpb_5_485 (
.data_in( data_in[489 : 485]),
.data_out(data_out_97)
);

xpb_5_490  u_xpb_5_490 (
.data_in( data_in[494 : 490]),
.data_out(data_out_98)
);

xpb_5_495  u_xpb_5_495 (
.data_in( data_in[499 : 495]),
.data_out(data_out_99)
);

xpb_5_500  u_xpb_5_500 (
.data_in( data_in[504 : 500]),
.data_out(data_out_100)
);

xpb_5_505  u_xpb_5_505 (
.data_in( data_in[509 : 505]),
.data_out(data_out_101)
);

xpb_5_510  u_xpb_5_510 (
.data_in( data_in[514 : 510]),
.data_out(data_out_102)
);

xpb_5_515  u_xpb_5_515 (
.data_in( data_in[519 : 515]),
.data_out(data_out_103)
);

xpb_5_520  u_xpb_5_520 (
.data_in( data_in[524 : 520]),
.data_out(data_out_104)
);

xpb_5_525  u_xpb_5_525 (
.data_in( data_in[529 : 525]),
.data_out(data_out_105)
);

xpb_5_530  u_xpb_5_530 (
.data_in( data_in[534 : 530]),
.data_out(data_out_106)
);

xpb_5_535  u_xpb_5_535 (
.data_in( data_in[539 : 535]),
.data_out(data_out_107)
);

xpb_5_540  u_xpb_5_540 (
.data_in( data_in[544 : 540]),
.data_out(data_out_108)
);

xpb_5_545  u_xpb_5_545 (
.data_in( data_in[549 : 545]),
.data_out(data_out_109)
);

xpb_5_550  u_xpb_5_550 (
.data_in( data_in[554 : 550]),
.data_out(data_out_110)
);

xpb_5_555  u_xpb_5_555 (
.data_in( data_in[559 : 555]),
.data_out(data_out_111)
);

xpb_5_560  u_xpb_5_560 (
.data_in( data_in[564 : 560]),
.data_out(data_out_112)
);

xpb_5_565  u_xpb_5_565 (
.data_in( data_in[569 : 565]),
.data_out(data_out_113)
);

xpb_5_570  u_xpb_5_570 (
.data_in( data_in[574 : 570]),
.data_out(data_out_114)
);

xpb_5_575  u_xpb_5_575 (
.data_in( data_in[579 : 575]),
.data_out(data_out_115)
);

xpb_5_580  u_xpb_5_580 (
.data_in( data_in[584 : 580]),
.data_out(data_out_116)
);

xpb_5_585  u_xpb_5_585 (
.data_in( data_in[589 : 585]),
.data_out(data_out_117)
);

xpb_5_590  u_xpb_5_590 (
.data_in( data_in[594 : 590]),
.data_out(data_out_118)
);

xpb_5_595  u_xpb_5_595 (
.data_in( data_in[599 : 595]),
.data_out(data_out_119)
);

xpb_5_600  u_xpb_5_600 (
.data_in( data_in[604 : 600]),
.data_out(data_out_120)
);

xpb_5_605  u_xpb_5_605 (
.data_in( data_in[609 : 605]),
.data_out(data_out_121)
);

xpb_5_610  u_xpb_5_610 (
.data_in( data_in[614 : 610]),
.data_out(data_out_122)
);

xpb_5_615  u_xpb_5_615 (
.data_in( data_in[619 : 615]),
.data_out(data_out_123)
);

xpb_5_620  u_xpb_5_620 (
.data_in( data_in[624 : 620]),
.data_out(data_out_124)
);

xpb_5_625  u_xpb_5_625 (
.data_in( data_in[629 : 625]),
.data_out(data_out_125)
);

xpb_5_630  u_xpb_5_630 (
.data_in( data_in[634 : 630]),
.data_out(data_out_126)
);

xpb_5_635  u_xpb_5_635 (
.data_in( data_in[639 : 635]),
.data_out(data_out_127)
);

xpb_5_640  u_xpb_5_640 (
.data_in( data_in[644 : 640]),
.data_out(data_out_128)
);

xpb_5_645  u_xpb_5_645 (
.data_in( data_in[649 : 645]),
.data_out(data_out_129)
);

xpb_5_650  u_xpb_5_650 (
.data_in( data_in[654 : 650]),
.data_out(data_out_130)
);

xpb_5_655  u_xpb_5_655 (
.data_in( data_in[659 : 655]),
.data_out(data_out_131)
);

xpb_5_660  u_xpb_5_660 (
.data_in( data_in[664 : 660]),
.data_out(data_out_132)
);

xpb_5_665  u_xpb_5_665 (
.data_in( data_in[669 : 665]),
.data_out(data_out_133)
);

xpb_5_670  u_xpb_5_670 (
.data_in( data_in[674 : 670]),
.data_out(data_out_134)
);

xpb_5_675  u_xpb_5_675 (
.data_in( data_in[679 : 675]),
.data_out(data_out_135)
);

xpb_5_680  u_xpb_5_680 (
.data_in( data_in[684 : 680]),
.data_out(data_out_136)
);

xpb_5_685  u_xpb_5_685 (
.data_in( data_in[689 : 685]),
.data_out(data_out_137)
);

xpb_5_690  u_xpb_5_690 (
.data_in( data_in[694 : 690]),
.data_out(data_out_138)
);

xpb_5_695  u_xpb_5_695 (
.data_in( data_in[699 : 695]),
.data_out(data_out_139)
);

xpb_5_700  u_xpb_5_700 (
.data_in( data_in[704 : 700]),
.data_out(data_out_140)
);

xpb_5_705  u_xpb_5_705 (
.data_in( data_in[709 : 705]),
.data_out(data_out_141)
);

xpb_5_710  u_xpb_5_710 (
.data_in( data_in[714 : 710]),
.data_out(data_out_142)
);

xpb_5_715  u_xpb_5_715 (
.data_in( data_in[719 : 715]),
.data_out(data_out_143)
);

xpb_5_720  u_xpb_5_720 (
.data_in( data_in[724 : 720]),
.data_out(data_out_144)
);

xpb_5_725  u_xpb_5_725 (
.data_in( data_in[729 : 725]),
.data_out(data_out_145)
);

xpb_5_730  u_xpb_5_730 (
.data_in( data_in[734 : 730]),
.data_out(data_out_146)
);

xpb_5_735  u_xpb_5_735 (
.data_in( data_in[739 : 735]),
.data_out(data_out_147)
);

xpb_5_740  u_xpb_5_740 (
.data_in( data_in[744 : 740]),
.data_out(data_out_148)
);

xpb_5_745  u_xpb_5_745 (
.data_in( data_in[749 : 745]),
.data_out(data_out_149)
);

xpb_5_750  u_xpb_5_750 (
.data_in( data_in[754 : 750]),
.data_out(data_out_150)
);

xpb_5_755  u_xpb_5_755 (
.data_in( data_in[759 : 755]),
.data_out(data_out_151)
);

xpb_5_760  u_xpb_5_760 (
.data_in( data_in[764 : 760]),
.data_out(data_out_152)
);

xpb_5_765  u_xpb_5_765 (
.data_in( data_in[769 : 765]),
.data_out(data_out_153)
);

xpb_5_770  u_xpb_5_770 (
.data_in( data_in[774 : 770]),
.data_out(data_out_154)
);

xpb_5_775  u_xpb_5_775 (
.data_in( data_in[779 : 775]),
.data_out(data_out_155)
);

xpb_5_780  u_xpb_5_780 (
.data_in( data_in[784 : 780]),
.data_out(data_out_156)
);

xpb_5_785  u_xpb_5_785 (
.data_in( data_in[789 : 785]),
.data_out(data_out_157)
);

xpb_5_790  u_xpb_5_790 (
.data_in( data_in[794 : 790]),
.data_out(data_out_158)
);

xpb_5_795  u_xpb_5_795 (
.data_in( data_in[799 : 795]),
.data_out(data_out_159)
);

xpb_5_800  u_xpb_5_800 (
.data_in( data_in[804 : 800]),
.data_out(data_out_160)
);

xpb_5_805  u_xpb_5_805 (
.data_in( data_in[809 : 805]),
.data_out(data_out_161)
);

xpb_5_810  u_xpb_5_810 (
.data_in( data_in[814 : 810]),
.data_out(data_out_162)
);

xpb_5_815  u_xpb_5_815 (
.data_in( data_in[819 : 815]),
.data_out(data_out_163)
);

xpb_5_820  u_xpb_5_820 (
.data_in( data_in[824 : 820]),
.data_out(data_out_164)
);

xpb_5_825  u_xpb_5_825 (
.data_in( data_in[829 : 825]),
.data_out(data_out_165)
);

xpb_5_830  u_xpb_5_830 (
.data_in( data_in[834 : 830]),
.data_out(data_out_166)
);

xpb_5_835  u_xpb_5_835 (
.data_in( data_in[839 : 835]),
.data_out(data_out_167)
);

xpb_5_840  u_xpb_5_840 (
.data_in( data_in[844 : 840]),
.data_out(data_out_168)
);

xpb_5_845  u_xpb_5_845 (
.data_in( data_in[849 : 845]),
.data_out(data_out_169)
);

xpb_5_850  u_xpb_5_850 (
.data_in( data_in[854 : 850]),
.data_out(data_out_170)
);

xpb_5_855  u_xpb_5_855 (
.data_in( data_in[859 : 855]),
.data_out(data_out_171)
);

xpb_5_860  u_xpb_5_860 (
.data_in( data_in[864 : 860]),
.data_out(data_out_172)
);

xpb_5_865  u_xpb_5_865 (
.data_in( data_in[869 : 865]),
.data_out(data_out_173)
);

xpb_5_870  u_xpb_5_870 (
.data_in( data_in[874 : 870]),
.data_out(data_out_174)
);

xpb_5_875  u_xpb_5_875 (
.data_in( data_in[879 : 875]),
.data_out(data_out_175)
);

xpb_5_880  u_xpb_5_880 (
.data_in( data_in[884 : 880]),
.data_out(data_out_176)
);

xpb_5_885  u_xpb_5_885 (
.data_in( data_in[889 : 885]),
.data_out(data_out_177)
);

xpb_5_890  u_xpb_5_890 (
.data_in( data_in[894 : 890]),
.data_out(data_out_178)
);

xpb_5_895  u_xpb_5_895 (
.data_in( data_in[899 : 895]),
.data_out(data_out_179)
);

xpb_5_900  u_xpb_5_900 (
.data_in( data_in[904 : 900]),
.data_out(data_out_180)
);

xpb_5_905  u_xpb_5_905 (
.data_in( data_in[909 : 905]),
.data_out(data_out_181)
);

xpb_5_910  u_xpb_5_910 (
.data_in( data_in[914 : 910]),
.data_out(data_out_182)
);

xpb_5_915  u_xpb_5_915 (
.data_in( data_in[919 : 915]),
.data_out(data_out_183)
);

xpb_5_920  u_xpb_5_920 (
.data_in( data_in[924 : 920]),
.data_out(data_out_184)
);

xpb_5_925  u_xpb_5_925 (
.data_in( data_in[929 : 925]),
.data_out(data_out_185)
);

xpb_5_930  u_xpb_5_930 (
.data_in( data_in[934 : 930]),
.data_out(data_out_186)
);

xpb_5_935  u_xpb_5_935 (
.data_in( data_in[939 : 935]),
.data_out(data_out_187)
);

xpb_5_940  u_xpb_5_940 (
.data_in( data_in[944 : 940]),
.data_out(data_out_188)
);

xpb_5_945  u_xpb_5_945 (
.data_in( data_in[949 : 945]),
.data_out(data_out_189)
);

xpb_5_950  u_xpb_5_950 (
.data_in( data_in[954 : 950]),
.data_out(data_out_190)
);

xpb_5_955  u_xpb_5_955 (
.data_in( data_in[959 : 955]),
.data_out(data_out_191)
);

xpb_5_960  u_xpb_5_960 (
.data_in( data_in[964 : 960]),
.data_out(data_out_192)
);

xpb_5_965  u_xpb_5_965 (
.data_in( data_in[969 : 965]),
.data_out(data_out_193)
);

xpb_5_970  u_xpb_5_970 (
.data_in( data_in[974 : 970]),
.data_out(data_out_194)
);

xpb_5_975  u_xpb_5_975 (
.data_in( data_in[979 : 975]),
.data_out(data_out_195)
);

xpb_5_980  u_xpb_5_980 (
.data_in( data_in[984 : 980]),
.data_out(data_out_196)
);

xpb_5_985  u_xpb_5_985 (
.data_in( data_in[989 : 985]),
.data_out(data_out_197)
);


xpb_5_990  u_xpb_5_990 (
.data_in( data_in[994 : 990]),
.data_out(data_out_198)
);

xpb_5_995  u_xpb_5_995 (
.data_in( data_in[999 : 995]),
.data_out(data_out_199)
);

xpb_5_1000  u_xpb_5_1000 (
.data_in( data_in[1004 : 1000]),
.data_out(data_out_200)
);

xpb_5_1005  u_xpb_5_1005 (
.data_in( data_in[1009 : 1005]),
.data_out(data_out_201)
);

xpb_5_1010  u_xpb_5_1010 (
.data_in( data_in[1014 : 1010]),
.data_out(data_out_202)
);

xpb_5_1015  u_xpb_5_1015 (
.data_in( data_in[1019 : 1015]),
.data_out(data_out_203)
);

xpb_4_1020  u_xpb_4_1020 (
.data_in( data_in[1023 : 1020]),
.data_out(data_out_204)
);

endmodule
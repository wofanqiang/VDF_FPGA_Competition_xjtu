module xpb_5_775
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6410ebc73fc41b38f6e7e6f7ee3643963b9d5c705b9a83f5c0bf5e5b1d7d5d3816d59ba4efff3e99a49077a184f2a1d65d050b1a649a90d40c546d0cfd0167397a07877fe96eb9fb6c233e3615cd94d30b8a8bb16ca60bdb824aff12bb9169719f4ceb9fa7baa561d76cad086f0d933d79e4f54e9d146a2a2ad7db57b66c8aee;
    5'b00010 : xpb = 1024'h17749238bd9a01a922ca5618cc123fdb05c4b5afe1bd677403a2036087f80d682a62b9d115d7fea4a9c2affc268732e255efee4ea682515c68099abbbf3059c17fbfda51234c76b1c5ac79c992bf657523101dca4cc5eaa64f096c2abcf830510f9245159eac523628197331e64b0051a4f00bbae9dd77240f403baae3f6af71;
    5'b00011 : xpb = 1024'h7b857dfffd5e1ce219b23d10ba488371416212203d57eb69c46161bba5756aa04138557605d73d3e4e53279dab79d4b8b2f4f9690b1ce230745e07c8bc31c0faf9c761d10cbb30ad31cfb7ffa88cfa482e9aa97bb96bf681d1546b3d788999c2aedf30b54666f797ff86203a5558938f1ed5010986f1e14e3a1817029a633a5f;
    5'b00100 : xpb = 1024'h2ee924717b3403524594ac3198247fb60b896b5fc37acee8074406c10ff01ad054c573a22baffd4953855ff84d0e65c4abdfdc9d4d04a2b8d01335777e60b382ff7fb4a24698ed638b58f393257ecaea46203b94998bd54c9e12d85579f060a21f248a2b3d58a46c5032e663cc9600a349e01775d3baee481e807755c7ed5ee2;
    5'b00101 : xpb = 1024'h92fa1038baf81e8b3c7c9329865ac34c4726c7d01f1552ddc803651c2d6d78086b9b0f471baf3be2f815d799d201079b08e4e7b7b19f338cdc67a2847b621abc79873c223007a75ef77c31c93b4c5fbd51aac7460631e128205dd7683581ca13be7175cae51349ce279f936c3ba393e0c3c50cc470cf5872495852ad7e59e9d0;
    5'b00110 : xpb = 1024'h465db6aa38ce04fb685f024a6436bf91114e210fa538365c0ae60a2197e828387f282d734187fbedfd480ff4739598a701cfcaebf386f415381cd0333d910d447f3f8ef369e5641551056d5cb83e305f6930595ee651bff2ed1c448036e890f32eb6cf40dc04f6a2784c5995b2e100f4eed02330bd98656c2dc0b300abe40e53;
    5'b00111 : xpb = 1024'haa6ea271789220345f46e942526d03274ceb7d8000d2ba51cba5687cb565857095fdc91831873a87a1d88795f8883a7d5ed4d606582184e944713d403a92747df947167353541e10bd28ab92ce0bc53274bae51052f7cbce6f674392f279fa64ce03bae083bf9c044fb9069e21ee943268b5187f5aaccf9658988e5862509941;
    5'b01000 : xpb = 1024'h5dd248e2f66806a48b2958633048ff6c1712d6bf86f59dd00e880d821fe035a0a98ae744575ffa92a70abff09a1ccb8957bfb93a9a094571a0266aeefcc16705feff69448d31dac716b1e7264afd95d48c4077293317aa993c25b0aaf3e0c1443e4914567ab148d8a065ccc7992c014693c02eeba775dc903d00eeab8fdabdc4;
    5'b01001 : xpb = 1024'h1135ef54743ded14b70bc7840e24fbb0e13a2fff0d18814e516ab2878a5ae5d0bd1805707d38ba9dac3cf84b3bb15c9550aa9c6edbf105f9fbdb989dbef0598e04b7bc15c70f977d703b22b9c7ef6676a3c609421337896408e41dc2f5478823ae8e6dcc71a2f5acf11292f110696e5abecb4557f43ee98a21694efebd64e247;
    5'b01010 : xpb = 1024'h7546db1bb402084dadf3ae7bfc5b3f471cd78c6f68b30544122a10e2a7d84308d3eda1156d37f93750cd6fecc0a3fe6badafa789408b96ce083005aabbf1c0c77ebf4395b07e5178dc5e60efddbcfb49af5094f37fdd953f8b2f1cd5b0d8f1954ddb596c195d9b0ec87f3ff97f77019838b03aa6915353b44c412a5673d16d35;
    5'b01011 : xpb = 1024'h28aa818d31d7eebdd9d61d9cda373b8be6fee5aeeed5e8c2550cb5e81252f338e77abf419310b94255ffa84762388f77a69a8abd8273575663e533597e20b34f84779666ea5c0e2f35e79c835aaecbebc6d6270c5ffd740a57ed89edb23fb874be20b2e2104f47e3192c0622f6b46eac63bb5112de1c60ae30a98aa9a15b91b8;
    5'b01100 : xpb = 1024'h8cbb6d54719c09f6d0be0494c86d7f22229c421f4a706cb815cc14432fd05070fe505ae6830ff7dbfa901fe8e72b314e039f95d7e70de82a7039a0667b221a88fe7f1de6d3cac82aa20adab9707c60bed260b2bdcca37fe5da3889006dd121e65d6d9e81b809ed44f098b32b65c201e9dda046617b30cad85b81660157c81ca6;
    5'b01101 : xpb = 1024'h401f13c5ef71f066fca073b5a6497b66ecc39b5ed093503658aeb9489a4b00a111dd7912a8e8b7e6ffc2584388bfc259fc8a790c28f5a8b2cbeece153d510d11043770b80da884e0fb94164ced6e3160e9e644d6acc35eb0a6f6f6186f37e8c5cdb2f7f7aefb9a1941457954dcff6efe08ab5ccdc7f9d7d23fe9c65485524129;
    5'b01110 : xpb = 1024'ha42fff8d2f360b9ff3885aad947fbefd2860f7cf2c2dd42c196e17a3b7c85dd928b314b798e7f680a452cfe50db26430598f84268d903986d8433b223a52744a7e3ef837f7173edc67b75483033bc633f570d08819696a8c2941f52b2ac952376cffe39756b63f7b18b2265d4c0d023b8290521c650e41fc6ac1a1ac3bbecc17;
    5'b01111 : xpb = 1024'h5793a5fead0bf2101f6ac9ce725bbb41f288510eb250b7aa5c50bca922430e093c4032e3bec0b68ba985083faf46f53c527a675acf77fa0f33f868d0fc8166d283f74b0930f4fb92c1409016802d96d60cf662a0f9894956f60062432c301916dd453d0d4da7ec4f695eec86c34a6f4fad9b6888b1d74ef64f2a01ff6948f09a;
    5'b10000 : xpb = 1024'haf74c702ae1d8804b4d38ef5037b786bcafaa4e38739b289f3361ae8cbdbe394fcd510fe4997696aeb7409a50db86484b654a8f115fba978fad967fbeb0595a89af9dda6ad2b8491ac9cba9fd1f6778247bf4b9d9a92821c2becf5b2d96dff64d8a968344999923ba0bb2b03a87dc63d8a67ef4fea05bf03392625296d3151d;
    5'b10001 : xpb = 1024'h6f0838376aa5f3b942351fe73e6dfb1cf84d06be940e1f1e5ff2c009aa3b1b7166a2ecb4d498b5305347b83bd5ce281ea86a55a975fa4b6b9c02038cbbb1c09403b7255a5441724486ed09e012ecfc4b3006806b464f33fd4509ce6de9284967ecd78222ec543e8591785fb8a9956fa1528b74439bb4c61a5e6a3daa4d3fa00b;
    5'b10010 : xpb = 1024'h226bdea8e87bda296e178f081c49f761c2745ffe1a31029ca2d5650f14b5cba17a300ae0fa71753b5879f0967762b92aa15538ddb7e20bf3f7b7313b7de0b31c096f782b8e1f2efae07645738fdecced478c1284266f12c811c83b85ea8f10475d1cdb98e345eb59e22525e220d2dcb57d968aafe87dd31442d29dfd7ac9c48e;
    5'b10011 : xpb = 1024'h867cca70283ff56264ff76000a803af7fe11bc6e75cb86926394c36a323328d99105a685ea70b3d4fd0a6837fc555b00fe5a43f81c7c9cc8040b9e487ae21a558376ffab778de8f64c9983a9a5ac61c053169e3593151ea394133a98a62079b8fc69c7388b0090bbb991d2ea8fe06ff2f77b7ffe85923d3e6daa795531364f7c;
    5'b10100 : xpb = 1024'h39e070e1a615dbd290e1e520e85c373cc83915adfbee6a10a677686f9cadd909a492c4b2104973e0023ca0929de9ec0cf745272c5e645d505fc0cbf73d110cdd892f527cb16ba5aca622bf3d229e32626a9c304e7334fd6e60d1a7b0a78740986caf20ae81f23d900a3e9914071ddd072286966ad25b4a385212d9a85ec073ff;
    5'b10101 : xpb = 1024'h9df15ca8e5d9f70b87c9cc18d6927ad303d6721e5788ee066736c6caba2b3641bb6860570048b279a6cd183422dc8de3544a3246c2feee246c1539043a1274170336d9fc9ada5fa81245fd73386bc7357626bbffdfdb0949e31ca6c36318aa0a0bfc0c4e29ace2f1e1ab461c762b70449c6b8bb96f6fb4627ceab500152cfeed;
    5'b10110 : xpb = 1024'h5155031a63afdd7bb3ac3b39b46e7717cdfdcb5dddabd184aa196bd024a5e671cef57e8326217284abff508ec4711eef4d35157b04e6aeacc7ca66b2fc41669f08ef2ccdd4b81c5e6bcf3906b55d97d78dac4e18bffae814afdb13db647f70e97c4165c4209e8fc632580c45ed68dd58c776a225bc38c15c6153155342b72370;
    5'b10111 : xpb = 1024'h4b8a98be185c3ebdf8eaa5a924a735c9825249d63ceb502ecfc10d58f2096a1e2829caf4bfa328fb13188e96605affb461ff8af46ce6f35237f9461be7059270ea77f9f0e95d914c558749a324f6879a531e031a01ac6df7c9980f365e637c8ec86bf3a17903c9a8304d26f64a64a6cf281b8920901ce5645bb75a6704147f3;
    5'b11000 : xpb = 1024'h68c995532149df24d67691528080b6f2d3c2810dbf6938f8adbb6f30ac9df3d9f95838543bf9712955c2008aeaf851d1a32503c9ab6900092fd4016ebb71c06088af071ef8049310317bb2d0481cfd4cb0bc6be30cc0d2bafee480062177a13a8bd3aad9bf4ae1fc5a717f77d3b3ddaa6c66ade0a6163880709350fe26add2e1;
    5'b11001 : xpb = 1024'h1c2d3bc49f1fc595025900735e5cb3379de9da4d458c1c76f09e14361718a40a0ce5568061d231345af438e58c8ce2dd9c0fe6fded50c0918b892f1d7da0b2e88e6759f031e24fc68b04ee63c50ecdeec841fdfbece0b185cba2ed1e22de6819fc19044fb63c8ed0ab1e45a14af14abe9771c44cf2df457a54fbb1515437f764;
    5'b11010 : xpb = 1024'h803e278bdee3e0cdf940e76b4c92f6cdd98736bda126a06cb15d72913496014223baf22551d16fcdff84b087117f84b3f914f21851eb516597dd9c2a7aa21a22086ee1701b5109c1f7282c99dadc62c1d3cc89ad5986bd614dedec30de6fd18b9b65efef5df73432828af2a9b9feddfc1156b99b8ff3afa47fd38ca90aa48252;
    5'b11011 : xpb = 1024'h33a1cdfd5cb9c73e2523568c2a6ef312a3ae8ffd274983eaf44017969f10b1723748105177aa2fd904b6e8e1b31415bff1ffd54c93d311edf392c9d93cd10caa0e273441552ec67850b1682d57ce3363eb521bc639a69c2c1aac5948dfd6986b0bab496554e8e106d337b8d3313c4b103c61d007dcbcbc9e643becfc382ea6d5;
    5'b11100 : xpb = 1024'h97b2b9c49c7de2771c0b3d8418a536a8df4bec6d82e407e0b4ff75f1bc8e0eaa4e1dabf667a96e72a94760833806b7964f04e066f86da2c1ffe736e639d273e3882ebbc13e9d8073bcd4a6636d9bc836f6dca777a64ca8079cf7585b9b6801dcaaf83504fca38668aaa465dba049de4db646c55679d126c88f13c853ee9b31c3;
    5'b11101 : xpb = 1024'h4b1660361a53c8e747edaca4f68132eda97345ad0906eb5ef7e21af72708beda61aaca228d822e7dae7998ddd99b48a247efc39b3a55634a5b9c6494fc01666b8de70e92787b3d2a165de1f6ea8d98d90e623990866c86d269b5c5739ccec8bc1b3d8e7af395333cfb512c0517874b61e151dbc2c69a33c2737c28a71c255646;
    5'b11110 : xpb = 1024'haf274bfd5a17e4203ed5939ce4b77683e510a21d64a16f54b8a1795244861c12788065c77d816d17530a107f5e8dea78a4f4ceb59eeff41e67f0d1a1f902cda507ee961261e9f7258281202d005b2dac19ecc541f31292adec00c4865860322dba8a7a1a9b4fd89ed2bdd90d8694de9f5b36d11163ae9dec9e5403fed291e134;
    5'b11111 : xpb = 1024'h628af26ed7edca906ab802bdc29372c8af37fb5ceac452d2fb841e57af00cc428c0d83f3a35a2d22583c48da00227b849ddfb1e9e0d7b4a6c3a5ff50bb31c02d0da6e8e39bc7b3dbdc0a5bc07d4cfe4e3172575ad3327178b8bf319e59c6f90d2acfd39092418573236a9f36fdd24bb38641e77db077aae682bc6452001c05b7;
    endcase
end

endmodule

module xpb_5_350
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h43abad172127c84c32460efd153d0e2bc9bface4acb6525c496e7c78245ce7deb50b306d4fe5b8c326ff03c338f9fd424d9889f9274f6efcd0791ba11b309893a7145a12ba95b191daa02f24a156e7acc5d79a9bed242ffddb10c3f21e6c8f446af7536f497d0011f108700fc1673005b6d14faf975114b0697a9d7d729531c5;
    5'b00010 : xpb = 1024'h87575a2e424f9098648c1dfa2a7a1c57937f59c9596ca4b892dcf8f048b9cfbd6a1660da9fcb71864dfe078671f3fa849b3113f24e9eddf9a0f23742366131274e28b425752b6323b5405e4942adcf598baf3537da485ffbb62187e43cd91e88d5eea6de92fa0023e210e01f82ce600b6da29f5f2ea22960d2f53afae52a638a;
    5'b00011 : xpb = 1024'h1a55c1efa189241bcbccb5202f5ce331ebc9037d30ab569d5e6ebc12ba140a941bd913cf258aabbad59ecc02c78fe6fc84af7605533b7caac0cc138516bf550980edd989803017707d468acb4b28f2d55d81d63b3ae662e8dba5b9dba11b0b3b11de68242bae07a84c5969504c6569e7d59a102c75a7e0e0f6005d73cedd2ee4;
    5'b00100 : xpb = 1024'h5e016f06c2b0ec67fe12c41d4499f15db588b061dd61a8f9a7dd388ade70f272d0e4443c7570647dfc9dcfc60089e43ed247fffe7a8aeba791452f2631efed9d2802339c3ac5c90257e6b9efec7fda82235970d7280a92e6b6b67dcdbf879a7f7cd5bb93752b07ba3d61d9600dcc99ed8c6b5fdc0cf8f5915f7afaf1417260a9;
    5'b00101 : xpb = 1024'ha1ad1c1de3d8b4b43058d31a59d6ff897f485d468a17fb55f14bb50302cdda5185ef74a9c5561d41239cd3893983e1811fe089f7a1da5aa461be4ac74d208630cf168daef55b7a943286e9148dd6c22ee9310b73152ec2e491c741bfddf429c3e7cd0f02bea807cc2e6a496fcf33c9f3433caf8ba44a0a41c8f5986eb407926e;
    5'b00110 : xpb = 1024'h34ab83df4312483797996a405eb9c663d79206fa6156ad3abcdd78257428152837b2279e4b155775ab3d98058f1fcdf9095eec0aa676f9558198270a2d7eaa1301dbb31300602ee0fa8d15969651e5aabb03ac7675ccc5d1b74b73b74236167623bcd048575c0f5098b2d2a098cad3cfab342058eb4fc1c1ec00bae79dba5dc8;
    5'b00111 : xpb = 1024'h785730f6643a1083c9df793d73f6d48fa151b3df0e0cff97064bf49d9884fd06ecbd580b9afb1038d23c9bc8c819cb3b56f77603cdc66852521142ab48af42a6a8f00d25baf5e072d52d44bb37a8cd5780db471262f0f5cf925c37a960a2a5ba8eb423b7a0d90f6289bb42b05a3203d56205700882a0d672557b5865104f8f8d;
    5'b01000 : xpb = 1024'hb5598b7c373a4073120106378d99b69f99b5d92e54bb17bd1ddb7c009df37dd9e800b0020ba4a6d59dd60451db5b7b34075d816d263070371eb1eee290d6688dbb53289c5fa94bf9d33713d4023f0d352ade815c38ef8bcb7e069a0c4e4926ccaa3e4fd398d16e6f403cbe123c90db1c9fce0d5c9a68df278867addfa025ae7;
    5'b01001 : xpb = 1024'h4f0145cee49b6c5363661f608e16a995c35b0a77920203d81b4c34382e3c1fbc538b3b6d70a0033080dc640856afb4f58e0e620ff9b2760042643a8f443dff1c82c98c9c8090465177d3a061e17ad880188582b1b0b328ba92f12d92e35121b1359b386c830a16f8e50c3bf0e5303db780ce308560f7a2a2e201185b6c978cac;
    5'b01010 : xpb = 1024'h92acf2e605c3349f95ac2e5da353b7c18d1ab75c3eb8563464bab0b05299079b08966bdac085bbf3a7db67cb8fa9b237dba6ec092101e4fd12dd56305f6e97b029dde6af3b25f7e35273cf8682d1c02cde5d1d4d9dd758b86e01f18501bdb0f5a0928bdbcc87170ad614ac00a6976dbd379f8034f848b7534b7bb5d8df2cbe71;
    5'b01011 : xpb = 1024'h25ab5aa764fcc822fcecc583a8367e9be564611015f70819304c73d2c3f34271ba591ecf4644f6282f7c2c47e5459eafc5254e1c259e83ae32b732733fccbb925ca30c13462aac301a79fc088b4ce3a8b02fbe50fe755ba59386237c65ff9da7dc824d21653b1e8f405d3531702e77999f96f1023f4e6ed36e86d851c8df89cb;
    5'b01100 : xpb = 1024'h695707be8624906f2f32d480bd738cc7af240df4c2ad5a7579baf04ae8502a506f644f3c962aaeeb567b300b1e3f9bf212bdd8154cedf2ab03304e145afd542603b7662600c05dc1f51a2b2d2ca3cb55760758eceb998ba36e96e76e846c2cec4779a090aeb81ea13165a5413195a79f566840b1d69f8383d80175cf3b74bb90;
    5'b01101 : xpb = 1024'had02b4d5a74c58bb6178e37dd2b09af378e3bad96f63acd1c3296cc30cad122f246f7fa9e61067ae7d7a33ce573999346056620e743d61a7d3a969b5762decb9aacbc038bb560f53cfba5a51cdfab3023bdef388d8bdbba149a7ab60a2d8bc30b270f3fff8351eb3226e1550f2fcd7a50d3990616df09834417c134cae09ed55;
    5'b01110 : xpb = 1024'h40011c970685ec3ec8b97aa3d79361cdd12d648d46a25eb68ebb2fe57e074d05d632329e6bcfa1e3051af84aacd585ac49d4c42178da0058f38345f8568c109bdd90e59cc65ac3a097c086d3d675d67e0db1948c395bbe8e6f2bdd58071aa8e2ee60b54590e926378cb69e81bc93e1817531012eb4f64fb4648735c597bcb8af;
    5'b01111 : xpb = 1024'h83acc9ae27adb48afaff89a0ecd06ff99aed1171f358b112d829ac5da26434e48b3d630bbbb55aa62c19fc0de5cf82ee976d4e1aa0296f55c3fc619971bca92f84a53faf80f075327260b5f877ccbe2ad3892f28267fee8c4a3ca14a25873827595808b4da6626497dbf0e917dfb11872c0250de4c476464ce01d3430a51ea74;
    5'b10000 : xpb = 1024'h16ab316f86e7480e624020c6f1b336d3f336bb25ca9762f7a3bb6f8013be6fbb3d001600417494dab3bac08a3b6b6f6680ebb02da4c60e06e3d63ddc521acd11b76a65138bf5297f3a66e27a8047e1a6a55bd02b871df1796fc0d34189c924d99547c9fa731a2dcde80797c247921b6393f9c1ab934d1be4f10cf5bbf404b5ce;
    5'b10001 : xpb = 1024'h5a56de86a80f105a94862fc406f044ffbcf6680a774db553ed29ebf8381b5799f20b466d915a4d9ddab9c44d74656ca8ce843a26cc157d03b44f597d6d4b65a55e7ebf26468adb111507119f219ec9536b336ac7744221774ad19733a835b41e003f1d69bc972ddfd91007d208f94b694acb115b2a9e30955a8793396699e793;
    5'b10010 : xpb = 1024'h9e028b9dc936d8a6c6cc3ec11c2d532b86b614ef240407b0369868705c783f78a71676dae140066101b8c810ad5f69eb1c1cc41ff364ec0084c8751e887bfe390593193901208ca2efa740c3c2f5b100310b05636166517525e25b25c6a243626b3670d906142df1ca1877e1ca607b6f019c610ac1ef4545c40230b6d92f1958;
    5'b10011 : xpb = 1024'h3100f35f28706c2a2e0cd5e721101a05deffbea2fb42b995022a2b92cdd27a4f58d929cf66ff409589598c8d02fb5663059b2632f8018ab1a4a2516168da221b38583e9d0c2540efb7ad6d45cb70d47c02dda666c20454624b668d1d2ae43014a726321e9ec835763461011293f7854b6993d1d808f4fcc5e70d532fc2e1e4b2;
    5'b10100 : xpb = 1024'h74aca076499834766052e4e4364d2831a8bf6b87a7f90bf14b98a80af22f622e0de45a3cb6e4f958b05890503bf553a55333b02c1f50f9ae751b6d02840abaaedf6c98afc6baf281924d9c6a6cc7bc28c8b54102af2884602677510f4950bf59121d858de845358825697122555eb55120652187a04611765087f0ad35771677;
    5'b10101 : xpb = 1024'h7ab0837a8d1c7f9c7937c0a3b2fef0c0109153b7f37bdd6172a6b2d63899d04bfa70d313ca4338d37f954cc9191401d3cb2123f23ed985f94f549456468de911231be13d1bfa6ce5a53c8ec7542dfa49a87e2060fc6874d4bfb8306ad92ac0b4e0d46d380f93d0c8fb1fa531ef5bf2d885c9254e74bc8f6739313261f29e1d1;
    5'b10110 : xpb = 1024'h4b56b54ec9f99045f9d98b07506cfd37cac8c2202bee10326098e7a587e684e374b23d9e8c89ec505ef8588fca8b3d5f8a4a9c384b3d075c656e64e67f997724b94618268c55586034f3f8111699c751605f7ca1fceab74b270c46f8cbff3b4fb9049a42ca763d1e80ba6a62e05cef333f2de2047e9cdda6dd0db0a391bf1396;
    5'b10111 : xpb = 1024'h8f026265eb2158922c1f9a0465aa0b6394886f04d8a4628eaa07641dac436cc229bd6e0bdc6fa51385f75c5303853aa1d7e32631728c765935e780879aca0fb8605a723946eb09f20f942735b7f0aefe2637173dea0ee749021d0aeaea6bca9423fbedb213f33d3071c2da72a1c41f38f5ff31b415edf25746884e210454455b;
    5'b11000 : xpb = 1024'h2200ca274a5aec159360312a6a8cd23decd218b8afe31473759927401d9da798db802100622edf480d9820cf59212719c16188447729150a55c15cca7b28339a931f979d51efbe3ed79a53b7c06bd279f809b8414aacea3627a13ce24eadb7465febaef7aca744b4dc0b63a36b5b29155df6a2815cf3a9d769937099ee0710b5;
    5'b11001 : xpb = 1024'h65ac773e6b82b461c5a640277fc9e069b691c59d5c9966cfbf07a3b841fa8f77908b516db214980b34972492921b245c0efa123d9e788407263a786b9658cc2e3a33f1b00c856fd0b23a82dc61c2ba26bde152dd37d11a3402b200d46d1a468acae30266f62444c6cd13d3b32cc2591b14c7f230f444be87d30e0e17609c427a;
    5'b11010 : xpb = 1024'ha95824558caa7cadf7ec4f249506ee9580517282094fb92c0876203066577756459681db01fa50ce5b962855cb15219e5c929c36c5c7f303f6b3940cb18964c1e1484bc2c71b21628cdab2010319a1d383b8ed7924f54a31ddc2c4c68b86d5cf35da55d63fa144d8be1c43c2ee298920cb9941e08b95d3383c88ab94d331743f;
    5'b11011 : xpb = 1024'h3c568c16ebe410315f2ce64a99e9b56fd89b1c35e08e6b10d407e352d7b1b22cf75934cf87b98b02e336ecd220b10e164610fe49ca6491b5168d704f91e788a4140d7126d21fd5af54e0de830b94c54f558b8e7c85934d1f0346f6bdefc8c28171ca171bd8554c5d2864ccf3b7c092fd3390b2add29b8ab85f93ce0dbce43f99;
    5'b11100 : xpb = 1024'h8002392e0d0bd87d9172f547af26c39ba25ac91a8d44bd6d1d765fcafc0e9a0bac64653cd79f43c60a35f09559ab0b5893a98842f1b400b1e7068bf0ad182137bb21cb398cb587412f810da7acebacfc1b63291872b77d1cde57bab00e3551c5dcc16a8b21d24c6f196d3d037927c302ea62025d69ec9f68c90e6b8b2f79715e;
    5'b11101 : xpb = 1024'h1300a0ef6c456c00f8b38c6db4098a75faa472ce64836f51e90822ed6d68d4e25e2718315d5e7dfa91d6b511af46f7d07d27ea55f6509f6306e068338d764519ede6f09d97ba3b8df7873a29b566d077ed35ca1bd355800a03dbeca772773e7818b12bd0ba8653f383b5c63442beccdf5259732ab0f256e8ec198e04192c3cb8;
    5'b11110 : xpb = 1024'h56ac4e068d6d344d2af99b6ac94698a1c4641fb31139c1ae32769f6591c5bcc11332489ead4436bdb8d5b8d4e840f512cac0744f1da00e5fd75983d4a8a6ddad94fb4ab0524fed1fd227694e56bdb824b30d64b7c079b007deecb09990e3cdbc83a87f400403540574be36440425fce5092ac2da48436b9955942b818bc16e7d;
    5'b11111 : xpb = 1024'h9a57fb1dae94fc995d3faa67de83a6cd8e23cc97bdf0140a7be51bddb622a49fc83d790bfd29ef80dfd4bc98213af2551858fe4844ef7d5ca7d29f75c3d776413c0fa4c30ce59eb1acc79872f8149fd178e4ff53ad9de005b9fd748baf505d00ee9fd2af4d80541765c6a653c58d2ceabffc1289df948049bf0ec8fefe56a042;
    endcase
end

endmodule

module xpb_5_95
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h460eceb48b03fbf5ba01a94cdbe1edfa3dfc84484c82bb233ea4eb304b785e1edd925aae5b49961da87d9c784dc6e07a3c43b8619573d4fd03fc4b180feb3b164cad317400907e06fd9a832605008952d8c1479f95c20d36670b60534453d5d06e65fbb016d35556c87f901458a78c938ebcfc8728e653ec2126b8fb0d1d02d4;
    5'b00010 : xpb = 1024'h8c1d9d691607f7eb74035299b7c3dbf47bf90890990576467d49d66096f0bc3dbb24b55cb6932c3b50fb38f09b8dc0f4788770c32ae7a9fa07f896301fd6762c995a62e80120fc0dfb35064c0a0112a5b1828f3f2b841a6cce16c0a688a7aba0dccbf7602da6aaad90ff2028b14f19271d79f90e51cca7d8424d71f61a3a05a8;
    5'b00011 : xpb = 1024'h217f26c7df1dbf1862ff840f834b829d487f89a8101090f23e12083b2f666d54956e929247b643ca5a1a962205f690a450b1013e9da8aeab5b55a1e9f4ef3c9171b85fad52207ccfe63586cf7625d7c7963edd4634bffa927f958eff12d0dedf1c2a60e693b10776d2bec95e12267f915d5d16b32a679e941d04afec9e74a211;
    5'b00100 : xpb = 1024'h678df57c6a21bb0e1d012d5c5f2d7097867c0df05c934c157cb6f36b7adecb737300ed40a2ffd9e80298329a53bd711e8cf4b9a0331c83a85f51ed0204da77a7be65912152b0fad6e3d009f57b26611a6f0024e5ca8207c8e6a0ef525724b4af8a905c96aa845ccd9b3e59726ace0c24ec1a133a534df2803e2b68e7ab91a4e5;
    5'b00101 : xpb = 1024'had9cc430f525b703d702d6a93b0f5e91c4789238a9160738bb5bde9bc6572992509347eefe497005ab15cf12a1845198c9387201c89058a5634e381a14c5b2be0b12c295534178dde16a8d1b8026ea6d47c16c85604414ff4dac4fa59b788a7ff8f65846c157b22463bde986c37598b87ad70fc17c34466c5f5221e2b8aea7b9;
    5'b00110 : xpb = 1024'h42fe4d8fbe3b7e30c5ff081f0697053a90ff1350202121e47c2410765eccdaa92add25248f6c8794b4352c440bed2148a162027d3b515d56b6ab43d3e9de7922e370bf5aa440f99fcc6b0d9eec4baf8f2c7dba8c697ff524ff2b1dfe25a1bdbe3854c1cd27620eeda57d92bc244cff22baba2d6654cf3d283a095fd93ce94422;
    5'b00111 : xpb = 1024'h890d1c44493f7a268000b16be278f334cefb97986ca3dd07bac8fba6aa4538c8086f7fd2eab61db25cb2c8bc59b401c2dda5baded0c53253baa78eebf9c9b439301df0cea4d177a6ca0590c4f14c38e2053f022bff42025b66367e5169f5938ea6babd7d3e3564446dfd22d07cf48bb6497729ed7db591145b3018d44a0646f6;
    5'b01000 : xpb = 1024'h1e6ea5a3125541536efce2e1ae0099dd9b8218afe3aef7b37b912d8142bae9dee2b95d087bd9354165d225edc41cd172b5cf4b5a438637050e049aa5cee27a9e087bed93f5d0f868b50611485d70fe03e9fb5033087de28117b54ca9f41ec6cce6192703a43fc10dafbccc05ddcbf220895a4792565087d035e756cace40e35f;
    5'b01001 : xpb = 1024'h647d74579d593d4928fe8c2e89e287d7d97e9cf83031b2d6ba3618b18e3347fdc04bb7b6d722cb5f0e4fc26611e3b1ecf21303bbd8fa0c021200e5bddecdb5b455291f07f661766fb2a0946e62718756c2bc97d29e3fefb77ec0acfd38729c9d547f22b3bb131664783c5c1a36737eb4181744197f36dbbc570e0fc5db5de633;
    5'b01010 : xpb = 1024'haa8c430c285d393ee300357b65c475d2177b21407cb46df9f8db03e1d9aba61c9dde1265326c617cb6cd5ede5faa92672e56bc1d6e6de0ff15fd30d5eeb8f0caa1d6507bf6f1f476b03b1794677210a99b7ddf723401fcede5cc0d507cc6726dc2e51e63d1e66bbb40bbec2e8f1b0b47a6d440a0a81d2fa87834c8c0e87ae907;
    5'b01011 : xpb = 1024'h3fedcc6af173006bd1fc66f1314c1c7ae401a257f3bf88a5b9a335bc722157337827ef9ac38f790bbfecbc0fca13621706804c98e12ee5b0695a3c8fc3d1b72f7a344d4147f175389b3b9817d396d5cb803a2d793d3ddd13974adba906efa5ac024387ea37f0c884827b9563eff271b1e6b75e4580b8266452ec06b76cb58570;
    5'b01100 : xpb = 1024'h85fc9b1f7c76fc618bfe103e0d2e0a7521fe26a0404243c8f84820ecbd99b55255ba4a491ed90f29686a588817da429142c404fa76a2baad6d5687a7d3bcf245c6e17eb54881f33f98d61b3dd8975f1e58fb7518d2ffea49fe563bfc4b437b7c70a9839a4ec41ddb4afb25784899fe4575745acca99e7a507412bfb279d28844;
    5'b01101 : xpb = 1024'h1b5e247e458cc38e7afa41b3d8b5b11dee84a7b7b74d5e74b91052c7560f66693004277eaffc26b87189b5b9824312411aed9575e963bf5ec0b39361a8d5b8aa9f3f7b7a9981740183d69bc144bc24403db7c31fdc3bca6fafd50a54d56caebab007ed20b4ce7aa48cbaceada97164afb55778718239710c4ec9fda8fe0d24ad;
    5'b01110 : xpb = 1024'h616cf332d090bf8434fbeb00b4979f182c812c0003d01997f7b53df7a187c4880d96822d0b45bcd61a075231d009f2bb57314dd77ed7945bc4afde79b8c0f3c0ebecacee9a11f20881711ee749bcad9316790abf71fdd7a616e06aa819c0848b1e6de8d0cba1cffb553a5ec20218f143441474f8ab1fc4f86ff0b6a40b2a2781;
    5'b01111 : xpb = 1024'ha77bc1e75b94bb79eefd944d90798d126a7db0485052d4bb365a2927ed0022a6eb28dcdb668f52f3c284eeaa1dd0d33593750639144b6958c8ac2991c8ac2ed73899de629aa2700f7f0ba20d4ebd36e5ef3a525f07bfe4dc7debcafb5e145a5b8cd3e480e27525521db9eed65ac07dd6d2d1717fd40618e491176f9f18472a55;
    5'b10000 : xpb = 1024'h3cdd4b4624aa82a6ddf9c5c35c0133bb3704315fc75def66f7225b028575d3bdc572ba10f7b26a82cba44bdb8839a2e56b9e96b4870c6e0a1c09354b9dc4f53c10f7db27eba1f0d16a0c2290bae1fc07d3f6a06610fbc5022f6a9953e83d8d99cc324e07487f821b5f79980bbb97e44112b48f24aca10fa06bcead959c81c6be;
    5'b10001 : xpb = 1024'h82ec19faafae7e9c97fb6f1037e321b57500b5a813e0aa8a35c74632d0ee31dca30514bf52fc00a07421e853d600835fa7e24f161c80430720058063adb030525da50c9bec326ed867a6a5b6bfe2855aacb7e805a6bdd2389675f9a72c91636a3a9849b75f52d77227f92820143f70d4a1718babd587638c8cf56690a99ec992;
    5'b10010 : xpb = 1024'h184da35978c445c986f7a086036ac85e418736bf8aebc535f68f780d6963e2f37d4ef1f4e41f182f7d4145854069530f800bdf918f4147b873628c1d82c8f6b7360309613d31ef9a52a7263a2c074a7c9174360caff9b25e47f4c7ffb6ba96a879f6b33dc55d343b69b8d1557516d73ee154a950ae225a4867aca4872dd965fb;
    5'b10011 : xpb = 1024'h5e5c720e03c841bf40f949d2df4cb6587f83bb07d76e80593534633db4dc41125ae14ca33f68ae4d25bee1fd8e303389bc4f97f324b51cb5775ed73592b431cd82b03ad53dc26da15041a9603107d3cf6a357dac45bbbf94af002852fb0e6c78e85caeeddc30899232386169cdbe63d27011a5d7d708ae3488d35d823af668cf;
    5'b10100 : xpb = 1024'ha46b40c28ecc3db4fafaf31fbb2ea452bd803f5023f13b7c73d94e6e00549f313873a7519ab2446ace3c7e75dbf71403f8935054ba28f1b27b5b224da29f6ce3cf5d6c493e52eba84ddc2c8636085d2242f6c54bdb7dcccb160b88a63f62424956c2aa9df303dee8fab7f17e2665f065fecea25effef0220a9fa167d48136ba3;
    5'b10101 : xpb = 1024'h39ccca2157e204e1e9f7249586b64afb8a06c0679afc562834a1804898ca504812bd84872bd55bf9d75bdba7465fe3b3d0bce0d02ce9f663ceb82e0777b83348a7bb690e8f526c6a38dcad09a22d224427b31352e4b9acf0c78a56fec98b758796211424590e3bb23c779ab3873d56d03eb1c003d889f8dc84b15473cc4e080c;
    5'b10110 : xpb = 1024'h7fdb98d5e2e600d7a3f8cde2629838f5c80344afe77f114b73466b78e442ae66f04fdf35871ef2177fd9781f9426c42e0d009931c25dcb60d2b4791f87a36e5ef4689a828fe2ea713677302fa72dab9700745af27a7bba272e95b7520ddf4b5804870fd46fe1910904f72ac7dfe4e363cd6ebc8b01704cc8a5d80d6ed96b0ae0;
    5'b10111 : xpb = 1024'h153d2234abfbc80492f4ff582e1fdf9e9489c5c75e8a2bf7340e9d537cb85f7dca99bc6b184209a688f8d550fe8f93dde52a29ad351ed012261184d95cbc34c3ccc69747e0e26b332177b0b3135270b8e530a8f983b79a4ce01485aa98087e9643e5795ad5ebedd246b6d3fd40bc49ce0d51da2fda0b4384808f4b655da5a749;
    5'b11000 : xpb = 1024'h5b4bf0e936ffc3fa4cf6a8a50a01cd98d2864a0fab0ce71a72b38883c830bd9ca82c1719738b9fc4317671c94c567458216de20eca92a50f2a0dcff16ca76fda1973c8bbe172e93a1f1233d91852fa0bbdf1f0991979a783471fe5fddc5c5466b24b750aecbf43290f3664119963d6619c0ed6b702f19770a1b604606ac2aa1d;
    5'b11001 : xpb = 1024'ha15abf9dc203bff006f851f1e5e3bb931082ce57f78fa23db15873b413a91bbb85be71c7ced535e1d9f40e419a1d54d25db19a7060067a0c2e0a1b097c92aaf06620fa2fe20367411cacb6ff1d53835e96b33838af3bb4b9ae2b465120b02a3720b170bb0392987fd7b5f425f20b62f52acbd33e2bd7eb5cc2dcbd5b77dfacf1;
    5'b11010 : xpb = 1024'h36bc48fc8b19871cf5f48367b16b623bdd094f6f6e9abce97220a58eac1eccd260084efd5ff84d70e3136b730486248235db2aebd2c77ebd816726c351ab71553e7ef6f53302e80307ad3782897848807b6f863fb87794df5faa14a9aad95d75600fda41699cf54919759d5b52e2c95f6aaef0e30472e2189d93fb51fc1a495a;
    5'b11011 : xpb = 1024'h7ccb17b1161d8312aff62cb48d4d50361b05d3b7bb1d780cb0c590bef7972af13d9aa9abbb41e38e8b9107eb524d04fc721ee34d683b53ba856371db6196ac6b8b2c28693393660a0547baa88e78d1d35430cddf4e39a215c6b574fcef2d3345ce75d5f180704a9fe1f52d6fab8a55f2f96bed6a2d593604bebab44d09374c2e;
    5'b11100 : xpb = 1024'h122ca10fdf334a3f9ef25e2a58d4f6dee78c54cf322892b8718dc299900cdc0817e486e14c64fb1d94b0651cbcb5d4ac4a4873c8dafc586bd8c07d9536af72d0638a252e8492e6cbf0483b2bfa9d96f538ed1be65775823b78344355795666840dd43f77e67aa76923b4d6a50c61bc5d394f0b0f05f42cc09971f2438d71e897;
    5'b11101 : xpb = 1024'h583b6fc46a37463558f4077734b6e4d92588d9177eab4ddbb032adc9db853a26f576e18fa7ae913b3d2e01950a7cb526868c2c2a70702d68dcbcc8ad469aade6b03756a2852364d2ede2be51ff9e204811ae6385ed378f71df3fa3a8bdaa3c547c3a3b27fd4dfcbfec3466b9650948f0c80c07962eda80acba98ab3e9a8eeb6b;
    5'b11110 : xpb = 1024'h9e4a3e78f53b422b12f5b0c41098d2d363855d5fcb2e08feeed798fa26fd9845d3093c3e02f82758e5ab9e0d584395a0c2cfe48c05e40265e0b913c55685e8fcfce4881685b3e2d9eb7d4178049ea99aea6fab2582f99ca8464b03fc01fe1224eaa036d814215216b4b3f6cdbdb0d58456c9041d57c0d498dbbf6439a7abee3f;
    5'b11111 : xpb = 1024'h33abc7d7be51095801f1e239dc20797c300bde77423923aaaf9fcad4bf73495cad531973941b3ee7eecafb3ec2ac65509af9750778a5071734161f7f2b9eaf61d54284dbd6b3639bd67dc1fb70c36ebccf2bf92c8c357ccdf7c9d2548c27456329fea05e7a2baedff673a0031e883bee96ac21c2305bcb54b676a2302be68aa8;
    endcase
end

endmodule

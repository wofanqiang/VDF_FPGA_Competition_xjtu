module xpb_5_685
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha144ce6f545dcfacff14da7b96d982c40bae2cd7a8f94b4c7e65c69ff1654f20f91e7efe752afe8531fbc8509c1ee79ef18844e6f9c0a7e3b89c656622524466d597b5457fe7857d8206c24c47d7787666e0af423465dd0a1643e887ae46151e5c75dbe13e63217b1dfc3fceb2cf5197757ed6bc330d83357b45c39e6e1419a9;
    5'b00010 : xpb = 1024'h91dc5788e6cd6a9133243d201d58be36a5e6567e7c7af6217eeed3ea2fc7f139eef48084202f7e7bc499515a54dfbe737ef661e7d0ce7f7bc0998b6e09d2141c36e035dc503e0db5f17381f5f6d32cbbd9bc64ebdc458d0376fb3f14a26187aa89e42598cbfd4a68b53898be6dce7d059c23ce9615cfa93ab01c0c385345cce7;
    5'b00011 : xpb = 1024'h8273e0a2793d057567339fc4a3d7f9a9401e80254ffca0f67f77e1346e2a9352e4ca8209cb33fe725736da640da095480c647ee8a7dc5713c896b175f151e3d19828b673209495ee60e0419fa5cee1014c981a9584253cfcd7b295a1967cfa36b7526f50599773564c74f1ae28cda873c2c8c66ff891cf3fe4f254d238778025;
    5'b00100 : xpb = 1024'h730b69bc0baca0599b4302692a57351bda56a9cc237e4bcb8000ee7eac8d356bdaa0838f76387e68e9d4636dc6616c1c99d29be97eea2eabd093d77dd8d1b386f9713709f0eb1e26d04d014954ca9546bf73d03f2c04ecf63869ec2e8a986cc2e4c0b907e7319c43e3b14a9de3ccd3e1e96dbe49db53f54519c89d6c1da93363;
    5'b00101 : xpb = 1024'h63a2f2d59e1c3b3dcf52650db0d6708e748ed372f6fff6a08089fbc8eaefd784d0768515213cfe5f7c71ec777f2242f12740b8ea55f80643d890fd85c051833c5ab9b7a0c141a65f3fb9c0f303c6498c324f85e8d3e49cef992142bb7eb3df4f122f02bf74cbc5317aeda38d9ecbff501012b623be161b4a4e9ee60602dae6a1;
    5'b00110 : xpb = 1024'h543a7bef308bd6220361c7b23755ac010ec6fd19ca81a175811309132952799dc64c869acc417e560f0f758137e319c5b4aed5eb2d05dddbe08e238da7d152f1bc02383791982e97af26809cb2c1fdd1a52b3b927bc44ce8f9d8994872cf51db3f9d4c770265ee1f1229fc7d59cb2abe36b7adfda0d8414f83752e9fe80c99df;
    5'b00111 : xpb = 1024'h44d20508c2fb710637712a56bdd4e773a8ff26c09e034c4a819c165d67b51bb6bc2288207745fe4ca1acfe8af0a3f09a421cf2ec0413b573e88b49958f5122a71d4ab8ce61eeb6d01e93404661bdb2171806f13c23a3fce25a8fefd566eac4676d0b962e9000170ca966556d14ca562c5d5ca5d7839a6754b84b7739cd3e4d1d;
    5'b01000 : xpb = 1024'h35698e22556b0bea6b808cfb445422e6433750677184f71f822523a7a617bdcfb1f889a6224a7e43344a8794a964c76ecf8b0fecdb218d0bf0886f9d76d0f25c7e93396532453f088dfffff010b9665c8ae2a6e5cb83acdbbb4746625b0636f39a79dfe61d9a3ffa40a2ae5ccfc9819a84019db1665c8d59ed21bfd3b270005b;
    5'b01001 : xpb = 1024'h2601173be7daa6ce9f8fef9fcad35e58dd6f7a0e4506a1f482ae30f1e47a5fe8a7ce8b2bcd4efe39c6e8109e62259e435cf92cedb22f64a3f88595a55e50c211dfdbb9fc029bc740fd6cbf99bfb51aa1fdbe5c8f73635cd51bfe9cef4f21a97fc7e8299dab3468e7d7df074c8ac8ad08aaa6958b491eb35f21f8086d97a1b399;
    5'b01010 : xpb = 1024'h1698a0557a4a41b2d39f5244515299cb77a7a3b518884cc983373e3c22dd02019da48cb178537e30598599a81ae67517ea6749ee893d3c3c0082bbad45d091c741243a92d2f24f796cd97f436eb0cee7709a12391b430cce7cb5f37c433d1c0bf556735538ce91d56f1b603c45c7d876d14b8d652be0d96456ce51077cd366d7;
    5'b01011 : xpb = 1024'h730296f0cb9dc9707aeb4e8d7d1d53e11dfcd5bec09f79e83c04b86613fa41a937a8e372357fe26ec2322b1d3a74bec77d566ef604b13d4087fe1b52d50617ca26cbb29a348d7b1dc463eed1dac832ce375c7e2c322bcc7dd6d4a0937588e9822c4bd0cc668bac30657b92c00c703e4f7f0853f0ea2ff698ba499a162051a15;
    5'b01100 : xpb = 1024'ha874f7de6117ac4406c38f646eab58021d8dfa33950342eb0226122652a4f33b8c990d359882fcac1e1eeb026fc6338b695dabd65a0bbbb7c11c471b4fa2a5e37804706f23305d2f5e4d01396583fba34a567724f78899d1f3b13290e59ea3b67f3a98ee04cbdc3e2453f8fab396557c6d6f5bfb41b0829f06ea5d3fd01933be;
    5'b01101 : xpb = 1024'h990c80f7f38747283ad2f208f52a9374b7c623da6884edc002af1f7091079554826f0ebb43877ca2b0bc740c28870a5ff6cbc8d73119934fc9196d2337227598d94cf105f386e567cdb9c0e3147fafe8bd322cce9f6849cb5468891dd9ba1642aca8e2a59266052bbb9051ea6e9580ea941453d52472a8a43bc0a5d9b54ae6fc;
    5'b01110 : xpb = 1024'h89a40a1185f6e20c6ee254ad7ba9cee751fe4d813c06989503382cbacf6a376d78451040ee8bfc994359fd15e147e1348439e5d808276ae7d116932b1ea2454e3a95719cc3dd6da03d26808cc37b642e300de2784747f9c4b51fdfaacdd588ceda172c5d20002e1952ccaada2994ac58bab94baf0734cea97096ee739a7c9a3a;
    5'b01111 : xpb = 1024'h7a3b932b18667cf0a2f1b75202290a59ec3677280f88436a03c13a050dccd9866e1b11c699907c8fd5f7861f9a08b80911a802d8df35427fd913b933062215039bddf2339433f5d8ac93403672771873a2e99821ef27a9be15d73637c1f0fb5b07857614ad9a5706ea0903c9e493d7c6e15e4388e9f6f4aea56d370d7fae4d78;
    5'b10000 : xpb = 1024'h6ad31c44aad617d4d70119f688a845cc866ea0cee309ee3f044a474f4c2f7b9f63f1134c4494fc8668950f2952c98edd9f161fd9b6431a17e110df3aeda1e4b8fd2672ca648a7e111bffffe02172ccb915c54dcb970759b7768e8cc4b60c6de734f3bfcc3b347ff481455cb99f93033508033b62ccb91ab3da437fa764e000b6;
    5'b10001 : xpb = 1024'h5b6aa55e3d45b2b90b107c9b0f27813f20a6ca75b68b991404d354998a921db859c714d1ef997c7cfb3298330b8a65b22c843cda8d50f1afe90e0542d521b46e5e6ef36134e106498b6cbf89d06e80fe88a103753ee709b0d745e351aa27e07362620983c8cea8e21881b5a95a922ea32ea8333caf7b40b90f19c8414a11b3f4;
    5'b10010 : xpb = 1024'h4c022e77cfb54d9d3f1fdf3f95a6bcb1badef41c8a0d43e9055c61e3c8f4bfd14f9d16579a9dfc738dd0213cc44b3c86b9f259db645ec947f10b2b4abca18423bfb773f805378e81fad97f337f6a3543fb7cb91ee6c6b9aa37fd39de9e4352ff8fd0533b5668d1cfafbe0e9915915a11554d2b16923d66be43f010db2f436732;
    5'b10011 : xpb = 1024'h3c99b7916224e881732f41e41c25f82455171dc35d8eeebe05e56f2e075761ea457317dd45a27c6a206daa467d0c135b476076dc3b6ca0dff9085152a42153d920fff48ed58e16ba6a463edd2e65e9896e586ec88ea669a398b4906b925ec58bbd3e9cf2e402fabd46fa6788d090857f7bf222f074ff8cc378c6597514751a70;
    5'b10100 : xpb = 1024'h2d3140aaf4948365a73ea488a2a53396ef4f476a31109993066e7c7845ba04033b491962f0a6fc60b30b335035ccea2fd4ce93dd127a78780105775a8ba1238e82487525a5e49ef2d9b2fe86dd619dcee13424723686199cf96be6f8867a3817eaace6aa719d23aade36c0788b8fb0eda2971aca57c1b2c8ad9ca20ef9a6cdae;
    5'b10101 : xpb = 1024'h1dc8c9c487041e49db4e072d29246f09898771110492446806f789c2841ca61c311f1ae89bab7c5745a8bc59ee8dc104623cb0dde988501009029d627320f343e390f5bc763b272b491fbe308c5d5214540fda1bde65c9965a233d857a95aaa4181b3061ff374c9875731968468edc5bc93c12a43a83d8cde272eaa8ded880ec;
    5'b10110 : xpb = 1024'he6052de1973b92e0f5d69d1afa3aa7c23bf9ab7d813ef3d0780970cc27f483526f51c6e46affc4dd8464563a74e97d8efaacddec09627a810ffc36a5aa0c2f944d976534691af63b88c7dda3b590659c6eb8fc58645798fbada94126eb11d3045897a198cd175860caf7258018e07c9efe10a7e1d45fed317493342c40a342a;
    5'b10111 : xpb = 1024'hafa5214d6dd188db0e72444d467d2d402f6dc78f810d3a8985e65dacb3e4975620139b6cbbdafad30a420db4436d7f77e13312c5ba56cf8bc99c28d07cf307601a712b98c67934e13a93402683307ed02dcc3f07baab5699d11e7c9a1cf7324ea1ff55facb3497012aabb226b45d5961655fe13a50538208928ef6e1321e4dd3;
    5'b11000 : xpb = 1024'ha03caa67004123bf4281a6f1ccfc68b2c9a5f136548ee55e866f6af6f247396f15e99cf266df7ac99cdf96bdfc2e564c6ea12fc69164a723d1994ed86472d7157bb9ac2f96cfbd19a9ffffd0322c3315a0a7f4b1628b069331d5d3271112a4dacf6d9fb258cebfeec1e80b166f5c84cf8c04d9143315a80dc7653f7b17500111;
    5'b11001 : xpb = 1024'h90d4338092b0bea376910996537ba42563de1add2810903386f8784130a9db880bbf9e7811e3fac02f7d1fc7b4ef2d20fc0f4cc768727ebbd99674e04bf2a6cadd022cc667264552196cbf79e127e75b1383aa5b0a6ab68c928d29b4052e1766fcdbe969e668e8dc592464062a5bb03db2a9d0ee15d7ce12fc3b8814fc81b44f;
    5'b11010 : xpb = 1024'h816bbc9a25205987aaa06c3ad9fadf97fe164483fb923b088781858b6f0c7da101959ffdbce87ab6c21aa8d16db003f5897d69c83f805653e1939ae8337276803e4aad5d377ccd8a88d97f2390239ba0865f6004b24a6685f3448040f94989f32a4a3321740311c9f060bcf5e55adbabd94ec8c7f899f4183111d0aee1b3678d;
    5'b11011 : xpb = 1024'h720345b3b78ff46bdeafcedf607a1b0a984e6e2acf13e5dd880a92d5ad6f1fb9f76ba18367ecfaad54b831db2670daca16eb86c9168e2debe990c0f01af246359f932df407d355c2f8463ecd3f1f4fe5f93b15ae5a2a167f53fbd6cded64fc7f57b87cd9019d3ab7879d15e5a05a0719fff3c0a1db5c1a1d65e81948c6e51acb;
    5'b11100 : xpb = 1024'h629acecd49ff8f5012bf3183e6f9567d328697d1a29590b28893a01febd1c1d2ed41a30912f17aa3e755bae4df31b19ea459a3c9ed9c0583f18de6f8027215eb00dbae8ad829ddfb67b2fe76ee1b042b6c16cb580209c678b4b32d5ae1806f0b8526c6908f3763a51ed96ed55b5932882698b87bbe1e40229abe61e2ac16ce09;
    5'b11101 : xpb = 1024'h533257e6dc6f2a3446ce94286d7891efccbec17876173b87891cad6a2a3463ebe317a48ebdf5fa9a79f343ee97f2887331c7c0cac4a9dd1bf98b0cffe9f1e5a062242f21a8806633d71fbe209d16b870def28101a9e97672156a83e7d59be197b29510481cd18c92b615c7c516585df64d3db055a0e06627cf94aa7c91488147;
    5'b11110 : xpb = 1024'h43c9e1006edec5187addf6ccf3f7cd6266f6eb1f4998e65c89a5bab468970604d8eda61468fa7a910c90ccf850b35f47bf35ddcb9bb7b4b401883307d171b555c36cafb878d6ee6c468c7dca4c126cb651ce36ab51c9266b7621da74c9b75423e00359ffaa6bb5804d5220b4d157896473e2a82f83a28c2d046af316767a3485;
    5'b11111 : xpb = 1024'h34616a1a014e5ffcaeed59717a7708d5012f14c61d1a91318a2ec7fea6f9a81dcec3a79a13fefa879f2e56020974361c4ca3facc72c58c4c0985590fb8f1850b24b5304f492d76a4b5f93d73fb0e20fbc4a9ec54f9a8d664d6d93101bdd2c6b00d71a3b73805de6de48e79a48c56b4d29a87a0096664b23239413bb05babe7c3;
    endcase
end

endmodule

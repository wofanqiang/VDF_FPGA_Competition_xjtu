module xpb_5_580
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha2734612eacc3045a103064b3061cf21c47846e2a3220122a59b8f65c1aaed8ecb927944bebf832a9d790d6ae876a6e95940dba126ff59bb42849eefad39afcafbcb8fdbe5e70e9e9f7ce06c93871bc8c883a54cd280b090cb5b431877cba5a8f09a2a36c25e5d2a161bc46da0b37f864845be9b7d0a8769ea52a72a2cd97e8f;
    5'b00010 : xpb = 1024'h943946d013aa2bc2770094bf506956f2177a8a9470cc61cdcd5a6575d0532e1593dc7510b35887c69b93db8eed8f3d084e678f5c2b4be32ad469fe811fa0eae48347eb091c3d1ff82c5fbe368e3273609d025101187b3410e129f436356ca8bfb22cc243d3f3c1c6a577a1fc4996d8e341b19e54a9c9b1a38e35d34fd0d096b3;
    5'b00011 : xpb = 1024'h85ff478d3c88273f4cfe23337070dec26a7cce463e76c278f5193b85defb6e9c5c2670dca7f18c6299aea9b2f2a7d327438e43172f986c9a664f5e12920825fe0ac4463652933151b9429c0088ddcaf87180fcb55e75b790f6f8a553f30dabd673bf5a50e589266334d37f8af27a32403b1d7e0dd688dbdd3218ff7574c7aed7;
    5'b00100 : xpb = 1024'h77c5484a656622bc22fbb1a790786692bd7f11f80c2123241cd81195eda3af2324706ca89c8a90fe97c977d6f7c0694638b4f6d233e4f609f834bda4046f61179240a16388e942ab462579ca8389229045ffa869a4703b110cc75671b0aeaeed3551f25df71e8affc42f5d199b5d8b9d34895dc703480616d5fc2b9b18bec6fb;
    5'b00101 : xpb = 1024'h698b49078e441e38f8f9401bb07fee63108155a9d9cb83cf4496e7a5fc4befa9ecba68749123959a95e445fafcd8ff652ddbaa8d38317f798a1a1d3576d69c3119bcfc90bf3f5404d30857947e347a281a7e541dea6abe912296078f6e4fb203f6e48a6b08b3ef9c538b3aa84440e4fa2df53d803007305079df57c0bcb5df1f;
    5'b00110 : xpb = 1024'h5b5149c4b72219b5cef6ce8fd08776336383995ba775e47a6c55bdb60af43030b504644085bc9a3693ff141f01f1958423025e483c7e08e91bff7cc6e93dd74aa13957bdf595655e5feb355e78dfd1bfeefcffd2306542113864b8ad2bf0b51ab87722781a495438e2e71836ed243e5727611d395cc65a8a1dc283e660acf743;
    5'b00111 : xpb = 1024'h4d174a81e0001532a4f45d03f08efe03b685dd0d75204525941493c6199c70b77d4e600c7a559ed29219e243070a2ba31829120340ca9258ade4dc585ba5126428b5b2eb2beb76b7ecce1328738b2957c37bab86765fc5914e3369cae991b8317a09ba852bdeb8d57242f5c5960797b420ccfcf2898584c3c1a5b00c04a40f67;
    5'b01000 : xpb = 1024'h3edd4b3f08de10af7af1eb78109685d4098820bf42caa5d0bbd369d62844b13e45985bd86eeea36e9034b0670c22c1c20d4fc5be45171bc83fca3be9ce0c4d7db0320e186241881179b0f0f26e3680ef97fa573abc5a491164021ae8a732bb483b9c52923d741d72019ed3543eeaf1111a38dcabb644aefd6588dc31a89b278b;
    5'b01001 : xpb = 1024'h30a34bfc31bc0c2c50ef79ec309e0da45c8a64711075067be3923fe636ecf1c50de257a46387a80a8e4f7e8b113b57e1027679794963a537d1af9b7b4073889737ae69459897996b0693cebc68e1d8876c7902ef0254cc9179d0cc0664d3be5efd2eea9f4f09820e90fab0e2e7ce4a6e13a4bc64e303d937096c08574c923faf;
    5'b01010 : xpb = 1024'h22694cb95a9a07a926ed086050a59574af8ca822de1f67270b5115f64595324bd62c53705820aca68c6a4caf1653edfff79d2d344db02ea76394fb0cb2dac3b0bf2ac472ceedaac49376ac86638d301f40f7aea3484f50118f9f7d242274c175bec182ac609ee6ab20568e7190b1a3cb0d109c1e0fc30370ad4f347cf08957d3;
    5'b01011 : xpb = 1024'h142f4d7683780325fcea96d470ad1d45028eebd4abc9c7d2330fec06543d72d29e764f3c4cb9b1428a851ad31b6c841eecc3e0ef51fcb816f57a5a9e2541feca46a71fa00543bc1e20598a505e3887b715765a578e49d391a56e2e41e015c48c80541ab972344b47afb26c003994fd28067c7bd73c822daa513260a294806ff7;
    5'b01100 : xpb = 1024'h5f54e33ac55fea2d2e8254890b4a51555912f867974287d5acec21662e5b35966c04b084152b5de889fe8f720851a3de1ea94aa56494186875fba2f97a939e3ce237acd3b99cd77ad3c681a58e3df4ee9f5060bd4445711bb3cdf5f9db6c7a341e6b2c683c9afe43f0e498ee2785684ffe85b90694157e3f5158cc83877881b;
    5'b01101 : xpb = 1024'ha868944697222ee873eb2b93c11674371a0976691c9629a0006a517c2490a0e83252c44d001239092618f66208fbc1273b2b704b7d489b41c9e4591f44e2e9aec9ef0aa92180dc164cb94886ec6afb17b278ab58a6c507a28698227815826d4c3280dcfd46280d0e552a0dfc832bd60b482e1a2be64bdf4ddf6833f2655106aa;
    5'b01110 : xpb = 1024'h9a2e9503c0002a6549e8ba07e11dfc076d0bba1aea408a4b2829278c3338e16efa9cc018f4ab3da52433c4860e14574630522406819524b15bc9b8b0b74a24c8516b65d657d6ed6fd99c2650e71652af86f7570cecbf8b229c66d395d3237062f413750a57bd71aae485eb8b2c0f2f684199f9e5130b0987834b601809481ece;
    5'b01111 : xpb = 1024'h8bf495c0e8de25e21fe6487c012583d7c00dfdccb7eaeaf64fe7fd9c41e121f5c2e6bbe4e9444241224e92aa132ced652578d7c185e1ae20edaf184229b15fe1d8e7c1038e2cfec9667f041ae1c1aa475b7602c132ba0ea2b23584b390c47379b5a60d176952d64773e1c919d4f288c53b05d99e3fca33c1272e8c3dad3f36f2;
    5'b10000 : xpb = 1024'h7dba967e11bc215ef5e3d6f0212d0ba81310417e85954ba177a6d3ac5089627c8b30b7b0dddd46dd206960ce184583841a9f8b7c8a2e37907f9477d39c189afb60641c30c4831022f361e1e4dc6d01df2ff4ae7578b49222c80435d14e6576907738a5247ae83ae4033da6a87dd5e2223471b9576c895dfacb11b86351364f16;
    5'b10001 : xpb = 1024'h6f80973b3a9a1cdbcbe165644134937866128530533fac4c9f65a9bc5f31a303537ab37cd2764b791e842ef21d5e19a30fc63f378e7ac1001179d7650e7fd614e7e0775dfad9217c8044bfaed718597704735a29beaf15a2ddd2e6ef0c0679a738cb3d318c7d9f809299843726b93b7f2ddd9910994888346ef4e488f52d673a;
    5'b10010 : xpb = 1024'h614697f863781858a1def3d8613c1b48b914c8e220ea0cf7c7247fcc6dd9e38a1bc4af48c70f50151c9efd162276afc204ecf2f292c74a6fa35f36f680e7112e6f5cd28b312f32d60d279d78d1c3b10ed8f205de04a99922f3a1980cc9a77cbdfa5dd53e9e13041d21f561c5cf9c94dc274978c9c607b26e12d810ae99247f5e;
    5'b10011 : xpb = 1024'h530c98b58c5613d577dc824c8143a3190c170c93ee946da2eee355dc7c822410e40eab14bba854b11ab9cb3a278f45e0fa13a6ad9713d3df35449687f34e4c47f6d92db86785442f9a0a7b42cc6f08a6ad70b1924aa41ca30970492a87487fd4bbf06d4bafa868b9b1513f54787fee3920b55882f2c6dca7b6bb3cd43d1b9782;
    5'b10100 : xpb = 1024'h44d29972b5340f524dda10c0a14b2ae95f195045bc3ece4e16a22bec8b2a6497ac58a6e0b041594d18d4995e2ca7dbffef3a5a689b605d4ec729f61965b587617e5588e59ddb558926ed590cc71a603e81ef5d46909ea0231f3efa4844e982eb7d830558c13dcd5640ad1ce3216347961a21383c1f8606e15a9e68f9e112afa6;
    5'b10101 : xpb = 1024'h36989a2fde120acf23d79f34c152b2b9b21b93f789e92ef93e6101fc99d2a51e74a2a2aca4da5de916ef678231c0721ee4610e239face6be590f55aad81cc27b05d1e412d43166e2b3d036d6c1c5b7d6566e08fad69923a3350dab66028a86023f159d65d2d331f2d008fa71ca46a0f3138d17f54c45311afe81951f8509c7ca;
    5'b10110 : xpb = 1024'h285e9aed06f0064bf9d52da8e15a3a8a051dd7a957938fa4661fd80ca87ae5a53cec9e7899736285150a35a636d9083dd987c1dea3f9702deaf4b53c4a83fd948d4e3f400a87783c40b314a0bc710f6e2aecb4af1c93a7234adc5c83c02b891900a83572e468968f5f64d8007329fa500cf8f7ae79045b54a264c1452900dfee;
    5'b10111 : xpb = 1024'h1a249baa2fce01c8cfd2bc1d0161c25a58201b5b253df04f8ddeae1cb723262c05369a448e0c6721132503ca3bf19e5cceae7599a845f99d7cda14cdbceb38ae14ca9a6d40dd8995cd95f26ab71c6705ff6b6063628e2aa360ab0da17dcc8c2fc23acd7ff5fdfb2beec0b58f1c0d53ad0664d767a5c3858e4647ed6accf7f812;
    5'b11000 : xpb = 1024'hbea9c6758abfd45a5d04a9121694a2aab225f0cf2e850fab59d842cc5cb66b2cd80961082a56bbd113fd1ee410a347bc3d52954ac92830d0ebf745f2f5273c79c46f59a77339aef5a78d034b1c7be9dd3ea0c17a888ae237679bebf3b6d8f4683cd658d07935fc87e1c931dc4f0ad09ffd0b720d282afc7ea2b199070ef1036;
    5'b11001 : xpb = 1024'hae5de27a43782d8b46d350dc51cb194c6f9aa5ef960a521d5b3913928776544199130f554164eee7aeb8df592980db651d1604f5d391dcc85144134edc8c2392981285765d1aa98df9f5b0a1454eda669c6db1647b095eb441d501d7b33934ef74678fc3c9f1bcf29438578b65a42c90481675bc4f8d3731d47dc0ba9dc88ec5;
    5'b11010 : xpb = 1024'ha023e3376c5629081cd0df5071d2a11cc29ce9a163b4b2c882f7e9a2961e94c8615d0b2135fdf383acd3ad7d2e997184123cb8b0d7de6637e32972e04ef35eac1f8ee0a39370bae786d88e6b3ffa31fe70ec5d18c103e23457a3b2f570da380635fa27d0db87218f2394351a0e8785ed418255757c4c616b7860ece041bfa6e9;
    5'b11011 : xpb = 1024'h91e9e3f495342484f2ce6dc491da28ed159f2d53315f1373aab6bfb2a4c6d54f29a706ed2a96f81faaee7ba133b207a307636c6bdc2aefa7750ed271c15a99c5a70b3bd0c9c6cc4113bb6c353aa58996456b08cd06fe65b46d7264132e7b3b1cf78cbfdded1c862bb2f012a8b76adf4a3aee352ea90b8ba51c441905e5b6bf0d;
    5'b11100 : xpb = 1024'h83afe4b1be122001c8cbfc38b1e1b0bd68a17104ff09741ed27595c2b36f15d5f1f102b91f2ffcbba90949c538ca9dc1fc8a2026e077791706f4320333c1d4df2e8796fe001cdd9aa09e49ff3550e12e19e9b4814cf8e93483411530ec1c3e33b91f57eafeb1eac8424bf037604e38a7345a14e7d5cab5dec027452b89add731;
    5'b11101 : xpb = 1024'h7575e56ee6f01b7e9ec98aacd1e9388dbba3b4b6ccb3d4c9fa346bd2c217565cba3afe8513c90157a72417e93de333e0f1b0d3e1e4c4028698d99194a6290ff8b603f22b3672eef42d8127c92ffc38c5ee68603592f36cb4990fc64ea9bd414a7ab1eff810474f64d1a7cdc6093192042dc5f4a10289e018640a71512da4ef55;
    5'b11110 : xpb = 1024'h673be62c0fce16fb74c71920f1f0c05e0ea5f8689a5e357521f341e2d0bf96e38284fa51086205f3a53ee60d42fbc9ffe6d7879ce9108bf62abef12618904b123d804d586cc9004dba6405932aa7905dc2e70be9d8edf034aede776c675e44613c44880521dcb4016103ab54b214eb612731d45a2f490a5207ed9d76d19c0779;
    5'b11111 : xpb = 1024'h5901e6e938ac12784ac4a79511f8482e61a83c1a6808962049b217f2df67d76a4acef61cfcfb0a8fa359b4314814601edbfe3b57ed5d1565bca450b78af7862bc4fca885a31f11a74746e35d2552e7f59765b79e1ee873b4c4ad288a24ff4777fdd720123372189df05f88e35af844be209db4135c08348babd0c99c75931f9d;
    endcase
end

endmodule

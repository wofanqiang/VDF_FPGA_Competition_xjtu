module xpb_5_660
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9b8b7fe2f2858e6ed0bbd40392e60879c3c6eeb2e06fbc53d6c94fb32c00f770d5271a7ea7f6e6d3b34d5b3e08eec22fff9499f7372eceaa2062f45a687bb701517f29fbc41ecdd6e9bb3b152d59c8a8d7bde65900afff9e962ac97665bf3f829f51479baad799bf1641ea8846be891bc24c0e03f0001b74434f593420bde7af;
    5'b00010 : xpb = 1024'h8669ba70231ce814d67230301571c9a21617da34eb67d8302fb5e610a4ff41d9a705b78485c74f18c73c77352e7f73959b0f0c084baacd089026a9569624f9512eaf1f48d8ac9e68c0dc7387c1d7cd20bb76d31974d9d22c76c900f21153dc730f9afd0da4e63af0a5c3ee3195acec0e35be3d258fb4d9b8402f3763b89968f3;
    5'b00011 : xpb = 1024'h7147f4fd53b441badc288c5c97fd8aca6868c5b6f65ff40c88a27c6e1dfd8c4278e4548a6397b75ddb2b932c541024fb36897e196026cb66ffea5e52c3ce3ba10bdf1495ed3a6efa97fdabfa5655d1989f2fbfd9e903a4ba5767386dbce879637fe4b27f9ef4dc223545f1dae49b4f00a9306c472f6997fc3d0f15935074ea37;
    5'b00100 : xpb = 1024'h5c262f8a844b9b60e1dee8891a894bf2bab9b13901580fe8e18f12cb96fbd6ab4ac2f19041681fa2ef1aaf2379a0d660d203f02a74a2c9c56fae134ef1777df0e90f09e301c83f8c6f1ee46cead3d61082e8ac9a5d2d774838056fe9687d1653f02e67f199037d53c4c7f5843389b1f31ca29b68cf1e564039eef3c2e8506b7b;
    5'b00101 : xpb = 1024'h47046a17b4e2f506e79544b59d150d1b0d0a9cbb0c502bc53a7ba9290ffa21141ca18e961f3887e80309cb1a9f3187c66d7e623b891ec823df71c84b1f20c040c63eff301656101e46401cdf7f51da8866a1995ad15749d618a3a7651411b34460781d6393121e855449f92d827814e59014ca8a6ed3148436ced1f2802becbf;
    5'b00110 : xpb = 1024'h31e2a4a4e57a4eaced4ba0e21fa0ce435f5b883d174847a193683f8688f86b7cee802b9bfd08f02d16f8e711c4c2392c08f8d44c9d9ac6824f357d474cca0290a36ef47d2ae3e0b01d61555213cfdf004a5a861b45811c63f941dee0bfa65034d0c1d2d58d20bfb6e3cbfcd6d16677d80386f9ac0e87d2c833aeb02218076e03;
    5'b00111 : xpb = 1024'h1cc0df321611a852f301fd0ea22c8f6bb1ac73bf2240637dec54d5e401f6b5e5c05ec8a1dad958722ae80308ea52ea91a473465db216c4e0bef932437a7344e0809ee9ca3f71b141f4828dc4a84de3782e1372dbb9aaeef1d9e0165c6b3aed25410b8847872f60e8734e00802054daca76f928cdae3c910c308e8e51afe2ef47;
    5'b01000 : xpb = 1024'h79f19bf46a901f8f8b8593b24b8509403fd5f412d387f5a45416c417af5004e923d65a7b8a9c0b73ed71f000fe39bf73fedb86ec692c33f2ebce73fa81c87305dcedf1753ff81d3cba3c6373ccbe7f011cc5f9c2dd4c17fba7e4dd816cf8a15b1553db9813e021a02d004296f433dbcea6b57ef4df14f502d6e6c8147be708b;
    5'b01001 : xpb = 1024'ha32a99a2392e9067c9742d3eb79e590dc7c44df40da83bae1c0abbf4a6f5f7bf6764802660a0a78af2247a3e18d25e273f825265fdc191e94f1fdb9a10983e31af4e0913181e4faab55f014c6a25b098e98a45f52e84c11e50a9174e7c8ec99850a685552c159bd91911eeb1b601c6d8acb765f33df16ac470bdc5b5687c583a;
    5'b01010 : xpb = 1024'h8e08d42f69c5ea0dcf2a896b3a2a1a361a15397618a0578a74f752521ff4422839431d2c3e710fd0061396353e630f8cdafcc477123d9047bee390963e4180818c7dfe602cac203c8c8039befea3b510cd4332b5a2ae93ac31474eca28236688c0f03ac726243d0aa893f25b04f029cb20299514dda629086d9da3e50057d97e;
    5'b01011 : xpb = 1024'h78e70ebc9a5d43b3d4e0e597bcb5db5e6c6624f823987366cde3e8af98f28c910b21ba321c4178151a02b22c63f3c0f27677368826b98ea62ea745926beac2d169adf3ad4139f0ce63a172319321b988b0fc1f7616d8663a11e58645d3b803793139f0392032de3c3815f60453de8cbd939bc4367d5ae74c6a7d821498335ac2;
    5'b01100 : xpb = 1024'h63c54949caf49d59da9741c43f419c86beb7107a2e908f4326d07f0d11f0d6f9dd005737fa11e05a2df1ce238984725811f1a8993b358d049e6afa8e9994052146dde8fa55c7c1603ac2aaa4279fbe0094b50c368b0238c7f283bdc17f4ca069a183a5ab1a417f6dc797f9ada2ccefb0070df3581d0fa590675d6044300edc06;
    5'b01101 : xpb = 1024'h4ea383d6fb8bf6ffe04d9df0c1cd5daf1107fbfc3988ab1f7fbd156a8aef2162aedef43dd7e2489f41e0ea1aaf1523bdad6c1aaa4fb18b630e2eaf8ac73d4771240dde476a5591f211e3e316bc1dc278786df8f6ff2c0b55d321f53d2ae13d5a11cd5b1d1450209f5719fd56f1bb52a27a802279bcc463d4643d3e73c7ea5d4a;
    5'b01110 : xpb = 1024'h3981be642c2350a5e603fa1d44591ed76358e77e4480c6fbd8a9abc803ed6bcb80bd9143b5b2b0e455d00611d4a5d52348e68cbb642d89c17df26486f4e689c1013dd3947ee36283e9051b89509bc6f05c26e5b77355dde3b3c02cb8d675da4a8217108f0e5ec1d0e69c010040a9b594edf2519b5c792218611d1ca35fc5de8e;
    5'b01111 : xpb = 1024'h245ff8f15cbaaa4bebba5649c6e4dfffb5a9d3004f78e2d8319642257cebb634529c2e499383192969bf2208fa368688e460fecc78a9881fedb61983228fcc10de6dc8e193713315c02653fbe519cb683fdfd277e77fb071945e6434820a773af260c601086d6302761e04a98f981887616480bcfc2de05c5dfcfad2f7a15fd2;
    5'b10000 : xpb = 1024'hf3e337e8d5203f1f170b2764970a12807fabe825a70feb48a82d882f5ea009d247acb4f7153816e7dae3e001fc737ee7fdb70dd8d25867e5d79ce7f50390e60bb9dbe2ea7ff03a797478c6e7997cfe02398bf385ba982ff74fc9bb02d9f142b62aa7b73027c043405a00852de867b79d4d6afde9be29ea05adcd9028f7ce116;
    5'b10001 : xpb = 1024'haac9b3617fd79260c22c8679dc56a9a1cbc1ad353ae0bb08614c283621eaf80df9a1e5ce194a684230fb993e28b5fa1e7f700ad4c45455287ddcc2d9b8b4c5620d1ce82a6c1dd17e8102c783a6f19888fb56a5915c59829e0b276526935e53ae01fbc30ead539df31be1f2db254504959722bde28be2ba149e2c3236b03ac8c5;
    5'b10010 : xpb = 1024'h95a7edeeb06eec06c7e2e2a65ee26aca1e1298b745d8d6e4ba38be939ae94276cb8082d3f71ad08744eab5354e46ab841aea7ce5d8d05386eda077d5e65e07b1ea4cdd7780aba2105823fff63b6f9d00df0f9251d083552bebc59ca23ef2f09e72457880a7623f24ab63f684743367880a94ed042b9778589b0c106648164a09;
    5'b10011 : xpb = 1024'h8086287be10645accd993ed2e16e2bf27063843950d0f2c1132554f113e78cdf9d5f1fd9d4eb38cc58d9d12c73d75ce9b664eef6ed4c51e55d642cd214074a01c77cd2c4953972a22f453868cfeda178c2c87f1244ad27b9cc63d41dea878d8ee28f2df2a170e0563ae5fa2dc321ca7a7e071c25cb4c369c97ebee95dff1cb4d;
    5'b10100 : xpb = 1024'h6b646309119d9f52d34f9aff63f9ed1ac2b46fbb5bc90e9d6c11eb4e8ce5d7486f3dbcdfb2bba1116cc8ed2399680e4f51df610801c85043cd27e1ce41b08c51a4acc811a9c74334066670db646ba5f0a6816bd2b8d6fa47ad020b99961c2a7f52d8e3649b7f8187ca67fdd712102d6cf1794b476b00f4e094cbccc577cd4c91;
    5'b10101 : xpb = 1024'h56429d964234f8f8d905f72be685ae4315055b3d66c12a79c4fe81ac05e421b1411c59e5908c095680b8091abef8bfb4ed59d31916444ea23ceb96ca6f59cea181dcbd5ebe5513c5dd87a94df8e9aa688a3a58932d00ccd58da0431541b0c76fc32298d6958e22b959ea018060fe905f64eb7a690ab5b32491abaaf50fa8cdd5;
    5'b10110 : xpb = 1024'h4120d82372cc529edebc535869116f6b675646bf71b946561deb18097ee26c1a12faf6eb6e5c719b94a72511e489711a88d4452a2ac04d00acaf4bc69d0310f15f0cb2abd2e2e457b4a8e1c08d67aee06df34553a12a9f636e3e7a90ed456460336c4e488f9cc3eae96c0529afecf351d85da98aaa6a71688e8b8924a7844f19;
    5'b10111 : xpb = 1024'h2bff12b0a363ac44e472af84eb9d3093b9a732417cb1623276d7ae66f7e0b682e4d993f14c2cd9e0a89641090a1a2280244eb73b3f3c4b5f1c7300c2caac53413c3ca7f8e770b4e98bca1a3321e5b35851ac3214155471f14edcb20c98da0150a3b603ba89ab651c78ee08d2fedb56444bcfd8ac4a1f2fac8b6b67543f5fd05d;
    5'b11000 : xpb = 1024'h16dd4d3dd3fb05eaea290bb16e28f1bc0bf81dc387a97e0ecfc444c470df00ebb6b830f729fd4225bc855d002faad3e5bfc9294c53b849bd8c36b5bef8559591196c9d45fbfe857b62eb52a5b663b7d035651ed4897e447f2f7ae988446e9e4113ffb92c83ba064e08700c7c4dc9b936bf4207cde9d3edf0884b4583d73b51a1;
    5'b11001 : xpb = 1024'h1bb87cb04925f90efdf67ddf0b4b2e45e49094592a199eb28b0db21e9dd4b548896cdfd07cdaa6ad07478f7553b854b5b439b5d6834481bfbfa6abb25fed7e0f69c9293108c560d3a0c8b184ae1bc48191e0b94fda8170d10192103f0033b3184496e9e7dc8a77f97f210259cb81c2932b436ef8988ac34852b23b36f16d2e5;
    5'b11010 : xpb = 1024'h9d4707adf717edffc09b3be1839abb5e220ff7f87311563eff7a2ad515de42c55dbde87bafc4913e83c1d4355e2a477b5ad835549f6316c61c5d5f158e7a8ee2481bbc8ed4ab23e423c7c62d783b84f0f0dbf1edfe5816aba643ea7a55c27ab4239ab63a28a0413eae33faade376a544f50044f37988c7a8c87a7ce78fd4ba94;
    5'b11011 : xpb = 1024'h8825423b27af47a5c651980e06267c867460e37a7e09721b5866c1328edc8d2e2f9c85818d94f98397b0f02c83baf8e0f652a765b3df15248c211411bc23d132254bb1dbe938f475fae8fea00cb98968d494deae7281e93986e221f6015717a493e46bac22aee2703db5fe573265083768727415193d85ecc55a5b1727b03bd8;
    5'b11100 : xpb = 1024'h73037cc85846a14bcc07f43a88b23daec6b1cefc89018df7b153579007dad797017b22876b6561c8aba00c23a94baa4691cd1976c85b1382fbe4c90de9cd1382027ba728fdc6c507d20a3712a1378de0b84dcb6ee6abbbc767805971acebb495042e211e1cbd83a1cd38020081536b29dbe4a336b8f24430c23a3946bf8bbd1c;
    5'b11101 : xpb = 1024'h5de1b75588ddfaf1d1be50670b3dfed71902ba7e93f9a9d40a3feded80d921ffd359bf8d4935ca0dbf8f281acedc5bac2d478b87dcd711e16ba87e0a177655d1dfab9c7612549599a92b6f8535b592589c06b82f5ad58e55481e90ed588051857477d69016cc24d35cba05a9d041ce1c4f56d25858a70274bf1a177657673e60;
    5'b11110 : xpb = 1024'h48bff1e2b9755497d774ac938dc9bfff6b53a6009ef1c5b0632c844af9d76c68a5385c9327063252d37e4411f46d0d11c8c1fd98f153103fdb6c3306451f9821bcdb91c326e2662b804ca7f7ca3396d07fbfa4efceff60e328bcc8690414ee75e4c18c0210dac604ec3c09531f30310ec2c90179f85bc0b8bbf9f5a5ef42bfa4;
    5'b11111 : xpb = 1024'h339e2c6fea0cae3ddd2b08c010558127bda49182a9e9e18cbc191aa872d5b6d17716f99904d69a97e76d600919fdbe77643c6faa05cf0e9e4b2fe80272c8da719a0b87103b7036bd576de06a5eb19b48637891b043293371095affe4afa98b66550b41740ae967367bbe0cfc6e1e9401363b309b98107efcb8d9d3d5871e40e8;
    endcase
end

endmodule

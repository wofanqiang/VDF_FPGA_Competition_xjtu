module xpb_5_85
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6f2e7c4e9c199031451cf0c8947fbf55b6eab722c8535c99eef779c9b1a78ce991c7fb7fa2b907fd39a46532b3119a4767838405d437d1f4d95525ed090256325fb8fb6e396a5367f27242490ba376851e2d514ad845d2dacfc72aa6c3e5e53363af5c6b243419265770d0163ef011e31f7ab46b76499f305754660c18d9a9aa;
    5'b00010 : xpb = 1024'h2dafb3477644eb99bf3469ba18a53759fc5f6b14bb2f18bc60123a3db04c6ccb204779867b4b916bd3ea8b1e82c523c46aece02585bcd39e020b0c7bd73237b34b22c22dc343a98ad24a81ef7e6b28d94855a8fd240578a4ea01c352cda127d4985726ac979f39bf2821b94d860ffd9cf01b89f49c47e13068395113a8d0ece9;
    5'b00011 : xpb = 1024'h9cde2f96125e7bcb04515a82ad24f6afb34a2237838275564f09b40761f3f9b4b20f75061e0499690d8ef05135d6be0bd270642b59f4a592db603268e0348de5aadbbd9bfcadfcf2c4bcc4388a0e9f5e6682fa47fc4b4b7fb9c8edf991870d07fc068317bbd352e57f928963c5000f800f963e6012918060bf8db71fc1aa9693;
    5'b00100 : xpb = 1024'h5b5f668eec89d7337e68d374314a6eb3f8bed629765e3178c024747b6098d996408ef30cf69722d7a7d5163d058a4788d5d9c04b0b79a73c041618f7ae646f669645845b86875315a49503defcd651b290ab51fa480af149d40386a59b424fa930ae4d592f3e737e5043729b0c1ffb39e03713e9388fc260d072a22751a1d9d2;
    5'b00101 : xpb = 1024'h19e09d87c6b5329bf8804c65b56fe6b83e338a1b6939ed9b313f34ef5f3db977cf0e7113cf29ac46421b3c28d53dd105d9431c6abcfea8e52ccbff867c9450e781af4b1b1060a938846d43856f9e0406bad3a9ac93ca9713ee3e1f51a4fd924a6556179aa2a9941720f45bd2533fe6f3b0d7e9725e8e0460e1578d2ee1991d11;
    5'b00110 : xpb = 1024'h890f19d662cec2cd3d9d3d2e49efa60df51e413e318d4a352036aeb910e5466160d66c9371e2b4437bbfa15b884f6b4d40c6a07091367ada062125738596a719e168468949cafca076df85ce7b417a8bd900faf76c1069eebe0549f868e3777dc9057405c6ddad3d78652be8922ff8d6d0529dddd4d7a39138abf33afa72c6bb;
    5'b00111 : xpb = 1024'h479050cf3cfa1e35b7b4b61fce151e123a92f5302469065791516f2d0f8a2642ef55ea9a4a753db21605c7475802f4ca442ffc9042bb7c832ed70c0253c6889accd20d48d3a452c356b7c574ee092ce0032952a9b7d00fb8d83fe2a4729eba1efdad3e473a48cdd64916151fd94fe490a0f37366fad5e5914990de428a6a09fa;
    5'b01000 : xpb = 1024'h61187c81725799e31cc2f11523a96168007a9221744c27a026c2fa10e2f06247dd568a12307c720b04bed3327b67e47479958aff4407e2c578cf29121f66a1bb83bd4085d7da8e63690051b60d0df342d51aa5c038fb582f27a7b507c59fcc032550888adb3ee6f19c6fe57206fd04a719448f020d427915a75c94a1a614d39;
    5'b01001 : xpb = 1024'h75400416b33f09cf76e91fd9e6ba556c36f26044df981f13f163a96abfd6930e0f9d6420c5c0cf1de9f05265dac8188eaf1cdcb5c878502130e2187e2af8c04e17f4cf7696e7fc4e290247646c7455b94b7efba6dbd5885dc241a5f7403fe1f3960464f3d1e807957137ce6d5f5fe22d910efd5b971dc6c1b1ca2f56333af6e3;
    5'b01010 : xpb = 1024'h33c13b0f8d6a6537f10098cb6adfcd707c671436d273db36627e69debe7b72ef9e1ce2279e53588c84367851aa7ba20bb28638d579fd51ca5997ff0cf928a1cf035e963620c1527108da870adf3c080d75a7535927952e27dc7c3ea349fb2494caac2f354553282e41e8b7a4a67fcde761afd2e4bd1c08c1c2af1a5dc3323a22;
    5'b01011 : xpb = 1024'ha2efb75e2983f569361d8993ff5f8cc63351cb599ac737d05175e3a87022ffd92fe4dda7410c6089bddadd845d8d3c531a09bcdb4e3523bf32ed24fa022af801631791a45a2ba5d8fb4cc953eadf7e9293d4a4a3ffdb0102ac43694a0de109c82e5b8ba069874154995987bae56fdfca812a87503365a7f21a038069dc0be3cc;
    5'b01100 : xpb = 1024'h6170ee5703af50d1b0350285838504ca78c67f4b8da2f3f2c290a41c6ec7dfbabe645bae199ee9f8582103702d40c5d01d7318faffba25685ba30b88d05ad9824e815863e404fbfbdb2508fa5da730e6bdfcfc564b9aa6ccc67e01f6179c4c69630355e1dcf261ed6a0a70f22c8fcb8451cb5cd95963e9f22ae86b716c03270b;
    5'b01101 : xpb = 1024'h1ff2254fdddaac3a2a4c7b7707aa7ccebe3b333d807eb01533ab64906d6cbf9c4ce3d9b4f2317366f267295bfcf44f4d20dc751ab13f27118458f2179e8abb0339eb1f236dde521ebafd48a0d06ee33ae8255408975a4c96e0b89aa221578f0a97ab2023505d82863abb5a2973afb73e226c32627f622bf23bcd5678fbfa6a4a;
    5'b01110 : xpb = 1024'h8f20a19e79f43c6b6f696c3f9c2a3c247525ea6048d20caf22a2de5a1f144c85deabd53494ea7b642c0b8e8eb005e994885ff9208576f9065dae1804a78d113599a41a91a748a586ad6f8ae9dc1259c00652a5536fa01f71b07fc548e53d743dfb5a7c8e74919bac922c2a3fb29fc92141e6e6cdf5abcb229321bc8514d413f4;
    5'b01111 : xpb = 1024'h4da1d897541f97d3e980e531204fb428ba9a9e523badc8d193bd9ece1db92c676d2b533b6d7d04d2c651b47a7fb973118bc9554036fbfaaf8663fe9375bcf2b6850de1513121fba98d47ca904eda0c14307afd05bb5fc53bcaba5df4eef8b6df300246cfe7fcbc4562dd1376f9bfb4db1287bc571baa0d22a406a78ca4cb5733;
    5'b10000 : xpb = 1024'hc230f902e4af33c63985e22a4752c2d000f52442e8984f404d85f421c5e0c48fbaad142460f8e416097da664f6cfc8e8f32b15fe880fc58af19e52243ecd4377077a810bafb51cc6d200a36c1a1be685aa354b8071f6b05e4f4f6a0f8b3f98064aa11115b67dcde338dfcae40dfa094e32891e041a84f22b4eb929434c29a72;
    5'b10001 : xpb = 1024'h7b518bdeca64836da8b54eeb38f4eb82b6fa0966f6dce18df3cfd90bce0599328d72ccc1e8c8963e9a3c3f99027e96d5f6b63565bcb8ce4d886f0b0f4cef2a69d030a37ef465a5345f924c7fcd4534ed78d0a602df653de0b4bc2147bc99deb3c8596d7c7f9bf6048afeccc47fcfb27802a3464bb7f1ee530c3ff8a04d9c441c;
    5'b10010 : xpb = 1024'h39d2c2d7a48fded622ccc7dcbd1a6386fc6ebd58e9b89db064ea997fccaa79141bf24ac8c15b1fad34826584d2322052fa1f91856e3dcff6b124f19e1b1f0beabb9a6a3e7e3efb573f6a8c26400ce741a2f8fdb52b24e3aacef6b9f3c6552154fd0137bdf307169d5bafb5fbc6ef9e31d3441bd4ddf030531d24e3a7dd93875b;
    5'b10011 : xpb = 1024'ha9013f2640a96f0767e9b8a5519a22dcb359747bb20bfa4a53e213497e5205fdadba4648641427aa6e26cab78543ba9a61a3158b4275a1eb8a7a178b2421621d1b5365acb7a94ebf31dcce6f4bb05dc6c1264f00036ab6859ebde49a8a3b068860b09429173b2fc3b320861205dfb014f2bed0405439cf83747949b3f66d3105;
    5'b10100 : xpb = 1024'h6782761f1ad4ca6fe2013196d5bf9ae0f8ce286da4e7b66cc4fcd3bd7cf6e5df3c39c44f3ca6b119086cf0a354f74417650c71aaf3faa394b32ffe19f251439e06bd2c6c4182a4e211b50e15be78101aeb4ea6b24f2a5c4fb8f87d4693f6492995585e6a8aa6505c83d16f494cff9bcec35fa5c97a381183855e34bb86647444;
    5'b10101 : xpb = 1024'h2603ad17f50025d85c18aa8859e512e53e42dc5f97c3728f361794317b9bc5c0cab9425615393a87a2b3168f24aacd946875cdcaa57fa53ddbe5e4a8c081251ef226f32bcb5bfb04f18d4dbc313fc26f1576fe649aea0219d33315f29db18bcaca0028abfe1170f554825880941f878894007b52a036538396431fc3165bb783;
    5'b10110 : xpb = 1024'h953229669119b609a1359b50ee64d23af52d93826016cf29250f0dfb2d4352aa5c813dd5b7f24284dc577bc1d7bc67dbcff951d079b77732b53b0a95c9837b5151dfee9a04c64e6ce3ff90053ce338f433a44faf732fd4f4a2fa4099619770fe2daf851722458a1babf32896d30f996bb37b2fbe167ff2b3ed9785cf2f35612d;
    5'b10111 : xpb = 1024'h53b3605f6b4511721b4d1442728a4a3f3aa2477452f28b4b9629ce6f2be8328beb00bbdc9084cbf3769da1ada76ff158d362adf02b3c78dbddf0f12497b35cd23d49b5598e9fa48fc3d7cfabafaaeb485dcca761beef7abebd34d9456b52b39f62574f5895b0aab47ca411ce1a2f8525841c05473c7e34b3fe7c70d6bf2ca46c;
    5'b11000 : xpb = 1024'h1234975845706cda95648d33f6afc2438016fb6645ce476e07448ee32a8d126d798039e36917556210e3c79977237ad5d6cc0a0fdcc17a8506a6d7b365e33e5328b37c191878fab2a3b00f5222729d9c87f4ff140aaf2088d76f71f1750df64096ff199a091bcb4d4d54fb05614f70df54bcdad0627c76b40f615bde4f23e7ab;
    5'b11001 : xpb = 1024'h816313a6e189fd0bda817dfc8b2f81993701b2890e21a407f63c08acdc349f570b4835630bd05d5f4a882ccc2a35151d3e4f8e15b0f94c79dffbfda06ee59485886c778751e34e1a9622519b2e161421a622505ee2f4f363a7369c9838f3db73faae76052d4fe473a4c5cb1ba03f82c274378f3bd8c615e466b5c1ea67fd9155;
    5'b11010 : xpb = 1024'h3fe44a9fbbb558745498f6ee0f54f99d7c76667b00fd602a6756c920dad97f3899c7b369e462e6cde4ce52b7f9e89e9a41b8ea35627e4e2308b1e42f3d15760673d63e46dbbca43d75fa9141a0ddc675d04aa8112eb4992dc171354442af1e152f564046a0bb050c7576b452e75f6e7c44d864c4fec457e4779aacf1f7f4d494;
    5'b11011 : xpb = 1024'haf12c6ee57cee8a599b5e7b6a3d4b8f333611d9dc950bcc4564e42ea8c810c222b8faee9871beecb1e72b7eaacfa38e1a93c6e3b36b62017e2070a1c4617cc38d38f39b51526f7a5686cd38aac813cfaee77f95c06fa6c0891385feb0695034893059cb1c4ef1e32cce78469264f805f64531930750df714ceef12fe10ce7e3e;
    5'b11100 : xpb = 1024'h6d93fde731fa440e13cd60a827fa30f778d5d18fbc2c78e6c769035e8b25ec03ba0f2cf05fae7839b8b8ddd67cadc25eaca5ca5ae83b21c10abcf0ab1447adb9bef900749f004dc8484513311f48ef4f18a0510e52ba11d2ab72f897105045e9c7ad66f3385a3ecb9d986da06d6f6c1934f3eeb99b0c3914dfd3fe05a0c5c17d;
    5'b11101 : xpb = 1024'h2c1534e00c259f768de4d999ac1fa8fbbe4a8581af0835093883c3d289cacbe5488eaaf7384101a852ff03c24c614bdbb00f267a99c0236a3372d739e2778f3aaa62c73428d9a3eb281d52d79210a1a342c8a8c09e79b79cc5ad91431a0b888afc553134abc55f646e4956d7b48f57d30594c442c10a7b14f0b8e90d30bd04bc;
    5'b11110 : xpb = 1024'h9b43b12ea83f2fa7d301ca62409f685175353ca4775b91a3277b3d9c3b7258ceda56a676dafa09a58ca368f4ff72e6231792aa806df7f55f0cc7fd26eb79e56d0a1bc2a26243f7531a8f95209db4182860f5fa0b76bf8a779574bbe9ddf16dbe60048d9fcff9788ac5ba26edf37f69b6250f78ae37541a45480d4f194996ae66;
    5'b11111 : xpb = 1024'h59c4e827826a8b104d194353c4c4e055baa9f0966a374dc59895fe103a1738b068d6247db38c931426e98ee0cf266fa01afc06a01f7cf708357de3b5b9a9c6edf5858961ec1d4d75fa67d4c7107bca7c8b1e51bdc27f3041afaf5495e7acb05f94ac57e143649923966b10253a9f556ff5b04e375d525c4558f23a20d98df1a5;
    endcase
end

endmodule

module xpb_5_125
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'heda7a3d1a34fef602a9dc01cab4cdb8999c21da7194f86028fd4ec11ae84ea9db661b6a0d2087c6b499240462d6255d33ffec8dece5dbe50ec33dcc4e8184ceca234ff66e226287e12228c155f568eeb1dcc414814d6c56524cde75dab436c07da0eeddcf829900220a8d5f26b98ea01c1a8a88310d494280e4e33c2de47caa;
    5'b00010 : xpb = 1024'h1db4f47a3469fdec0553b80395699b71333843b4e329f0c051fa9d8235d09d53b6cc36d41a410f8d69324808c5ac4aba67ffd91bd9cbb7ca1d867b989d03099d94469fecdc44c50fc2445182abead1dd63b98829029ad8aca499bcebb5686d80fb41ddbb9f05320044151abe4d731d4038351510621a928501c9c6785bc8f954;
    5'b00011 : xpb = 1024'h2c8f6eb74e9efce207fd9405601e6929ccd4658f54bee9207af7ec4350b8ebfd9232523e276197541dcb6c0d288270179bffc5a9c6b193af2c49b964eb848e6c5e69efe34a672797a3667a4401e03acc15964c3d83e84502f6e69b61901ca44178e2cc996e87cb00661fa81d742cabe0544f9f989327dbc782aea9b489ad75fe;
    5'b00100 : xpb = 1024'h3b69e8f468d3fbd80aa770072ad336e266708769c653e180a3f53b046ba13aa76d986da834821f1ad26490118b589574cfffb237b3976f943b0cf7313a06133b288d3fd9b8898a1f8488a30557d5a3bac77310520535b159493379d76ad0db01f683bb773e0a6400882a357c9ae63a80706a2a20c435250a03938cf0b791f2a8;
    5'b00101 : xpb = 1024'h4a4463318308face0d514c08f588049b000ca94437e8d9e0ccf289c58689895148fe891241a2a6e186fdb415ee2ebad203ff9ec5a07d4b7949d034fd88879809f2b08fd026abeca765aacbc6adcb0ca9794fd46686831daf9b80584d458511c27424aa550d8cfd00aa34c2dbc19fc9208c84b4a8f5426e4c8478702ce5766f52;
    5'b00110 : xpb = 1024'h591edd6e9d3df9c40ffb280ac03cd25399a8cb1ea97dd240f5efd886a171d7fb2464a47c4ec32ea83b96d81a5104e02f37ff8b538d63275e589372c9d7091cd8bcd3dfc694ce4f2f46ccf48803c075982b2c987b07d08a05edcd36c320394882f1c59932dd0f9600cc3f503ae85957c0a89f3f31264fb78f055d5369135aebfc;
    5'b00111 : xpb = 1024'h67f957abb772f8ba12a5040c8af1a00c3344ecf91b12caa11eed2747bc5a26a4ffcabfe65be3b66ef02ffc1eb3db058c6bff77e17a4903436756b096258aa1a786f72fbd02f0b1b727ef1d4959b5de86dd095c8f891df65c401a1538faed7f436f668810ac922f00ee49dd9a0f12e660c4b9c9b9575d00d1864236a5413f68a6;
    5'b01000 : xpb = 1024'h76d3d1e8d1a7f7b0154ee00e55a66dc4cce10ed38ca7c30147ea7608d742754edb30db5069043e35a4c9202316b12ae99fff646f672edf287619ee62740c2676511a7fb37113143f0911460aafab47758ee620a40a6b62b29266f3aed5a1b603ed0776ee7c14c80110546af935cc7500e0d45441886a4a14072719e16f23e550;
    5'b01001 : xpb = 1024'h85ae4c25ebdcf6a617f8bc10205b3b7d667d30adfe3cbb6170e7c4c9f22ac3f8b696f6ba7624c5fc5962442779875046d3ff50fd5414bb0d84dd2c2ec28dab451b3dcfa9df3576c6ea336ecc05a0b06440c2e4b88bb8cf08e4b3d224b055ecc46aa865cc4b976101325ef8585c8603a0fceedec9b9779356880bfd1d9d0861fa;
    5'b01010 : xpb = 1024'h9488c6630611f59c1aa29811eb100936001952886fd1b3c199e5138b0d1312a291fd122483454dc30dfb682bdc5d75a407ff3d8b40fa96f293a069fb110f3013e5611fa04d57d94ecb55978d5b961952f29fa8cd0d063b5f3700b09a8b0a2384e84954aa1b19fa01546985b7833f924119096951ea84dc9908f0e059caecdea4;
    5'b01011 : xpb = 1024'ha36340a02046f4921d4c7413b5c4d6ee99b57462e166ac21c2e2624c27fb614c6d632d8e9065d589c2948c303f339b013bff2a192de072d7a263a7c75f90b4e2af846f96bb7a3bd6ac77c04eb18b8241a47c6ce18e53a7b5894d8f1065be5a4565ea4387ea9c930176741316a9f920e13523f3da1b9225db89d5c395f8d15b4e;
    5'b01100 : xpb = 1024'h1907587788dbebf54f0d83e701f5d55c1db930c7d84040a6e02f7b78fe102ee4580cb7fd35fdec1d7cf70edbeabaf940be4eec0f8137e710087a635733fc50005588ade7a0ba1197affe66d6ea526ff6254375d831ae6fb260ddb8b8647ee73b483a03c0956337411beb996d8e2895802649f7ffc5411edc44b2bcd9dd3718d;
    5'b01101 : xpb = 1024'h106aefc492c2bdb5579ab4403ad42b0e5b77b4e6ef18fc6a97004678aac9519820e6e6e9e08066888c6894f22181d4f13fe4db4ee4f95a560f4ae401c1c149cecf7bdad4e82e03a15c220f2ec49a8fee1430fb7204685351785aba0160fc253432248f19d8d8cc7433c946f5ff9c17f81e7f2a082d615b3045300f09cbb7ee37;
    5'b01110 : xpb = 1024'h1f456a01acf7bcab5a4490420588f8c6f513d6c160adf4cabffd9539c5b1a041fc4d0253eda0ee4f4101b8f68457fa4e73e4c7dcd1df363b1e0e21ce1042ce9d999f2acb565066293d4437f01a8ff8dcc60dbf8685b5bfa7caa798773bb05bf4afc57df7a85b657455d3d4552655a6983a99b4905e6ea472c614f245f99c6ae1;
    5'b01111 : xpb = 1024'h2e1fe43ec72cbba15cee6c43d03dc67f8eaff89bd242ed2ae8fae3fae099eeebd7b31dbdfac17615f59adcfae72e1faba7e4b46abec512202cd15f9a5ec4536c63c27ac1c472c8b11e6660b1708561cb77ea839b07032bfe1cf476ed166492b52d666cd577ddfe7477de61b44d0f353856b43f188f7bedb546f9d5822780e78b;
    5'b10000 : xpb = 1024'h3cfa5e7be161ba975f9848459af29438284c1a7643d7e58b11f832bbfb823d95b319392807e1fddcaa3400ff4a044508dbe4a0f8abaaee053b949d66ad45d83b2de5cab832952b38ff888972c67acaba29c747af885098546f415562f118c975ab075bb34760977499e8ef1373c8c3d872cec9a0c08936f7c7deb8be55656435;
    5'b10001 : xpb = 1024'h4bd4d8b8fb96b98d6242244765a761f0c1e83c50b56cddeb3af5817d166a8c3f8e7f5492150285a35ecd2503acda6a660fe48d869890c9ea4a57db32fbc75d09f8091aaea0b78dc0e0aab2341c7033a8dba40bc4099e04aac18e33d8cbcd003628a84a9116e33074bbf37c729a8252788ee95428f196803a48c39bfa8349e0df;
    5'b10010 : xpb = 1024'h5aaf52f615cbb88364ec0049305c2fa95b845e2b2701d64b63f2d03e3152dae969e56ffc22230d6a136649080fb08fc343e47a148576a5cf591b18ff4a48e1d8c22c6aa50ed9f048c1ccdaf572659c978d80cfd88aeb710113db124ea68136f6a649396ee665c974ddfe09d1c13be118ab03deb122a3c97cc9a87f36b12e5d89;
    5'b10011 : xpb = 1024'h6989cd333000b7796795dc4afb10fd61f52080059896ceab8cf01eff4c3b2993454b8b662f439530c7ff6d0c7286b52077e466a2725c81b467de56cb98ca66a78c4fba9b7cfc52d0a2ef03b6c85b05863f5d93ed0c38dd576627f0c481356db723ea284cb5e8627500089730e7f56fb8c71e693953b112bf4a8d6272df12da33;
    5'b10100 : xpb = 1024'h786447704a35b66f6a3fb84cc5c5cb1a8ebca1e00a2bc70bb5ed6dc06723783d20b1a6d03c641cf77c989110d55cda7dabe453305f425d9976a19497e74beb7656730a91eb1eb55884112c781e506e74f13a58018d8649adb874cf3a5be9a477a18b172a856afb75221324900eaefe58e338f3c184be5c01cb7245af0cf756dd;
    5'b10101 : xpb = 1024'h873ec1ad646ab5656ce9944e907a98d32858c3ba7bc0bf6bdeeabc81820bc6e6fc17c23a4984a4be3131b5153832ffdadfe43fbe4c28397e8564d26435cd704520965a88594117e0653355397445d763a3171c160ed3b6040ac1adb0369ddb381f2c060854ed9475441db1ef35688cf8ff537e49b5cba5444c5728eb3adbd387;
    5'b10110 : xpb = 1024'h96193bea7e9fb45b6f9370505b2f668bc1f4e594ed55b7cc07e80b429cf41590d77ddda456a52c84e5cad9199b09253813e42c4c390e156394281030844ef513eab9aa7ec7637a6846557dfaca3b405254f3e02a9021225a5d0e8c26115211f89cccf4e624702d7566283f4e5c221b991b6e08d1e6d8ee86cd3c0c2768c05031;
    5'b10111 : xpb = 1024'ha4f3b62798d4b351723d4c5225e434445b91076f5eeab02c30e55a03b7dc643ab2e3f90e63c5b44b9a63fd1dfddf4a9547e418da25f3f148a2eb4dfcd2d079e2b4dcfa753585dcf02777a6bc2030a94106d0a43f116e8eb0af5b6a9bec0648b91a6de3c3f3f2c6758832ccad82dbaa393788935a17e637c94e20ef6396a4ccdb;
    5'b11000 : xpb = 1024'h320eb0ef11b7d7ea9e1b07ce03ebaab83b72618fb080814dc05ef6f1fc205dc8b0196ffa6bfbd83af9ee1db7d575f2817c9dd81f026fce2010f4c6ae67f8a000ab115bcf4174232f5ffccdadd4a4dfec4a86ebb0635cdf64c1bb7170c8fdce76907407812ac66e8237d732db1c512b004c93efff8a823db8896579b3ba6e31a;
    5'b11001 : xpb = 1024'h11fb654c0b507c74ac8b8c7eaaf388641d5347f36c9d007505033e303aaa54866667b269b3e0454a643805dfe02d84854bc9ca0fdd0cd8c70fd28a3735010eced4d465b36239a4bad721f59c333fb6ed768532cf87833a4c9e68958ce74413a7e6a82f55e22effe84588008cd87ea15020e3c98829b56d1e097b3ad7698b5fc4;
    5'b11010 : xpb = 1024'h20d5df8925857b6aaf35688075a8561cb6ef69cdde31f8d52e008cf15592a33041cdcdd3c100cd1118d129e44303a9e27fc9b69dc9f2b4ac1e95c8038382939d9ef7b5a9d05c0742b8441e5d89351fdc2861f6e408d0a6a2f0b57402c1f84a6864491e33b1b198e867928debff382ff03cfe54105ac2b6608a601e13976fdc6e;
    5'b11011 : xpb = 1024'h2fb059c63fba7a60b1df4482405d23d5508b8ba84fc6f13556fddbb2707af1da1d33e93dce2154d7cd6a4de8a5d9cf3fb3c9a32bb6d890912d5905cfd204186c691b05a03e7e69ca9966471edf2a88cada3ebaf88a1e12f9430252789cac8128e1ea0d11813431e8899d1b4b25f1be905918de988bcfffa30b45014fc5545918;
    5'b11100 : xpb = 1024'h3e8ad40359ef7956b48920840b11f18dea27ad82c15be9957ffb2a738b634083f89a04a7db41dc9e820371ed08aff49ce7c98fb9a3be6c763c1c439c20859d3b333e5596aca0cc527a886fe0351ff1b98c1b7f0d0b6b7f4f954f30ee7760b7e95f8afbef50b6cae8aba7a8aa4cab4d3075336920bcdd48e58c29e48bf338d5c2;
    5'b11101 : xpb = 1024'h4d654e407424784cb732fc85d5c6bf4683c3cf5d32f0e1f5a8f87934a64b8f2dd4002011e8626465369c95f16b8619fa1bc97c4790a4485b4adf81686f072209fd61a58d1ac32eda5baa98a18b155aa83df843218cb8eba5e79c0f645214eea9dd2beacd203963e8cdb236097364dbd0914df3a8edea92280d0ec7c8211d526c;
    5'b11110 : xpb = 1024'h5c3fc87d8e597742b9dcd887a07b8cff1d5ff137a485da55d1f5c7f5c133ddd7af663b7bf582ec2beb35b9f5ce5c3f574fc968d57d8a244059a2bf34bd88a6d8c784f58388e591623cccc162e10ac396efd507360e0657fc39e8edda2cc9256a5accd9aaefbbfce8efbcc3689a1e6a70ad687e311ef7db6a8df3ab044f01cf16;
    5'b11111 : xpb = 1024'h6b1a42baa88e7638bc86b4896b305ab7b6fc1312161ad2b5faf316b6dc1c2c818acc56e602a373f29fceddfa313264b483c955636a7000256865fd010c0a2ba791a84579f707f3ea1deeea2437002c85a1b1cb4a8f53c4528c35cc50077d5c2ad86dc888bf3e95e911c750c7c0d7f910c98308b9500524ad0ed88e407ce64bc0;
    endcase
end

endmodule

module first_reduction_data
(
    input clk,
    input [1023:0] partial_product_high0,
    input [1023:0] partial_product_high1,
    input [1032:0] partial_product_low0,
    input [1032:0] partial_product_low1,

    output [511:0] col_out_0,
    output [511:0] col_out_1,
    output [511:0] col_out_2,
    output [511:0] col_out_3,
    output [511:0] col_out_4,
    output [511:0] col_out_5,
    output [511:0] col_out_6,
    output [511:0] col_out_7,
    output [511:0] col_out_8,
    output [511:0] col_out_9,
    output [511:0] col_out_10,
    output [511:0] col_out_11,
    output [511:0] col_out_12,
    output [511:0] col_out_13,
    output [511:0] col_out_14,
    output [511:0] col_out_15,
    output [511:0] col_out_16,
    output [511:0] col_out_17,
    output [511:0] col_out_18,
    output [511:0] col_out_19,
    output [511:0] col_out_20,
    output [511:0] col_out_21,
    output [511:0] col_out_22,
    output [511:0] col_out_23,
    output [511:0] col_out_24,
    output [511:0] col_out_25,
    output [511:0] col_out_26,
    output [511:0] col_out_27,
    output [511:0] col_out_28,
    output [511:0] col_out_29,
    output [511:0] col_out_30,
    output [511:0] col_out_31,
    output [511:0] col_out_32,
    output [511:0] col_out_33,
    output [511:0] col_out_34,
    output [511:0] col_out_35,
    output [511:0] col_out_36,
    output [511:0] col_out_37,
    output [511:0] col_out_38,
    output [511:0] col_out_39,
    output [511:0] col_out_40,
    output [511:0] col_out_41,
    output [511:0] col_out_42,
    output [511:0] col_out_43,
    output [511:0] col_out_44,
    output [511:0] col_out_45,
    output [511:0] col_out_46,
    output [511:0] col_out_47,
    output [511:0] col_out_48,
    output [511:0] col_out_49,
    output [511:0] col_out_50,
    output [511:0] col_out_51,
    output [511:0] col_out_52,
    output [511:0] col_out_53,
    output [511:0] col_out_54,
    output [511:0] col_out_55,
    output [511:0] col_out_56,
    output [511:0] col_out_57,
    output [511:0] col_out_58,
    output [511:0] col_out_59,
    output [511:0] col_out_60,
    output [511:0] col_out_61,
    output [511:0] col_out_62,
    output [511:0] col_out_63,
    output [511:0] col_out_64,
    output [511:0] col_out_65,
    output [511:0] col_out_66,
    output [511:0] col_out_67,
    output [511:0] col_out_68,
    output [511:0] col_out_69,
    output [511:0] col_out_70,
    output [511:0] col_out_71,
    output [511:0] col_out_72,
    output [511:0] col_out_73,
    output [511:0] col_out_74,
    output [511:0] col_out_75,
    output [511:0] col_out_76,
    output [511:0] col_out_77,
    output [511:0] col_out_78,
    output [511:0] col_out_79,
    output [511:0] col_out_80,
    output [511:0] col_out_81,
    output [511:0] col_out_82,
    output [511:0] col_out_83,
    output [511:0] col_out_84,
    output [511:0] col_out_85,
    output [511:0] col_out_86,
    output [511:0] col_out_87,
    output [511:0] col_out_88,
    output [511:0] col_out_89,
    output [511:0] col_out_90,
    output [511:0] col_out_91,
    output [511:0] col_out_92,
    output [511:0] col_out_93,
    output [511:0] col_out_94,
    output [511:0] col_out_95,
    output [511:0] col_out_96,
    output [511:0] col_out_97,
    output [511:0] col_out_98,
    output [511:0] col_out_99,
    output [511:0] col_out_100,
    output [511:0] col_out_101,
    output [511:0] col_out_102,
    output [511:0] col_out_103,
    output [511:0] col_out_104,
    output [511:0] col_out_105,
    output [511:0] col_out_106,
    output [511:0] col_out_107,
    output [511:0] col_out_108,
    output [511:0] col_out_109,
    output [511:0] col_out_110,
    output [511:0] col_out_111,
    output [511:0] col_out_112,
    output [511:0] col_out_113,
    output [511:0] col_out_114,
    output [511:0] col_out_115,
    output [511:0] col_out_116,
    output [511:0] col_out_117,
    output [511:0] col_out_118,
    output [511:0] col_out_119,
    output [511:0] col_out_120,
    output [511:0] col_out_121,
    output [511:0] col_out_122,
    output [511:0] col_out_123,
    output [511:0] col_out_124,
    output [511:0] col_out_125,
    output [511:0] col_out_126,
    output [511:0] col_out_127,
    output [511:0] col_out_128,
    output [511:0] col_out_129,
    output [511:0] col_out_130,
    output [511:0] col_out_131,
    output [511:0] col_out_132,
    output [511:0] col_out_133,
    output [511:0] col_out_134,
    output [511:0] col_out_135,
    output [511:0] col_out_136,
    output [511:0] col_out_137,
    output [511:0] col_out_138,
    output [511:0] col_out_139,
    output [511:0] col_out_140,
    output [511:0] col_out_141,
    output [511:0] col_out_142,
    output [511:0] col_out_143,
    output [511:0] col_out_144,
    output [511:0] col_out_145,
    output [511:0] col_out_146,
    output [511:0] col_out_147,
    output [511:0] col_out_148,
    output [511:0] col_out_149,
    output [511:0] col_out_150,
    output [511:0] col_out_151,
    output [511:0] col_out_152,
    output [511:0] col_out_153,
    output [511:0] col_out_154,
    output [511:0] col_out_155,
    output [511:0] col_out_156,
    output [511:0] col_out_157,
    output [511:0] col_out_158,
    output [511:0] col_out_159,
    output [511:0] col_out_160,
    output [511:0] col_out_161,
    output [511:0] col_out_162,
    output [511:0] col_out_163,
    output [511:0] col_out_164,
    output [511:0] col_out_165,
    output [511:0] col_out_166,
    output [511:0] col_out_167,
    output [511:0] col_out_168,
    output [511:0] col_out_169,
    output [511:0] col_out_170,
    output [511:0] col_out_171,
    output [511:0] col_out_172,
    output [511:0] col_out_173,
    output [511:0] col_out_174,
    output [511:0] col_out_175,
    output [511:0] col_out_176,
    output [511:0] col_out_177,
    output [511:0] col_out_178,
    output [511:0] col_out_179,
    output [511:0] col_out_180,
    output [511:0] col_out_181,
    output [511:0] col_out_182,
    output [511:0] col_out_183,
    output [511:0] col_out_184,
    output [511:0] col_out_185,
    output [511:0] col_out_186,
    output [511:0] col_out_187,
    output [511:0] col_out_188,
    output [511:0] col_out_189,
    output [511:0] col_out_190,
    output [511:0] col_out_191,
    output [511:0] col_out_192,
    output [511:0] col_out_193,
    output [511:0] col_out_194,
    output [511:0] col_out_195,
    output [511:0] col_out_196,
    output [511:0] col_out_197,
    output [511:0] col_out_198,
    output [511:0] col_out_199,
    output [511:0] col_out_200,
    output [511:0] col_out_201,
    output [511:0] col_out_202,
    output [511:0] col_out_203,
    output [511:0] col_out_204,
    output [511:0] col_out_205,
    output [511:0] col_out_206,
    output [511:0] col_out_207,
    output [511:0] col_out_208,
    output [511:0] col_out_209,
    output [511:0] col_out_210,
    output [511:0] col_out_211,
    output [511:0] col_out_212,
    output [511:0] col_out_213,
    output [511:0] col_out_214,
    output [511:0] col_out_215,
    output [511:0] col_out_216,
    output [511:0] col_out_217,
    output [511:0] col_out_218,
    output [511:0] col_out_219,
    output [511:0] col_out_220,
    output [511:0] col_out_221,
    output [511:0] col_out_222,
    output [511:0] col_out_223,
    output [511:0] col_out_224,
    output [511:0] col_out_225,
    output [511:0] col_out_226,
    output [511:0] col_out_227,
    output [511:0] col_out_228,
    output [511:0] col_out_229,
    output [511:0] col_out_230,
    output [511:0] col_out_231,
    output [511:0] col_out_232,
    output [511:0] col_out_233,
    output [511:0] col_out_234,
    output [511:0] col_out_235,
    output [511:0] col_out_236,
    output [511:0] col_out_237,
    output [511:0] col_out_238,
    output [511:0] col_out_239,
    output [511:0] col_out_240,
    output [511:0] col_out_241,
    output [511:0] col_out_242,
    output [511:0] col_out_243,
    output [511:0] col_out_244,
    output [511:0] col_out_245,
    output [511:0] col_out_246,
    output [511:0] col_out_247,
    output [511:0] col_out_248,
    output [511:0] col_out_249,
    output [511:0] col_out_250,
    output [511:0] col_out_251,
    output [511:0] col_out_252,
    output [511:0] col_out_253,
    output [511:0] col_out_254,
    output [511:0] col_out_255,
    output [511:0] col_out_256,
    output [511:0] col_out_257,
    output [511:0] col_out_258,
    output [511:0] col_out_259,
    output [511:0] col_out_260,
    output [511:0] col_out_261,
    output [511:0] col_out_262,
    output [511:0] col_out_263,
    output [511:0] col_out_264,
    output [511:0] col_out_265,
    output [511:0] col_out_266,
    output [511:0] col_out_267,
    output [511:0] col_out_268,
    output [511:0] col_out_269,
    output [511:0] col_out_270,
    output [511:0] col_out_271,
    output [511:0] col_out_272,
    output [511:0] col_out_273,
    output [511:0] col_out_274,
    output [511:0] col_out_275,
    output [511:0] col_out_276,
    output [511:0] col_out_277,
    output [511:0] col_out_278,
    output [511:0] col_out_279,
    output [511:0] col_out_280,
    output [511:0] col_out_281,
    output [511:0] col_out_282,
    output [511:0] col_out_283,
    output [511:0] col_out_284,
    output [511:0] col_out_285,
    output [511:0] col_out_286,
    output [511:0] col_out_287,
    output [511:0] col_out_288,
    output [511:0] col_out_289,
    output [511:0] col_out_290,
    output [511:0] col_out_291,
    output [511:0] col_out_292,
    output [511:0] col_out_293,
    output [511:0] col_out_294,
    output [511:0] col_out_295,
    output [511:0] col_out_296,
    output [511:0] col_out_297,
    output [511:0] col_out_298,
    output [511:0] col_out_299,
    output [511:0] col_out_300,
    output [511:0] col_out_301,
    output [511:0] col_out_302,
    output [511:0] col_out_303,
    output [511:0] col_out_304,
    output [511:0] col_out_305,
    output [511:0] col_out_306,
    output [511:0] col_out_307,
    output [511:0] col_out_308,
    output [511:0] col_out_309,
    output [511:0] col_out_310,
    output [511:0] col_out_311,
    output [511:0] col_out_312,
    output [511:0] col_out_313,
    output [511:0] col_out_314,
    output [511:0] col_out_315,
    output [511:0] col_out_316,
    output [511:0] col_out_317,
    output [511:0] col_out_318,
    output [511:0] col_out_319,
    output [511:0] col_out_320,
    output [511:0] col_out_321,
    output [511:0] col_out_322,
    output [511:0] col_out_323,
    output [511:0] col_out_324,
    output [511:0] col_out_325,
    output [511:0] col_out_326,
    output [511:0] col_out_327,
    output [511:0] col_out_328,
    output [511:0] col_out_329,
    output [511:0] col_out_330,
    output [511:0] col_out_331,
    output [511:0] col_out_332,
    output [511:0] col_out_333,
    output [511:0] col_out_334,
    output [511:0] col_out_335,
    output [511:0] col_out_336,
    output [511:0] col_out_337,
    output [511:0] col_out_338,
    output [511:0] col_out_339,
    output [511:0] col_out_340,
    output [511:0] col_out_341,
    output [511:0] col_out_342,
    output [511:0] col_out_343,
    output [511:0] col_out_344,
    output [511:0] col_out_345,
    output [511:0] col_out_346,
    output [511:0] col_out_347,
    output [511:0] col_out_348,
    output [511:0] col_out_349,
    output [511:0] col_out_350,
    output [511:0] col_out_351,
    output [511:0] col_out_352,
    output [511:0] col_out_353,
    output [511:0] col_out_354,
    output [511:0] col_out_355,
    output [511:0] col_out_356,
    output [511:0] col_out_357,
    output [511:0] col_out_358,
    output [511:0] col_out_359,
    output [511:0] col_out_360,
    output [511:0] col_out_361,
    output [511:0] col_out_362,
    output [511:0] col_out_363,
    output [511:0] col_out_364,
    output [511:0] col_out_365,
    output [511:0] col_out_366,
    output [511:0] col_out_367,
    output [511:0] col_out_368,
    output [511:0] col_out_369,
    output [511:0] col_out_370,
    output [511:0] col_out_371,
    output [511:0] col_out_372,
    output [511:0] col_out_373,
    output [511:0] col_out_374,
    output [511:0] col_out_375,
    output [511:0] col_out_376,
    output [511:0] col_out_377,
    output [511:0] col_out_378,
    output [511:0] col_out_379,
    output [511:0] col_out_380,
    output [511:0] col_out_381,
    output [511:0] col_out_382,
    output [511:0] col_out_383,
    output [511:0] col_out_384,
    output [511:0] col_out_385,
    output [511:0] col_out_386,
    output [511:0] col_out_387,
    output [511:0] col_out_388,
    output [511:0] col_out_389,
    output [511:0] col_out_390,
    output [511:0] col_out_391,
    output [511:0] col_out_392,
    output [511:0] col_out_393,
    output [511:0] col_out_394,
    output [511:0] col_out_395,
    output [511:0] col_out_396,
    output [511:0] col_out_397,
    output [511:0] col_out_398,
    output [511:0] col_out_399,
    output [511:0] col_out_400,
    output [511:0] col_out_401,
    output [511:0] col_out_402,
    output [511:0] col_out_403,
    output [511:0] col_out_404,
    output [511:0] col_out_405,
    output [511:0] col_out_406,
    output [511:0] col_out_407,
    output [511:0] col_out_408,
    output [511:0] col_out_409,
    output [511:0] col_out_410,
    output [511:0] col_out_411,
    output [511:0] col_out_412,
    output [511:0] col_out_413,
    output [511:0] col_out_414,
    output [511:0] col_out_415,
    output [511:0] col_out_416,
    output [511:0] col_out_417,
    output [511:0] col_out_418,
    output [511:0] col_out_419,
    output [511:0] col_out_420,
    output [511:0] col_out_421,
    output [511:0] col_out_422,
    output [511:0] col_out_423,
    output [511:0] col_out_424,
    output [511:0] col_out_425,
    output [511:0] col_out_426,
    output [511:0] col_out_427,
    output [511:0] col_out_428,
    output [511:0] col_out_429,
    output [511:0] col_out_430,
    output [511:0] col_out_431,
    output [511:0] col_out_432,
    output [511:0] col_out_433,
    output [511:0] col_out_434,
    output [511:0] col_out_435,
    output [511:0] col_out_436,
    output [511:0] col_out_437,
    output [511:0] col_out_438,
    output [511:0] col_out_439,
    output [511:0] col_out_440,
    output [511:0] col_out_441,
    output [511:0] col_out_442,
    output [511:0] col_out_443,
    output [511:0] col_out_444,
    output [511:0] col_out_445,
    output [511:0] col_out_446,
    output [511:0] col_out_447,
    output [511:0] col_out_448,
    output [511:0] col_out_449,
    output [511:0] col_out_450,
    output [511:0] col_out_451,
    output [511:0] col_out_452,
    output [511:0] col_out_453,
    output [511:0] col_out_454,
    output [511:0] col_out_455,
    output [511:0] col_out_456,
    output [511:0] col_out_457,
    output [511:0] col_out_458,
    output [511:0] col_out_459,
    output [511:0] col_out_460,
    output [511:0] col_out_461,
    output [511:0] col_out_462,
    output [511:0] col_out_463,
    output [511:0] col_out_464,
    output [511:0] col_out_465,
    output [511:0] col_out_466,
    output [511:0] col_out_467,
    output [511:0] col_out_468,
    output [511:0] col_out_469,
    output [511:0] col_out_470,
    output [511:0] col_out_471,
    output [511:0] col_out_472,
    output [511:0] col_out_473,
    output [511:0] col_out_474,
    output [511:0] col_out_475,
    output [511:0] col_out_476,
    output [511:0] col_out_477,
    output [511:0] col_out_478,
    output [511:0] col_out_479,
    output [511:0] col_out_480,
    output [511:0] col_out_481,
    output [511:0] col_out_482,
    output [511:0] col_out_483,
    output [511:0] col_out_484,
    output [511:0] col_out_485,
    output [511:0] col_out_486,
    output [511:0] col_out_487,
    output [511:0] col_out_488,
    output [511:0] col_out_489,
    output [511:0] col_out_490,
    output [511:0] col_out_491,
    output [511:0] col_out_492,
    output [511:0] col_out_493,
    output [511:0] col_out_494,
    output [511:0] col_out_495,
    output [511:0] col_out_496,
    output [511:0] col_out_497,
    output [511:0] col_out_498,
    output [511:0] col_out_499,
    output [511:0] col_out_500,
    output [511:0] col_out_501,
    output [511:0] col_out_502,
    output [511:0] col_out_503,
    output [511:0] col_out_504,
    output [511:0] col_out_505,
    output [511:0] col_out_506,
    output [511:0] col_out_507,
    output [511:0] col_out_508,
    output [511:0] col_out_509,
    output [511:0] col_out_510,
    output [511:0] col_out_511,
    output [511:0] col_out_512,
    output [511:0] col_out_513,
    output [511:0] col_out_514,
    output [511:0] col_out_515,
    output [511:0] col_out_516,
    output [511:0] col_out_517,
    output [511:0] col_out_518,
    output [511:0] col_out_519,
    output [511:0] col_out_520,
    output [511:0] col_out_521,
    output [511:0] col_out_522,
    output [511:0] col_out_523,
    output [511:0] col_out_524,
    output [511:0] col_out_525,
    output [511:0] col_out_526,
    output [511:0] col_out_527,
    output [511:0] col_out_528,
    output [511:0] col_out_529,
    output [511:0] col_out_530,
    output [511:0] col_out_531,
    output [511:0] col_out_532,
    output [511:0] col_out_533,
    output [511:0] col_out_534,
    output [511:0] col_out_535,
    output [511:0] col_out_536,
    output [511:0] col_out_537,
    output [511:0] col_out_538,
    output [511:0] col_out_539,
    output [511:0] col_out_540,
    output [511:0] col_out_541,
    output [511:0] col_out_542,
    output [511:0] col_out_543,
    output [511:0] col_out_544,
    output [511:0] col_out_545,
    output [511:0] col_out_546,
    output [511:0] col_out_547,
    output [511:0] col_out_548,
    output [511:0] col_out_549,
    output [511:0] col_out_550,
    output [511:0] col_out_551,
    output [511:0] col_out_552,
    output [511:0] col_out_553,
    output [511:0] col_out_554,
    output [511:0] col_out_555,
    output [511:0] col_out_556,
    output [511:0] col_out_557,
    output [511:0] col_out_558,
    output [511:0] col_out_559,
    output [511:0] col_out_560,
    output [511:0] col_out_561,
    output [511:0] col_out_562,
    output [511:0] col_out_563,
    output [511:0] col_out_564,
    output [511:0] col_out_565,
    output [511:0] col_out_566,
    output [511:0] col_out_567,
    output [511:0] col_out_568,
    output [511:0] col_out_569,
    output [511:0] col_out_570,
    output [511:0] col_out_571,
    output [511:0] col_out_572,
    output [511:0] col_out_573,
    output [511:0] col_out_574,
    output [511:0] col_out_575,
    output [511:0] col_out_576,
    output [511:0] col_out_577,
    output [511:0] col_out_578,
    output [511:0] col_out_579,
    output [511:0] col_out_580,
    output [511:0] col_out_581,
    output [511:0] col_out_582,
    output [511:0] col_out_583,
    output [511:0] col_out_584,
    output [511:0] col_out_585,
    output [511:0] col_out_586,
    output [511:0] col_out_587,
    output [511:0] col_out_588,
    output [511:0] col_out_589,
    output [511:0] col_out_590,
    output [511:0] col_out_591,
    output [511:0] col_out_592,
    output [511:0] col_out_593,
    output [511:0] col_out_594,
    output [511:0] col_out_595,
    output [511:0] col_out_596,
    output [511:0] col_out_597,
    output [511:0] col_out_598,
    output [511:0] col_out_599,
    output [511:0] col_out_600,
    output [511:0] col_out_601,
    output [511:0] col_out_602,
    output [511:0] col_out_603,
    output [511:0] col_out_604,
    output [511:0] col_out_605,
    output [511:0] col_out_606,
    output [511:0] col_out_607,
    output [511:0] col_out_608,
    output [511:0] col_out_609,
    output [511:0] col_out_610,
    output [511:0] col_out_611,
    output [511:0] col_out_612,
    output [511:0] col_out_613,
    output [511:0] col_out_614,
    output [511:0] col_out_615,
    output [511:0] col_out_616,
    output [511:0] col_out_617,
    output [511:0] col_out_618,
    output [511:0] col_out_619,
    output [511:0] col_out_620,
    output [511:0] col_out_621,
    output [511:0] col_out_622,
    output [511:0] col_out_623,
    output [511:0] col_out_624,
    output [511:0] col_out_625,
    output [511:0] col_out_626,
    output [511:0] col_out_627,
    output [511:0] col_out_628,
    output [511:0] col_out_629,
    output [511:0] col_out_630,
    output [511:0] col_out_631,
    output [511:0] col_out_632,
    output [511:0] col_out_633,
    output [511:0] col_out_634,
    output [511:0] col_out_635,
    output [511:0] col_out_636,
    output [511:0] col_out_637,
    output [511:0] col_out_638,
    output [511:0] col_out_639,
    output [511:0] col_out_640,
    output [511:0] col_out_641,
    output [511:0] col_out_642,
    output [511:0] col_out_643,
    output [511:0] col_out_644,
    output [511:0] col_out_645,
    output [511:0] col_out_646,
    output [511:0] col_out_647,
    output [511:0] col_out_648,
    output [511:0] col_out_649,
    output [511:0] col_out_650,
    output [511:0] col_out_651,
    output [511:0] col_out_652,
    output [511:0] col_out_653,
    output [511:0] col_out_654,
    output [511:0] col_out_655,
    output [511:0] col_out_656,
    output [511:0] col_out_657,
    output [511:0] col_out_658,
    output [511:0] col_out_659,
    output [511:0] col_out_660,
    output [511:0] col_out_661,
    output [511:0] col_out_662,
    output [511:0] col_out_663,
    output [511:0] col_out_664,
    output [511:0] col_out_665,
    output [511:0] col_out_666,
    output [511:0] col_out_667,
    output [511:0] col_out_668,
    output [511:0] col_out_669,
    output [511:0] col_out_670,
    output [511:0] col_out_671,
    output [511:0] col_out_672,
    output [511:0] col_out_673,
    output [511:0] col_out_674,
    output [511:0] col_out_675,
    output [511:0] col_out_676,
    output [511:0] col_out_677,
    output [511:0] col_out_678,
    output [511:0] col_out_679,
    output [511:0] col_out_680,
    output [511:0] col_out_681,
    output [511:0] col_out_682,
    output [511:0] col_out_683,
    output [511:0] col_out_684,
    output [511:0] col_out_685,
    output [511:0] col_out_686,
    output [511:0] col_out_687,
    output [511:0] col_out_688,
    output [511:0] col_out_689,
    output [511:0] col_out_690,
    output [511:0] col_out_691,
    output [511:0] col_out_692,
    output [511:0] col_out_693,
    output [511:0] col_out_694,
    output [511:0] col_out_695,
    output [511:0] col_out_696,
    output [511:0] col_out_697,
    output [511:0] col_out_698,
    output [511:0] col_out_699,
    output [511:0] col_out_700,
    output [511:0] col_out_701,
    output [511:0] col_out_702,
    output [511:0] col_out_703,
    output [511:0] col_out_704,
    output [511:0] col_out_705,
    output [511:0] col_out_706,
    output [511:0] col_out_707,
    output [511:0] col_out_708,
    output [511:0] col_out_709,
    output [511:0] col_out_710,
    output [511:0] col_out_711,
    output [511:0] col_out_712,
    output [511:0] col_out_713,
    output [511:0] col_out_714,
    output [511:0] col_out_715,
    output [511:0] col_out_716,
    output [511:0] col_out_717,
    output [511:0] col_out_718,
    output [511:0] col_out_719,
    output [511:0] col_out_720,
    output [511:0] col_out_721,
    output [511:0] col_out_722,
    output [511:0] col_out_723,
    output [511:0] col_out_724,
    output [511:0] col_out_725,
    output [511:0] col_out_726,
    output [511:0] col_out_727,
    output [511:0] col_out_728,
    output [511:0] col_out_729,
    output [511:0] col_out_730,
    output [511:0] col_out_731,
    output [511:0] col_out_732,
    output [511:0] col_out_733,
    output [511:0] col_out_734,
    output [511:0] col_out_735,
    output [511:0] col_out_736,
    output [511:0] col_out_737,
    output [511:0] col_out_738,
    output [511:0] col_out_739,
    output [511:0] col_out_740,
    output [511:0] col_out_741,
    output [511:0] col_out_742,
    output [511:0] col_out_743,
    output [511:0] col_out_744,
    output [511:0] col_out_745,
    output [511:0] col_out_746,
    output [511:0] col_out_747,
    output [511:0] col_out_748,
    output [511:0] col_out_749,
    output [511:0] col_out_750,
    output [511:0] col_out_751,
    output [511:0] col_out_752,
    output [511:0] col_out_753,
    output [511:0] col_out_754,
    output [511:0] col_out_755,
    output [511:0] col_out_756,
    output [511:0] col_out_757,
    output [511:0] col_out_758,
    output [511:0] col_out_759,
    output [511:0] col_out_760,
    output [511:0] col_out_761,
    output [511:0] col_out_762,
    output [511:0] col_out_763,
    output [511:0] col_out_764,
    output [511:0] col_out_765,
    output [511:0] col_out_766,
    output [511:0] col_out_767,
    output [511:0] col_out_768,
    output [511:0] col_out_769,
    output [511:0] col_out_770,
    output [511:0] col_out_771,
    output [511:0] col_out_772,
    output [511:0] col_out_773,
    output [511:0] col_out_774,
    output [511:0] col_out_775,
    output [511:0] col_out_776,
    output [511:0] col_out_777,
    output [511:0] col_out_778,
    output [511:0] col_out_779,
    output [511:0] col_out_780,
    output [511:0] col_out_781,
    output [511:0] col_out_782,
    output [511:0] col_out_783,
    output [511:0] col_out_784,
    output [511:0] col_out_785,
    output [511:0] col_out_786,
    output [511:0] col_out_787,
    output [511:0] col_out_788,
    output [511:0] col_out_789,
    output [511:0] col_out_790,
    output [511:0] col_out_791,
    output [511:0] col_out_792,
    output [511:0] col_out_793,
    output [511:0] col_out_794,
    output [511:0] col_out_795,
    output [511:0] col_out_796,
    output [511:0] col_out_797,
    output [511:0] col_out_798,
    output [511:0] col_out_799,
    output [511:0] col_out_800,
    output [511:0] col_out_801,
    output [511:0] col_out_802,
    output [511:0] col_out_803,
    output [511:0] col_out_804,
    output [511:0] col_out_805,
    output [511:0] col_out_806,
    output [511:0] col_out_807,
    output [511:0] col_out_808,
    output [511:0] col_out_809,
    output [511:0] col_out_810,
    output [511:0] col_out_811,
    output [511:0] col_out_812,
    output [511:0] col_out_813,
    output [511:0] col_out_814,
    output [511:0] col_out_815,
    output [511:0] col_out_816,
    output [511:0] col_out_817,
    output [511:0] col_out_818,
    output [511:0] col_out_819,
    output [511:0] col_out_820,
    output [511:0] col_out_821,
    output [511:0] col_out_822,
    output [511:0] col_out_823,
    output [511:0] col_out_824,
    output [511:0] col_out_825,
    output [511:0] col_out_826,
    output [511:0] col_out_827,
    output [511:0] col_out_828,
    output [511:0] col_out_829,
    output [511:0] col_out_830,
    output [511:0] col_out_831,
    output [511:0] col_out_832,
    output [511:0] col_out_833,
    output [511:0] col_out_834,
    output [511:0] col_out_835,
    output [511:0] col_out_836,
    output [511:0] col_out_837,
    output [511:0] col_out_838,
    output [511:0] col_out_839,
    output [511:0] col_out_840,
    output [511:0] col_out_841,
    output [511:0] col_out_842,
    output [511:0] col_out_843,
    output [511:0] col_out_844,
    output [511:0] col_out_845,
    output [511:0] col_out_846,
    output [511:0] col_out_847,
    output [511:0] col_out_848,
    output [511:0] col_out_849,
    output [511:0] col_out_850,
    output [511:0] col_out_851,
    output [511:0] col_out_852,
    output [511:0] col_out_853,
    output [511:0] col_out_854,
    output [511:0] col_out_855,
    output [511:0] col_out_856,
    output [511:0] col_out_857,
    output [511:0] col_out_858,
    output [511:0] col_out_859,
    output [511:0] col_out_860,
    output [511:0] col_out_861,
    output [511:0] col_out_862,
    output [511:0] col_out_863,
    output [511:0] col_out_864,
    output [511:0] col_out_865,
    output [511:0] col_out_866,
    output [511:0] col_out_867,
    output [511:0] col_out_868,
    output [511:0] col_out_869,
    output [511:0] col_out_870,
    output [511:0] col_out_871,
    output [511:0] col_out_872,
    output [511:0] col_out_873,
    output [511:0] col_out_874,
    output [511:0] col_out_875,
    output [511:0] col_out_876,
    output [511:0] col_out_877,
    output [511:0] col_out_878,
    output [511:0] col_out_879,
    output [511:0] col_out_880,
    output [511:0] col_out_881,
    output [511:0] col_out_882,
    output [511:0] col_out_883,
    output [511:0] col_out_884,
    output [511:0] col_out_885,
    output [511:0] col_out_886,
    output [511:0] col_out_887,
    output [511:0] col_out_888,
    output [511:0] col_out_889,
    output [511:0] col_out_890,
    output [511:0] col_out_891,
    output [511:0] col_out_892,
    output [511:0] col_out_893,
    output [511:0] col_out_894,
    output [511:0] col_out_895,
    output [511:0] col_out_896,
    output [511:0] col_out_897,
    output [511:0] col_out_898,
    output [511:0] col_out_899,
    output [511:0] col_out_900,
    output [511:0] col_out_901,
    output [511:0] col_out_902,
    output [511:0] col_out_903,
    output [511:0] col_out_904,
    output [511:0] col_out_905,
    output [511:0] col_out_906,
    output [511:0] col_out_907,
    output [511:0] col_out_908,
    output [511:0] col_out_909,
    output [511:0] col_out_910,
    output [511:0] col_out_911,
    output [511:0] col_out_912,
    output [511:0] col_out_913,
    output [511:0] col_out_914,
    output [511:0] col_out_915,
    output [511:0] col_out_916,
    output [511:0] col_out_917,
    output [511:0] col_out_918,
    output [511:0] col_out_919,
    output [511:0] col_out_920,
    output [511:0] col_out_921,
    output [511:0] col_out_922,
    output [511:0] col_out_923,
    output [511:0] col_out_924,
    output [511:0] col_out_925,
    output [511:0] col_out_926,
    output [511:0] col_out_927,
    output [511:0] col_out_928,
    output [511:0] col_out_929,
    output [511:0] col_out_930,
    output [511:0] col_out_931,
    output [511:0] col_out_932,
    output [511:0] col_out_933,
    output [511:0] col_out_934,
    output [511:0] col_out_935,
    output [511:0] col_out_936,
    output [511:0] col_out_937,
    output [511:0] col_out_938,
    output [511:0] col_out_939,
    output [511:0] col_out_940,
    output [511:0] col_out_941,
    output [511:0] col_out_942,
    output [511:0] col_out_943,
    output [511:0] col_out_944,
    output [511:0] col_out_945,
    output [511:0] col_out_946,
    output [511:0] col_out_947,
    output [511:0] col_out_948,
    output [511:0] col_out_949,
    output [511:0] col_out_950,
    output [511:0] col_out_951,
    output [511:0] col_out_952,
    output [511:0] col_out_953,
    output [511:0] col_out_954,
    output [511:0] col_out_955,
    output [511:0] col_out_956,
    output [511:0] col_out_957,
    output [511:0] col_out_958,
    output [511:0] col_out_959,
    output [511:0] col_out_960,
    output [511:0] col_out_961,
    output [511:0] col_out_962,
    output [511:0] col_out_963,
    output [511:0] col_out_964,
    output [511:0] col_out_965,
    output [511:0] col_out_966,
    output [511:0] col_out_967,
    output [511:0] col_out_968,
    output [511:0] col_out_969,
    output [511:0] col_out_970,
    output [511:0] col_out_971,
    output [511:0] col_out_972,
    output [511:0] col_out_973,
    output [511:0] col_out_974,
    output [511:0] col_out_975,
    output [511:0] col_out_976,
    output [511:0] col_out_977,
    output [511:0] col_out_978,
    output [511:0] col_out_979,
    output [511:0] col_out_980,
    output [511:0] col_out_981,
    output [511:0] col_out_982,
    output [511:0] col_out_983,
    output [511:0] col_out_984,
    output [511:0] col_out_985,
    output [511:0] col_out_986,
    output [511:0] col_out_987,
    output [511:0] col_out_988,
    output [511:0] col_out_989,
    output [511:0] col_out_990,
    output [511:0] col_out_991,
    output [511:0] col_out_992,
    output [511:0] col_out_993,
    output [511:0] col_out_994,
    output [511:0] col_out_995,
    output [511:0] col_out_996,
    output [511:0] col_out_997,
    output [511:0] col_out_998,
    output [511:0] col_out_999,
    output [511:0] col_out_1000,
    output [511:0] col_out_1001,
    output [511:0] col_out_1002,
    output [511:0] col_out_1003,
    output [511:0] col_out_1004,
    output [511:0] col_out_1005,
    output [511:0] col_out_1006,
    output [511:0] col_out_1007,
    output [511:0] col_out_1008,
    output [511:0] col_out_1009,
    output [511:0] col_out_1010,
    output [511:0] col_out_1011,
    output [511:0] col_out_1012,
    output [511:0] col_out_1013,
    output [511:0] col_out_1014,
    output [511:0] col_out_1015,
    output [511:0] col_out_1016,
    output [511:0] col_out_1017,
    output [511:0] col_out_1018,
    output [511:0] col_out_1019,
    output [511:0] col_out_1020,
    output [511:0] col_out_1021,
    output [511:0] col_out_1022,
    output [511:0] col_out_1023
);




// xpb_2018_col Outputs
wire  [409:0]  u0_col_out_0;
wire  [409:0]  u0_col_out_1;
wire  [409:0]  u0_col_out_2;
wire  [409:0]  u0_col_out_3;
wire  [409:0]  u0_col_out_4;
wire  [409:0]  u0_col_out_5;
wire  [409:0]  u0_col_out_6;
wire  [409:0]  u0_col_out_7;
wire  [409:0]  u0_col_out_8;
wire  [409:0]  u0_col_out_9;
wire  [409:0]  u0_col_out_10;
wire  [409:0]  u0_col_out_11;
wire  [409:0]  u0_col_out_12;
wire  [409:0]  u0_col_out_13;
wire  [409:0]  u0_col_out_14;
wire  [409:0]  u0_col_out_15;
wire  [409:0]  u0_col_out_16;
wire  [409:0]  u0_col_out_17;
wire  [409:0]  u0_col_out_18;
wire  [409:0]  u0_col_out_19;
wire  [409:0]  u0_col_out_20;
wire  [409:0]  u0_col_out_21;
wire  [409:0]  u0_col_out_22;
wire  [409:0]  u0_col_out_23;
wire  [409:0]  u0_col_out_24;
wire  [409:0]  u0_col_out_25;
wire  [409:0]  u0_col_out_26;
wire  [409:0]  u0_col_out_27;
wire  [409:0]  u0_col_out_28;
wire  [409:0]  u0_col_out_29;
wire  [409:0]  u0_col_out_30;
wire  [409:0]  u0_col_out_31;
wire  [409:0]  u0_col_out_32;
wire  [409:0]  u0_col_out_33;
wire  [409:0]  u0_col_out_34;
wire  [409:0]  u0_col_out_35;
wire  [409:0]  u0_col_out_36;
wire  [409:0]  u0_col_out_37;
wire  [409:0]  u0_col_out_38;
wire  [409:0]  u0_col_out_39;
wire  [409:0]  u0_col_out_40;
wire  [409:0]  u0_col_out_41;
wire  [409:0]  u0_col_out_42;
wire  [409:0]  u0_col_out_43;
wire  [409:0]  u0_col_out_44;
wire  [409:0]  u0_col_out_45;
wire  [409:0]  u0_col_out_46;
wire  [409:0]  u0_col_out_47;
wire  [409:0]  u0_col_out_48;
wire  [409:0]  u0_col_out_49;
wire  [409:0]  u0_col_out_50;
wire  [409:0]  u0_col_out_51;
wire  [409:0]  u0_col_out_52;
wire  [409:0]  u0_col_out_53;
wire  [409:0]  u0_col_out_54;
wire  [409:0]  u0_col_out_55;
wire  [409:0]  u0_col_out_56;
wire  [409:0]  u0_col_out_57;
wire  [409:0]  u0_col_out_58;
wire  [409:0]  u0_col_out_59;
wire  [409:0]  u0_col_out_60;
wire  [409:0]  u0_col_out_61;
wire  [409:0]  u0_col_out_62;
wire  [409:0]  u0_col_out_63;
wire  [409:0]  u0_col_out_64;
wire  [409:0]  u0_col_out_65;
wire  [409:0]  u0_col_out_66;
wire  [409:0]  u0_col_out_67;
wire  [409:0]  u0_col_out_68;
wire  [409:0]  u0_col_out_69;
wire  [409:0]  u0_col_out_70;
wire  [409:0]  u0_col_out_71;
wire  [409:0]  u0_col_out_72;
wire  [409:0]  u0_col_out_73;
wire  [409:0]  u0_col_out_74;
wire  [409:0]  u0_col_out_75;
wire  [409:0]  u0_col_out_76;
wire  [409:0]  u0_col_out_77;
wire  [409:0]  u0_col_out_78;
wire  [409:0]  u0_col_out_79;
wire  [409:0]  u0_col_out_80;
wire  [409:0]  u0_col_out_81;
wire  [409:0]  u0_col_out_82;
wire  [409:0]  u0_col_out_83;
wire  [409:0]  u0_col_out_84;
wire  [409:0]  u0_col_out_85;
wire  [409:0]  u0_col_out_86;
wire  [409:0]  u0_col_out_87;
wire  [409:0]  u0_col_out_88;
wire  [409:0]  u0_col_out_89;
wire  [409:0]  u0_col_out_90;
wire  [409:0]  u0_col_out_91;
wire  [409:0]  u0_col_out_92;
wire  [409:0]  u0_col_out_93;
wire  [409:0]  u0_col_out_94;
wire  [409:0]  u0_col_out_95;
wire  [409:0]  u0_col_out_96;
wire  [409:0]  u0_col_out_97;
wire  [409:0]  u0_col_out_98;
wire  [409:0]  u0_col_out_99;
wire  [409:0]  u0_col_out_100;
wire  [409:0]  u0_col_out_101;
wire  [409:0]  u0_col_out_102;
wire  [409:0]  u0_col_out_103;
wire  [409:0]  u0_col_out_104;
wire  [409:0]  u0_col_out_105;
wire  [409:0]  u0_col_out_106;
wire  [409:0]  u0_col_out_107;
wire  [409:0]  u0_col_out_108;
wire  [409:0]  u0_col_out_109;
wire  [409:0]  u0_col_out_110;
wire  [409:0]  u0_col_out_111;
wire  [409:0]  u0_col_out_112;
wire  [409:0]  u0_col_out_113;
wire  [409:0]  u0_col_out_114;
wire  [409:0]  u0_col_out_115;
wire  [409:0]  u0_col_out_116;
wire  [409:0]  u0_col_out_117;
wire  [409:0]  u0_col_out_118;
wire  [409:0]  u0_col_out_119;
wire  [409:0]  u0_col_out_120;
wire  [409:0]  u0_col_out_121;
wire  [409:0]  u0_col_out_122;
wire  [409:0]  u0_col_out_123;
wire  [409:0]  u0_col_out_124;
wire  [409:0]  u0_col_out_125;
wire  [409:0]  u0_col_out_126;
wire  [409:0]  u0_col_out_127;
wire  [409:0]  u0_col_out_128;
wire  [409:0]  u0_col_out_129;
wire  [409:0]  u0_col_out_130;
wire  [409:0]  u0_col_out_131;
wire  [409:0]  u0_col_out_132;
wire  [409:0]  u0_col_out_133;
wire  [409:0]  u0_col_out_134;
wire  [409:0]  u0_col_out_135;
wire  [409:0]  u0_col_out_136;
wire  [409:0]  u0_col_out_137;
wire  [409:0]  u0_col_out_138;
wire  [409:0]  u0_col_out_139;
wire  [409:0]  u0_col_out_140;
wire  [409:0]  u0_col_out_141;
wire  [409:0]  u0_col_out_142;
wire  [409:0]  u0_col_out_143;
wire  [409:0]  u0_col_out_144;
wire  [409:0]  u0_col_out_145;
wire  [409:0]  u0_col_out_146;
wire  [409:0]  u0_col_out_147;
wire  [409:0]  u0_col_out_148;
wire  [409:0]  u0_col_out_149;
wire  [409:0]  u0_col_out_150;
wire  [409:0]  u0_col_out_151;
wire  [409:0]  u0_col_out_152;
wire  [409:0]  u0_col_out_153;
wire  [409:0]  u0_col_out_154;
wire  [409:0]  u0_col_out_155;
wire  [409:0]  u0_col_out_156;
wire  [409:0]  u0_col_out_157;
wire  [409:0]  u0_col_out_158;
wire  [409:0]  u0_col_out_159;
wire  [409:0]  u0_col_out_160;
wire  [409:0]  u0_col_out_161;
wire  [409:0]  u0_col_out_162;
wire  [409:0]  u0_col_out_163;
wire  [409:0]  u0_col_out_164;
wire  [409:0]  u0_col_out_165;
wire  [409:0]  u0_col_out_166;
wire  [409:0]  u0_col_out_167;
wire  [409:0]  u0_col_out_168;
wire  [409:0]  u0_col_out_169;
wire  [409:0]  u0_col_out_170;
wire  [409:0]  u0_col_out_171;
wire  [409:0]  u0_col_out_172;
wire  [409:0]  u0_col_out_173;
wire  [409:0]  u0_col_out_174;
wire  [409:0]  u0_col_out_175;
wire  [409:0]  u0_col_out_176;
wire  [409:0]  u0_col_out_177;
wire  [409:0]  u0_col_out_178;
wire  [409:0]  u0_col_out_179;
wire  [409:0]  u0_col_out_180;
wire  [409:0]  u0_col_out_181;
wire  [409:0]  u0_col_out_182;
wire  [409:0]  u0_col_out_183;
wire  [409:0]  u0_col_out_184;
wire  [409:0]  u0_col_out_185;
wire  [409:0]  u0_col_out_186;
wire  [409:0]  u0_col_out_187;
wire  [409:0]  u0_col_out_188;
wire  [409:0]  u0_col_out_189;
wire  [409:0]  u0_col_out_190;
wire  [409:0]  u0_col_out_191;
wire  [409:0]  u0_col_out_192;
wire  [409:0]  u0_col_out_193;
wire  [409:0]  u0_col_out_194;
wire  [409:0]  u0_col_out_195;
wire  [409:0]  u0_col_out_196;
wire  [409:0]  u0_col_out_197;
wire  [409:0]  u0_col_out_198;
wire  [409:0]  u0_col_out_199;
wire  [409:0]  u0_col_out_200;
wire  [409:0]  u0_col_out_201;
wire  [409:0]  u0_col_out_202;
wire  [409:0]  u0_col_out_203;
wire  [409:0]  u0_col_out_204;
wire  [409:0]  u0_col_out_205;
wire  [409:0]  u0_col_out_206;
wire  [409:0]  u0_col_out_207;
wire  [409:0]  u0_col_out_208;
wire  [409:0]  u0_col_out_209;
wire  [409:0]  u0_col_out_210;
wire  [409:0]  u0_col_out_211;
wire  [409:0]  u0_col_out_212;
wire  [409:0]  u0_col_out_213;
wire  [409:0]  u0_col_out_214;
wire  [409:0]  u0_col_out_215;
wire  [409:0]  u0_col_out_216;
wire  [409:0]  u0_col_out_217;
wire  [409:0]  u0_col_out_218;
wire  [409:0]  u0_col_out_219;
wire  [409:0]  u0_col_out_220;
wire  [409:0]  u0_col_out_221;
wire  [409:0]  u0_col_out_222;
wire  [409:0]  u0_col_out_223;
wire  [409:0]  u0_col_out_224;
wire  [409:0]  u0_col_out_225;
wire  [409:0]  u0_col_out_226;
wire  [409:0]  u0_col_out_227;
wire  [409:0]  u0_col_out_228;
wire  [409:0]  u0_col_out_229;
wire  [409:0]  u0_col_out_230;
wire  [409:0]  u0_col_out_231;
wire  [409:0]  u0_col_out_232;
wire  [409:0]  u0_col_out_233;
wire  [409:0]  u0_col_out_234;
wire  [409:0]  u0_col_out_235;
wire  [409:0]  u0_col_out_236;
wire  [409:0]  u0_col_out_237;
wire  [409:0]  u0_col_out_238;
wire  [409:0]  u0_col_out_239;
wire  [409:0]  u0_col_out_240;
wire  [409:0]  u0_col_out_241;
wire  [409:0]  u0_col_out_242;
wire  [409:0]  u0_col_out_243;
wire  [409:0]  u0_col_out_244;
wire  [409:0]  u0_col_out_245;
wire  [409:0]  u0_col_out_246;
wire  [409:0]  u0_col_out_247;
wire  [409:0]  u0_col_out_248;
wire  [409:0]  u0_col_out_249;
wire  [409:0]  u0_col_out_250;
wire  [409:0]  u0_col_out_251;
wire  [409:0]  u0_col_out_252;
wire  [409:0]  u0_col_out_253;
wire  [409:0]  u0_col_out_254;
wire  [409:0]  u0_col_out_255;
wire  [409:0]  u0_col_out_256;
wire  [409:0]  u0_col_out_257;
wire  [409:0]  u0_col_out_258;
wire  [409:0]  u0_col_out_259;
wire  [409:0]  u0_col_out_260;
wire  [409:0]  u0_col_out_261;
wire  [409:0]  u0_col_out_262;
wire  [409:0]  u0_col_out_263;
wire  [409:0]  u0_col_out_264;
wire  [409:0]  u0_col_out_265;
wire  [409:0]  u0_col_out_266;
wire  [409:0]  u0_col_out_267;
wire  [409:0]  u0_col_out_268;
wire  [409:0]  u0_col_out_269;
wire  [409:0]  u0_col_out_270;
wire  [409:0]  u0_col_out_271;
wire  [409:0]  u0_col_out_272;
wire  [409:0]  u0_col_out_273;
wire  [409:0]  u0_col_out_274;
wire  [409:0]  u0_col_out_275;
wire  [409:0]  u0_col_out_276;
wire  [409:0]  u0_col_out_277;
wire  [409:0]  u0_col_out_278;
wire  [409:0]  u0_col_out_279;
wire  [409:0]  u0_col_out_280;
wire  [409:0]  u0_col_out_281;
wire  [409:0]  u0_col_out_282;
wire  [409:0]  u0_col_out_283;
wire  [409:0]  u0_col_out_284;
wire  [409:0]  u0_col_out_285;
wire  [409:0]  u0_col_out_286;
wire  [409:0]  u0_col_out_287;
wire  [409:0]  u0_col_out_288;
wire  [409:0]  u0_col_out_289;
wire  [409:0]  u0_col_out_290;
wire  [409:0]  u0_col_out_291;
wire  [409:0]  u0_col_out_292;
wire  [409:0]  u0_col_out_293;
wire  [409:0]  u0_col_out_294;
wire  [409:0]  u0_col_out_295;
wire  [409:0]  u0_col_out_296;
wire  [409:0]  u0_col_out_297;
wire  [409:0]  u0_col_out_298;
wire  [409:0]  u0_col_out_299;
wire  [409:0]  u0_col_out_300;
wire  [409:0]  u0_col_out_301;
wire  [409:0]  u0_col_out_302;
wire  [409:0]  u0_col_out_303;
wire  [409:0]  u0_col_out_304;
wire  [409:0]  u0_col_out_305;
wire  [409:0]  u0_col_out_306;
wire  [409:0]  u0_col_out_307;
wire  [409:0]  u0_col_out_308;
wire  [409:0]  u0_col_out_309;
wire  [409:0]  u0_col_out_310;
wire  [409:0]  u0_col_out_311;
wire  [409:0]  u0_col_out_312;
wire  [409:0]  u0_col_out_313;
wire  [409:0]  u0_col_out_314;
wire  [409:0]  u0_col_out_315;
wire  [409:0]  u0_col_out_316;
wire  [409:0]  u0_col_out_317;
wire  [409:0]  u0_col_out_318;
wire  [409:0]  u0_col_out_319;
wire  [409:0]  u0_col_out_320;
wire  [409:0]  u0_col_out_321;
wire  [409:0]  u0_col_out_322;
wire  [409:0]  u0_col_out_323;
wire  [409:0]  u0_col_out_324;
wire  [409:0]  u0_col_out_325;
wire  [409:0]  u0_col_out_326;
wire  [409:0]  u0_col_out_327;
wire  [409:0]  u0_col_out_328;
wire  [409:0]  u0_col_out_329;
wire  [409:0]  u0_col_out_330;
wire  [409:0]  u0_col_out_331;
wire  [409:0]  u0_col_out_332;
wire  [409:0]  u0_col_out_333;
wire  [409:0]  u0_col_out_334;
wire  [409:0]  u0_col_out_335;
wire  [409:0]  u0_col_out_336;
wire  [409:0]  u0_col_out_337;
wire  [409:0]  u0_col_out_338;
wire  [409:0]  u0_col_out_339;
wire  [409:0]  u0_col_out_340;
wire  [409:0]  u0_col_out_341;
wire  [409:0]  u0_col_out_342;
wire  [409:0]  u0_col_out_343;
wire  [409:0]  u0_col_out_344;
wire  [409:0]  u0_col_out_345;
wire  [409:0]  u0_col_out_346;
wire  [409:0]  u0_col_out_347;
wire  [409:0]  u0_col_out_348;
wire  [409:0]  u0_col_out_349;
wire  [409:0]  u0_col_out_350;
wire  [409:0]  u0_col_out_351;
wire  [409:0]  u0_col_out_352;
wire  [409:0]  u0_col_out_353;
wire  [409:0]  u0_col_out_354;
wire  [409:0]  u0_col_out_355;
wire  [409:0]  u0_col_out_356;
wire  [409:0]  u0_col_out_357;
wire  [409:0]  u0_col_out_358;
wire  [409:0]  u0_col_out_359;
wire  [409:0]  u0_col_out_360;
wire  [409:0]  u0_col_out_361;
wire  [409:0]  u0_col_out_362;
wire  [409:0]  u0_col_out_363;
wire  [409:0]  u0_col_out_364;
wire  [409:0]  u0_col_out_365;
wire  [409:0]  u0_col_out_366;
wire  [409:0]  u0_col_out_367;
wire  [409:0]  u0_col_out_368;
wire  [409:0]  u0_col_out_369;
wire  [409:0]  u0_col_out_370;
wire  [409:0]  u0_col_out_371;
wire  [409:0]  u0_col_out_372;
wire  [409:0]  u0_col_out_373;
wire  [409:0]  u0_col_out_374;
wire  [409:0]  u0_col_out_375;
wire  [409:0]  u0_col_out_376;
wire  [409:0]  u0_col_out_377;
wire  [409:0]  u0_col_out_378;
wire  [409:0]  u0_col_out_379;
wire  [409:0]  u0_col_out_380;
wire  [409:0]  u0_col_out_381;
wire  [409:0]  u0_col_out_382;
wire  [409:0]  u0_col_out_383;
wire  [409:0]  u0_col_out_384;
wire  [409:0]  u0_col_out_385;
wire  [409:0]  u0_col_out_386;
wire  [409:0]  u0_col_out_387;
wire  [409:0]  u0_col_out_388;
wire  [409:0]  u0_col_out_389;
wire  [409:0]  u0_col_out_390;
wire  [409:0]  u0_col_out_391;
wire  [409:0]  u0_col_out_392;
wire  [409:0]  u0_col_out_393;
wire  [409:0]  u0_col_out_394;
wire  [409:0]  u0_col_out_395;
wire  [409:0]  u0_col_out_396;
wire  [409:0]  u0_col_out_397;
wire  [409:0]  u0_col_out_398;
wire  [409:0]  u0_col_out_399;
wire  [409:0]  u0_col_out_400;
wire  [409:0]  u0_col_out_401;
wire  [409:0]  u0_col_out_402;
wire  [409:0]  u0_col_out_403;
wire  [409:0]  u0_col_out_404;
wire  [409:0]  u0_col_out_405;
wire  [409:0]  u0_col_out_406;
wire  [409:0]  u0_col_out_407;
wire  [409:0]  u0_col_out_408;
wire  [409:0]  u0_col_out_409;
wire  [409:0]  u0_col_out_410;
wire  [409:0]  u0_col_out_411;
wire  [409:0]  u0_col_out_412;
wire  [409:0]  u0_col_out_413;
wire  [409:0]  u0_col_out_414;
wire  [409:0]  u0_col_out_415;
wire  [409:0]  u0_col_out_416;
wire  [409:0]  u0_col_out_417;
wire  [409:0]  u0_col_out_418;
wire  [409:0]  u0_col_out_419;
wire  [409:0]  u0_col_out_420;
wire  [409:0]  u0_col_out_421;
wire  [409:0]  u0_col_out_422;
wire  [409:0]  u0_col_out_423;
wire  [409:0]  u0_col_out_424;
wire  [409:0]  u0_col_out_425;
wire  [409:0]  u0_col_out_426;
wire  [409:0]  u0_col_out_427;
wire  [409:0]  u0_col_out_428;
wire  [409:0]  u0_col_out_429;
wire  [409:0]  u0_col_out_430;
wire  [409:0]  u0_col_out_431;
wire  [409:0]  u0_col_out_432;
wire  [409:0]  u0_col_out_433;
wire  [409:0]  u0_col_out_434;
wire  [409:0]  u0_col_out_435;
wire  [409:0]  u0_col_out_436;
wire  [409:0]  u0_col_out_437;
wire  [409:0]  u0_col_out_438;
wire  [409:0]  u0_col_out_439;
wire  [409:0]  u0_col_out_440;
wire  [409:0]  u0_col_out_441;
wire  [409:0]  u0_col_out_442;
wire  [409:0]  u0_col_out_443;
wire  [409:0]  u0_col_out_444;
wire  [409:0]  u0_col_out_445;
wire  [409:0]  u0_col_out_446;
wire  [409:0]  u0_col_out_447;
wire  [409:0]  u0_col_out_448;
wire  [409:0]  u0_col_out_449;
wire  [409:0]  u0_col_out_450;
wire  [409:0]  u0_col_out_451;
wire  [409:0]  u0_col_out_452;
wire  [409:0]  u0_col_out_453;
wire  [409:0]  u0_col_out_454;
wire  [409:0]  u0_col_out_455;
wire  [409:0]  u0_col_out_456;
wire  [409:0]  u0_col_out_457;
wire  [409:0]  u0_col_out_458;
wire  [409:0]  u0_col_out_459;
wire  [409:0]  u0_col_out_460;
wire  [409:0]  u0_col_out_461;
wire  [409:0]  u0_col_out_462;
wire  [409:0]  u0_col_out_463;
wire  [409:0]  u0_col_out_464;
wire  [409:0]  u0_col_out_465;
wire  [409:0]  u0_col_out_466;
wire  [409:0]  u0_col_out_467;
wire  [409:0]  u0_col_out_468;
wire  [409:0]  u0_col_out_469;
wire  [409:0]  u0_col_out_470;
wire  [409:0]  u0_col_out_471;
wire  [409:0]  u0_col_out_472;
wire  [409:0]  u0_col_out_473;
wire  [409:0]  u0_col_out_474;
wire  [409:0]  u0_col_out_475;
wire  [409:0]  u0_col_out_476;
wire  [409:0]  u0_col_out_477;
wire  [409:0]  u0_col_out_478;
wire  [409:0]  u0_col_out_479;
wire  [409:0]  u0_col_out_480;
wire  [409:0]  u0_col_out_481;
wire  [409:0]  u0_col_out_482;
wire  [409:0]  u0_col_out_483;
wire  [409:0]  u0_col_out_484;
wire  [409:0]  u0_col_out_485;
wire  [409:0]  u0_col_out_486;
wire  [409:0]  u0_col_out_487;
wire  [409:0]  u0_col_out_488;
wire  [409:0]  u0_col_out_489;
wire  [409:0]  u0_col_out_490;
wire  [409:0]  u0_col_out_491;
wire  [409:0]  u0_col_out_492;
wire  [409:0]  u0_col_out_493;
wire  [409:0]  u0_col_out_494;
wire  [409:0]  u0_col_out_495;
wire  [409:0]  u0_col_out_496;
wire  [409:0]  u0_col_out_497;
wire  [409:0]  u0_col_out_498;
wire  [409:0]  u0_col_out_499;
wire  [409:0]  u0_col_out_500;
wire  [409:0]  u0_col_out_501;
wire  [409:0]  u0_col_out_502;
wire  [409:0]  u0_col_out_503;
wire  [409:0]  u0_col_out_504;
wire  [409:0]  u0_col_out_505;
wire  [409:0]  u0_col_out_506;
wire  [409:0]  u0_col_out_507;
wire  [409:0]  u0_col_out_508;
wire  [409:0]  u0_col_out_509;
wire  [409:0]  u0_col_out_510;
wire  [409:0]  u0_col_out_511;
wire  [409:0]  u0_col_out_512;
wire  [409:0]  u0_col_out_513;
wire  [409:0]  u0_col_out_514;
wire  [409:0]  u0_col_out_515;
wire  [409:0]  u0_col_out_516;
wire  [409:0]  u0_col_out_517;
wire  [409:0]  u0_col_out_518;
wire  [409:0]  u0_col_out_519;
wire  [409:0]  u0_col_out_520;
wire  [409:0]  u0_col_out_521;
wire  [409:0]  u0_col_out_522;
wire  [409:0]  u0_col_out_523;
wire  [409:0]  u0_col_out_524;
wire  [409:0]  u0_col_out_525;
wire  [409:0]  u0_col_out_526;
wire  [409:0]  u0_col_out_527;
wire  [409:0]  u0_col_out_528;
wire  [409:0]  u0_col_out_529;
wire  [409:0]  u0_col_out_530;
wire  [409:0]  u0_col_out_531;
wire  [409:0]  u0_col_out_532;
wire  [409:0]  u0_col_out_533;
wire  [409:0]  u0_col_out_534;
wire  [409:0]  u0_col_out_535;
wire  [409:0]  u0_col_out_536;
wire  [409:0]  u0_col_out_537;
wire  [409:0]  u0_col_out_538;
wire  [409:0]  u0_col_out_539;
wire  [409:0]  u0_col_out_540;
wire  [409:0]  u0_col_out_541;
wire  [409:0]  u0_col_out_542;
wire  [409:0]  u0_col_out_543;
wire  [409:0]  u0_col_out_544;
wire  [409:0]  u0_col_out_545;
wire  [409:0]  u0_col_out_546;
wire  [409:0]  u0_col_out_547;
wire  [409:0]  u0_col_out_548;
wire  [409:0]  u0_col_out_549;
wire  [409:0]  u0_col_out_550;
wire  [409:0]  u0_col_out_551;
wire  [409:0]  u0_col_out_552;
wire  [409:0]  u0_col_out_553;
wire  [409:0]  u0_col_out_554;
wire  [409:0]  u0_col_out_555;
wire  [409:0]  u0_col_out_556;
wire  [409:0]  u0_col_out_557;
wire  [409:0]  u0_col_out_558;
wire  [409:0]  u0_col_out_559;
wire  [409:0]  u0_col_out_560;
wire  [409:0]  u0_col_out_561;
wire  [409:0]  u0_col_out_562;
wire  [409:0]  u0_col_out_563;
wire  [409:0]  u0_col_out_564;
wire  [409:0]  u0_col_out_565;
wire  [409:0]  u0_col_out_566;
wire  [409:0]  u0_col_out_567;
wire  [409:0]  u0_col_out_568;
wire  [409:0]  u0_col_out_569;
wire  [409:0]  u0_col_out_570;
wire  [409:0]  u0_col_out_571;
wire  [409:0]  u0_col_out_572;
wire  [409:0]  u0_col_out_573;
wire  [409:0]  u0_col_out_574;
wire  [409:0]  u0_col_out_575;
wire  [409:0]  u0_col_out_576;
wire  [409:0]  u0_col_out_577;
wire  [409:0]  u0_col_out_578;
wire  [409:0]  u0_col_out_579;
wire  [409:0]  u0_col_out_580;
wire  [409:0]  u0_col_out_581;
wire  [409:0]  u0_col_out_582;
wire  [409:0]  u0_col_out_583;
wire  [409:0]  u0_col_out_584;
wire  [409:0]  u0_col_out_585;
wire  [409:0]  u0_col_out_586;
wire  [409:0]  u0_col_out_587;
wire  [409:0]  u0_col_out_588;
wire  [409:0]  u0_col_out_589;
wire  [409:0]  u0_col_out_590;
wire  [409:0]  u0_col_out_591;
wire  [409:0]  u0_col_out_592;
wire  [409:0]  u0_col_out_593;
wire  [409:0]  u0_col_out_594;
wire  [409:0]  u0_col_out_595;
wire  [409:0]  u0_col_out_596;
wire  [409:0]  u0_col_out_597;
wire  [409:0]  u0_col_out_598;
wire  [409:0]  u0_col_out_599;
wire  [409:0]  u0_col_out_600;
wire  [409:0]  u0_col_out_601;
wire  [409:0]  u0_col_out_602;
wire  [409:0]  u0_col_out_603;
wire  [409:0]  u0_col_out_604;
wire  [409:0]  u0_col_out_605;
wire  [409:0]  u0_col_out_606;
wire  [409:0]  u0_col_out_607;
wire  [409:0]  u0_col_out_608;
wire  [409:0]  u0_col_out_609;
wire  [409:0]  u0_col_out_610;
wire  [409:0]  u0_col_out_611;
wire  [409:0]  u0_col_out_612;
wire  [409:0]  u0_col_out_613;
wire  [409:0]  u0_col_out_614;
wire  [409:0]  u0_col_out_615;
wire  [409:0]  u0_col_out_616;
wire  [409:0]  u0_col_out_617;
wire  [409:0]  u0_col_out_618;
wire  [409:0]  u0_col_out_619;
wire  [409:0]  u0_col_out_620;
wire  [409:0]  u0_col_out_621;
wire  [409:0]  u0_col_out_622;
wire  [409:0]  u0_col_out_623;
wire  [409:0]  u0_col_out_624;
wire  [409:0]  u0_col_out_625;
wire  [409:0]  u0_col_out_626;
wire  [409:0]  u0_col_out_627;
wire  [409:0]  u0_col_out_628;
wire  [409:0]  u0_col_out_629;
wire  [409:0]  u0_col_out_630;
wire  [409:0]  u0_col_out_631;
wire  [409:0]  u0_col_out_632;
wire  [409:0]  u0_col_out_633;
wire  [409:0]  u0_col_out_634;
wire  [409:0]  u0_col_out_635;
wire  [409:0]  u0_col_out_636;
wire  [409:0]  u0_col_out_637;
wire  [409:0]  u0_col_out_638;
wire  [409:0]  u0_col_out_639;
wire  [409:0]  u0_col_out_640;
wire  [409:0]  u0_col_out_641;
wire  [409:0]  u0_col_out_642;
wire  [409:0]  u0_col_out_643;
wire  [409:0]  u0_col_out_644;
wire  [409:0]  u0_col_out_645;
wire  [409:0]  u0_col_out_646;
wire  [409:0]  u0_col_out_647;
wire  [409:0]  u0_col_out_648;
wire  [409:0]  u0_col_out_649;
wire  [409:0]  u0_col_out_650;
wire  [409:0]  u0_col_out_651;
wire  [409:0]  u0_col_out_652;
wire  [409:0]  u0_col_out_653;
wire  [409:0]  u0_col_out_654;
wire  [409:0]  u0_col_out_655;
wire  [409:0]  u0_col_out_656;
wire  [409:0]  u0_col_out_657;
wire  [409:0]  u0_col_out_658;
wire  [409:0]  u0_col_out_659;
wire  [409:0]  u0_col_out_660;
wire  [409:0]  u0_col_out_661;
wire  [409:0]  u0_col_out_662;
wire  [409:0]  u0_col_out_663;
wire  [409:0]  u0_col_out_664;
wire  [409:0]  u0_col_out_665;
wire  [409:0]  u0_col_out_666;
wire  [409:0]  u0_col_out_667;
wire  [409:0]  u0_col_out_668;
wire  [409:0]  u0_col_out_669;
wire  [409:0]  u0_col_out_670;
wire  [409:0]  u0_col_out_671;
wire  [409:0]  u0_col_out_672;
wire  [409:0]  u0_col_out_673;
wire  [409:0]  u0_col_out_674;
wire  [409:0]  u0_col_out_675;
wire  [409:0]  u0_col_out_676;
wire  [409:0]  u0_col_out_677;
wire  [409:0]  u0_col_out_678;
wire  [409:0]  u0_col_out_679;
wire  [409:0]  u0_col_out_680;
wire  [409:0]  u0_col_out_681;
wire  [409:0]  u0_col_out_682;
wire  [409:0]  u0_col_out_683;
wire  [409:0]  u0_col_out_684;
wire  [409:0]  u0_col_out_685;
wire  [409:0]  u0_col_out_686;
wire  [409:0]  u0_col_out_687;
wire  [409:0]  u0_col_out_688;
wire  [409:0]  u0_col_out_689;
wire  [409:0]  u0_col_out_690;
wire  [409:0]  u0_col_out_691;
wire  [409:0]  u0_col_out_692;
wire  [409:0]  u0_col_out_693;
wire  [409:0]  u0_col_out_694;
wire  [409:0]  u0_col_out_695;
wire  [409:0]  u0_col_out_696;
wire  [409:0]  u0_col_out_697;
wire  [409:0]  u0_col_out_698;
wire  [409:0]  u0_col_out_699;
wire  [409:0]  u0_col_out_700;
wire  [409:0]  u0_col_out_701;
wire  [409:0]  u0_col_out_702;
wire  [409:0]  u0_col_out_703;
wire  [409:0]  u0_col_out_704;
wire  [409:0]  u0_col_out_705;
wire  [409:0]  u0_col_out_706;
wire  [409:0]  u0_col_out_707;
wire  [409:0]  u0_col_out_708;
wire  [409:0]  u0_col_out_709;
wire  [409:0]  u0_col_out_710;
wire  [409:0]  u0_col_out_711;
wire  [409:0]  u0_col_out_712;
wire  [409:0]  u0_col_out_713;
wire  [409:0]  u0_col_out_714;
wire  [409:0]  u0_col_out_715;
wire  [409:0]  u0_col_out_716;
wire  [409:0]  u0_col_out_717;
wire  [409:0]  u0_col_out_718;
wire  [409:0]  u0_col_out_719;
wire  [409:0]  u0_col_out_720;
wire  [409:0]  u0_col_out_721;
wire  [409:0]  u0_col_out_722;
wire  [409:0]  u0_col_out_723;
wire  [409:0]  u0_col_out_724;
wire  [409:0]  u0_col_out_725;
wire  [409:0]  u0_col_out_726;
wire  [409:0]  u0_col_out_727;
wire  [409:0]  u0_col_out_728;
wire  [409:0]  u0_col_out_729;
wire  [409:0]  u0_col_out_730;
wire  [409:0]  u0_col_out_731;
wire  [409:0]  u0_col_out_732;
wire  [409:0]  u0_col_out_733;
wire  [409:0]  u0_col_out_734;
wire  [409:0]  u0_col_out_735;
wire  [409:0]  u0_col_out_736;
wire  [409:0]  u0_col_out_737;
wire  [409:0]  u0_col_out_738;
wire  [409:0]  u0_col_out_739;
wire  [409:0]  u0_col_out_740;
wire  [409:0]  u0_col_out_741;
wire  [409:0]  u0_col_out_742;
wire  [409:0]  u0_col_out_743;
wire  [409:0]  u0_col_out_744;
wire  [409:0]  u0_col_out_745;
wire  [409:0]  u0_col_out_746;
wire  [409:0]  u0_col_out_747;
wire  [409:0]  u0_col_out_748;
wire  [409:0]  u0_col_out_749;
wire  [409:0]  u0_col_out_750;
wire  [409:0]  u0_col_out_751;
wire  [409:0]  u0_col_out_752;
wire  [409:0]  u0_col_out_753;
wire  [409:0]  u0_col_out_754;
wire  [409:0]  u0_col_out_755;
wire  [409:0]  u0_col_out_756;
wire  [409:0]  u0_col_out_757;
wire  [409:0]  u0_col_out_758;
wire  [409:0]  u0_col_out_759;
wire  [409:0]  u0_col_out_760;
wire  [409:0]  u0_col_out_761;
wire  [409:0]  u0_col_out_762;
wire  [409:0]  u0_col_out_763;
wire  [409:0]  u0_col_out_764;
wire  [409:0]  u0_col_out_765;
wire  [409:0]  u0_col_out_766;
wire  [409:0]  u0_col_out_767;
wire  [409:0]  u0_col_out_768;
wire  [409:0]  u0_col_out_769;
wire  [409:0]  u0_col_out_770;
wire  [409:0]  u0_col_out_771;
wire  [409:0]  u0_col_out_772;
wire  [409:0]  u0_col_out_773;
wire  [409:0]  u0_col_out_774;
wire  [409:0]  u0_col_out_775;
wire  [409:0]  u0_col_out_776;
wire  [409:0]  u0_col_out_777;
wire  [409:0]  u0_col_out_778;
wire  [409:0]  u0_col_out_779;
wire  [409:0]  u0_col_out_780;
wire  [409:0]  u0_col_out_781;
wire  [409:0]  u0_col_out_782;
wire  [409:0]  u0_col_out_783;
wire  [409:0]  u0_col_out_784;
wire  [409:0]  u0_col_out_785;
wire  [409:0]  u0_col_out_786;
wire  [409:0]  u0_col_out_787;
wire  [409:0]  u0_col_out_788;
wire  [409:0]  u0_col_out_789;
wire  [409:0]  u0_col_out_790;
wire  [409:0]  u0_col_out_791;
wire  [409:0]  u0_col_out_792;
wire  [409:0]  u0_col_out_793;
wire  [409:0]  u0_col_out_794;
wire  [409:0]  u0_col_out_795;
wire  [409:0]  u0_col_out_796;
wire  [409:0]  u0_col_out_797;
wire  [409:0]  u0_col_out_798;
wire  [409:0]  u0_col_out_799;
wire  [409:0]  u0_col_out_800;
wire  [409:0]  u0_col_out_801;
wire  [409:0]  u0_col_out_802;
wire  [409:0]  u0_col_out_803;
wire  [409:0]  u0_col_out_804;
wire  [409:0]  u0_col_out_805;
wire  [409:0]  u0_col_out_806;
wire  [409:0]  u0_col_out_807;
wire  [409:0]  u0_col_out_808;
wire  [409:0]  u0_col_out_809;
wire  [409:0]  u0_col_out_810;
wire  [409:0]  u0_col_out_811;
wire  [409:0]  u0_col_out_812;
wire  [409:0]  u0_col_out_813;
wire  [409:0]  u0_col_out_814;
wire  [409:0]  u0_col_out_815;
wire  [409:0]  u0_col_out_816;
wire  [409:0]  u0_col_out_817;
wire  [409:0]  u0_col_out_818;
wire  [409:0]  u0_col_out_819;
wire  [409:0]  u0_col_out_820;
wire  [409:0]  u0_col_out_821;
wire  [409:0]  u0_col_out_822;
wire  [409:0]  u0_col_out_823;
wire  [409:0]  u0_col_out_824;
wire  [409:0]  u0_col_out_825;
wire  [409:0]  u0_col_out_826;
wire  [409:0]  u0_col_out_827;
wire  [409:0]  u0_col_out_828;
wire  [409:0]  u0_col_out_829;
wire  [409:0]  u0_col_out_830;
wire  [409:0]  u0_col_out_831;
wire  [409:0]  u0_col_out_832;
wire  [409:0]  u0_col_out_833;
wire  [409:0]  u0_col_out_834;
wire  [409:0]  u0_col_out_835;
wire  [409:0]  u0_col_out_836;
wire  [409:0]  u0_col_out_837;
wire  [409:0]  u0_col_out_838;
wire  [409:0]  u0_col_out_839;
wire  [409:0]  u0_col_out_840;
wire  [409:0]  u0_col_out_841;
wire  [409:0]  u0_col_out_842;
wire  [409:0]  u0_col_out_843;
wire  [409:0]  u0_col_out_844;
wire  [409:0]  u0_col_out_845;
wire  [409:0]  u0_col_out_846;
wire  [409:0]  u0_col_out_847;
wire  [409:0]  u0_col_out_848;
wire  [409:0]  u0_col_out_849;
wire  [409:0]  u0_col_out_850;
wire  [409:0]  u0_col_out_851;
wire  [409:0]  u0_col_out_852;
wire  [409:0]  u0_col_out_853;
wire  [409:0]  u0_col_out_854;
wire  [409:0]  u0_col_out_855;
wire  [409:0]  u0_col_out_856;
wire  [409:0]  u0_col_out_857;
wire  [409:0]  u0_col_out_858;
wire  [409:0]  u0_col_out_859;
wire  [409:0]  u0_col_out_860;
wire  [409:0]  u0_col_out_861;
wire  [409:0]  u0_col_out_862;
wire  [409:0]  u0_col_out_863;
wire  [409:0]  u0_col_out_864;
wire  [409:0]  u0_col_out_865;
wire  [409:0]  u0_col_out_866;
wire  [409:0]  u0_col_out_867;
wire  [409:0]  u0_col_out_868;
wire  [409:0]  u0_col_out_869;
wire  [409:0]  u0_col_out_870;
wire  [409:0]  u0_col_out_871;
wire  [409:0]  u0_col_out_872;
wire  [409:0]  u0_col_out_873;
wire  [409:0]  u0_col_out_874;
wire  [409:0]  u0_col_out_875;
wire  [409:0]  u0_col_out_876;
wire  [409:0]  u0_col_out_877;
wire  [409:0]  u0_col_out_878;
wire  [409:0]  u0_col_out_879;
wire  [409:0]  u0_col_out_880;
wire  [409:0]  u0_col_out_881;
wire  [409:0]  u0_col_out_882;
wire  [409:0]  u0_col_out_883;
wire  [409:0]  u0_col_out_884;
wire  [409:0]  u0_col_out_885;
wire  [409:0]  u0_col_out_886;
wire  [409:0]  u0_col_out_887;
wire  [409:0]  u0_col_out_888;
wire  [409:0]  u0_col_out_889;
wire  [409:0]  u0_col_out_890;
wire  [409:0]  u0_col_out_891;
wire  [409:0]  u0_col_out_892;
wire  [409:0]  u0_col_out_893;
wire  [409:0]  u0_col_out_894;
wire  [409:0]  u0_col_out_895;
wire  [409:0]  u0_col_out_896;
wire  [409:0]  u0_col_out_897;
wire  [409:0]  u0_col_out_898;
wire  [409:0]  u0_col_out_899;
wire  [409:0]  u0_col_out_900;
wire  [409:0]  u0_col_out_901;
wire  [409:0]  u0_col_out_902;
wire  [409:0]  u0_col_out_903;
wire  [409:0]  u0_col_out_904;
wire  [409:0]  u0_col_out_905;
wire  [409:0]  u0_col_out_906;
wire  [409:0]  u0_col_out_907;
wire  [409:0]  u0_col_out_908;
wire  [409:0]  u0_col_out_909;
wire  [409:0]  u0_col_out_910;
wire  [409:0]  u0_col_out_911;
wire  [409:0]  u0_col_out_912;
wire  [409:0]  u0_col_out_913;
wire  [409:0]  u0_col_out_914;
wire  [409:0]  u0_col_out_915;
wire  [409:0]  u0_col_out_916;
wire  [409:0]  u0_col_out_917;
wire  [409:0]  u0_col_out_918;
wire  [409:0]  u0_col_out_919;
wire  [409:0]  u0_col_out_920;
wire  [409:0]  u0_col_out_921;
wire  [409:0]  u0_col_out_922;
wire  [409:0]  u0_col_out_923;
wire  [409:0]  u0_col_out_924;
wire  [409:0]  u0_col_out_925;
wire  [409:0]  u0_col_out_926;
wire  [409:0]  u0_col_out_927;
wire  [409:0]  u0_col_out_928;
wire  [409:0]  u0_col_out_929;
wire  [409:0]  u0_col_out_930;
wire  [409:0]  u0_col_out_931;
wire  [409:0]  u0_col_out_932;
wire  [409:0]  u0_col_out_933;
wire  [409:0]  u0_col_out_934;
wire  [409:0]  u0_col_out_935;
wire  [409:0]  u0_col_out_936;
wire  [409:0]  u0_col_out_937;
wire  [409:0]  u0_col_out_938;
wire  [409:0]  u0_col_out_939;
wire  [409:0]  u0_col_out_940;
wire  [409:0]  u0_col_out_941;
wire  [409:0]  u0_col_out_942;
wire  [409:0]  u0_col_out_943;
wire  [409:0]  u0_col_out_944;
wire  [409:0]  u0_col_out_945;
wire  [409:0]  u0_col_out_946;
wire  [409:0]  u0_col_out_947;
wire  [409:0]  u0_col_out_948;
wire  [409:0]  u0_col_out_949;
wire  [409:0]  u0_col_out_950;
wire  [409:0]  u0_col_out_951;
wire  [409:0]  u0_col_out_952;
wire  [409:0]  u0_col_out_953;
wire  [409:0]  u0_col_out_954;
wire  [409:0]  u0_col_out_955;
wire  [409:0]  u0_col_out_956;
wire  [409:0]  u0_col_out_957;
wire  [409:0]  u0_col_out_958;
wire  [409:0]  u0_col_out_959;
wire  [409:0]  u0_col_out_960;
wire  [409:0]  u0_col_out_961;
wire  [409:0]  u0_col_out_962;
wire  [409:0]  u0_col_out_963;
wire  [409:0]  u0_col_out_964;
wire  [409:0]  u0_col_out_965;
wire  [409:0]  u0_col_out_966;
wire  [409:0]  u0_col_out_967;
wire  [409:0]  u0_col_out_968;
wire  [409:0]  u0_col_out_969;
wire  [409:0]  u0_col_out_970;
wire  [409:0]  u0_col_out_971;
wire  [409:0]  u0_col_out_972;
wire  [409:0]  u0_col_out_973;
wire  [409:0]  u0_col_out_974;
wire  [409:0]  u0_col_out_975;
wire  [409:0]  u0_col_out_976;
wire  [409:0]  u0_col_out_977;
wire  [409:0]  u0_col_out_978;
wire  [409:0]  u0_col_out_979;
wire  [409:0]  u0_col_out_980;
wire  [409:0]  u0_col_out_981;
wire  [409:0]  u0_col_out_982;
wire  [409:0]  u0_col_out_983;
wire  [409:0]  u0_col_out_984;
wire  [409:0]  u0_col_out_985;
wire  [409:0]  u0_col_out_986;
wire  [409:0]  u0_col_out_987;
wire  [409:0]  u0_col_out_988;
wire  [409:0]  u0_col_out_989;
wire  [409:0]  u0_col_out_990;
wire  [409:0]  u0_col_out_991;
wire  [409:0]  u0_col_out_992;
wire  [409:0]  u0_col_out_993;
wire  [409:0]  u0_col_out_994;
wire  [409:0]  u0_col_out_995;
wire  [409:0]  u0_col_out_996;
wire  [409:0]  u0_col_out_997;
wire  [409:0]  u0_col_out_998;
wire  [409:0]  u0_col_out_999;
wire  [409:0]  u0_col_out_1000;
wire  [409:0]  u0_col_out_1001;
wire  [409:0]  u0_col_out_1002;
wire  [409:0]  u0_col_out_1003;
wire  [409:0]  u0_col_out_1004;
wire  [409:0]  u0_col_out_1005;
wire  [409:0]  u0_col_out_1006;
wire  [409:0]  u0_col_out_1007;
wire  [409:0]  u0_col_out_1008;
wire  [409:0]  u0_col_out_1009;
wire  [409:0]  u0_col_out_1010;
wire  [409:0]  u0_col_out_1011;
wire  [409:0]  u0_col_out_1012;
wire  [409:0]  u0_col_out_1013;
wire  [409:0]  u0_col_out_1014;
wire  [409:0]  u0_col_out_1015;
wire  [409:0]  u0_col_out_1016;
wire  [409:0]  u0_col_out_1017;
wire  [409:0]  u0_col_out_1018;
wire  [409:0]  u0_col_out_1019;
wire  [409:0]  u0_col_out_1020;
wire  [409:0]  u0_col_out_1021;
wire  [409:0]  u0_col_out_1022;
wire  [409:0]  u0_col_out_1023;

xpb_2018_col  u0_xpb_2018_col (
    .clk(clk),
    .data_in0                ( partial_product_high0       ),
    .data_in1                ( partial_product_high1       ),

    .col_out_0               ( u0_col_out_0[409:0]      ),
    .col_out_1               ( u0_col_out_1[409:0]      ),
    .col_out_2               ( u0_col_out_2[409:0]      ),
    .col_out_3               ( u0_col_out_3[409:0]      ),
    .col_out_4               ( u0_col_out_4[409:0]      ),
    .col_out_5               ( u0_col_out_5[409:0]      ),
    .col_out_6               ( u0_col_out_6[409:0]      ),
    .col_out_7               ( u0_col_out_7[409:0]      ),
    .col_out_8               ( u0_col_out_8[409:0]      ),
    .col_out_9               ( u0_col_out_9[409:0]      ),
    .col_out_10              ( u0_col_out_10[409:0]     ),
    .col_out_11              ( u0_col_out_11[409:0]     ),
    .col_out_12              ( u0_col_out_12[409:0]     ),
    .col_out_13              ( u0_col_out_13[409:0]     ),
    .col_out_14              ( u0_col_out_14[409:0]     ),
    .col_out_15              ( u0_col_out_15[409:0]     ),
    .col_out_16              ( u0_col_out_16[409:0]     ),
    .col_out_17              ( u0_col_out_17[409:0]     ),
    .col_out_18              ( u0_col_out_18[409:0]     ),
    .col_out_19              ( u0_col_out_19[409:0]     ),
    .col_out_20              ( u0_col_out_20[409:0]     ),
    .col_out_21              ( u0_col_out_21[409:0]     ),
    .col_out_22              ( u0_col_out_22[409:0]     ),
    .col_out_23              ( u0_col_out_23[409:0]     ),
    .col_out_24              ( u0_col_out_24[409:0]     ),
    .col_out_25              ( u0_col_out_25[409:0]     ),
    .col_out_26              ( u0_col_out_26[409:0]     ),
    .col_out_27              ( u0_col_out_27[409:0]     ),
    .col_out_28              ( u0_col_out_28[409:0]     ),
    .col_out_29              ( u0_col_out_29[409:0]     ),
    .col_out_30              ( u0_col_out_30[409:0]     ),
    .col_out_31              ( u0_col_out_31[409:0]     ),
    .col_out_32              ( u0_col_out_32[409:0]     ),
    .col_out_33              ( u0_col_out_33[409:0]     ),
    .col_out_34              ( u0_col_out_34[409:0]     ),
    .col_out_35              ( u0_col_out_35[409:0]     ),
    .col_out_36              ( u0_col_out_36[409:0]     ),
    .col_out_37              ( u0_col_out_37[409:0]     ),
    .col_out_38              ( u0_col_out_38[409:0]     ),
    .col_out_39              ( u0_col_out_39[409:0]     ),
    .col_out_40              ( u0_col_out_40[409:0]     ),
    .col_out_41              ( u0_col_out_41[409:0]     ),
    .col_out_42              ( u0_col_out_42[409:0]     ),
    .col_out_43              ( u0_col_out_43[409:0]     ),
    .col_out_44              ( u0_col_out_44[409:0]     ),
    .col_out_45              ( u0_col_out_45[409:0]     ),
    .col_out_46              ( u0_col_out_46[409:0]     ),
    .col_out_47              ( u0_col_out_47[409:0]     ),
    .col_out_48              ( u0_col_out_48[409:0]     ),
    .col_out_49              ( u0_col_out_49[409:0]     ),
    .col_out_50              ( u0_col_out_50[409:0]     ),
    .col_out_51              ( u0_col_out_51[409:0]     ),
    .col_out_52              ( u0_col_out_52[409:0]     ),
    .col_out_53              ( u0_col_out_53[409:0]     ),
    .col_out_54              ( u0_col_out_54[409:0]     ),
    .col_out_55              ( u0_col_out_55[409:0]     ),
    .col_out_56              ( u0_col_out_56[409:0]     ),
    .col_out_57              ( u0_col_out_57[409:0]     ),
    .col_out_58              ( u0_col_out_58[409:0]     ),
    .col_out_59              ( u0_col_out_59[409:0]     ),
    .col_out_60              ( u0_col_out_60[409:0]     ),
    .col_out_61              ( u0_col_out_61[409:0]     ),
    .col_out_62              ( u0_col_out_62[409:0]     ),
    .col_out_63              ( u0_col_out_63[409:0]     ),
    .col_out_64              ( u0_col_out_64[409:0]     ),
    .col_out_65              ( u0_col_out_65[409:0]     ),
    .col_out_66              ( u0_col_out_66[409:0]     ),
    .col_out_67              ( u0_col_out_67[409:0]     ),
    .col_out_68              ( u0_col_out_68[409:0]     ),
    .col_out_69              ( u0_col_out_69[409:0]     ),
    .col_out_70              ( u0_col_out_70[409:0]     ),
    .col_out_71              ( u0_col_out_71[409:0]     ),
    .col_out_72              ( u0_col_out_72[409:0]     ),
    .col_out_73              ( u0_col_out_73[409:0]     ),
    .col_out_74              ( u0_col_out_74[409:0]     ),
    .col_out_75              ( u0_col_out_75[409:0]     ),
    .col_out_76              ( u0_col_out_76[409:0]     ),
    .col_out_77              ( u0_col_out_77[409:0]     ),
    .col_out_78              ( u0_col_out_78[409:0]     ),
    .col_out_79              ( u0_col_out_79[409:0]     ),
    .col_out_80              ( u0_col_out_80[409:0]     ),
    .col_out_81              ( u0_col_out_81[409:0]     ),
    .col_out_82              ( u0_col_out_82[409:0]     ),
    .col_out_83              ( u0_col_out_83[409:0]     ),
    .col_out_84              ( u0_col_out_84[409:0]     ),
    .col_out_85              ( u0_col_out_85[409:0]     ),
    .col_out_86              ( u0_col_out_86[409:0]     ),
    .col_out_87              ( u0_col_out_87[409:0]     ),
    .col_out_88              ( u0_col_out_88[409:0]     ),
    .col_out_89              ( u0_col_out_89[409:0]     ),
    .col_out_90              ( u0_col_out_90[409:0]     ),
    .col_out_91              ( u0_col_out_91[409:0]     ),
    .col_out_92              ( u0_col_out_92[409:0]     ),
    .col_out_93              ( u0_col_out_93[409:0]     ),
    .col_out_94              ( u0_col_out_94[409:0]     ),
    .col_out_95              ( u0_col_out_95[409:0]     ),
    .col_out_96              ( u0_col_out_96[409:0]     ),
    .col_out_97              ( u0_col_out_97[409:0]     ),
    .col_out_98              ( u0_col_out_98[409:0]     ),
    .col_out_99              ( u0_col_out_99[409:0]     ),
    .col_out_100             ( u0_col_out_100[409:0]    ),
    .col_out_101             ( u0_col_out_101[409:0]    ),
    .col_out_102             ( u0_col_out_102[409:0]    ),
    .col_out_103             ( u0_col_out_103[409:0]    ),
    .col_out_104             ( u0_col_out_104[409:0]    ),
    .col_out_105             ( u0_col_out_105[409:0]    ),
    .col_out_106             ( u0_col_out_106[409:0]    ),
    .col_out_107             ( u0_col_out_107[409:0]    ),
    .col_out_108             ( u0_col_out_108[409:0]    ),
    .col_out_109             ( u0_col_out_109[409:0]    ),
    .col_out_110             ( u0_col_out_110[409:0]    ),
    .col_out_111             ( u0_col_out_111[409:0]    ),
    .col_out_112             ( u0_col_out_112[409:0]    ),
    .col_out_113             ( u0_col_out_113[409:0]    ),
    .col_out_114             ( u0_col_out_114[409:0]    ),
    .col_out_115             ( u0_col_out_115[409:0]    ),
    .col_out_116             ( u0_col_out_116[409:0]    ),
    .col_out_117             ( u0_col_out_117[409:0]    ),
    .col_out_118             ( u0_col_out_118[409:0]    ),
    .col_out_119             ( u0_col_out_119[409:0]    ),
    .col_out_120             ( u0_col_out_120[409:0]    ),
    .col_out_121             ( u0_col_out_121[409:0]    ),
    .col_out_122             ( u0_col_out_122[409:0]    ),
    .col_out_123             ( u0_col_out_123[409:0]    ),
    .col_out_124             ( u0_col_out_124[409:0]    ),
    .col_out_125             ( u0_col_out_125[409:0]    ),
    .col_out_126             ( u0_col_out_126[409:0]    ),
    .col_out_127             ( u0_col_out_127[409:0]    ),
    .col_out_128             ( u0_col_out_128[409:0]    ),
    .col_out_129             ( u0_col_out_129[409:0]    ),
    .col_out_130             ( u0_col_out_130[409:0]    ),
    .col_out_131             ( u0_col_out_131[409:0]    ),
    .col_out_132             ( u0_col_out_132[409:0]    ),
    .col_out_133             ( u0_col_out_133[409:0]    ),
    .col_out_134             ( u0_col_out_134[409:0]    ),
    .col_out_135             ( u0_col_out_135[409:0]    ),
    .col_out_136             ( u0_col_out_136[409:0]    ),
    .col_out_137             ( u0_col_out_137[409:0]    ),
    .col_out_138             ( u0_col_out_138[409:0]    ),
    .col_out_139             ( u0_col_out_139[409:0]    ),
    .col_out_140             ( u0_col_out_140[409:0]    ),
    .col_out_141             ( u0_col_out_141[409:0]    ),
    .col_out_142             ( u0_col_out_142[409:0]    ),
    .col_out_143             ( u0_col_out_143[409:0]    ),
    .col_out_144             ( u0_col_out_144[409:0]    ),
    .col_out_145             ( u0_col_out_145[409:0]    ),
    .col_out_146             ( u0_col_out_146[409:0]    ),
    .col_out_147             ( u0_col_out_147[409:0]    ),
    .col_out_148             ( u0_col_out_148[409:0]    ),
    .col_out_149             ( u0_col_out_149[409:0]    ),
    .col_out_150             ( u0_col_out_150[409:0]    ),
    .col_out_151             ( u0_col_out_151[409:0]    ),
    .col_out_152             ( u0_col_out_152[409:0]    ),
    .col_out_153             ( u0_col_out_153[409:0]    ),
    .col_out_154             ( u0_col_out_154[409:0]    ),
    .col_out_155             ( u0_col_out_155[409:0]    ),
    .col_out_156             ( u0_col_out_156[409:0]    ),
    .col_out_157             ( u0_col_out_157[409:0]    ),
    .col_out_158             ( u0_col_out_158[409:0]    ),
    .col_out_159             ( u0_col_out_159[409:0]    ),
    .col_out_160             ( u0_col_out_160[409:0]    ),
    .col_out_161             ( u0_col_out_161[409:0]    ),
    .col_out_162             ( u0_col_out_162[409:0]    ),
    .col_out_163             ( u0_col_out_163[409:0]    ),
    .col_out_164             ( u0_col_out_164[409:0]    ),
    .col_out_165             ( u0_col_out_165[409:0]    ),
    .col_out_166             ( u0_col_out_166[409:0]    ),
    .col_out_167             ( u0_col_out_167[409:0]    ),
    .col_out_168             ( u0_col_out_168[409:0]    ),
    .col_out_169             ( u0_col_out_169[409:0]    ),
    .col_out_170             ( u0_col_out_170[409:0]    ),
    .col_out_171             ( u0_col_out_171[409:0]    ),
    .col_out_172             ( u0_col_out_172[409:0]    ),
    .col_out_173             ( u0_col_out_173[409:0]    ),
    .col_out_174             ( u0_col_out_174[409:0]    ),
    .col_out_175             ( u0_col_out_175[409:0]    ),
    .col_out_176             ( u0_col_out_176[409:0]    ),
    .col_out_177             ( u0_col_out_177[409:0]    ),
    .col_out_178             ( u0_col_out_178[409:0]    ),
    .col_out_179             ( u0_col_out_179[409:0]    ),
    .col_out_180             ( u0_col_out_180[409:0]    ),
    .col_out_181             ( u0_col_out_181[409:0]    ),
    .col_out_182             ( u0_col_out_182[409:0]    ),
    .col_out_183             ( u0_col_out_183[409:0]    ),
    .col_out_184             ( u0_col_out_184[409:0]    ),
    .col_out_185             ( u0_col_out_185[409:0]    ),
    .col_out_186             ( u0_col_out_186[409:0]    ),
    .col_out_187             ( u0_col_out_187[409:0]    ),
    .col_out_188             ( u0_col_out_188[409:0]    ),
    .col_out_189             ( u0_col_out_189[409:0]    ),
    .col_out_190             ( u0_col_out_190[409:0]    ),
    .col_out_191             ( u0_col_out_191[409:0]    ),
    .col_out_192             ( u0_col_out_192[409:0]    ),
    .col_out_193             ( u0_col_out_193[409:0]    ),
    .col_out_194             ( u0_col_out_194[409:0]    ),
    .col_out_195             ( u0_col_out_195[409:0]    ),
    .col_out_196             ( u0_col_out_196[409:0]    ),
    .col_out_197             ( u0_col_out_197[409:0]    ),
    .col_out_198             ( u0_col_out_198[409:0]    ),
    .col_out_199             ( u0_col_out_199[409:0]    ),
    .col_out_200             ( u0_col_out_200[409:0]    ),
    .col_out_201             ( u0_col_out_201[409:0]    ),
    .col_out_202             ( u0_col_out_202[409:0]    ),
    .col_out_203             ( u0_col_out_203[409:0]    ),
    .col_out_204             ( u0_col_out_204[409:0]    ),
    .col_out_205             ( u0_col_out_205[409:0]    ),
    .col_out_206             ( u0_col_out_206[409:0]    ),
    .col_out_207             ( u0_col_out_207[409:0]    ),
    .col_out_208             ( u0_col_out_208[409:0]    ),
    .col_out_209             ( u0_col_out_209[409:0]    ),
    .col_out_210             ( u0_col_out_210[409:0]    ),
    .col_out_211             ( u0_col_out_211[409:0]    ),
    .col_out_212             ( u0_col_out_212[409:0]    ),
    .col_out_213             ( u0_col_out_213[409:0]    ),
    .col_out_214             ( u0_col_out_214[409:0]    ),
    .col_out_215             ( u0_col_out_215[409:0]    ),
    .col_out_216             ( u0_col_out_216[409:0]    ),
    .col_out_217             ( u0_col_out_217[409:0]    ),
    .col_out_218             ( u0_col_out_218[409:0]    ),
    .col_out_219             ( u0_col_out_219[409:0]    ),
    .col_out_220             ( u0_col_out_220[409:0]    ),
    .col_out_221             ( u0_col_out_221[409:0]    ),
    .col_out_222             ( u0_col_out_222[409:0]    ),
    .col_out_223             ( u0_col_out_223[409:0]    ),
    .col_out_224             ( u0_col_out_224[409:0]    ),
    .col_out_225             ( u0_col_out_225[409:0]    ),
    .col_out_226             ( u0_col_out_226[409:0]    ),
    .col_out_227             ( u0_col_out_227[409:0]    ),
    .col_out_228             ( u0_col_out_228[409:0]    ),
    .col_out_229             ( u0_col_out_229[409:0]    ),
    .col_out_230             ( u0_col_out_230[409:0]    ),
    .col_out_231             ( u0_col_out_231[409:0]    ),
    .col_out_232             ( u0_col_out_232[409:0]    ),
    .col_out_233             ( u0_col_out_233[409:0]    ),
    .col_out_234             ( u0_col_out_234[409:0]    ),
    .col_out_235             ( u0_col_out_235[409:0]    ),
    .col_out_236             ( u0_col_out_236[409:0]    ),
    .col_out_237             ( u0_col_out_237[409:0]    ),
    .col_out_238             ( u0_col_out_238[409:0]    ),
    .col_out_239             ( u0_col_out_239[409:0]    ),
    .col_out_240             ( u0_col_out_240[409:0]    ),
    .col_out_241             ( u0_col_out_241[409:0]    ),
    .col_out_242             ( u0_col_out_242[409:0]    ),
    .col_out_243             ( u0_col_out_243[409:0]    ),
    .col_out_244             ( u0_col_out_244[409:0]    ),
    .col_out_245             ( u0_col_out_245[409:0]    ),
    .col_out_246             ( u0_col_out_246[409:0]    ),
    .col_out_247             ( u0_col_out_247[409:0]    ),
    .col_out_248             ( u0_col_out_248[409:0]    ),
    .col_out_249             ( u0_col_out_249[409:0]    ),
    .col_out_250             ( u0_col_out_250[409:0]    ),
    .col_out_251             ( u0_col_out_251[409:0]    ),
    .col_out_252             ( u0_col_out_252[409:0]    ),
    .col_out_253             ( u0_col_out_253[409:0]    ),
    .col_out_254             ( u0_col_out_254[409:0]    ),
    .col_out_255             ( u0_col_out_255[409:0]    ),
    .col_out_256             ( u0_col_out_256[409:0]    ),
    .col_out_257             ( u0_col_out_257[409:0]    ),
    .col_out_258             ( u0_col_out_258[409:0]    ),
    .col_out_259             ( u0_col_out_259[409:0]    ),
    .col_out_260             ( u0_col_out_260[409:0]    ),
    .col_out_261             ( u0_col_out_261[409:0]    ),
    .col_out_262             ( u0_col_out_262[409:0]    ),
    .col_out_263             ( u0_col_out_263[409:0]    ),
    .col_out_264             ( u0_col_out_264[409:0]    ),
    .col_out_265             ( u0_col_out_265[409:0]    ),
    .col_out_266             ( u0_col_out_266[409:0]    ),
    .col_out_267             ( u0_col_out_267[409:0]    ),
    .col_out_268             ( u0_col_out_268[409:0]    ),
    .col_out_269             ( u0_col_out_269[409:0]    ),
    .col_out_270             ( u0_col_out_270[409:0]    ),
    .col_out_271             ( u0_col_out_271[409:0]    ),
    .col_out_272             ( u0_col_out_272[409:0]    ),
    .col_out_273             ( u0_col_out_273[409:0]    ),
    .col_out_274             ( u0_col_out_274[409:0]    ),
    .col_out_275             ( u0_col_out_275[409:0]    ),
    .col_out_276             ( u0_col_out_276[409:0]    ),
    .col_out_277             ( u0_col_out_277[409:0]    ),
    .col_out_278             ( u0_col_out_278[409:0]    ),
    .col_out_279             ( u0_col_out_279[409:0]    ),
    .col_out_280             ( u0_col_out_280[409:0]    ),
    .col_out_281             ( u0_col_out_281[409:0]    ),
    .col_out_282             ( u0_col_out_282[409:0]    ),
    .col_out_283             ( u0_col_out_283[409:0]    ),
    .col_out_284             ( u0_col_out_284[409:0]    ),
    .col_out_285             ( u0_col_out_285[409:0]    ),
    .col_out_286             ( u0_col_out_286[409:0]    ),
    .col_out_287             ( u0_col_out_287[409:0]    ),
    .col_out_288             ( u0_col_out_288[409:0]    ),
    .col_out_289             ( u0_col_out_289[409:0]    ),
    .col_out_290             ( u0_col_out_290[409:0]    ),
    .col_out_291             ( u0_col_out_291[409:0]    ),
    .col_out_292             ( u0_col_out_292[409:0]    ),
    .col_out_293             ( u0_col_out_293[409:0]    ),
    .col_out_294             ( u0_col_out_294[409:0]    ),
    .col_out_295             ( u0_col_out_295[409:0]    ),
    .col_out_296             ( u0_col_out_296[409:0]    ),
    .col_out_297             ( u0_col_out_297[409:0]    ),
    .col_out_298             ( u0_col_out_298[409:0]    ),
    .col_out_299             ( u0_col_out_299[409:0]    ),
    .col_out_300             ( u0_col_out_300[409:0]    ),
    .col_out_301             ( u0_col_out_301[409:0]    ),
    .col_out_302             ( u0_col_out_302[409:0]    ),
    .col_out_303             ( u0_col_out_303[409:0]    ),
    .col_out_304             ( u0_col_out_304[409:0]    ),
    .col_out_305             ( u0_col_out_305[409:0]    ),
    .col_out_306             ( u0_col_out_306[409:0]    ),
    .col_out_307             ( u0_col_out_307[409:0]    ),
    .col_out_308             ( u0_col_out_308[409:0]    ),
    .col_out_309             ( u0_col_out_309[409:0]    ),
    .col_out_310             ( u0_col_out_310[409:0]    ),
    .col_out_311             ( u0_col_out_311[409:0]    ),
    .col_out_312             ( u0_col_out_312[409:0]    ),
    .col_out_313             ( u0_col_out_313[409:0]    ),
    .col_out_314             ( u0_col_out_314[409:0]    ),
    .col_out_315             ( u0_col_out_315[409:0]    ),
    .col_out_316             ( u0_col_out_316[409:0]    ),
    .col_out_317             ( u0_col_out_317[409:0]    ),
    .col_out_318             ( u0_col_out_318[409:0]    ),
    .col_out_319             ( u0_col_out_319[409:0]    ),
    .col_out_320             ( u0_col_out_320[409:0]    ),
    .col_out_321             ( u0_col_out_321[409:0]    ),
    .col_out_322             ( u0_col_out_322[409:0]    ),
    .col_out_323             ( u0_col_out_323[409:0]    ),
    .col_out_324             ( u0_col_out_324[409:0]    ),
    .col_out_325             ( u0_col_out_325[409:0]    ),
    .col_out_326             ( u0_col_out_326[409:0]    ),
    .col_out_327             ( u0_col_out_327[409:0]    ),
    .col_out_328             ( u0_col_out_328[409:0]    ),
    .col_out_329             ( u0_col_out_329[409:0]    ),
    .col_out_330             ( u0_col_out_330[409:0]    ),
    .col_out_331             ( u0_col_out_331[409:0]    ),
    .col_out_332             ( u0_col_out_332[409:0]    ),
    .col_out_333             ( u0_col_out_333[409:0]    ),
    .col_out_334             ( u0_col_out_334[409:0]    ),
    .col_out_335             ( u0_col_out_335[409:0]    ),
    .col_out_336             ( u0_col_out_336[409:0]    ),
    .col_out_337             ( u0_col_out_337[409:0]    ),
    .col_out_338             ( u0_col_out_338[409:0]    ),
    .col_out_339             ( u0_col_out_339[409:0]    ),
    .col_out_340             ( u0_col_out_340[409:0]    ),
    .col_out_341             ( u0_col_out_341[409:0]    ),
    .col_out_342             ( u0_col_out_342[409:0]    ),
    .col_out_343             ( u0_col_out_343[409:0]    ),
    .col_out_344             ( u0_col_out_344[409:0]    ),
    .col_out_345             ( u0_col_out_345[409:0]    ),
    .col_out_346             ( u0_col_out_346[409:0]    ),
    .col_out_347             ( u0_col_out_347[409:0]    ),
    .col_out_348             ( u0_col_out_348[409:0]    ),
    .col_out_349             ( u0_col_out_349[409:0]    ),
    .col_out_350             ( u0_col_out_350[409:0]    ),
    .col_out_351             ( u0_col_out_351[409:0]    ),
    .col_out_352             ( u0_col_out_352[409:0]    ),
    .col_out_353             ( u0_col_out_353[409:0]    ),
    .col_out_354             ( u0_col_out_354[409:0]    ),
    .col_out_355             ( u0_col_out_355[409:0]    ),
    .col_out_356             ( u0_col_out_356[409:0]    ),
    .col_out_357             ( u0_col_out_357[409:0]    ),
    .col_out_358             ( u0_col_out_358[409:0]    ),
    .col_out_359             ( u0_col_out_359[409:0]    ),
    .col_out_360             ( u0_col_out_360[409:0]    ),
    .col_out_361             ( u0_col_out_361[409:0]    ),
    .col_out_362             ( u0_col_out_362[409:0]    ),
    .col_out_363             ( u0_col_out_363[409:0]    ),
    .col_out_364             ( u0_col_out_364[409:0]    ),
    .col_out_365             ( u0_col_out_365[409:0]    ),
    .col_out_366             ( u0_col_out_366[409:0]    ),
    .col_out_367             ( u0_col_out_367[409:0]    ),
    .col_out_368             ( u0_col_out_368[409:0]    ),
    .col_out_369             ( u0_col_out_369[409:0]    ),
    .col_out_370             ( u0_col_out_370[409:0]    ),
    .col_out_371             ( u0_col_out_371[409:0]    ),
    .col_out_372             ( u0_col_out_372[409:0]    ),
    .col_out_373             ( u0_col_out_373[409:0]    ),
    .col_out_374             ( u0_col_out_374[409:0]    ),
    .col_out_375             ( u0_col_out_375[409:0]    ),
    .col_out_376             ( u0_col_out_376[409:0]    ),
    .col_out_377             ( u0_col_out_377[409:0]    ),
    .col_out_378             ( u0_col_out_378[409:0]    ),
    .col_out_379             ( u0_col_out_379[409:0]    ),
    .col_out_380             ( u0_col_out_380[409:0]    ),
    .col_out_381             ( u0_col_out_381[409:0]    ),
    .col_out_382             ( u0_col_out_382[409:0]    ),
    .col_out_383             ( u0_col_out_383[409:0]    ),
    .col_out_384             ( u0_col_out_384[409:0]    ),
    .col_out_385             ( u0_col_out_385[409:0]    ),
    .col_out_386             ( u0_col_out_386[409:0]    ),
    .col_out_387             ( u0_col_out_387[409:0]    ),
    .col_out_388             ( u0_col_out_388[409:0]    ),
    .col_out_389             ( u0_col_out_389[409:0]    ),
    .col_out_390             ( u0_col_out_390[409:0]    ),
    .col_out_391             ( u0_col_out_391[409:0]    ),
    .col_out_392             ( u0_col_out_392[409:0]    ),
    .col_out_393             ( u0_col_out_393[409:0]    ),
    .col_out_394             ( u0_col_out_394[409:0]    ),
    .col_out_395             ( u0_col_out_395[409:0]    ),
    .col_out_396             ( u0_col_out_396[409:0]    ),
    .col_out_397             ( u0_col_out_397[409:0]    ),
    .col_out_398             ( u0_col_out_398[409:0]    ),
    .col_out_399             ( u0_col_out_399[409:0]    ),
    .col_out_400             ( u0_col_out_400[409:0]    ),
    .col_out_401             ( u0_col_out_401[409:0]    ),
    .col_out_402             ( u0_col_out_402[409:0]    ),
    .col_out_403             ( u0_col_out_403[409:0]    ),
    .col_out_404             ( u0_col_out_404[409:0]    ),
    .col_out_405             ( u0_col_out_405[409:0]    ),
    .col_out_406             ( u0_col_out_406[409:0]    ),
    .col_out_407             ( u0_col_out_407[409:0]    ),
    .col_out_408             ( u0_col_out_408[409:0]    ),
    .col_out_409             ( u0_col_out_409[409:0]    ),
    .col_out_410             ( u0_col_out_410[409:0]    ),
    .col_out_411             ( u0_col_out_411[409:0]    ),
    .col_out_412             ( u0_col_out_412[409:0]    ),
    .col_out_413             ( u0_col_out_413[409:0]    ),
    .col_out_414             ( u0_col_out_414[409:0]    ),
    .col_out_415             ( u0_col_out_415[409:0]    ),
    .col_out_416             ( u0_col_out_416[409:0]    ),
    .col_out_417             ( u0_col_out_417[409:0]    ),
    .col_out_418             ( u0_col_out_418[409:0]    ),
    .col_out_419             ( u0_col_out_419[409:0]    ),
    .col_out_420             ( u0_col_out_420[409:0]    ),
    .col_out_421             ( u0_col_out_421[409:0]    ),
    .col_out_422             ( u0_col_out_422[409:0]    ),
    .col_out_423             ( u0_col_out_423[409:0]    ),
    .col_out_424             ( u0_col_out_424[409:0]    ),
    .col_out_425             ( u0_col_out_425[409:0]    ),
    .col_out_426             ( u0_col_out_426[409:0]    ),
    .col_out_427             ( u0_col_out_427[409:0]    ),
    .col_out_428             ( u0_col_out_428[409:0]    ),
    .col_out_429             ( u0_col_out_429[409:0]    ),
    .col_out_430             ( u0_col_out_430[409:0]    ),
    .col_out_431             ( u0_col_out_431[409:0]    ),
    .col_out_432             ( u0_col_out_432[409:0]    ),
    .col_out_433             ( u0_col_out_433[409:0]    ),
    .col_out_434             ( u0_col_out_434[409:0]    ),
    .col_out_435             ( u0_col_out_435[409:0]    ),
    .col_out_436             ( u0_col_out_436[409:0]    ),
    .col_out_437             ( u0_col_out_437[409:0]    ),
    .col_out_438             ( u0_col_out_438[409:0]    ),
    .col_out_439             ( u0_col_out_439[409:0]    ),
    .col_out_440             ( u0_col_out_440[409:0]    ),
    .col_out_441             ( u0_col_out_441[409:0]    ),
    .col_out_442             ( u0_col_out_442[409:0]    ),
    .col_out_443             ( u0_col_out_443[409:0]    ),
    .col_out_444             ( u0_col_out_444[409:0]    ),
    .col_out_445             ( u0_col_out_445[409:0]    ),
    .col_out_446             ( u0_col_out_446[409:0]    ),
    .col_out_447             ( u0_col_out_447[409:0]    ),
    .col_out_448             ( u0_col_out_448[409:0]    ),
    .col_out_449             ( u0_col_out_449[409:0]    ),
    .col_out_450             ( u0_col_out_450[409:0]    ),
    .col_out_451             ( u0_col_out_451[409:0]    ),
    .col_out_452             ( u0_col_out_452[409:0]    ),
    .col_out_453             ( u0_col_out_453[409:0]    ),
    .col_out_454             ( u0_col_out_454[409:0]    ),
    .col_out_455             ( u0_col_out_455[409:0]    ),
    .col_out_456             ( u0_col_out_456[409:0]    ),
    .col_out_457             ( u0_col_out_457[409:0]    ),
    .col_out_458             ( u0_col_out_458[409:0]    ),
    .col_out_459             ( u0_col_out_459[409:0]    ),
    .col_out_460             ( u0_col_out_460[409:0]    ),
    .col_out_461             ( u0_col_out_461[409:0]    ),
    .col_out_462             ( u0_col_out_462[409:0]    ),
    .col_out_463             ( u0_col_out_463[409:0]    ),
    .col_out_464             ( u0_col_out_464[409:0]    ),
    .col_out_465             ( u0_col_out_465[409:0]    ),
    .col_out_466             ( u0_col_out_466[409:0]    ),
    .col_out_467             ( u0_col_out_467[409:0]    ),
    .col_out_468             ( u0_col_out_468[409:0]    ),
    .col_out_469             ( u0_col_out_469[409:0]    ),
    .col_out_470             ( u0_col_out_470[409:0]    ),
    .col_out_471             ( u0_col_out_471[409:0]    ),
    .col_out_472             ( u0_col_out_472[409:0]    ),
    .col_out_473             ( u0_col_out_473[409:0]    ),
    .col_out_474             ( u0_col_out_474[409:0]    ),
    .col_out_475             ( u0_col_out_475[409:0]    ),
    .col_out_476             ( u0_col_out_476[409:0]    ),
    .col_out_477             ( u0_col_out_477[409:0]    ),
    .col_out_478             ( u0_col_out_478[409:0]    ),
    .col_out_479             ( u0_col_out_479[409:0]    ),
    .col_out_480             ( u0_col_out_480[409:0]    ),
    .col_out_481             ( u0_col_out_481[409:0]    ),
    .col_out_482             ( u0_col_out_482[409:0]    ),
    .col_out_483             ( u0_col_out_483[409:0]    ),
    .col_out_484             ( u0_col_out_484[409:0]    ),
    .col_out_485             ( u0_col_out_485[409:0]    ),
    .col_out_486             ( u0_col_out_486[409:0]    ),
    .col_out_487             ( u0_col_out_487[409:0]    ),
    .col_out_488             ( u0_col_out_488[409:0]    ),
    .col_out_489             ( u0_col_out_489[409:0]    ),
    .col_out_490             ( u0_col_out_490[409:0]    ),
    .col_out_491             ( u0_col_out_491[409:0]    ),
    .col_out_492             ( u0_col_out_492[409:0]    ),
    .col_out_493             ( u0_col_out_493[409:0]    ),
    .col_out_494             ( u0_col_out_494[409:0]    ),
    .col_out_495             ( u0_col_out_495[409:0]    ),
    .col_out_496             ( u0_col_out_496[409:0]    ),
    .col_out_497             ( u0_col_out_497[409:0]    ),
    .col_out_498             ( u0_col_out_498[409:0]    ),
    .col_out_499             ( u0_col_out_499[409:0]    ),
    .col_out_500             ( u0_col_out_500[409:0]    ),
    .col_out_501             ( u0_col_out_501[409:0]    ),
    .col_out_502             ( u0_col_out_502[409:0]    ),
    .col_out_503             ( u0_col_out_503[409:0]    ),
    .col_out_504             ( u0_col_out_504[409:0]    ),
    .col_out_505             ( u0_col_out_505[409:0]    ),
    .col_out_506             ( u0_col_out_506[409:0]    ),
    .col_out_507             ( u0_col_out_507[409:0]    ),
    .col_out_508             ( u0_col_out_508[409:0]    ),
    .col_out_509             ( u0_col_out_509[409:0]    ),
    .col_out_510             ( u0_col_out_510[409:0]    ),
    .col_out_511             ( u0_col_out_511[409:0]    ),
    .col_out_512             ( u0_col_out_512[409:0]    ),
    .col_out_513             ( u0_col_out_513[409:0]    ),
    .col_out_514             ( u0_col_out_514[409:0]    ),
    .col_out_515             ( u0_col_out_515[409:0]    ),
    .col_out_516             ( u0_col_out_516[409:0]    ),
    .col_out_517             ( u0_col_out_517[409:0]    ),
    .col_out_518             ( u0_col_out_518[409:0]    ),
    .col_out_519             ( u0_col_out_519[409:0]    ),
    .col_out_520             ( u0_col_out_520[409:0]    ),
    .col_out_521             ( u0_col_out_521[409:0]    ),
    .col_out_522             ( u0_col_out_522[409:0]    ),
    .col_out_523             ( u0_col_out_523[409:0]    ),
    .col_out_524             ( u0_col_out_524[409:0]    ),
    .col_out_525             ( u0_col_out_525[409:0]    ),
    .col_out_526             ( u0_col_out_526[409:0]    ),
    .col_out_527             ( u0_col_out_527[409:0]    ),
    .col_out_528             ( u0_col_out_528[409:0]    ),
    .col_out_529             ( u0_col_out_529[409:0]    ),
    .col_out_530             ( u0_col_out_530[409:0]    ),
    .col_out_531             ( u0_col_out_531[409:0]    ),
    .col_out_532             ( u0_col_out_532[409:0]    ),
    .col_out_533             ( u0_col_out_533[409:0]    ),
    .col_out_534             ( u0_col_out_534[409:0]    ),
    .col_out_535             ( u0_col_out_535[409:0]    ),
    .col_out_536             ( u0_col_out_536[409:0]    ),
    .col_out_537             ( u0_col_out_537[409:0]    ),
    .col_out_538             ( u0_col_out_538[409:0]    ),
    .col_out_539             ( u0_col_out_539[409:0]    ),
    .col_out_540             ( u0_col_out_540[409:0]    ),
    .col_out_541             ( u0_col_out_541[409:0]    ),
    .col_out_542             ( u0_col_out_542[409:0]    ),
    .col_out_543             ( u0_col_out_543[409:0]    ),
    .col_out_544             ( u0_col_out_544[409:0]    ),
    .col_out_545             ( u0_col_out_545[409:0]    ),
    .col_out_546             ( u0_col_out_546[409:0]    ),
    .col_out_547             ( u0_col_out_547[409:0]    ),
    .col_out_548             ( u0_col_out_548[409:0]    ),
    .col_out_549             ( u0_col_out_549[409:0]    ),
    .col_out_550             ( u0_col_out_550[409:0]    ),
    .col_out_551             ( u0_col_out_551[409:0]    ),
    .col_out_552             ( u0_col_out_552[409:0]    ),
    .col_out_553             ( u0_col_out_553[409:0]    ),
    .col_out_554             ( u0_col_out_554[409:0]    ),
    .col_out_555             ( u0_col_out_555[409:0]    ),
    .col_out_556             ( u0_col_out_556[409:0]    ),
    .col_out_557             ( u0_col_out_557[409:0]    ),
    .col_out_558             ( u0_col_out_558[409:0]    ),
    .col_out_559             ( u0_col_out_559[409:0]    ),
    .col_out_560             ( u0_col_out_560[409:0]    ),
    .col_out_561             ( u0_col_out_561[409:0]    ),
    .col_out_562             ( u0_col_out_562[409:0]    ),
    .col_out_563             ( u0_col_out_563[409:0]    ),
    .col_out_564             ( u0_col_out_564[409:0]    ),
    .col_out_565             ( u0_col_out_565[409:0]    ),
    .col_out_566             ( u0_col_out_566[409:0]    ),
    .col_out_567             ( u0_col_out_567[409:0]    ),
    .col_out_568             ( u0_col_out_568[409:0]    ),
    .col_out_569             ( u0_col_out_569[409:0]    ),
    .col_out_570             ( u0_col_out_570[409:0]    ),
    .col_out_571             ( u0_col_out_571[409:0]    ),
    .col_out_572             ( u0_col_out_572[409:0]    ),
    .col_out_573             ( u0_col_out_573[409:0]    ),
    .col_out_574             ( u0_col_out_574[409:0]    ),
    .col_out_575             ( u0_col_out_575[409:0]    ),
    .col_out_576             ( u0_col_out_576[409:0]    ),
    .col_out_577             ( u0_col_out_577[409:0]    ),
    .col_out_578             ( u0_col_out_578[409:0]    ),
    .col_out_579             ( u0_col_out_579[409:0]    ),
    .col_out_580             ( u0_col_out_580[409:0]    ),
    .col_out_581             ( u0_col_out_581[409:0]    ),
    .col_out_582             ( u0_col_out_582[409:0]    ),
    .col_out_583             ( u0_col_out_583[409:0]    ),
    .col_out_584             ( u0_col_out_584[409:0]    ),
    .col_out_585             ( u0_col_out_585[409:0]    ),
    .col_out_586             ( u0_col_out_586[409:0]    ),
    .col_out_587             ( u0_col_out_587[409:0]    ),
    .col_out_588             ( u0_col_out_588[409:0]    ),
    .col_out_589             ( u0_col_out_589[409:0]    ),
    .col_out_590             ( u0_col_out_590[409:0]    ),
    .col_out_591             ( u0_col_out_591[409:0]    ),
    .col_out_592             ( u0_col_out_592[409:0]    ),
    .col_out_593             ( u0_col_out_593[409:0]    ),
    .col_out_594             ( u0_col_out_594[409:0]    ),
    .col_out_595             ( u0_col_out_595[409:0]    ),
    .col_out_596             ( u0_col_out_596[409:0]    ),
    .col_out_597             ( u0_col_out_597[409:0]    ),
    .col_out_598             ( u0_col_out_598[409:0]    ),
    .col_out_599             ( u0_col_out_599[409:0]    ),
    .col_out_600             ( u0_col_out_600[409:0]    ),
    .col_out_601             ( u0_col_out_601[409:0]    ),
    .col_out_602             ( u0_col_out_602[409:0]    ),
    .col_out_603             ( u0_col_out_603[409:0]    ),
    .col_out_604             ( u0_col_out_604[409:0]    ),
    .col_out_605             ( u0_col_out_605[409:0]    ),
    .col_out_606             ( u0_col_out_606[409:0]    ),
    .col_out_607             ( u0_col_out_607[409:0]    ),
    .col_out_608             ( u0_col_out_608[409:0]    ),
    .col_out_609             ( u0_col_out_609[409:0]    ),
    .col_out_610             ( u0_col_out_610[409:0]    ),
    .col_out_611             ( u0_col_out_611[409:0]    ),
    .col_out_612             ( u0_col_out_612[409:0]    ),
    .col_out_613             ( u0_col_out_613[409:0]    ),
    .col_out_614             ( u0_col_out_614[409:0]    ),
    .col_out_615             ( u0_col_out_615[409:0]    ),
    .col_out_616             ( u0_col_out_616[409:0]    ),
    .col_out_617             ( u0_col_out_617[409:0]    ),
    .col_out_618             ( u0_col_out_618[409:0]    ),
    .col_out_619             ( u0_col_out_619[409:0]    ),
    .col_out_620             ( u0_col_out_620[409:0]    ),
    .col_out_621             ( u0_col_out_621[409:0]    ),
    .col_out_622             ( u0_col_out_622[409:0]    ),
    .col_out_623             ( u0_col_out_623[409:0]    ),
    .col_out_624             ( u0_col_out_624[409:0]    ),
    .col_out_625             ( u0_col_out_625[409:0]    ),
    .col_out_626             ( u0_col_out_626[409:0]    ),
    .col_out_627             ( u0_col_out_627[409:0]    ),
    .col_out_628             ( u0_col_out_628[409:0]    ),
    .col_out_629             ( u0_col_out_629[409:0]    ),
    .col_out_630             ( u0_col_out_630[409:0]    ),
    .col_out_631             ( u0_col_out_631[409:0]    ),
    .col_out_632             ( u0_col_out_632[409:0]    ),
    .col_out_633             ( u0_col_out_633[409:0]    ),
    .col_out_634             ( u0_col_out_634[409:0]    ),
    .col_out_635             ( u0_col_out_635[409:0]    ),
    .col_out_636             ( u0_col_out_636[409:0]    ),
    .col_out_637             ( u0_col_out_637[409:0]    ),
    .col_out_638             ( u0_col_out_638[409:0]    ),
    .col_out_639             ( u0_col_out_639[409:0]    ),
    .col_out_640             ( u0_col_out_640[409:0]    ),
    .col_out_641             ( u0_col_out_641[409:0]    ),
    .col_out_642             ( u0_col_out_642[409:0]    ),
    .col_out_643             ( u0_col_out_643[409:0]    ),
    .col_out_644             ( u0_col_out_644[409:0]    ),
    .col_out_645             ( u0_col_out_645[409:0]    ),
    .col_out_646             ( u0_col_out_646[409:0]    ),
    .col_out_647             ( u0_col_out_647[409:0]    ),
    .col_out_648             ( u0_col_out_648[409:0]    ),
    .col_out_649             ( u0_col_out_649[409:0]    ),
    .col_out_650             ( u0_col_out_650[409:0]    ),
    .col_out_651             ( u0_col_out_651[409:0]    ),
    .col_out_652             ( u0_col_out_652[409:0]    ),
    .col_out_653             ( u0_col_out_653[409:0]    ),
    .col_out_654             ( u0_col_out_654[409:0]    ),
    .col_out_655             ( u0_col_out_655[409:0]    ),
    .col_out_656             ( u0_col_out_656[409:0]    ),
    .col_out_657             ( u0_col_out_657[409:0]    ),
    .col_out_658             ( u0_col_out_658[409:0]    ),
    .col_out_659             ( u0_col_out_659[409:0]    ),
    .col_out_660             ( u0_col_out_660[409:0]    ),
    .col_out_661             ( u0_col_out_661[409:0]    ),
    .col_out_662             ( u0_col_out_662[409:0]    ),
    .col_out_663             ( u0_col_out_663[409:0]    ),
    .col_out_664             ( u0_col_out_664[409:0]    ),
    .col_out_665             ( u0_col_out_665[409:0]    ),
    .col_out_666             ( u0_col_out_666[409:0]    ),
    .col_out_667             ( u0_col_out_667[409:0]    ),
    .col_out_668             ( u0_col_out_668[409:0]    ),
    .col_out_669             ( u0_col_out_669[409:0]    ),
    .col_out_670             ( u0_col_out_670[409:0]    ),
    .col_out_671             ( u0_col_out_671[409:0]    ),
    .col_out_672             ( u0_col_out_672[409:0]    ),
    .col_out_673             ( u0_col_out_673[409:0]    ),
    .col_out_674             ( u0_col_out_674[409:0]    ),
    .col_out_675             ( u0_col_out_675[409:0]    ),
    .col_out_676             ( u0_col_out_676[409:0]    ),
    .col_out_677             ( u0_col_out_677[409:0]    ),
    .col_out_678             ( u0_col_out_678[409:0]    ),
    .col_out_679             ( u0_col_out_679[409:0]    ),
    .col_out_680             ( u0_col_out_680[409:0]    ),
    .col_out_681             ( u0_col_out_681[409:0]    ),
    .col_out_682             ( u0_col_out_682[409:0]    ),
    .col_out_683             ( u0_col_out_683[409:0]    ),
    .col_out_684             ( u0_col_out_684[409:0]    ),
    .col_out_685             ( u0_col_out_685[409:0]    ),
    .col_out_686             ( u0_col_out_686[409:0]    ),
    .col_out_687             ( u0_col_out_687[409:0]    ),
    .col_out_688             ( u0_col_out_688[409:0]    ),
    .col_out_689             ( u0_col_out_689[409:0]    ),
    .col_out_690             ( u0_col_out_690[409:0]    ),
    .col_out_691             ( u0_col_out_691[409:0]    ),
    .col_out_692             ( u0_col_out_692[409:0]    ),
    .col_out_693             ( u0_col_out_693[409:0]    ),
    .col_out_694             ( u0_col_out_694[409:0]    ),
    .col_out_695             ( u0_col_out_695[409:0]    ),
    .col_out_696             ( u0_col_out_696[409:0]    ),
    .col_out_697             ( u0_col_out_697[409:0]    ),
    .col_out_698             ( u0_col_out_698[409:0]    ),
    .col_out_699             ( u0_col_out_699[409:0]    ),
    .col_out_700             ( u0_col_out_700[409:0]    ),
    .col_out_701             ( u0_col_out_701[409:0]    ),
    .col_out_702             ( u0_col_out_702[409:0]    ),
    .col_out_703             ( u0_col_out_703[409:0]    ),
    .col_out_704             ( u0_col_out_704[409:0]    ),
    .col_out_705             ( u0_col_out_705[409:0]    ),
    .col_out_706             ( u0_col_out_706[409:0]    ),
    .col_out_707             ( u0_col_out_707[409:0]    ),
    .col_out_708             ( u0_col_out_708[409:0]    ),
    .col_out_709             ( u0_col_out_709[409:0]    ),
    .col_out_710             ( u0_col_out_710[409:0]    ),
    .col_out_711             ( u0_col_out_711[409:0]    ),
    .col_out_712             ( u0_col_out_712[409:0]    ),
    .col_out_713             ( u0_col_out_713[409:0]    ),
    .col_out_714             ( u0_col_out_714[409:0]    ),
    .col_out_715             ( u0_col_out_715[409:0]    ),
    .col_out_716             ( u0_col_out_716[409:0]    ),
    .col_out_717             ( u0_col_out_717[409:0]    ),
    .col_out_718             ( u0_col_out_718[409:0]    ),
    .col_out_719             ( u0_col_out_719[409:0]    ),
    .col_out_720             ( u0_col_out_720[409:0]    ),
    .col_out_721             ( u0_col_out_721[409:0]    ),
    .col_out_722             ( u0_col_out_722[409:0]    ),
    .col_out_723             ( u0_col_out_723[409:0]    ),
    .col_out_724             ( u0_col_out_724[409:0]    ),
    .col_out_725             ( u0_col_out_725[409:0]    ),
    .col_out_726             ( u0_col_out_726[409:0]    ),
    .col_out_727             ( u0_col_out_727[409:0]    ),
    .col_out_728             ( u0_col_out_728[409:0]    ),
    .col_out_729             ( u0_col_out_729[409:0]    ),
    .col_out_730             ( u0_col_out_730[409:0]    ),
    .col_out_731             ( u0_col_out_731[409:0]    ),
    .col_out_732             ( u0_col_out_732[409:0]    ),
    .col_out_733             ( u0_col_out_733[409:0]    ),
    .col_out_734             ( u0_col_out_734[409:0]    ),
    .col_out_735             ( u0_col_out_735[409:0]    ),
    .col_out_736             ( u0_col_out_736[409:0]    ),
    .col_out_737             ( u0_col_out_737[409:0]    ),
    .col_out_738             ( u0_col_out_738[409:0]    ),
    .col_out_739             ( u0_col_out_739[409:0]    ),
    .col_out_740             ( u0_col_out_740[409:0]    ),
    .col_out_741             ( u0_col_out_741[409:0]    ),
    .col_out_742             ( u0_col_out_742[409:0]    ),
    .col_out_743             ( u0_col_out_743[409:0]    ),
    .col_out_744             ( u0_col_out_744[409:0]    ),
    .col_out_745             ( u0_col_out_745[409:0]    ),
    .col_out_746             ( u0_col_out_746[409:0]    ),
    .col_out_747             ( u0_col_out_747[409:0]    ),
    .col_out_748             ( u0_col_out_748[409:0]    ),
    .col_out_749             ( u0_col_out_749[409:0]    ),
    .col_out_750             ( u0_col_out_750[409:0]    ),
    .col_out_751             ( u0_col_out_751[409:0]    ),
    .col_out_752             ( u0_col_out_752[409:0]    ),
    .col_out_753             ( u0_col_out_753[409:0]    ),
    .col_out_754             ( u0_col_out_754[409:0]    ),
    .col_out_755             ( u0_col_out_755[409:0]    ),
    .col_out_756             ( u0_col_out_756[409:0]    ),
    .col_out_757             ( u0_col_out_757[409:0]    ),
    .col_out_758             ( u0_col_out_758[409:0]    ),
    .col_out_759             ( u0_col_out_759[409:0]    ),
    .col_out_760             ( u0_col_out_760[409:0]    ),
    .col_out_761             ( u0_col_out_761[409:0]    ),
    .col_out_762             ( u0_col_out_762[409:0]    ),
    .col_out_763             ( u0_col_out_763[409:0]    ),
    .col_out_764             ( u0_col_out_764[409:0]    ),
    .col_out_765             ( u0_col_out_765[409:0]    ),
    .col_out_766             ( u0_col_out_766[409:0]    ),
    .col_out_767             ( u0_col_out_767[409:0]    ),
    .col_out_768             ( u0_col_out_768[409:0]    ),
    .col_out_769             ( u0_col_out_769[409:0]    ),
    .col_out_770             ( u0_col_out_770[409:0]    ),
    .col_out_771             ( u0_col_out_771[409:0]    ),
    .col_out_772             ( u0_col_out_772[409:0]    ),
    .col_out_773             ( u0_col_out_773[409:0]    ),
    .col_out_774             ( u0_col_out_774[409:0]    ),
    .col_out_775             ( u0_col_out_775[409:0]    ),
    .col_out_776             ( u0_col_out_776[409:0]    ),
    .col_out_777             ( u0_col_out_777[409:0]    ),
    .col_out_778             ( u0_col_out_778[409:0]    ),
    .col_out_779             ( u0_col_out_779[409:0]    ),
    .col_out_780             ( u0_col_out_780[409:0]    ),
    .col_out_781             ( u0_col_out_781[409:0]    ),
    .col_out_782             ( u0_col_out_782[409:0]    ),
    .col_out_783             ( u0_col_out_783[409:0]    ),
    .col_out_784             ( u0_col_out_784[409:0]    ),
    .col_out_785             ( u0_col_out_785[409:0]    ),
    .col_out_786             ( u0_col_out_786[409:0]    ),
    .col_out_787             ( u0_col_out_787[409:0]    ),
    .col_out_788             ( u0_col_out_788[409:0]    ),
    .col_out_789             ( u0_col_out_789[409:0]    ),
    .col_out_790             ( u0_col_out_790[409:0]    ),
    .col_out_791             ( u0_col_out_791[409:0]    ),
    .col_out_792             ( u0_col_out_792[409:0]    ),
    .col_out_793             ( u0_col_out_793[409:0]    ),
    .col_out_794             ( u0_col_out_794[409:0]    ),
    .col_out_795             ( u0_col_out_795[409:0]    ),
    .col_out_796             ( u0_col_out_796[409:0]    ),
    .col_out_797             ( u0_col_out_797[409:0]    ),
    .col_out_798             ( u0_col_out_798[409:0]    ),
    .col_out_799             ( u0_col_out_799[409:0]    ),
    .col_out_800             ( u0_col_out_800[409:0]    ),
    .col_out_801             ( u0_col_out_801[409:0]    ),
    .col_out_802             ( u0_col_out_802[409:0]    ),
    .col_out_803             ( u0_col_out_803[409:0]    ),
    .col_out_804             ( u0_col_out_804[409:0]    ),
    .col_out_805             ( u0_col_out_805[409:0]    ),
    .col_out_806             ( u0_col_out_806[409:0]    ),
    .col_out_807             ( u0_col_out_807[409:0]    ),
    .col_out_808             ( u0_col_out_808[409:0]    ),
    .col_out_809             ( u0_col_out_809[409:0]    ),
    .col_out_810             ( u0_col_out_810[409:0]    ),
    .col_out_811             ( u0_col_out_811[409:0]    ),
    .col_out_812             ( u0_col_out_812[409:0]    ),
    .col_out_813             ( u0_col_out_813[409:0]    ),
    .col_out_814             ( u0_col_out_814[409:0]    ),
    .col_out_815             ( u0_col_out_815[409:0]    ),
    .col_out_816             ( u0_col_out_816[409:0]    ),
    .col_out_817             ( u0_col_out_817[409:0]    ),
    .col_out_818             ( u0_col_out_818[409:0]    ),
    .col_out_819             ( u0_col_out_819[409:0]    ),
    .col_out_820             ( u0_col_out_820[409:0]    ),
    .col_out_821             ( u0_col_out_821[409:0]    ),
    .col_out_822             ( u0_col_out_822[409:0]    ),
    .col_out_823             ( u0_col_out_823[409:0]    ),
    .col_out_824             ( u0_col_out_824[409:0]    ),
    .col_out_825             ( u0_col_out_825[409:0]    ),
    .col_out_826             ( u0_col_out_826[409:0]    ),
    .col_out_827             ( u0_col_out_827[409:0]    ),
    .col_out_828             ( u0_col_out_828[409:0]    ),
    .col_out_829             ( u0_col_out_829[409:0]    ),
    .col_out_830             ( u0_col_out_830[409:0]    ),
    .col_out_831             ( u0_col_out_831[409:0]    ),
    .col_out_832             ( u0_col_out_832[409:0]    ),
    .col_out_833             ( u0_col_out_833[409:0]    ),
    .col_out_834             ( u0_col_out_834[409:0]    ),
    .col_out_835             ( u0_col_out_835[409:0]    ),
    .col_out_836             ( u0_col_out_836[409:0]    ),
    .col_out_837             ( u0_col_out_837[409:0]    ),
    .col_out_838             ( u0_col_out_838[409:0]    ),
    .col_out_839             ( u0_col_out_839[409:0]    ),
    .col_out_840             ( u0_col_out_840[409:0]    ),
    .col_out_841             ( u0_col_out_841[409:0]    ),
    .col_out_842             ( u0_col_out_842[409:0]    ),
    .col_out_843             ( u0_col_out_843[409:0]    ),
    .col_out_844             ( u0_col_out_844[409:0]    ),
    .col_out_845             ( u0_col_out_845[409:0]    ),
    .col_out_846             ( u0_col_out_846[409:0]    ),
    .col_out_847             ( u0_col_out_847[409:0]    ),
    .col_out_848             ( u0_col_out_848[409:0]    ),
    .col_out_849             ( u0_col_out_849[409:0]    ),
    .col_out_850             ( u0_col_out_850[409:0]    ),
    .col_out_851             ( u0_col_out_851[409:0]    ),
    .col_out_852             ( u0_col_out_852[409:0]    ),
    .col_out_853             ( u0_col_out_853[409:0]    ),
    .col_out_854             ( u0_col_out_854[409:0]    ),
    .col_out_855             ( u0_col_out_855[409:0]    ),
    .col_out_856             ( u0_col_out_856[409:0]    ),
    .col_out_857             ( u0_col_out_857[409:0]    ),
    .col_out_858             ( u0_col_out_858[409:0]    ),
    .col_out_859             ( u0_col_out_859[409:0]    ),
    .col_out_860             ( u0_col_out_860[409:0]    ),
    .col_out_861             ( u0_col_out_861[409:0]    ),
    .col_out_862             ( u0_col_out_862[409:0]    ),
    .col_out_863             ( u0_col_out_863[409:0]    ),
    .col_out_864             ( u0_col_out_864[409:0]    ),
    .col_out_865             ( u0_col_out_865[409:0]    ),
    .col_out_866             ( u0_col_out_866[409:0]    ),
    .col_out_867             ( u0_col_out_867[409:0]    ),
    .col_out_868             ( u0_col_out_868[409:0]    ),
    .col_out_869             ( u0_col_out_869[409:0]    ),
    .col_out_870             ( u0_col_out_870[409:0]    ),
    .col_out_871             ( u0_col_out_871[409:0]    ),
    .col_out_872             ( u0_col_out_872[409:0]    ),
    .col_out_873             ( u0_col_out_873[409:0]    ),
    .col_out_874             ( u0_col_out_874[409:0]    ),
    .col_out_875             ( u0_col_out_875[409:0]    ),
    .col_out_876             ( u0_col_out_876[409:0]    ),
    .col_out_877             ( u0_col_out_877[409:0]    ),
    .col_out_878             ( u0_col_out_878[409:0]    ),
    .col_out_879             ( u0_col_out_879[409:0]    ),
    .col_out_880             ( u0_col_out_880[409:0]    ),
    .col_out_881             ( u0_col_out_881[409:0]    ),
    .col_out_882             ( u0_col_out_882[409:0]    ),
    .col_out_883             ( u0_col_out_883[409:0]    ),
    .col_out_884             ( u0_col_out_884[409:0]    ),
    .col_out_885             ( u0_col_out_885[409:0]    ),
    .col_out_886             ( u0_col_out_886[409:0]    ),
    .col_out_887             ( u0_col_out_887[409:0]    ),
    .col_out_888             ( u0_col_out_888[409:0]    ),
    .col_out_889             ( u0_col_out_889[409:0]    ),
    .col_out_890             ( u0_col_out_890[409:0]    ),
    .col_out_891             ( u0_col_out_891[409:0]    ),
    .col_out_892             ( u0_col_out_892[409:0]    ),
    .col_out_893             ( u0_col_out_893[409:0]    ),
    .col_out_894             ( u0_col_out_894[409:0]    ),
    .col_out_895             ( u0_col_out_895[409:0]    ),
    .col_out_896             ( u0_col_out_896[409:0]    ),
    .col_out_897             ( u0_col_out_897[409:0]    ),
    .col_out_898             ( u0_col_out_898[409:0]    ),
    .col_out_899             ( u0_col_out_899[409:0]    ),
    .col_out_900             ( u0_col_out_900[409:0]    ),
    .col_out_901             ( u0_col_out_901[409:0]    ),
    .col_out_902             ( u0_col_out_902[409:0]    ),
    .col_out_903             ( u0_col_out_903[409:0]    ),
    .col_out_904             ( u0_col_out_904[409:0]    ),
    .col_out_905             ( u0_col_out_905[409:0]    ),
    .col_out_906             ( u0_col_out_906[409:0]    ),
    .col_out_907             ( u0_col_out_907[409:0]    ),
    .col_out_908             ( u0_col_out_908[409:0]    ),
    .col_out_909             ( u0_col_out_909[409:0]    ),
    .col_out_910             ( u0_col_out_910[409:0]    ),
    .col_out_911             ( u0_col_out_911[409:0]    ),
    .col_out_912             ( u0_col_out_912[409:0]    ),
    .col_out_913             ( u0_col_out_913[409:0]    ),
    .col_out_914             ( u0_col_out_914[409:0]    ),
    .col_out_915             ( u0_col_out_915[409:0]    ),
    .col_out_916             ( u0_col_out_916[409:0]    ),
    .col_out_917             ( u0_col_out_917[409:0]    ),
    .col_out_918             ( u0_col_out_918[409:0]    ),
    .col_out_919             ( u0_col_out_919[409:0]    ),
    .col_out_920             ( u0_col_out_920[409:0]    ),
    .col_out_921             ( u0_col_out_921[409:0]    ),
    .col_out_922             ( u0_col_out_922[409:0]    ),
    .col_out_923             ( u0_col_out_923[409:0]    ),
    .col_out_924             ( u0_col_out_924[409:0]    ),
    .col_out_925             ( u0_col_out_925[409:0]    ),
    .col_out_926             ( u0_col_out_926[409:0]    ),
    .col_out_927             ( u0_col_out_927[409:0]    ),
    .col_out_928             ( u0_col_out_928[409:0]    ),
    .col_out_929             ( u0_col_out_929[409:0]    ),
    .col_out_930             ( u0_col_out_930[409:0]    ),
    .col_out_931             ( u0_col_out_931[409:0]    ),
    .col_out_932             ( u0_col_out_932[409:0]    ),
    .col_out_933             ( u0_col_out_933[409:0]    ),
    .col_out_934             ( u0_col_out_934[409:0]    ),
    .col_out_935             ( u0_col_out_935[409:0]    ),
    .col_out_936             ( u0_col_out_936[409:0]    ),
    .col_out_937             ( u0_col_out_937[409:0]    ),
    .col_out_938             ( u0_col_out_938[409:0]    ),
    .col_out_939             ( u0_col_out_939[409:0]    ),
    .col_out_940             ( u0_col_out_940[409:0]    ),
    .col_out_941             ( u0_col_out_941[409:0]    ),
    .col_out_942             ( u0_col_out_942[409:0]    ),
    .col_out_943             ( u0_col_out_943[409:0]    ),
    .col_out_944             ( u0_col_out_944[409:0]    ),
    .col_out_945             ( u0_col_out_945[409:0]    ),
    .col_out_946             ( u0_col_out_946[409:0]    ),
    .col_out_947             ( u0_col_out_947[409:0]    ),
    .col_out_948             ( u0_col_out_948[409:0]    ),
    .col_out_949             ( u0_col_out_949[409:0]    ),
    .col_out_950             ( u0_col_out_950[409:0]    ),
    .col_out_951             ( u0_col_out_951[409:0]    ),
    .col_out_952             ( u0_col_out_952[409:0]    ),
    .col_out_953             ( u0_col_out_953[409:0]    ),
    .col_out_954             ( u0_col_out_954[409:0]    ),
    .col_out_955             ( u0_col_out_955[409:0]    ),
    .col_out_956             ( u0_col_out_956[409:0]    ),
    .col_out_957             ( u0_col_out_957[409:0]    ),
    .col_out_958             ( u0_col_out_958[409:0]    ),
    .col_out_959             ( u0_col_out_959[409:0]    ),
    .col_out_960             ( u0_col_out_960[409:0]    ),
    .col_out_961             ( u0_col_out_961[409:0]    ),
    .col_out_962             ( u0_col_out_962[409:0]    ),
    .col_out_963             ( u0_col_out_963[409:0]    ),
    .col_out_964             ( u0_col_out_964[409:0]    ),
    .col_out_965             ( u0_col_out_965[409:0]    ),
    .col_out_966             ( u0_col_out_966[409:0]    ),
    .col_out_967             ( u0_col_out_967[409:0]    ),
    .col_out_968             ( u0_col_out_968[409:0]    ),
    .col_out_969             ( u0_col_out_969[409:0]    ),
    .col_out_970             ( u0_col_out_970[409:0]    ),
    .col_out_971             ( u0_col_out_971[409:0]    ),
    .col_out_972             ( u0_col_out_972[409:0]    ),
    .col_out_973             ( u0_col_out_973[409:0]    ),
    .col_out_974             ( u0_col_out_974[409:0]    ),
    .col_out_975             ( u0_col_out_975[409:0]    ),
    .col_out_976             ( u0_col_out_976[409:0]    ),
    .col_out_977             ( u0_col_out_977[409:0]    ),
    .col_out_978             ( u0_col_out_978[409:0]    ),
    .col_out_979             ( u0_col_out_979[409:0]    ),
    .col_out_980             ( u0_col_out_980[409:0]    ),
    .col_out_981             ( u0_col_out_981[409:0]    ),
    .col_out_982             ( u0_col_out_982[409:0]    ),
    .col_out_983             ( u0_col_out_983[409:0]    ),
    .col_out_984             ( u0_col_out_984[409:0]    ),
    .col_out_985             ( u0_col_out_985[409:0]    ),
    .col_out_986             ( u0_col_out_986[409:0]    ),
    .col_out_987             ( u0_col_out_987[409:0]    ),
    .col_out_988             ( u0_col_out_988[409:0]    ),
    .col_out_989             ( u0_col_out_989[409:0]    ),
    .col_out_990             ( u0_col_out_990[409:0]    ),
    .col_out_991             ( u0_col_out_991[409:0]    ),
    .col_out_992             ( u0_col_out_992[409:0]    ),
    .col_out_993             ( u0_col_out_993[409:0]    ),
    .col_out_994             ( u0_col_out_994[409:0]    ),
    .col_out_995             ( u0_col_out_995[409:0]    ),
    .col_out_996             ( u0_col_out_996[409:0]    ),
    .col_out_997             ( u0_col_out_997[409:0]    ),
    .col_out_998             ( u0_col_out_998[409:0]    ),
    .col_out_999             ( u0_col_out_999[409:0]    ),
    .col_out_1000            ( u0_col_out_1000[409:0]   ),
    .col_out_1001            ( u0_col_out_1001[409:0]   ),
    .col_out_1002            ( u0_col_out_1002[409:0]   ),
    .col_out_1003            ( u0_col_out_1003[409:0]   ),
    .col_out_1004            ( u0_col_out_1004[409:0]   ),
    .col_out_1005            ( u0_col_out_1005[409:0]   ),
    .col_out_1006            ( u0_col_out_1006[409:0]   ),
    .col_out_1007            ( u0_col_out_1007[409:0]   ),
    .col_out_1008            ( u0_col_out_1008[409:0]   ),
    .col_out_1009            ( u0_col_out_1009[409:0]   ),
    .col_out_1010            ( u0_col_out_1010[409:0]   ),
    .col_out_1011            ( u0_col_out_1011[409:0]   ),
    .col_out_1012            ( u0_col_out_1012[409:0]   ),
    .col_out_1013            ( u0_col_out_1013[409:0]   ),
    .col_out_1014            ( u0_col_out_1014[409:0]   ),
    .col_out_1015            ( u0_col_out_1015[409:0]   ),
    .col_out_1016            ( u0_col_out_1016[409:0]   ),
    .col_out_1017            ( u0_col_out_1017[409:0]   ),
    .col_out_1018            ( u0_col_out_1018[409:0]   ),
    .col_out_1019            ( u0_col_out_1019[409:0]   ),
    .col_out_1020            ( u0_col_out_1020[409:0]   ),
    .col_out_1021            ( u0_col_out_1021[409:0]   ),
    .col_out_1022            ( u0_col_out_1022[409:0]   ),
    .col_out_1023            ( u0_col_out_1023[409:0]   )
);




// xpb_18 Outputs
wire  [1023:0]  u1_data_out_0;
wire  [1023:0]  u1_data_out_1;
wire  [1023:0]  u1_data_out_2;
wire  [1023:0]  u1_data_out_3;

xpb_18  u1_xpb_18 (
    .data_in0                ( partial_product_low0[1032:1024]     ),
    .data_in1                ( partial_product_low1[1032:1024]      ),

    .data_out_0              ( u1_data_out_0   ),
    .data_out_1              ( u1_data_out_1   ),
    .data_out_2              ( u1_data_out_2   ),
    .data_out_3              ( u1_data_out_3   )
);






assign col_out_0 = {u0_col_out_0,u1_data_out_0[0],u1_data_out_1[0],u1_data_out_2[0],u1_data_out_3[0],partial_product_low0[0],partial_product_low1[0],96'b0};
assign col_out_1 = {u0_col_out_1,u1_data_out_0[1],u1_data_out_1[1],u1_data_out_2[1],u1_data_out_3[1],partial_product_low0[1],partial_product_low1[1],96'b0};
assign col_out_2 = {u0_col_out_2,u1_data_out_0[2],u1_data_out_1[2],u1_data_out_2[2],u1_data_out_3[2],partial_product_low0[2],partial_product_low1[2],96'b0};
assign col_out_3 = {u0_col_out_3,u1_data_out_0[3],u1_data_out_1[3],u1_data_out_2[3],u1_data_out_3[3],partial_product_low0[3],partial_product_low1[3],96'b0};
assign col_out_4 = {u0_col_out_4,u1_data_out_0[4],u1_data_out_1[4],u1_data_out_2[4],u1_data_out_3[4],partial_product_low0[4],partial_product_low1[4],96'b0};
assign col_out_5 = {u0_col_out_5,u1_data_out_0[5],u1_data_out_1[5],u1_data_out_2[5],u1_data_out_3[5],partial_product_low0[5],partial_product_low1[5],96'b0};
assign col_out_6 = {u0_col_out_6,u1_data_out_0[6],u1_data_out_1[6],u1_data_out_2[6],u1_data_out_3[6],partial_product_low0[6],partial_product_low1[6],96'b0};
assign col_out_7 = {u0_col_out_7,u1_data_out_0[7],u1_data_out_1[7],u1_data_out_2[7],u1_data_out_3[7],partial_product_low0[7],partial_product_low1[7],96'b0};
assign col_out_8 = {u0_col_out_8,u1_data_out_0[8],u1_data_out_1[8],u1_data_out_2[8],u1_data_out_3[8],partial_product_low0[8],partial_product_low1[8],96'b0};
assign col_out_9 = {u0_col_out_9,u1_data_out_0[9],u1_data_out_1[9],u1_data_out_2[9],u1_data_out_3[9],partial_product_low0[9],partial_product_low1[9],96'b0};
assign col_out_10 = {u0_col_out_10,u1_data_out_0[10],u1_data_out_1[10],u1_data_out_2[10],u1_data_out_3[10],partial_product_low0[10],partial_product_low1[10],96'b0};
assign col_out_11 = {u0_col_out_11,u1_data_out_0[11],u1_data_out_1[11],u1_data_out_2[11],u1_data_out_3[11],partial_product_low0[11],partial_product_low1[11],96'b0};
assign col_out_12 = {u0_col_out_12,u1_data_out_0[12],u1_data_out_1[12],u1_data_out_2[12],u1_data_out_3[12],partial_product_low0[12],partial_product_low1[12],96'b0};
assign col_out_13 = {u0_col_out_13,u1_data_out_0[13],u1_data_out_1[13],u1_data_out_2[13],u1_data_out_3[13],partial_product_low0[13],partial_product_low1[13],96'b0};
assign col_out_14 = {u0_col_out_14,u1_data_out_0[14],u1_data_out_1[14],u1_data_out_2[14],u1_data_out_3[14],partial_product_low0[14],partial_product_low1[14],96'b0};
assign col_out_15 = {u0_col_out_15,u1_data_out_0[15],u1_data_out_1[15],u1_data_out_2[15],u1_data_out_3[15],partial_product_low0[15],partial_product_low1[15],96'b0};
assign col_out_16 = {u0_col_out_16,u1_data_out_0[16],u1_data_out_1[16],u1_data_out_2[16],u1_data_out_3[16],partial_product_low0[16],partial_product_low1[16],96'b0};
assign col_out_17 = {u0_col_out_17,u1_data_out_0[17],u1_data_out_1[17],u1_data_out_2[17],u1_data_out_3[17],partial_product_low0[17],partial_product_low1[17],96'b0};
assign col_out_18 = {u0_col_out_18,u1_data_out_0[18],u1_data_out_1[18],u1_data_out_2[18],u1_data_out_3[18],partial_product_low0[18],partial_product_low1[18],96'b0};
assign col_out_19 = {u0_col_out_19,u1_data_out_0[19],u1_data_out_1[19],u1_data_out_2[19],u1_data_out_3[19],partial_product_low0[19],partial_product_low1[19],96'b0};
assign col_out_20 = {u0_col_out_20,u1_data_out_0[20],u1_data_out_1[20],u1_data_out_2[20],u1_data_out_3[20],partial_product_low0[20],partial_product_low1[20],96'b0};
assign col_out_21 = {u0_col_out_21,u1_data_out_0[21],u1_data_out_1[21],u1_data_out_2[21],u1_data_out_3[21],partial_product_low0[21],partial_product_low1[21],96'b0};
assign col_out_22 = {u0_col_out_22,u1_data_out_0[22],u1_data_out_1[22],u1_data_out_2[22],u1_data_out_3[22],partial_product_low0[22],partial_product_low1[22],96'b0};
assign col_out_23 = {u0_col_out_23,u1_data_out_0[23],u1_data_out_1[23],u1_data_out_2[23],u1_data_out_3[23],partial_product_low0[23],partial_product_low1[23],96'b0};
assign col_out_24 = {u0_col_out_24,u1_data_out_0[24],u1_data_out_1[24],u1_data_out_2[24],u1_data_out_3[24],partial_product_low0[24],partial_product_low1[24],96'b0};
assign col_out_25 = {u0_col_out_25,u1_data_out_0[25],u1_data_out_1[25],u1_data_out_2[25],u1_data_out_3[25],partial_product_low0[25],partial_product_low1[25],96'b0};
assign col_out_26 = {u0_col_out_26,u1_data_out_0[26],u1_data_out_1[26],u1_data_out_2[26],u1_data_out_3[26],partial_product_low0[26],partial_product_low1[26],96'b0};
assign col_out_27 = {u0_col_out_27,u1_data_out_0[27],u1_data_out_1[27],u1_data_out_2[27],u1_data_out_3[27],partial_product_low0[27],partial_product_low1[27],96'b0};
assign col_out_28 = {u0_col_out_28,u1_data_out_0[28],u1_data_out_1[28],u1_data_out_2[28],u1_data_out_3[28],partial_product_low0[28],partial_product_low1[28],96'b0};
assign col_out_29 = {u0_col_out_29,u1_data_out_0[29],u1_data_out_1[29],u1_data_out_2[29],u1_data_out_3[29],partial_product_low0[29],partial_product_low1[29],96'b0};
assign col_out_30 = {u0_col_out_30,u1_data_out_0[30],u1_data_out_1[30],u1_data_out_2[30],u1_data_out_3[30],partial_product_low0[30],partial_product_low1[30],96'b0};
assign col_out_31 = {u0_col_out_31,u1_data_out_0[31],u1_data_out_1[31],u1_data_out_2[31],u1_data_out_3[31],partial_product_low0[31],partial_product_low1[31],96'b0};
assign col_out_32 = {u0_col_out_32,u1_data_out_0[32],u1_data_out_1[32],u1_data_out_2[32],u1_data_out_3[32],partial_product_low0[32],partial_product_low1[32],96'b0};
assign col_out_33 = {u0_col_out_33,u1_data_out_0[33],u1_data_out_1[33],u1_data_out_2[33],u1_data_out_3[33],partial_product_low0[33],partial_product_low1[33],96'b0};
assign col_out_34 = {u0_col_out_34,u1_data_out_0[34],u1_data_out_1[34],u1_data_out_2[34],u1_data_out_3[34],partial_product_low0[34],partial_product_low1[34],96'b0};
assign col_out_35 = {u0_col_out_35,u1_data_out_0[35],u1_data_out_1[35],u1_data_out_2[35],u1_data_out_3[35],partial_product_low0[35],partial_product_low1[35],96'b0};
assign col_out_36 = {u0_col_out_36,u1_data_out_0[36],u1_data_out_1[36],u1_data_out_2[36],u1_data_out_3[36],partial_product_low0[36],partial_product_low1[36],96'b0};
assign col_out_37 = {u0_col_out_37,u1_data_out_0[37],u1_data_out_1[37],u1_data_out_2[37],u1_data_out_3[37],partial_product_low0[37],partial_product_low1[37],96'b0};
assign col_out_38 = {u0_col_out_38,u1_data_out_0[38],u1_data_out_1[38],u1_data_out_2[38],u1_data_out_3[38],partial_product_low0[38],partial_product_low1[38],96'b0};
assign col_out_39 = {u0_col_out_39,u1_data_out_0[39],u1_data_out_1[39],u1_data_out_2[39],u1_data_out_3[39],partial_product_low0[39],partial_product_low1[39],96'b0};
assign col_out_40 = {u0_col_out_40,u1_data_out_0[40],u1_data_out_1[40],u1_data_out_2[40],u1_data_out_3[40],partial_product_low0[40],partial_product_low1[40],96'b0};
assign col_out_41 = {u0_col_out_41,u1_data_out_0[41],u1_data_out_1[41],u1_data_out_2[41],u1_data_out_3[41],partial_product_low0[41],partial_product_low1[41],96'b0};
assign col_out_42 = {u0_col_out_42,u1_data_out_0[42],u1_data_out_1[42],u1_data_out_2[42],u1_data_out_3[42],partial_product_low0[42],partial_product_low1[42],96'b0};
assign col_out_43 = {u0_col_out_43,u1_data_out_0[43],u1_data_out_1[43],u1_data_out_2[43],u1_data_out_3[43],partial_product_low0[43],partial_product_low1[43],96'b0};
assign col_out_44 = {u0_col_out_44,u1_data_out_0[44],u1_data_out_1[44],u1_data_out_2[44],u1_data_out_3[44],partial_product_low0[44],partial_product_low1[44],96'b0};
assign col_out_45 = {u0_col_out_45,u1_data_out_0[45],u1_data_out_1[45],u1_data_out_2[45],u1_data_out_3[45],partial_product_low0[45],partial_product_low1[45],96'b0};
assign col_out_46 = {u0_col_out_46,u1_data_out_0[46],u1_data_out_1[46],u1_data_out_2[46],u1_data_out_3[46],partial_product_low0[46],partial_product_low1[46],96'b0};
assign col_out_47 = {u0_col_out_47,u1_data_out_0[47],u1_data_out_1[47],u1_data_out_2[47],u1_data_out_3[47],partial_product_low0[47],partial_product_low1[47],96'b0};
assign col_out_48 = {u0_col_out_48,u1_data_out_0[48],u1_data_out_1[48],u1_data_out_2[48],u1_data_out_3[48],partial_product_low0[48],partial_product_low1[48],96'b0};
assign col_out_49 = {u0_col_out_49,u1_data_out_0[49],u1_data_out_1[49],u1_data_out_2[49],u1_data_out_3[49],partial_product_low0[49],partial_product_low1[49],96'b0};
assign col_out_50 = {u0_col_out_50,u1_data_out_0[50],u1_data_out_1[50],u1_data_out_2[50],u1_data_out_3[50],partial_product_low0[50],partial_product_low1[50],96'b0};
assign col_out_51 = {u0_col_out_51,u1_data_out_0[51],u1_data_out_1[51],u1_data_out_2[51],u1_data_out_3[51],partial_product_low0[51],partial_product_low1[51],96'b0};
assign col_out_52 = {u0_col_out_52,u1_data_out_0[52],u1_data_out_1[52],u1_data_out_2[52],u1_data_out_3[52],partial_product_low0[52],partial_product_low1[52],96'b0};
assign col_out_53 = {u0_col_out_53,u1_data_out_0[53],u1_data_out_1[53],u1_data_out_2[53],u1_data_out_3[53],partial_product_low0[53],partial_product_low1[53],96'b0};
assign col_out_54 = {u0_col_out_54,u1_data_out_0[54],u1_data_out_1[54],u1_data_out_2[54],u1_data_out_3[54],partial_product_low0[54],partial_product_low1[54],96'b0};
assign col_out_55 = {u0_col_out_55,u1_data_out_0[55],u1_data_out_1[55],u1_data_out_2[55],u1_data_out_3[55],partial_product_low0[55],partial_product_low1[55],96'b0};
assign col_out_56 = {u0_col_out_56,u1_data_out_0[56],u1_data_out_1[56],u1_data_out_2[56],u1_data_out_3[56],partial_product_low0[56],partial_product_low1[56],96'b0};
assign col_out_57 = {u0_col_out_57,u1_data_out_0[57],u1_data_out_1[57],u1_data_out_2[57],u1_data_out_3[57],partial_product_low0[57],partial_product_low1[57],96'b0};
assign col_out_58 = {u0_col_out_58,u1_data_out_0[58],u1_data_out_1[58],u1_data_out_2[58],u1_data_out_3[58],partial_product_low0[58],partial_product_low1[58],96'b0};
assign col_out_59 = {u0_col_out_59,u1_data_out_0[59],u1_data_out_1[59],u1_data_out_2[59],u1_data_out_3[59],partial_product_low0[59],partial_product_low1[59],96'b0};
assign col_out_60 = {u0_col_out_60,u1_data_out_0[60],u1_data_out_1[60],u1_data_out_2[60],u1_data_out_3[60],partial_product_low0[60],partial_product_low1[60],96'b0};
assign col_out_61 = {u0_col_out_61,u1_data_out_0[61],u1_data_out_1[61],u1_data_out_2[61],u1_data_out_3[61],partial_product_low0[61],partial_product_low1[61],96'b0};
assign col_out_62 = {u0_col_out_62,u1_data_out_0[62],u1_data_out_1[62],u1_data_out_2[62],u1_data_out_3[62],partial_product_low0[62],partial_product_low1[62],96'b0};
assign col_out_63 = {u0_col_out_63,u1_data_out_0[63],u1_data_out_1[63],u1_data_out_2[63],u1_data_out_3[63],partial_product_low0[63],partial_product_low1[63],96'b0};
assign col_out_64 = {u0_col_out_64,u1_data_out_0[64],u1_data_out_1[64],u1_data_out_2[64],u1_data_out_3[64],partial_product_low0[64],partial_product_low1[64],96'b0};
assign col_out_65 = {u0_col_out_65,u1_data_out_0[65],u1_data_out_1[65],u1_data_out_2[65],u1_data_out_3[65],partial_product_low0[65],partial_product_low1[65],96'b0};
assign col_out_66 = {u0_col_out_66,u1_data_out_0[66],u1_data_out_1[66],u1_data_out_2[66],u1_data_out_3[66],partial_product_low0[66],partial_product_low1[66],96'b0};
assign col_out_67 = {u0_col_out_67,u1_data_out_0[67],u1_data_out_1[67],u1_data_out_2[67],u1_data_out_3[67],partial_product_low0[67],partial_product_low1[67],96'b0};
assign col_out_68 = {u0_col_out_68,u1_data_out_0[68],u1_data_out_1[68],u1_data_out_2[68],u1_data_out_3[68],partial_product_low0[68],partial_product_low1[68],96'b0};
assign col_out_69 = {u0_col_out_69,u1_data_out_0[69],u1_data_out_1[69],u1_data_out_2[69],u1_data_out_3[69],partial_product_low0[69],partial_product_low1[69],96'b0};
assign col_out_70 = {u0_col_out_70,u1_data_out_0[70],u1_data_out_1[70],u1_data_out_2[70],u1_data_out_3[70],partial_product_low0[70],partial_product_low1[70],96'b0};
assign col_out_71 = {u0_col_out_71,u1_data_out_0[71],u1_data_out_1[71],u1_data_out_2[71],u1_data_out_3[71],partial_product_low0[71],partial_product_low1[71],96'b0};
assign col_out_72 = {u0_col_out_72,u1_data_out_0[72],u1_data_out_1[72],u1_data_out_2[72],u1_data_out_3[72],partial_product_low0[72],partial_product_low1[72],96'b0};
assign col_out_73 = {u0_col_out_73,u1_data_out_0[73],u1_data_out_1[73],u1_data_out_2[73],u1_data_out_3[73],partial_product_low0[73],partial_product_low1[73],96'b0};
assign col_out_74 = {u0_col_out_74,u1_data_out_0[74],u1_data_out_1[74],u1_data_out_2[74],u1_data_out_3[74],partial_product_low0[74],partial_product_low1[74],96'b0};
assign col_out_75 = {u0_col_out_75,u1_data_out_0[75],u1_data_out_1[75],u1_data_out_2[75],u1_data_out_3[75],partial_product_low0[75],partial_product_low1[75],96'b0};
assign col_out_76 = {u0_col_out_76,u1_data_out_0[76],u1_data_out_1[76],u1_data_out_2[76],u1_data_out_3[76],partial_product_low0[76],partial_product_low1[76],96'b0};
assign col_out_77 = {u0_col_out_77,u1_data_out_0[77],u1_data_out_1[77],u1_data_out_2[77],u1_data_out_3[77],partial_product_low0[77],partial_product_low1[77],96'b0};
assign col_out_78 = {u0_col_out_78,u1_data_out_0[78],u1_data_out_1[78],u1_data_out_2[78],u1_data_out_3[78],partial_product_low0[78],partial_product_low1[78],96'b0};
assign col_out_79 = {u0_col_out_79,u1_data_out_0[79],u1_data_out_1[79],u1_data_out_2[79],u1_data_out_3[79],partial_product_low0[79],partial_product_low1[79],96'b0};
assign col_out_80 = {u0_col_out_80,u1_data_out_0[80],u1_data_out_1[80],u1_data_out_2[80],u1_data_out_3[80],partial_product_low0[80],partial_product_low1[80],96'b0};
assign col_out_81 = {u0_col_out_81,u1_data_out_0[81],u1_data_out_1[81],u1_data_out_2[81],u1_data_out_3[81],partial_product_low0[81],partial_product_low1[81],96'b0};
assign col_out_82 = {u0_col_out_82,u1_data_out_0[82],u1_data_out_1[82],u1_data_out_2[82],u1_data_out_3[82],partial_product_low0[82],partial_product_low1[82],96'b0};
assign col_out_83 = {u0_col_out_83,u1_data_out_0[83],u1_data_out_1[83],u1_data_out_2[83],u1_data_out_3[83],partial_product_low0[83],partial_product_low1[83],96'b0};
assign col_out_84 = {u0_col_out_84,u1_data_out_0[84],u1_data_out_1[84],u1_data_out_2[84],u1_data_out_3[84],partial_product_low0[84],partial_product_low1[84],96'b0};
assign col_out_85 = {u0_col_out_85,u1_data_out_0[85],u1_data_out_1[85],u1_data_out_2[85],u1_data_out_3[85],partial_product_low0[85],partial_product_low1[85],96'b0};
assign col_out_86 = {u0_col_out_86,u1_data_out_0[86],u1_data_out_1[86],u1_data_out_2[86],u1_data_out_3[86],partial_product_low0[86],partial_product_low1[86],96'b0};
assign col_out_87 = {u0_col_out_87,u1_data_out_0[87],u1_data_out_1[87],u1_data_out_2[87],u1_data_out_3[87],partial_product_low0[87],partial_product_low1[87],96'b0};
assign col_out_88 = {u0_col_out_88,u1_data_out_0[88],u1_data_out_1[88],u1_data_out_2[88],u1_data_out_3[88],partial_product_low0[88],partial_product_low1[88],96'b0};
assign col_out_89 = {u0_col_out_89,u1_data_out_0[89],u1_data_out_1[89],u1_data_out_2[89],u1_data_out_3[89],partial_product_low0[89],partial_product_low1[89],96'b0};
assign col_out_90 = {u0_col_out_90,u1_data_out_0[90],u1_data_out_1[90],u1_data_out_2[90],u1_data_out_3[90],partial_product_low0[90],partial_product_low1[90],96'b0};
assign col_out_91 = {u0_col_out_91,u1_data_out_0[91],u1_data_out_1[91],u1_data_out_2[91],u1_data_out_3[91],partial_product_low0[91],partial_product_low1[91],96'b0};
assign col_out_92 = {u0_col_out_92,u1_data_out_0[92],u1_data_out_1[92],u1_data_out_2[92],u1_data_out_3[92],partial_product_low0[92],partial_product_low1[92],96'b0};
assign col_out_93 = {u0_col_out_93,u1_data_out_0[93],u1_data_out_1[93],u1_data_out_2[93],u1_data_out_3[93],partial_product_low0[93],partial_product_low1[93],96'b0};
assign col_out_94 = {u0_col_out_94,u1_data_out_0[94],u1_data_out_1[94],u1_data_out_2[94],u1_data_out_3[94],partial_product_low0[94],partial_product_low1[94],96'b0};
assign col_out_95 = {u0_col_out_95,u1_data_out_0[95],u1_data_out_1[95],u1_data_out_2[95],u1_data_out_3[95],partial_product_low0[95],partial_product_low1[95],96'b0};
assign col_out_96 = {u0_col_out_96,u1_data_out_0[96],u1_data_out_1[96],u1_data_out_2[96],u1_data_out_3[96],partial_product_low0[96],partial_product_low1[96],96'b0};
assign col_out_97 = {u0_col_out_97,u1_data_out_0[97],u1_data_out_1[97],u1_data_out_2[97],u1_data_out_3[97],partial_product_low0[97],partial_product_low1[97],96'b0};
assign col_out_98 = {u0_col_out_98,u1_data_out_0[98],u1_data_out_1[98],u1_data_out_2[98],u1_data_out_3[98],partial_product_low0[98],partial_product_low1[98],96'b0};
assign col_out_99 = {u0_col_out_99,u1_data_out_0[99],u1_data_out_1[99],u1_data_out_2[99],u1_data_out_3[99],partial_product_low0[99],partial_product_low1[99],96'b0};
assign col_out_100 = {u0_col_out_100,u1_data_out_0[100],u1_data_out_1[100],u1_data_out_2[100],u1_data_out_3[100],partial_product_low0[100],partial_product_low1[100],96'b0};
assign col_out_101 = {u0_col_out_101,u1_data_out_0[101],u1_data_out_1[101],u1_data_out_2[101],u1_data_out_3[101],partial_product_low0[101],partial_product_low1[101],96'b0};
assign col_out_102 = {u0_col_out_102,u1_data_out_0[102],u1_data_out_1[102],u1_data_out_2[102],u1_data_out_3[102],partial_product_low0[102],partial_product_low1[102],96'b0};
assign col_out_103 = {u0_col_out_103,u1_data_out_0[103],u1_data_out_1[103],u1_data_out_2[103],u1_data_out_3[103],partial_product_low0[103],partial_product_low1[103],96'b0};
assign col_out_104 = {u0_col_out_104,u1_data_out_0[104],u1_data_out_1[104],u1_data_out_2[104],u1_data_out_3[104],partial_product_low0[104],partial_product_low1[104],96'b0};
assign col_out_105 = {u0_col_out_105,u1_data_out_0[105],u1_data_out_1[105],u1_data_out_2[105],u1_data_out_3[105],partial_product_low0[105],partial_product_low1[105],96'b0};
assign col_out_106 = {u0_col_out_106,u1_data_out_0[106],u1_data_out_1[106],u1_data_out_2[106],u1_data_out_3[106],partial_product_low0[106],partial_product_low1[106],96'b0};
assign col_out_107 = {u0_col_out_107,u1_data_out_0[107],u1_data_out_1[107],u1_data_out_2[107],u1_data_out_3[107],partial_product_low0[107],partial_product_low1[107],96'b0};
assign col_out_108 = {u0_col_out_108,u1_data_out_0[108],u1_data_out_1[108],u1_data_out_2[108],u1_data_out_3[108],partial_product_low0[108],partial_product_low1[108],96'b0};
assign col_out_109 = {u0_col_out_109,u1_data_out_0[109],u1_data_out_1[109],u1_data_out_2[109],u1_data_out_3[109],partial_product_low0[109],partial_product_low1[109],96'b0};
assign col_out_110 = {u0_col_out_110,u1_data_out_0[110],u1_data_out_1[110],u1_data_out_2[110],u1_data_out_3[110],partial_product_low0[110],partial_product_low1[110],96'b0};
assign col_out_111 = {u0_col_out_111,u1_data_out_0[111],u1_data_out_1[111],u1_data_out_2[111],u1_data_out_3[111],partial_product_low0[111],partial_product_low1[111],96'b0};
assign col_out_112 = {u0_col_out_112,u1_data_out_0[112],u1_data_out_1[112],u1_data_out_2[112],u1_data_out_3[112],partial_product_low0[112],partial_product_low1[112],96'b0};
assign col_out_113 = {u0_col_out_113,u1_data_out_0[113],u1_data_out_1[113],u1_data_out_2[113],u1_data_out_3[113],partial_product_low0[113],partial_product_low1[113],96'b0};
assign col_out_114 = {u0_col_out_114,u1_data_out_0[114],u1_data_out_1[114],u1_data_out_2[114],u1_data_out_3[114],partial_product_low0[114],partial_product_low1[114],96'b0};
assign col_out_115 = {u0_col_out_115,u1_data_out_0[115],u1_data_out_1[115],u1_data_out_2[115],u1_data_out_3[115],partial_product_low0[115],partial_product_low1[115],96'b0};
assign col_out_116 = {u0_col_out_116,u1_data_out_0[116],u1_data_out_1[116],u1_data_out_2[116],u1_data_out_3[116],partial_product_low0[116],partial_product_low1[116],96'b0};
assign col_out_117 = {u0_col_out_117,u1_data_out_0[117],u1_data_out_1[117],u1_data_out_2[117],u1_data_out_3[117],partial_product_low0[117],partial_product_low1[117],96'b0};
assign col_out_118 = {u0_col_out_118,u1_data_out_0[118],u1_data_out_1[118],u1_data_out_2[118],u1_data_out_3[118],partial_product_low0[118],partial_product_low1[118],96'b0};
assign col_out_119 = {u0_col_out_119,u1_data_out_0[119],u1_data_out_1[119],u1_data_out_2[119],u1_data_out_3[119],partial_product_low0[119],partial_product_low1[119],96'b0};
assign col_out_120 = {u0_col_out_120,u1_data_out_0[120],u1_data_out_1[120],u1_data_out_2[120],u1_data_out_3[120],partial_product_low0[120],partial_product_low1[120],96'b0};
assign col_out_121 = {u0_col_out_121,u1_data_out_0[121],u1_data_out_1[121],u1_data_out_2[121],u1_data_out_3[121],partial_product_low0[121],partial_product_low1[121],96'b0};
assign col_out_122 = {u0_col_out_122,u1_data_out_0[122],u1_data_out_1[122],u1_data_out_2[122],u1_data_out_3[122],partial_product_low0[122],partial_product_low1[122],96'b0};
assign col_out_123 = {u0_col_out_123,u1_data_out_0[123],u1_data_out_1[123],u1_data_out_2[123],u1_data_out_3[123],partial_product_low0[123],partial_product_low1[123],96'b0};
assign col_out_124 = {u0_col_out_124,u1_data_out_0[124],u1_data_out_1[124],u1_data_out_2[124],u1_data_out_3[124],partial_product_low0[124],partial_product_low1[124],96'b0};
assign col_out_125 = {u0_col_out_125,u1_data_out_0[125],u1_data_out_1[125],u1_data_out_2[125],u1_data_out_3[125],partial_product_low0[125],partial_product_low1[125],96'b0};
assign col_out_126 = {u0_col_out_126,u1_data_out_0[126],u1_data_out_1[126],u1_data_out_2[126],u1_data_out_3[126],partial_product_low0[126],partial_product_low1[126],96'b0};
assign col_out_127 = {u0_col_out_127,u1_data_out_0[127],u1_data_out_1[127],u1_data_out_2[127],u1_data_out_3[127],partial_product_low0[127],partial_product_low1[127],96'b0};
assign col_out_128 = {u0_col_out_128,u1_data_out_0[128],u1_data_out_1[128],u1_data_out_2[128],u1_data_out_3[128],partial_product_low0[128],partial_product_low1[128],96'b0};
assign col_out_129 = {u0_col_out_129,u1_data_out_0[129],u1_data_out_1[129],u1_data_out_2[129],u1_data_out_3[129],partial_product_low0[129],partial_product_low1[129],96'b0};
assign col_out_130 = {u0_col_out_130,u1_data_out_0[130],u1_data_out_1[130],u1_data_out_2[130],u1_data_out_3[130],partial_product_low0[130],partial_product_low1[130],96'b0};
assign col_out_131 = {u0_col_out_131,u1_data_out_0[131],u1_data_out_1[131],u1_data_out_2[131],u1_data_out_3[131],partial_product_low0[131],partial_product_low1[131],96'b0};
assign col_out_132 = {u0_col_out_132,u1_data_out_0[132],u1_data_out_1[132],u1_data_out_2[132],u1_data_out_3[132],partial_product_low0[132],partial_product_low1[132],96'b0};
assign col_out_133 = {u0_col_out_133,u1_data_out_0[133],u1_data_out_1[133],u1_data_out_2[133],u1_data_out_3[133],partial_product_low0[133],partial_product_low1[133],96'b0};
assign col_out_134 = {u0_col_out_134,u1_data_out_0[134],u1_data_out_1[134],u1_data_out_2[134],u1_data_out_3[134],partial_product_low0[134],partial_product_low1[134],96'b0};
assign col_out_135 = {u0_col_out_135,u1_data_out_0[135],u1_data_out_1[135],u1_data_out_2[135],u1_data_out_3[135],partial_product_low0[135],partial_product_low1[135],96'b0};
assign col_out_136 = {u0_col_out_136,u1_data_out_0[136],u1_data_out_1[136],u1_data_out_2[136],u1_data_out_3[136],partial_product_low0[136],partial_product_low1[136],96'b0};
assign col_out_137 = {u0_col_out_137,u1_data_out_0[137],u1_data_out_1[137],u1_data_out_2[137],u1_data_out_3[137],partial_product_low0[137],partial_product_low1[137],96'b0};
assign col_out_138 = {u0_col_out_138,u1_data_out_0[138],u1_data_out_1[138],u1_data_out_2[138],u1_data_out_3[138],partial_product_low0[138],partial_product_low1[138],96'b0};
assign col_out_139 = {u0_col_out_139,u1_data_out_0[139],u1_data_out_1[139],u1_data_out_2[139],u1_data_out_3[139],partial_product_low0[139],partial_product_low1[139],96'b0};
assign col_out_140 = {u0_col_out_140,u1_data_out_0[140],u1_data_out_1[140],u1_data_out_2[140],u1_data_out_3[140],partial_product_low0[140],partial_product_low1[140],96'b0};
assign col_out_141 = {u0_col_out_141,u1_data_out_0[141],u1_data_out_1[141],u1_data_out_2[141],u1_data_out_3[141],partial_product_low0[141],partial_product_low1[141],96'b0};
assign col_out_142 = {u0_col_out_142,u1_data_out_0[142],u1_data_out_1[142],u1_data_out_2[142],u1_data_out_3[142],partial_product_low0[142],partial_product_low1[142],96'b0};
assign col_out_143 = {u0_col_out_143,u1_data_out_0[143],u1_data_out_1[143],u1_data_out_2[143],u1_data_out_3[143],partial_product_low0[143],partial_product_low1[143],96'b0};
assign col_out_144 = {u0_col_out_144,u1_data_out_0[144],u1_data_out_1[144],u1_data_out_2[144],u1_data_out_3[144],partial_product_low0[144],partial_product_low1[144],96'b0};
assign col_out_145 = {u0_col_out_145,u1_data_out_0[145],u1_data_out_1[145],u1_data_out_2[145],u1_data_out_3[145],partial_product_low0[145],partial_product_low1[145],96'b0};
assign col_out_146 = {u0_col_out_146,u1_data_out_0[146],u1_data_out_1[146],u1_data_out_2[146],u1_data_out_3[146],partial_product_low0[146],partial_product_low1[146],96'b0};
assign col_out_147 = {u0_col_out_147,u1_data_out_0[147],u1_data_out_1[147],u1_data_out_2[147],u1_data_out_3[147],partial_product_low0[147],partial_product_low1[147],96'b0};
assign col_out_148 = {u0_col_out_148,u1_data_out_0[148],u1_data_out_1[148],u1_data_out_2[148],u1_data_out_3[148],partial_product_low0[148],partial_product_low1[148],96'b0};
assign col_out_149 = {u0_col_out_149,u1_data_out_0[149],u1_data_out_1[149],u1_data_out_2[149],u1_data_out_3[149],partial_product_low0[149],partial_product_low1[149],96'b0};
assign col_out_150 = {u0_col_out_150,u1_data_out_0[150],u1_data_out_1[150],u1_data_out_2[150],u1_data_out_3[150],partial_product_low0[150],partial_product_low1[150],96'b0};
assign col_out_151 = {u0_col_out_151,u1_data_out_0[151],u1_data_out_1[151],u1_data_out_2[151],u1_data_out_3[151],partial_product_low0[151],partial_product_low1[151],96'b0};
assign col_out_152 = {u0_col_out_152,u1_data_out_0[152],u1_data_out_1[152],u1_data_out_2[152],u1_data_out_3[152],partial_product_low0[152],partial_product_low1[152],96'b0};
assign col_out_153 = {u0_col_out_153,u1_data_out_0[153],u1_data_out_1[153],u1_data_out_2[153],u1_data_out_3[153],partial_product_low0[153],partial_product_low1[153],96'b0};
assign col_out_154 = {u0_col_out_154,u1_data_out_0[154],u1_data_out_1[154],u1_data_out_2[154],u1_data_out_3[154],partial_product_low0[154],partial_product_low1[154],96'b0};
assign col_out_155 = {u0_col_out_155,u1_data_out_0[155],u1_data_out_1[155],u1_data_out_2[155],u1_data_out_3[155],partial_product_low0[155],partial_product_low1[155],96'b0};
assign col_out_156 = {u0_col_out_156,u1_data_out_0[156],u1_data_out_1[156],u1_data_out_2[156],u1_data_out_3[156],partial_product_low0[156],partial_product_low1[156],96'b0};
assign col_out_157 = {u0_col_out_157,u1_data_out_0[157],u1_data_out_1[157],u1_data_out_2[157],u1_data_out_3[157],partial_product_low0[157],partial_product_low1[157],96'b0};
assign col_out_158 = {u0_col_out_158,u1_data_out_0[158],u1_data_out_1[158],u1_data_out_2[158],u1_data_out_3[158],partial_product_low0[158],partial_product_low1[158],96'b0};
assign col_out_159 = {u0_col_out_159,u1_data_out_0[159],u1_data_out_1[159],u1_data_out_2[159],u1_data_out_3[159],partial_product_low0[159],partial_product_low1[159],96'b0};
assign col_out_160 = {u0_col_out_160,u1_data_out_0[160],u1_data_out_1[160],u1_data_out_2[160],u1_data_out_3[160],partial_product_low0[160],partial_product_low1[160],96'b0};
assign col_out_161 = {u0_col_out_161,u1_data_out_0[161],u1_data_out_1[161],u1_data_out_2[161],u1_data_out_3[161],partial_product_low0[161],partial_product_low1[161],96'b0};
assign col_out_162 = {u0_col_out_162,u1_data_out_0[162],u1_data_out_1[162],u1_data_out_2[162],u1_data_out_3[162],partial_product_low0[162],partial_product_low1[162],96'b0};
assign col_out_163 = {u0_col_out_163,u1_data_out_0[163],u1_data_out_1[163],u1_data_out_2[163],u1_data_out_3[163],partial_product_low0[163],partial_product_low1[163],96'b0};
assign col_out_164 = {u0_col_out_164,u1_data_out_0[164],u1_data_out_1[164],u1_data_out_2[164],u1_data_out_3[164],partial_product_low0[164],partial_product_low1[164],96'b0};
assign col_out_165 = {u0_col_out_165,u1_data_out_0[165],u1_data_out_1[165],u1_data_out_2[165],u1_data_out_3[165],partial_product_low0[165],partial_product_low1[165],96'b0};
assign col_out_166 = {u0_col_out_166,u1_data_out_0[166],u1_data_out_1[166],u1_data_out_2[166],u1_data_out_3[166],partial_product_low0[166],partial_product_low1[166],96'b0};
assign col_out_167 = {u0_col_out_167,u1_data_out_0[167],u1_data_out_1[167],u1_data_out_2[167],u1_data_out_3[167],partial_product_low0[167],partial_product_low1[167],96'b0};
assign col_out_168 = {u0_col_out_168,u1_data_out_0[168],u1_data_out_1[168],u1_data_out_2[168],u1_data_out_3[168],partial_product_low0[168],partial_product_low1[168],96'b0};
assign col_out_169 = {u0_col_out_169,u1_data_out_0[169],u1_data_out_1[169],u1_data_out_2[169],u1_data_out_3[169],partial_product_low0[169],partial_product_low1[169],96'b0};
assign col_out_170 = {u0_col_out_170,u1_data_out_0[170],u1_data_out_1[170],u1_data_out_2[170],u1_data_out_3[170],partial_product_low0[170],partial_product_low1[170],96'b0};
assign col_out_171 = {u0_col_out_171,u1_data_out_0[171],u1_data_out_1[171],u1_data_out_2[171],u1_data_out_3[171],partial_product_low0[171],partial_product_low1[171],96'b0};
assign col_out_172 = {u0_col_out_172,u1_data_out_0[172],u1_data_out_1[172],u1_data_out_2[172],u1_data_out_3[172],partial_product_low0[172],partial_product_low1[172],96'b0};
assign col_out_173 = {u0_col_out_173,u1_data_out_0[173],u1_data_out_1[173],u1_data_out_2[173],u1_data_out_3[173],partial_product_low0[173],partial_product_low1[173],96'b0};
assign col_out_174 = {u0_col_out_174,u1_data_out_0[174],u1_data_out_1[174],u1_data_out_2[174],u1_data_out_3[174],partial_product_low0[174],partial_product_low1[174],96'b0};
assign col_out_175 = {u0_col_out_175,u1_data_out_0[175],u1_data_out_1[175],u1_data_out_2[175],u1_data_out_3[175],partial_product_low0[175],partial_product_low1[175],96'b0};
assign col_out_176 = {u0_col_out_176,u1_data_out_0[176],u1_data_out_1[176],u1_data_out_2[176],u1_data_out_3[176],partial_product_low0[176],partial_product_low1[176],96'b0};
assign col_out_177 = {u0_col_out_177,u1_data_out_0[177],u1_data_out_1[177],u1_data_out_2[177],u1_data_out_3[177],partial_product_low0[177],partial_product_low1[177],96'b0};
assign col_out_178 = {u0_col_out_178,u1_data_out_0[178],u1_data_out_1[178],u1_data_out_2[178],u1_data_out_3[178],partial_product_low0[178],partial_product_low1[178],96'b0};
assign col_out_179 = {u0_col_out_179,u1_data_out_0[179],u1_data_out_1[179],u1_data_out_2[179],u1_data_out_3[179],partial_product_low0[179],partial_product_low1[179],96'b0};
assign col_out_180 = {u0_col_out_180,u1_data_out_0[180],u1_data_out_1[180],u1_data_out_2[180],u1_data_out_3[180],partial_product_low0[180],partial_product_low1[180],96'b0};
assign col_out_181 = {u0_col_out_181,u1_data_out_0[181],u1_data_out_1[181],u1_data_out_2[181],u1_data_out_3[181],partial_product_low0[181],partial_product_low1[181],96'b0};
assign col_out_182 = {u0_col_out_182,u1_data_out_0[182],u1_data_out_1[182],u1_data_out_2[182],u1_data_out_3[182],partial_product_low0[182],partial_product_low1[182],96'b0};
assign col_out_183 = {u0_col_out_183,u1_data_out_0[183],u1_data_out_1[183],u1_data_out_2[183],u1_data_out_3[183],partial_product_low0[183],partial_product_low1[183],96'b0};
assign col_out_184 = {u0_col_out_184,u1_data_out_0[184],u1_data_out_1[184],u1_data_out_2[184],u1_data_out_3[184],partial_product_low0[184],partial_product_low1[184],96'b0};
assign col_out_185 = {u0_col_out_185,u1_data_out_0[185],u1_data_out_1[185],u1_data_out_2[185],u1_data_out_3[185],partial_product_low0[185],partial_product_low1[185],96'b0};
assign col_out_186 = {u0_col_out_186,u1_data_out_0[186],u1_data_out_1[186],u1_data_out_2[186],u1_data_out_3[186],partial_product_low0[186],partial_product_low1[186],96'b0};
assign col_out_187 = {u0_col_out_187,u1_data_out_0[187],u1_data_out_1[187],u1_data_out_2[187],u1_data_out_3[187],partial_product_low0[187],partial_product_low1[187],96'b0};
assign col_out_188 = {u0_col_out_188,u1_data_out_0[188],u1_data_out_1[188],u1_data_out_2[188],u1_data_out_3[188],partial_product_low0[188],partial_product_low1[188],96'b0};
assign col_out_189 = {u0_col_out_189,u1_data_out_0[189],u1_data_out_1[189],u1_data_out_2[189],u1_data_out_3[189],partial_product_low0[189],partial_product_low1[189],96'b0};
assign col_out_190 = {u0_col_out_190,u1_data_out_0[190],u1_data_out_1[190],u1_data_out_2[190],u1_data_out_3[190],partial_product_low0[190],partial_product_low1[190],96'b0};
assign col_out_191 = {u0_col_out_191,u1_data_out_0[191],u1_data_out_1[191],u1_data_out_2[191],u1_data_out_3[191],partial_product_low0[191],partial_product_low1[191],96'b0};
assign col_out_192 = {u0_col_out_192,u1_data_out_0[192],u1_data_out_1[192],u1_data_out_2[192],u1_data_out_3[192],partial_product_low0[192],partial_product_low1[192],96'b0};
assign col_out_193 = {u0_col_out_193,u1_data_out_0[193],u1_data_out_1[193],u1_data_out_2[193],u1_data_out_3[193],partial_product_low0[193],partial_product_low1[193],96'b0};
assign col_out_194 = {u0_col_out_194,u1_data_out_0[194],u1_data_out_1[194],u1_data_out_2[194],u1_data_out_3[194],partial_product_low0[194],partial_product_low1[194],96'b0};
assign col_out_195 = {u0_col_out_195,u1_data_out_0[195],u1_data_out_1[195],u1_data_out_2[195],u1_data_out_3[195],partial_product_low0[195],partial_product_low1[195],96'b0};
assign col_out_196 = {u0_col_out_196,u1_data_out_0[196],u1_data_out_1[196],u1_data_out_2[196],u1_data_out_3[196],partial_product_low0[196],partial_product_low1[196],96'b0};
assign col_out_197 = {u0_col_out_197,u1_data_out_0[197],u1_data_out_1[197],u1_data_out_2[197],u1_data_out_3[197],partial_product_low0[197],partial_product_low1[197],96'b0};
assign col_out_198 = {u0_col_out_198,u1_data_out_0[198],u1_data_out_1[198],u1_data_out_2[198],u1_data_out_3[198],partial_product_low0[198],partial_product_low1[198],96'b0};
assign col_out_199 = {u0_col_out_199,u1_data_out_0[199],u1_data_out_1[199],u1_data_out_2[199],u1_data_out_3[199],partial_product_low0[199],partial_product_low1[199],96'b0};
assign col_out_200 = {u0_col_out_200,u1_data_out_0[200],u1_data_out_1[200],u1_data_out_2[200],u1_data_out_3[200],partial_product_low0[200],partial_product_low1[200],96'b0};
assign col_out_201 = {u0_col_out_201,u1_data_out_0[201],u1_data_out_1[201],u1_data_out_2[201],u1_data_out_3[201],partial_product_low0[201],partial_product_low1[201],96'b0};
assign col_out_202 = {u0_col_out_202,u1_data_out_0[202],u1_data_out_1[202],u1_data_out_2[202],u1_data_out_3[202],partial_product_low0[202],partial_product_low1[202],96'b0};
assign col_out_203 = {u0_col_out_203,u1_data_out_0[203],u1_data_out_1[203],u1_data_out_2[203],u1_data_out_3[203],partial_product_low0[203],partial_product_low1[203],96'b0};
assign col_out_204 = {u0_col_out_204,u1_data_out_0[204],u1_data_out_1[204],u1_data_out_2[204],u1_data_out_3[204],partial_product_low0[204],partial_product_low1[204],96'b0};
assign col_out_205 = {u0_col_out_205,u1_data_out_0[205],u1_data_out_1[205],u1_data_out_2[205],u1_data_out_3[205],partial_product_low0[205],partial_product_low1[205],96'b0};
assign col_out_206 = {u0_col_out_206,u1_data_out_0[206],u1_data_out_1[206],u1_data_out_2[206],u1_data_out_3[206],partial_product_low0[206],partial_product_low1[206],96'b0};
assign col_out_207 = {u0_col_out_207,u1_data_out_0[207],u1_data_out_1[207],u1_data_out_2[207],u1_data_out_3[207],partial_product_low0[207],partial_product_low1[207],96'b0};
assign col_out_208 = {u0_col_out_208,u1_data_out_0[208],u1_data_out_1[208],u1_data_out_2[208],u1_data_out_3[208],partial_product_low0[208],partial_product_low1[208],96'b0};
assign col_out_209 = {u0_col_out_209,u1_data_out_0[209],u1_data_out_1[209],u1_data_out_2[209],u1_data_out_3[209],partial_product_low0[209],partial_product_low1[209],96'b0};
assign col_out_210 = {u0_col_out_210,u1_data_out_0[210],u1_data_out_1[210],u1_data_out_2[210],u1_data_out_3[210],partial_product_low0[210],partial_product_low1[210],96'b0};
assign col_out_211 = {u0_col_out_211,u1_data_out_0[211],u1_data_out_1[211],u1_data_out_2[211],u1_data_out_3[211],partial_product_low0[211],partial_product_low1[211],96'b0};
assign col_out_212 = {u0_col_out_212,u1_data_out_0[212],u1_data_out_1[212],u1_data_out_2[212],u1_data_out_3[212],partial_product_low0[212],partial_product_low1[212],96'b0};
assign col_out_213 = {u0_col_out_213,u1_data_out_0[213],u1_data_out_1[213],u1_data_out_2[213],u1_data_out_3[213],partial_product_low0[213],partial_product_low1[213],96'b0};
assign col_out_214 = {u0_col_out_214,u1_data_out_0[214],u1_data_out_1[214],u1_data_out_2[214],u1_data_out_3[214],partial_product_low0[214],partial_product_low1[214],96'b0};
assign col_out_215 = {u0_col_out_215,u1_data_out_0[215],u1_data_out_1[215],u1_data_out_2[215],u1_data_out_3[215],partial_product_low0[215],partial_product_low1[215],96'b0};
assign col_out_216 = {u0_col_out_216,u1_data_out_0[216],u1_data_out_1[216],u1_data_out_2[216],u1_data_out_3[216],partial_product_low0[216],partial_product_low1[216],96'b0};
assign col_out_217 = {u0_col_out_217,u1_data_out_0[217],u1_data_out_1[217],u1_data_out_2[217],u1_data_out_3[217],partial_product_low0[217],partial_product_low1[217],96'b0};
assign col_out_218 = {u0_col_out_218,u1_data_out_0[218],u1_data_out_1[218],u1_data_out_2[218],u1_data_out_3[218],partial_product_low0[218],partial_product_low1[218],96'b0};
assign col_out_219 = {u0_col_out_219,u1_data_out_0[219],u1_data_out_1[219],u1_data_out_2[219],u1_data_out_3[219],partial_product_low0[219],partial_product_low1[219],96'b0};
assign col_out_220 = {u0_col_out_220,u1_data_out_0[220],u1_data_out_1[220],u1_data_out_2[220],u1_data_out_3[220],partial_product_low0[220],partial_product_low1[220],96'b0};
assign col_out_221 = {u0_col_out_221,u1_data_out_0[221],u1_data_out_1[221],u1_data_out_2[221],u1_data_out_3[221],partial_product_low0[221],partial_product_low1[221],96'b0};
assign col_out_222 = {u0_col_out_222,u1_data_out_0[222],u1_data_out_1[222],u1_data_out_2[222],u1_data_out_3[222],partial_product_low0[222],partial_product_low1[222],96'b0};
assign col_out_223 = {u0_col_out_223,u1_data_out_0[223],u1_data_out_1[223],u1_data_out_2[223],u1_data_out_3[223],partial_product_low0[223],partial_product_low1[223],96'b0};
assign col_out_224 = {u0_col_out_224,u1_data_out_0[224],u1_data_out_1[224],u1_data_out_2[224],u1_data_out_3[224],partial_product_low0[224],partial_product_low1[224],96'b0};
assign col_out_225 = {u0_col_out_225,u1_data_out_0[225],u1_data_out_1[225],u1_data_out_2[225],u1_data_out_3[225],partial_product_low0[225],partial_product_low1[225],96'b0};
assign col_out_226 = {u0_col_out_226,u1_data_out_0[226],u1_data_out_1[226],u1_data_out_2[226],u1_data_out_3[226],partial_product_low0[226],partial_product_low1[226],96'b0};
assign col_out_227 = {u0_col_out_227,u1_data_out_0[227],u1_data_out_1[227],u1_data_out_2[227],u1_data_out_3[227],partial_product_low0[227],partial_product_low1[227],96'b0};
assign col_out_228 = {u0_col_out_228,u1_data_out_0[228],u1_data_out_1[228],u1_data_out_2[228],u1_data_out_3[228],partial_product_low0[228],partial_product_low1[228],96'b0};
assign col_out_229 = {u0_col_out_229,u1_data_out_0[229],u1_data_out_1[229],u1_data_out_2[229],u1_data_out_3[229],partial_product_low0[229],partial_product_low1[229],96'b0};
assign col_out_230 = {u0_col_out_230,u1_data_out_0[230],u1_data_out_1[230],u1_data_out_2[230],u1_data_out_3[230],partial_product_low0[230],partial_product_low1[230],96'b0};
assign col_out_231 = {u0_col_out_231,u1_data_out_0[231],u1_data_out_1[231],u1_data_out_2[231],u1_data_out_3[231],partial_product_low0[231],partial_product_low1[231],96'b0};
assign col_out_232 = {u0_col_out_232,u1_data_out_0[232],u1_data_out_1[232],u1_data_out_2[232],u1_data_out_3[232],partial_product_low0[232],partial_product_low1[232],96'b0};
assign col_out_233 = {u0_col_out_233,u1_data_out_0[233],u1_data_out_1[233],u1_data_out_2[233],u1_data_out_3[233],partial_product_low0[233],partial_product_low1[233],96'b0};
assign col_out_234 = {u0_col_out_234,u1_data_out_0[234],u1_data_out_1[234],u1_data_out_2[234],u1_data_out_3[234],partial_product_low0[234],partial_product_low1[234],96'b0};
assign col_out_235 = {u0_col_out_235,u1_data_out_0[235],u1_data_out_1[235],u1_data_out_2[235],u1_data_out_3[235],partial_product_low0[235],partial_product_low1[235],96'b0};
assign col_out_236 = {u0_col_out_236,u1_data_out_0[236],u1_data_out_1[236],u1_data_out_2[236],u1_data_out_3[236],partial_product_low0[236],partial_product_low1[236],96'b0};
assign col_out_237 = {u0_col_out_237,u1_data_out_0[237],u1_data_out_1[237],u1_data_out_2[237],u1_data_out_3[237],partial_product_low0[237],partial_product_low1[237],96'b0};
assign col_out_238 = {u0_col_out_238,u1_data_out_0[238],u1_data_out_1[238],u1_data_out_2[238],u1_data_out_3[238],partial_product_low0[238],partial_product_low1[238],96'b0};
assign col_out_239 = {u0_col_out_239,u1_data_out_0[239],u1_data_out_1[239],u1_data_out_2[239],u1_data_out_3[239],partial_product_low0[239],partial_product_low1[239],96'b0};
assign col_out_240 = {u0_col_out_240,u1_data_out_0[240],u1_data_out_1[240],u1_data_out_2[240],u1_data_out_3[240],partial_product_low0[240],partial_product_low1[240],96'b0};
assign col_out_241 = {u0_col_out_241,u1_data_out_0[241],u1_data_out_1[241],u1_data_out_2[241],u1_data_out_3[241],partial_product_low0[241],partial_product_low1[241],96'b0};
assign col_out_242 = {u0_col_out_242,u1_data_out_0[242],u1_data_out_1[242],u1_data_out_2[242],u1_data_out_3[242],partial_product_low0[242],partial_product_low1[242],96'b0};
assign col_out_243 = {u0_col_out_243,u1_data_out_0[243],u1_data_out_1[243],u1_data_out_2[243],u1_data_out_3[243],partial_product_low0[243],partial_product_low1[243],96'b0};
assign col_out_244 = {u0_col_out_244,u1_data_out_0[244],u1_data_out_1[244],u1_data_out_2[244],u1_data_out_3[244],partial_product_low0[244],partial_product_low1[244],96'b0};
assign col_out_245 = {u0_col_out_245,u1_data_out_0[245],u1_data_out_1[245],u1_data_out_2[245],u1_data_out_3[245],partial_product_low0[245],partial_product_low1[245],96'b0};
assign col_out_246 = {u0_col_out_246,u1_data_out_0[246],u1_data_out_1[246],u1_data_out_2[246],u1_data_out_3[246],partial_product_low0[246],partial_product_low1[246],96'b0};
assign col_out_247 = {u0_col_out_247,u1_data_out_0[247],u1_data_out_1[247],u1_data_out_2[247],u1_data_out_3[247],partial_product_low0[247],partial_product_low1[247],96'b0};
assign col_out_248 = {u0_col_out_248,u1_data_out_0[248],u1_data_out_1[248],u1_data_out_2[248],u1_data_out_3[248],partial_product_low0[248],partial_product_low1[248],96'b0};
assign col_out_249 = {u0_col_out_249,u1_data_out_0[249],u1_data_out_1[249],u1_data_out_2[249],u1_data_out_3[249],partial_product_low0[249],partial_product_low1[249],96'b0};
assign col_out_250 = {u0_col_out_250,u1_data_out_0[250],u1_data_out_1[250],u1_data_out_2[250],u1_data_out_3[250],partial_product_low0[250],partial_product_low1[250],96'b0};
assign col_out_251 = {u0_col_out_251,u1_data_out_0[251],u1_data_out_1[251],u1_data_out_2[251],u1_data_out_3[251],partial_product_low0[251],partial_product_low1[251],96'b0};
assign col_out_252 = {u0_col_out_252,u1_data_out_0[252],u1_data_out_1[252],u1_data_out_2[252],u1_data_out_3[252],partial_product_low0[252],partial_product_low1[252],96'b0};
assign col_out_253 = {u0_col_out_253,u1_data_out_0[253],u1_data_out_1[253],u1_data_out_2[253],u1_data_out_3[253],partial_product_low0[253],partial_product_low1[253],96'b0};
assign col_out_254 = {u0_col_out_254,u1_data_out_0[254],u1_data_out_1[254],u1_data_out_2[254],u1_data_out_3[254],partial_product_low0[254],partial_product_low1[254],96'b0};
assign col_out_255 = {u0_col_out_255,u1_data_out_0[255],u1_data_out_1[255],u1_data_out_2[255],u1_data_out_3[255],partial_product_low0[255],partial_product_low1[255],96'b0};
assign col_out_256 = {u0_col_out_256,u1_data_out_0[256],u1_data_out_1[256],u1_data_out_2[256],u1_data_out_3[256],partial_product_low0[256],partial_product_low1[256],96'b0};
assign col_out_257 = {u0_col_out_257,u1_data_out_0[257],u1_data_out_1[257],u1_data_out_2[257],u1_data_out_3[257],partial_product_low0[257],partial_product_low1[257],96'b0};
assign col_out_258 = {u0_col_out_258,u1_data_out_0[258],u1_data_out_1[258],u1_data_out_2[258],u1_data_out_3[258],partial_product_low0[258],partial_product_low1[258],96'b0};
assign col_out_259 = {u0_col_out_259,u1_data_out_0[259],u1_data_out_1[259],u1_data_out_2[259],u1_data_out_3[259],partial_product_low0[259],partial_product_low1[259],96'b0};
assign col_out_260 = {u0_col_out_260,u1_data_out_0[260],u1_data_out_1[260],u1_data_out_2[260],u1_data_out_3[260],partial_product_low0[260],partial_product_low1[260],96'b0};
assign col_out_261 = {u0_col_out_261,u1_data_out_0[261],u1_data_out_1[261],u1_data_out_2[261],u1_data_out_3[261],partial_product_low0[261],partial_product_low1[261],96'b0};
assign col_out_262 = {u0_col_out_262,u1_data_out_0[262],u1_data_out_1[262],u1_data_out_2[262],u1_data_out_3[262],partial_product_low0[262],partial_product_low1[262],96'b0};
assign col_out_263 = {u0_col_out_263,u1_data_out_0[263],u1_data_out_1[263],u1_data_out_2[263],u1_data_out_3[263],partial_product_low0[263],partial_product_low1[263],96'b0};
assign col_out_264 = {u0_col_out_264,u1_data_out_0[264],u1_data_out_1[264],u1_data_out_2[264],u1_data_out_3[264],partial_product_low0[264],partial_product_low1[264],96'b0};
assign col_out_265 = {u0_col_out_265,u1_data_out_0[265],u1_data_out_1[265],u1_data_out_2[265],u1_data_out_3[265],partial_product_low0[265],partial_product_low1[265],96'b0};
assign col_out_266 = {u0_col_out_266,u1_data_out_0[266],u1_data_out_1[266],u1_data_out_2[266],u1_data_out_3[266],partial_product_low0[266],partial_product_low1[266],96'b0};
assign col_out_267 = {u0_col_out_267,u1_data_out_0[267],u1_data_out_1[267],u1_data_out_2[267],u1_data_out_3[267],partial_product_low0[267],partial_product_low1[267],96'b0};
assign col_out_268 = {u0_col_out_268,u1_data_out_0[268],u1_data_out_1[268],u1_data_out_2[268],u1_data_out_3[268],partial_product_low0[268],partial_product_low1[268],96'b0};
assign col_out_269 = {u0_col_out_269,u1_data_out_0[269],u1_data_out_1[269],u1_data_out_2[269],u1_data_out_3[269],partial_product_low0[269],partial_product_low1[269],96'b0};
assign col_out_270 = {u0_col_out_270,u1_data_out_0[270],u1_data_out_1[270],u1_data_out_2[270],u1_data_out_3[270],partial_product_low0[270],partial_product_low1[270],96'b0};
assign col_out_271 = {u0_col_out_271,u1_data_out_0[271],u1_data_out_1[271],u1_data_out_2[271],u1_data_out_3[271],partial_product_low0[271],partial_product_low1[271],96'b0};
assign col_out_272 = {u0_col_out_272,u1_data_out_0[272],u1_data_out_1[272],u1_data_out_2[272],u1_data_out_3[272],partial_product_low0[272],partial_product_low1[272],96'b0};
assign col_out_273 = {u0_col_out_273,u1_data_out_0[273],u1_data_out_1[273],u1_data_out_2[273],u1_data_out_3[273],partial_product_low0[273],partial_product_low1[273],96'b0};
assign col_out_274 = {u0_col_out_274,u1_data_out_0[274],u1_data_out_1[274],u1_data_out_2[274],u1_data_out_3[274],partial_product_low0[274],partial_product_low1[274],96'b0};
assign col_out_275 = {u0_col_out_275,u1_data_out_0[275],u1_data_out_1[275],u1_data_out_2[275],u1_data_out_3[275],partial_product_low0[275],partial_product_low1[275],96'b0};
assign col_out_276 = {u0_col_out_276,u1_data_out_0[276],u1_data_out_1[276],u1_data_out_2[276],u1_data_out_3[276],partial_product_low0[276],partial_product_low1[276],96'b0};
assign col_out_277 = {u0_col_out_277,u1_data_out_0[277],u1_data_out_1[277],u1_data_out_2[277],u1_data_out_3[277],partial_product_low0[277],partial_product_low1[277],96'b0};
assign col_out_278 = {u0_col_out_278,u1_data_out_0[278],u1_data_out_1[278],u1_data_out_2[278],u1_data_out_3[278],partial_product_low0[278],partial_product_low1[278],96'b0};
assign col_out_279 = {u0_col_out_279,u1_data_out_0[279],u1_data_out_1[279],u1_data_out_2[279],u1_data_out_3[279],partial_product_low0[279],partial_product_low1[279],96'b0};
assign col_out_280 = {u0_col_out_280,u1_data_out_0[280],u1_data_out_1[280],u1_data_out_2[280],u1_data_out_3[280],partial_product_low0[280],partial_product_low1[280],96'b0};
assign col_out_281 = {u0_col_out_281,u1_data_out_0[281],u1_data_out_1[281],u1_data_out_2[281],u1_data_out_3[281],partial_product_low0[281],partial_product_low1[281],96'b0};
assign col_out_282 = {u0_col_out_282,u1_data_out_0[282],u1_data_out_1[282],u1_data_out_2[282],u1_data_out_3[282],partial_product_low0[282],partial_product_low1[282],96'b0};
assign col_out_283 = {u0_col_out_283,u1_data_out_0[283],u1_data_out_1[283],u1_data_out_2[283],u1_data_out_3[283],partial_product_low0[283],partial_product_low1[283],96'b0};
assign col_out_284 = {u0_col_out_284,u1_data_out_0[284],u1_data_out_1[284],u1_data_out_2[284],u1_data_out_3[284],partial_product_low0[284],partial_product_low1[284],96'b0};
assign col_out_285 = {u0_col_out_285,u1_data_out_0[285],u1_data_out_1[285],u1_data_out_2[285],u1_data_out_3[285],partial_product_low0[285],partial_product_low1[285],96'b0};
assign col_out_286 = {u0_col_out_286,u1_data_out_0[286],u1_data_out_1[286],u1_data_out_2[286],u1_data_out_3[286],partial_product_low0[286],partial_product_low1[286],96'b0};
assign col_out_287 = {u0_col_out_287,u1_data_out_0[287],u1_data_out_1[287],u1_data_out_2[287],u1_data_out_3[287],partial_product_low0[287],partial_product_low1[287],96'b0};
assign col_out_288 = {u0_col_out_288,u1_data_out_0[288],u1_data_out_1[288],u1_data_out_2[288],u1_data_out_3[288],partial_product_low0[288],partial_product_low1[288],96'b0};
assign col_out_289 = {u0_col_out_289,u1_data_out_0[289],u1_data_out_1[289],u1_data_out_2[289],u1_data_out_3[289],partial_product_low0[289],partial_product_low1[289],96'b0};
assign col_out_290 = {u0_col_out_290,u1_data_out_0[290],u1_data_out_1[290],u1_data_out_2[290],u1_data_out_3[290],partial_product_low0[290],partial_product_low1[290],96'b0};
assign col_out_291 = {u0_col_out_291,u1_data_out_0[291],u1_data_out_1[291],u1_data_out_2[291],u1_data_out_3[291],partial_product_low0[291],partial_product_low1[291],96'b0};
assign col_out_292 = {u0_col_out_292,u1_data_out_0[292],u1_data_out_1[292],u1_data_out_2[292],u1_data_out_3[292],partial_product_low0[292],partial_product_low1[292],96'b0};
assign col_out_293 = {u0_col_out_293,u1_data_out_0[293],u1_data_out_1[293],u1_data_out_2[293],u1_data_out_3[293],partial_product_low0[293],partial_product_low1[293],96'b0};
assign col_out_294 = {u0_col_out_294,u1_data_out_0[294],u1_data_out_1[294],u1_data_out_2[294],u1_data_out_3[294],partial_product_low0[294],partial_product_low1[294],96'b0};
assign col_out_295 = {u0_col_out_295,u1_data_out_0[295],u1_data_out_1[295],u1_data_out_2[295],u1_data_out_3[295],partial_product_low0[295],partial_product_low1[295],96'b0};
assign col_out_296 = {u0_col_out_296,u1_data_out_0[296],u1_data_out_1[296],u1_data_out_2[296],u1_data_out_3[296],partial_product_low0[296],partial_product_low1[296],96'b0};
assign col_out_297 = {u0_col_out_297,u1_data_out_0[297],u1_data_out_1[297],u1_data_out_2[297],u1_data_out_3[297],partial_product_low0[297],partial_product_low1[297],96'b0};
assign col_out_298 = {u0_col_out_298,u1_data_out_0[298],u1_data_out_1[298],u1_data_out_2[298],u1_data_out_3[298],partial_product_low0[298],partial_product_low1[298],96'b0};
assign col_out_299 = {u0_col_out_299,u1_data_out_0[299],u1_data_out_1[299],u1_data_out_2[299],u1_data_out_3[299],partial_product_low0[299],partial_product_low1[299],96'b0};
assign col_out_300 = {u0_col_out_300,u1_data_out_0[300],u1_data_out_1[300],u1_data_out_2[300],u1_data_out_3[300],partial_product_low0[300],partial_product_low1[300],96'b0};
assign col_out_301 = {u0_col_out_301,u1_data_out_0[301],u1_data_out_1[301],u1_data_out_2[301],u1_data_out_3[301],partial_product_low0[301],partial_product_low1[301],96'b0};
assign col_out_302 = {u0_col_out_302,u1_data_out_0[302],u1_data_out_1[302],u1_data_out_2[302],u1_data_out_3[302],partial_product_low0[302],partial_product_low1[302],96'b0};
assign col_out_303 = {u0_col_out_303,u1_data_out_0[303],u1_data_out_1[303],u1_data_out_2[303],u1_data_out_3[303],partial_product_low0[303],partial_product_low1[303],96'b0};
assign col_out_304 = {u0_col_out_304,u1_data_out_0[304],u1_data_out_1[304],u1_data_out_2[304],u1_data_out_3[304],partial_product_low0[304],partial_product_low1[304],96'b0};
assign col_out_305 = {u0_col_out_305,u1_data_out_0[305],u1_data_out_1[305],u1_data_out_2[305],u1_data_out_3[305],partial_product_low0[305],partial_product_low1[305],96'b0};
assign col_out_306 = {u0_col_out_306,u1_data_out_0[306],u1_data_out_1[306],u1_data_out_2[306],u1_data_out_3[306],partial_product_low0[306],partial_product_low1[306],96'b0};
assign col_out_307 = {u0_col_out_307,u1_data_out_0[307],u1_data_out_1[307],u1_data_out_2[307],u1_data_out_3[307],partial_product_low0[307],partial_product_low1[307],96'b0};
assign col_out_308 = {u0_col_out_308,u1_data_out_0[308],u1_data_out_1[308],u1_data_out_2[308],u1_data_out_3[308],partial_product_low0[308],partial_product_low1[308],96'b0};
assign col_out_309 = {u0_col_out_309,u1_data_out_0[309],u1_data_out_1[309],u1_data_out_2[309],u1_data_out_3[309],partial_product_low0[309],partial_product_low1[309],96'b0};
assign col_out_310 = {u0_col_out_310,u1_data_out_0[310],u1_data_out_1[310],u1_data_out_2[310],u1_data_out_3[310],partial_product_low0[310],partial_product_low1[310],96'b0};
assign col_out_311 = {u0_col_out_311,u1_data_out_0[311],u1_data_out_1[311],u1_data_out_2[311],u1_data_out_3[311],partial_product_low0[311],partial_product_low1[311],96'b0};
assign col_out_312 = {u0_col_out_312,u1_data_out_0[312],u1_data_out_1[312],u1_data_out_2[312],u1_data_out_3[312],partial_product_low0[312],partial_product_low1[312],96'b0};
assign col_out_313 = {u0_col_out_313,u1_data_out_0[313],u1_data_out_1[313],u1_data_out_2[313],u1_data_out_3[313],partial_product_low0[313],partial_product_low1[313],96'b0};
assign col_out_314 = {u0_col_out_314,u1_data_out_0[314],u1_data_out_1[314],u1_data_out_2[314],u1_data_out_3[314],partial_product_low0[314],partial_product_low1[314],96'b0};
assign col_out_315 = {u0_col_out_315,u1_data_out_0[315],u1_data_out_1[315],u1_data_out_2[315],u1_data_out_3[315],partial_product_low0[315],partial_product_low1[315],96'b0};
assign col_out_316 = {u0_col_out_316,u1_data_out_0[316],u1_data_out_1[316],u1_data_out_2[316],u1_data_out_3[316],partial_product_low0[316],partial_product_low1[316],96'b0};
assign col_out_317 = {u0_col_out_317,u1_data_out_0[317],u1_data_out_1[317],u1_data_out_2[317],u1_data_out_3[317],partial_product_low0[317],partial_product_low1[317],96'b0};
assign col_out_318 = {u0_col_out_318,u1_data_out_0[318],u1_data_out_1[318],u1_data_out_2[318],u1_data_out_3[318],partial_product_low0[318],partial_product_low1[318],96'b0};
assign col_out_319 = {u0_col_out_319,u1_data_out_0[319],u1_data_out_1[319],u1_data_out_2[319],u1_data_out_3[319],partial_product_low0[319],partial_product_low1[319],96'b0};
assign col_out_320 = {u0_col_out_320,u1_data_out_0[320],u1_data_out_1[320],u1_data_out_2[320],u1_data_out_3[320],partial_product_low0[320],partial_product_low1[320],96'b0};
assign col_out_321 = {u0_col_out_321,u1_data_out_0[321],u1_data_out_1[321],u1_data_out_2[321],u1_data_out_3[321],partial_product_low0[321],partial_product_low1[321],96'b0};
assign col_out_322 = {u0_col_out_322,u1_data_out_0[322],u1_data_out_1[322],u1_data_out_2[322],u1_data_out_3[322],partial_product_low0[322],partial_product_low1[322],96'b0};
assign col_out_323 = {u0_col_out_323,u1_data_out_0[323],u1_data_out_1[323],u1_data_out_2[323],u1_data_out_3[323],partial_product_low0[323],partial_product_low1[323],96'b0};
assign col_out_324 = {u0_col_out_324,u1_data_out_0[324],u1_data_out_1[324],u1_data_out_2[324],u1_data_out_3[324],partial_product_low0[324],partial_product_low1[324],96'b0};
assign col_out_325 = {u0_col_out_325,u1_data_out_0[325],u1_data_out_1[325],u1_data_out_2[325],u1_data_out_3[325],partial_product_low0[325],partial_product_low1[325],96'b0};
assign col_out_326 = {u0_col_out_326,u1_data_out_0[326],u1_data_out_1[326],u1_data_out_2[326],u1_data_out_3[326],partial_product_low0[326],partial_product_low1[326],96'b0};
assign col_out_327 = {u0_col_out_327,u1_data_out_0[327],u1_data_out_1[327],u1_data_out_2[327],u1_data_out_3[327],partial_product_low0[327],partial_product_low1[327],96'b0};
assign col_out_328 = {u0_col_out_328,u1_data_out_0[328],u1_data_out_1[328],u1_data_out_2[328],u1_data_out_3[328],partial_product_low0[328],partial_product_low1[328],96'b0};
assign col_out_329 = {u0_col_out_329,u1_data_out_0[329],u1_data_out_1[329],u1_data_out_2[329],u1_data_out_3[329],partial_product_low0[329],partial_product_low1[329],96'b0};
assign col_out_330 = {u0_col_out_330,u1_data_out_0[330],u1_data_out_1[330],u1_data_out_2[330],u1_data_out_3[330],partial_product_low0[330],partial_product_low1[330],96'b0};
assign col_out_331 = {u0_col_out_331,u1_data_out_0[331],u1_data_out_1[331],u1_data_out_2[331],u1_data_out_3[331],partial_product_low0[331],partial_product_low1[331],96'b0};
assign col_out_332 = {u0_col_out_332,u1_data_out_0[332],u1_data_out_1[332],u1_data_out_2[332],u1_data_out_3[332],partial_product_low0[332],partial_product_low1[332],96'b0};
assign col_out_333 = {u0_col_out_333,u1_data_out_0[333],u1_data_out_1[333],u1_data_out_2[333],u1_data_out_3[333],partial_product_low0[333],partial_product_low1[333],96'b0};
assign col_out_334 = {u0_col_out_334,u1_data_out_0[334],u1_data_out_1[334],u1_data_out_2[334],u1_data_out_3[334],partial_product_low0[334],partial_product_low1[334],96'b0};
assign col_out_335 = {u0_col_out_335,u1_data_out_0[335],u1_data_out_1[335],u1_data_out_2[335],u1_data_out_3[335],partial_product_low0[335],partial_product_low1[335],96'b0};
assign col_out_336 = {u0_col_out_336,u1_data_out_0[336],u1_data_out_1[336],u1_data_out_2[336],u1_data_out_3[336],partial_product_low0[336],partial_product_low1[336],96'b0};
assign col_out_337 = {u0_col_out_337,u1_data_out_0[337],u1_data_out_1[337],u1_data_out_2[337],u1_data_out_3[337],partial_product_low0[337],partial_product_low1[337],96'b0};
assign col_out_338 = {u0_col_out_338,u1_data_out_0[338],u1_data_out_1[338],u1_data_out_2[338],u1_data_out_3[338],partial_product_low0[338],partial_product_low1[338],96'b0};
assign col_out_339 = {u0_col_out_339,u1_data_out_0[339],u1_data_out_1[339],u1_data_out_2[339],u1_data_out_3[339],partial_product_low0[339],partial_product_low1[339],96'b0};
assign col_out_340 = {u0_col_out_340,u1_data_out_0[340],u1_data_out_1[340],u1_data_out_2[340],u1_data_out_3[340],partial_product_low0[340],partial_product_low1[340],96'b0};
assign col_out_341 = {u0_col_out_341,u1_data_out_0[341],u1_data_out_1[341],u1_data_out_2[341],u1_data_out_3[341],partial_product_low0[341],partial_product_low1[341],96'b0};
assign col_out_342 = {u0_col_out_342,u1_data_out_0[342],u1_data_out_1[342],u1_data_out_2[342],u1_data_out_3[342],partial_product_low0[342],partial_product_low1[342],96'b0};
assign col_out_343 = {u0_col_out_343,u1_data_out_0[343],u1_data_out_1[343],u1_data_out_2[343],u1_data_out_3[343],partial_product_low0[343],partial_product_low1[343],96'b0};
assign col_out_344 = {u0_col_out_344,u1_data_out_0[344],u1_data_out_1[344],u1_data_out_2[344],u1_data_out_3[344],partial_product_low0[344],partial_product_low1[344],96'b0};
assign col_out_345 = {u0_col_out_345,u1_data_out_0[345],u1_data_out_1[345],u1_data_out_2[345],u1_data_out_3[345],partial_product_low0[345],partial_product_low1[345],96'b0};
assign col_out_346 = {u0_col_out_346,u1_data_out_0[346],u1_data_out_1[346],u1_data_out_2[346],u1_data_out_3[346],partial_product_low0[346],partial_product_low1[346],96'b0};
assign col_out_347 = {u0_col_out_347,u1_data_out_0[347],u1_data_out_1[347],u1_data_out_2[347],u1_data_out_3[347],partial_product_low0[347],partial_product_low1[347],96'b0};
assign col_out_348 = {u0_col_out_348,u1_data_out_0[348],u1_data_out_1[348],u1_data_out_2[348],u1_data_out_3[348],partial_product_low0[348],partial_product_low1[348],96'b0};
assign col_out_349 = {u0_col_out_349,u1_data_out_0[349],u1_data_out_1[349],u1_data_out_2[349],u1_data_out_3[349],partial_product_low0[349],partial_product_low1[349],96'b0};
assign col_out_350 = {u0_col_out_350,u1_data_out_0[350],u1_data_out_1[350],u1_data_out_2[350],u1_data_out_3[350],partial_product_low0[350],partial_product_low1[350],96'b0};
assign col_out_351 = {u0_col_out_351,u1_data_out_0[351],u1_data_out_1[351],u1_data_out_2[351],u1_data_out_3[351],partial_product_low0[351],partial_product_low1[351],96'b0};
assign col_out_352 = {u0_col_out_352,u1_data_out_0[352],u1_data_out_1[352],u1_data_out_2[352],u1_data_out_3[352],partial_product_low0[352],partial_product_low1[352],96'b0};
assign col_out_353 = {u0_col_out_353,u1_data_out_0[353],u1_data_out_1[353],u1_data_out_2[353],u1_data_out_3[353],partial_product_low0[353],partial_product_low1[353],96'b0};
assign col_out_354 = {u0_col_out_354,u1_data_out_0[354],u1_data_out_1[354],u1_data_out_2[354],u1_data_out_3[354],partial_product_low0[354],partial_product_low1[354],96'b0};
assign col_out_355 = {u0_col_out_355,u1_data_out_0[355],u1_data_out_1[355],u1_data_out_2[355],u1_data_out_3[355],partial_product_low0[355],partial_product_low1[355],96'b0};
assign col_out_356 = {u0_col_out_356,u1_data_out_0[356],u1_data_out_1[356],u1_data_out_2[356],u1_data_out_3[356],partial_product_low0[356],partial_product_low1[356],96'b0};
assign col_out_357 = {u0_col_out_357,u1_data_out_0[357],u1_data_out_1[357],u1_data_out_2[357],u1_data_out_3[357],partial_product_low0[357],partial_product_low1[357],96'b0};
assign col_out_358 = {u0_col_out_358,u1_data_out_0[358],u1_data_out_1[358],u1_data_out_2[358],u1_data_out_3[358],partial_product_low0[358],partial_product_low1[358],96'b0};
assign col_out_359 = {u0_col_out_359,u1_data_out_0[359],u1_data_out_1[359],u1_data_out_2[359],u1_data_out_3[359],partial_product_low0[359],partial_product_low1[359],96'b0};
assign col_out_360 = {u0_col_out_360,u1_data_out_0[360],u1_data_out_1[360],u1_data_out_2[360],u1_data_out_3[360],partial_product_low0[360],partial_product_low1[360],96'b0};
assign col_out_361 = {u0_col_out_361,u1_data_out_0[361],u1_data_out_1[361],u1_data_out_2[361],u1_data_out_3[361],partial_product_low0[361],partial_product_low1[361],96'b0};
assign col_out_362 = {u0_col_out_362,u1_data_out_0[362],u1_data_out_1[362],u1_data_out_2[362],u1_data_out_3[362],partial_product_low0[362],partial_product_low1[362],96'b0};
assign col_out_363 = {u0_col_out_363,u1_data_out_0[363],u1_data_out_1[363],u1_data_out_2[363],u1_data_out_3[363],partial_product_low0[363],partial_product_low1[363],96'b0};
assign col_out_364 = {u0_col_out_364,u1_data_out_0[364],u1_data_out_1[364],u1_data_out_2[364],u1_data_out_3[364],partial_product_low0[364],partial_product_low1[364],96'b0};
assign col_out_365 = {u0_col_out_365,u1_data_out_0[365],u1_data_out_1[365],u1_data_out_2[365],u1_data_out_3[365],partial_product_low0[365],partial_product_low1[365],96'b0};
assign col_out_366 = {u0_col_out_366,u1_data_out_0[366],u1_data_out_1[366],u1_data_out_2[366],u1_data_out_3[366],partial_product_low0[366],partial_product_low1[366],96'b0};
assign col_out_367 = {u0_col_out_367,u1_data_out_0[367],u1_data_out_1[367],u1_data_out_2[367],u1_data_out_3[367],partial_product_low0[367],partial_product_low1[367],96'b0};
assign col_out_368 = {u0_col_out_368,u1_data_out_0[368],u1_data_out_1[368],u1_data_out_2[368],u1_data_out_3[368],partial_product_low0[368],partial_product_low1[368],96'b0};
assign col_out_369 = {u0_col_out_369,u1_data_out_0[369],u1_data_out_1[369],u1_data_out_2[369],u1_data_out_3[369],partial_product_low0[369],partial_product_low1[369],96'b0};
assign col_out_370 = {u0_col_out_370,u1_data_out_0[370],u1_data_out_1[370],u1_data_out_2[370],u1_data_out_3[370],partial_product_low0[370],partial_product_low1[370],96'b0};
assign col_out_371 = {u0_col_out_371,u1_data_out_0[371],u1_data_out_1[371],u1_data_out_2[371],u1_data_out_3[371],partial_product_low0[371],partial_product_low1[371],96'b0};
assign col_out_372 = {u0_col_out_372,u1_data_out_0[372],u1_data_out_1[372],u1_data_out_2[372],u1_data_out_3[372],partial_product_low0[372],partial_product_low1[372],96'b0};
assign col_out_373 = {u0_col_out_373,u1_data_out_0[373],u1_data_out_1[373],u1_data_out_2[373],u1_data_out_3[373],partial_product_low0[373],partial_product_low1[373],96'b0};
assign col_out_374 = {u0_col_out_374,u1_data_out_0[374],u1_data_out_1[374],u1_data_out_2[374],u1_data_out_3[374],partial_product_low0[374],partial_product_low1[374],96'b0};
assign col_out_375 = {u0_col_out_375,u1_data_out_0[375],u1_data_out_1[375],u1_data_out_2[375],u1_data_out_3[375],partial_product_low0[375],partial_product_low1[375],96'b0};
assign col_out_376 = {u0_col_out_376,u1_data_out_0[376],u1_data_out_1[376],u1_data_out_2[376],u1_data_out_3[376],partial_product_low0[376],partial_product_low1[376],96'b0};
assign col_out_377 = {u0_col_out_377,u1_data_out_0[377],u1_data_out_1[377],u1_data_out_2[377],u1_data_out_3[377],partial_product_low0[377],partial_product_low1[377],96'b0};
assign col_out_378 = {u0_col_out_378,u1_data_out_0[378],u1_data_out_1[378],u1_data_out_2[378],u1_data_out_3[378],partial_product_low0[378],partial_product_low1[378],96'b0};
assign col_out_379 = {u0_col_out_379,u1_data_out_0[379],u1_data_out_1[379],u1_data_out_2[379],u1_data_out_3[379],partial_product_low0[379],partial_product_low1[379],96'b0};
assign col_out_380 = {u0_col_out_380,u1_data_out_0[380],u1_data_out_1[380],u1_data_out_2[380],u1_data_out_3[380],partial_product_low0[380],partial_product_low1[380],96'b0};
assign col_out_381 = {u0_col_out_381,u1_data_out_0[381],u1_data_out_1[381],u1_data_out_2[381],u1_data_out_3[381],partial_product_low0[381],partial_product_low1[381],96'b0};
assign col_out_382 = {u0_col_out_382,u1_data_out_0[382],u1_data_out_1[382],u1_data_out_2[382],u1_data_out_3[382],partial_product_low0[382],partial_product_low1[382],96'b0};
assign col_out_383 = {u0_col_out_383,u1_data_out_0[383],u1_data_out_1[383],u1_data_out_2[383],u1_data_out_3[383],partial_product_low0[383],partial_product_low1[383],96'b0};
assign col_out_384 = {u0_col_out_384,u1_data_out_0[384],u1_data_out_1[384],u1_data_out_2[384],u1_data_out_3[384],partial_product_low0[384],partial_product_low1[384],96'b0};
assign col_out_385 = {u0_col_out_385,u1_data_out_0[385],u1_data_out_1[385],u1_data_out_2[385],u1_data_out_3[385],partial_product_low0[385],partial_product_low1[385],96'b0};
assign col_out_386 = {u0_col_out_386,u1_data_out_0[386],u1_data_out_1[386],u1_data_out_2[386],u1_data_out_3[386],partial_product_low0[386],partial_product_low1[386],96'b0};
assign col_out_387 = {u0_col_out_387,u1_data_out_0[387],u1_data_out_1[387],u1_data_out_2[387],u1_data_out_3[387],partial_product_low0[387],partial_product_low1[387],96'b0};
assign col_out_388 = {u0_col_out_388,u1_data_out_0[388],u1_data_out_1[388],u1_data_out_2[388],u1_data_out_3[388],partial_product_low0[388],partial_product_low1[388],96'b0};
assign col_out_389 = {u0_col_out_389,u1_data_out_0[389],u1_data_out_1[389],u1_data_out_2[389],u1_data_out_3[389],partial_product_low0[389],partial_product_low1[389],96'b0};
assign col_out_390 = {u0_col_out_390,u1_data_out_0[390],u1_data_out_1[390],u1_data_out_2[390],u1_data_out_3[390],partial_product_low0[390],partial_product_low1[390],96'b0};
assign col_out_391 = {u0_col_out_391,u1_data_out_0[391],u1_data_out_1[391],u1_data_out_2[391],u1_data_out_3[391],partial_product_low0[391],partial_product_low1[391],96'b0};
assign col_out_392 = {u0_col_out_392,u1_data_out_0[392],u1_data_out_1[392],u1_data_out_2[392],u1_data_out_3[392],partial_product_low0[392],partial_product_low1[392],96'b0};
assign col_out_393 = {u0_col_out_393,u1_data_out_0[393],u1_data_out_1[393],u1_data_out_2[393],u1_data_out_3[393],partial_product_low0[393],partial_product_low1[393],96'b0};
assign col_out_394 = {u0_col_out_394,u1_data_out_0[394],u1_data_out_1[394],u1_data_out_2[394],u1_data_out_3[394],partial_product_low0[394],partial_product_low1[394],96'b0};
assign col_out_395 = {u0_col_out_395,u1_data_out_0[395],u1_data_out_1[395],u1_data_out_2[395],u1_data_out_3[395],partial_product_low0[395],partial_product_low1[395],96'b0};
assign col_out_396 = {u0_col_out_396,u1_data_out_0[396],u1_data_out_1[396],u1_data_out_2[396],u1_data_out_3[396],partial_product_low0[396],partial_product_low1[396],96'b0};
assign col_out_397 = {u0_col_out_397,u1_data_out_0[397],u1_data_out_1[397],u1_data_out_2[397],u1_data_out_3[397],partial_product_low0[397],partial_product_low1[397],96'b0};
assign col_out_398 = {u0_col_out_398,u1_data_out_0[398],u1_data_out_1[398],u1_data_out_2[398],u1_data_out_3[398],partial_product_low0[398],partial_product_low1[398],96'b0};
assign col_out_399 = {u0_col_out_399,u1_data_out_0[399],u1_data_out_1[399],u1_data_out_2[399],u1_data_out_3[399],partial_product_low0[399],partial_product_low1[399],96'b0};
assign col_out_400 = {u0_col_out_400,u1_data_out_0[400],u1_data_out_1[400],u1_data_out_2[400],u1_data_out_3[400],partial_product_low0[400],partial_product_low1[400],96'b0};
assign col_out_401 = {u0_col_out_401,u1_data_out_0[401],u1_data_out_1[401],u1_data_out_2[401],u1_data_out_3[401],partial_product_low0[401],partial_product_low1[401],96'b0};
assign col_out_402 = {u0_col_out_402,u1_data_out_0[402],u1_data_out_1[402],u1_data_out_2[402],u1_data_out_3[402],partial_product_low0[402],partial_product_low1[402],96'b0};
assign col_out_403 = {u0_col_out_403,u1_data_out_0[403],u1_data_out_1[403],u1_data_out_2[403],u1_data_out_3[403],partial_product_low0[403],partial_product_low1[403],96'b0};
assign col_out_404 = {u0_col_out_404,u1_data_out_0[404],u1_data_out_1[404],u1_data_out_2[404],u1_data_out_3[404],partial_product_low0[404],partial_product_low1[404],96'b0};
assign col_out_405 = {u0_col_out_405,u1_data_out_0[405],u1_data_out_1[405],u1_data_out_2[405],u1_data_out_3[405],partial_product_low0[405],partial_product_low1[405],96'b0};
assign col_out_406 = {u0_col_out_406,u1_data_out_0[406],u1_data_out_1[406],u1_data_out_2[406],u1_data_out_3[406],partial_product_low0[406],partial_product_low1[406],96'b0};
assign col_out_407 = {u0_col_out_407,u1_data_out_0[407],u1_data_out_1[407],u1_data_out_2[407],u1_data_out_3[407],partial_product_low0[407],partial_product_low1[407],96'b0};
assign col_out_408 = {u0_col_out_408,u1_data_out_0[408],u1_data_out_1[408],u1_data_out_2[408],u1_data_out_3[408],partial_product_low0[408],partial_product_low1[408],96'b0};
assign col_out_409 = {u0_col_out_409,u1_data_out_0[409],u1_data_out_1[409],u1_data_out_2[409],u1_data_out_3[409],partial_product_low0[409],partial_product_low1[409],96'b0};
assign col_out_410 = {u0_col_out_410,u1_data_out_0[410],u1_data_out_1[410],u1_data_out_2[410],u1_data_out_3[410],partial_product_low0[410],partial_product_low1[410],96'b0};
assign col_out_411 = {u0_col_out_411,u1_data_out_0[411],u1_data_out_1[411],u1_data_out_2[411],u1_data_out_3[411],partial_product_low0[411],partial_product_low1[411],96'b0};
assign col_out_412 = {u0_col_out_412,u1_data_out_0[412],u1_data_out_1[412],u1_data_out_2[412],u1_data_out_3[412],partial_product_low0[412],partial_product_low1[412],96'b0};
assign col_out_413 = {u0_col_out_413,u1_data_out_0[413],u1_data_out_1[413],u1_data_out_2[413],u1_data_out_3[413],partial_product_low0[413],partial_product_low1[413],96'b0};
assign col_out_414 = {u0_col_out_414,u1_data_out_0[414],u1_data_out_1[414],u1_data_out_2[414],u1_data_out_3[414],partial_product_low0[414],partial_product_low1[414],96'b0};
assign col_out_415 = {u0_col_out_415,u1_data_out_0[415],u1_data_out_1[415],u1_data_out_2[415],u1_data_out_3[415],partial_product_low0[415],partial_product_low1[415],96'b0};
assign col_out_416 = {u0_col_out_416,u1_data_out_0[416],u1_data_out_1[416],u1_data_out_2[416],u1_data_out_3[416],partial_product_low0[416],partial_product_low1[416],96'b0};
assign col_out_417 = {u0_col_out_417,u1_data_out_0[417],u1_data_out_1[417],u1_data_out_2[417],u1_data_out_3[417],partial_product_low0[417],partial_product_low1[417],96'b0};
assign col_out_418 = {u0_col_out_418,u1_data_out_0[418],u1_data_out_1[418],u1_data_out_2[418],u1_data_out_3[418],partial_product_low0[418],partial_product_low1[418],96'b0};
assign col_out_419 = {u0_col_out_419,u1_data_out_0[419],u1_data_out_1[419],u1_data_out_2[419],u1_data_out_3[419],partial_product_low0[419],partial_product_low1[419],96'b0};
assign col_out_420 = {u0_col_out_420,u1_data_out_0[420],u1_data_out_1[420],u1_data_out_2[420],u1_data_out_3[420],partial_product_low0[420],partial_product_low1[420],96'b0};
assign col_out_421 = {u0_col_out_421,u1_data_out_0[421],u1_data_out_1[421],u1_data_out_2[421],u1_data_out_3[421],partial_product_low0[421],partial_product_low1[421],96'b0};
assign col_out_422 = {u0_col_out_422,u1_data_out_0[422],u1_data_out_1[422],u1_data_out_2[422],u1_data_out_3[422],partial_product_low0[422],partial_product_low1[422],96'b0};
assign col_out_423 = {u0_col_out_423,u1_data_out_0[423],u1_data_out_1[423],u1_data_out_2[423],u1_data_out_3[423],partial_product_low0[423],partial_product_low1[423],96'b0};
assign col_out_424 = {u0_col_out_424,u1_data_out_0[424],u1_data_out_1[424],u1_data_out_2[424],u1_data_out_3[424],partial_product_low0[424],partial_product_low1[424],96'b0};
assign col_out_425 = {u0_col_out_425,u1_data_out_0[425],u1_data_out_1[425],u1_data_out_2[425],u1_data_out_3[425],partial_product_low0[425],partial_product_low1[425],96'b0};
assign col_out_426 = {u0_col_out_426,u1_data_out_0[426],u1_data_out_1[426],u1_data_out_2[426],u1_data_out_3[426],partial_product_low0[426],partial_product_low1[426],96'b0};
assign col_out_427 = {u0_col_out_427,u1_data_out_0[427],u1_data_out_1[427],u1_data_out_2[427],u1_data_out_3[427],partial_product_low0[427],partial_product_low1[427],96'b0};
assign col_out_428 = {u0_col_out_428,u1_data_out_0[428],u1_data_out_1[428],u1_data_out_2[428],u1_data_out_3[428],partial_product_low0[428],partial_product_low1[428],96'b0};
assign col_out_429 = {u0_col_out_429,u1_data_out_0[429],u1_data_out_1[429],u1_data_out_2[429],u1_data_out_3[429],partial_product_low0[429],partial_product_low1[429],96'b0};
assign col_out_430 = {u0_col_out_430,u1_data_out_0[430],u1_data_out_1[430],u1_data_out_2[430],u1_data_out_3[430],partial_product_low0[430],partial_product_low1[430],96'b0};
assign col_out_431 = {u0_col_out_431,u1_data_out_0[431],u1_data_out_1[431],u1_data_out_2[431],u1_data_out_3[431],partial_product_low0[431],partial_product_low1[431],96'b0};
assign col_out_432 = {u0_col_out_432,u1_data_out_0[432],u1_data_out_1[432],u1_data_out_2[432],u1_data_out_3[432],partial_product_low0[432],partial_product_low1[432],96'b0};
assign col_out_433 = {u0_col_out_433,u1_data_out_0[433],u1_data_out_1[433],u1_data_out_2[433],u1_data_out_3[433],partial_product_low0[433],partial_product_low1[433],96'b0};
assign col_out_434 = {u0_col_out_434,u1_data_out_0[434],u1_data_out_1[434],u1_data_out_2[434],u1_data_out_3[434],partial_product_low0[434],partial_product_low1[434],96'b0};
assign col_out_435 = {u0_col_out_435,u1_data_out_0[435],u1_data_out_1[435],u1_data_out_2[435],u1_data_out_3[435],partial_product_low0[435],partial_product_low1[435],96'b0};
assign col_out_436 = {u0_col_out_436,u1_data_out_0[436],u1_data_out_1[436],u1_data_out_2[436],u1_data_out_3[436],partial_product_low0[436],partial_product_low1[436],96'b0};
assign col_out_437 = {u0_col_out_437,u1_data_out_0[437],u1_data_out_1[437],u1_data_out_2[437],u1_data_out_3[437],partial_product_low0[437],partial_product_low1[437],96'b0};
assign col_out_438 = {u0_col_out_438,u1_data_out_0[438],u1_data_out_1[438],u1_data_out_2[438],u1_data_out_3[438],partial_product_low0[438],partial_product_low1[438],96'b0};
assign col_out_439 = {u0_col_out_439,u1_data_out_0[439],u1_data_out_1[439],u1_data_out_2[439],u1_data_out_3[439],partial_product_low0[439],partial_product_low1[439],96'b0};
assign col_out_440 = {u0_col_out_440,u1_data_out_0[440],u1_data_out_1[440],u1_data_out_2[440],u1_data_out_3[440],partial_product_low0[440],partial_product_low1[440],96'b0};
assign col_out_441 = {u0_col_out_441,u1_data_out_0[441],u1_data_out_1[441],u1_data_out_2[441],u1_data_out_3[441],partial_product_low0[441],partial_product_low1[441],96'b0};
assign col_out_442 = {u0_col_out_442,u1_data_out_0[442],u1_data_out_1[442],u1_data_out_2[442],u1_data_out_3[442],partial_product_low0[442],partial_product_low1[442],96'b0};
assign col_out_443 = {u0_col_out_443,u1_data_out_0[443],u1_data_out_1[443],u1_data_out_2[443],u1_data_out_3[443],partial_product_low0[443],partial_product_low1[443],96'b0};
assign col_out_444 = {u0_col_out_444,u1_data_out_0[444],u1_data_out_1[444],u1_data_out_2[444],u1_data_out_3[444],partial_product_low0[444],partial_product_low1[444],96'b0};
assign col_out_445 = {u0_col_out_445,u1_data_out_0[445],u1_data_out_1[445],u1_data_out_2[445],u1_data_out_3[445],partial_product_low0[445],partial_product_low1[445],96'b0};
assign col_out_446 = {u0_col_out_446,u1_data_out_0[446],u1_data_out_1[446],u1_data_out_2[446],u1_data_out_3[446],partial_product_low0[446],partial_product_low1[446],96'b0};
assign col_out_447 = {u0_col_out_447,u1_data_out_0[447],u1_data_out_1[447],u1_data_out_2[447],u1_data_out_3[447],partial_product_low0[447],partial_product_low1[447],96'b0};
assign col_out_448 = {u0_col_out_448,u1_data_out_0[448],u1_data_out_1[448],u1_data_out_2[448],u1_data_out_3[448],partial_product_low0[448],partial_product_low1[448],96'b0};
assign col_out_449 = {u0_col_out_449,u1_data_out_0[449],u1_data_out_1[449],u1_data_out_2[449],u1_data_out_3[449],partial_product_low0[449],partial_product_low1[449],96'b0};
assign col_out_450 = {u0_col_out_450,u1_data_out_0[450],u1_data_out_1[450],u1_data_out_2[450],u1_data_out_3[450],partial_product_low0[450],partial_product_low1[450],96'b0};
assign col_out_451 = {u0_col_out_451,u1_data_out_0[451],u1_data_out_1[451],u1_data_out_2[451],u1_data_out_3[451],partial_product_low0[451],partial_product_low1[451],96'b0};
assign col_out_452 = {u0_col_out_452,u1_data_out_0[452],u1_data_out_1[452],u1_data_out_2[452],u1_data_out_3[452],partial_product_low0[452],partial_product_low1[452],96'b0};
assign col_out_453 = {u0_col_out_453,u1_data_out_0[453],u1_data_out_1[453],u1_data_out_2[453],u1_data_out_3[453],partial_product_low0[453],partial_product_low1[453],96'b0};
assign col_out_454 = {u0_col_out_454,u1_data_out_0[454],u1_data_out_1[454],u1_data_out_2[454],u1_data_out_3[454],partial_product_low0[454],partial_product_low1[454],96'b0};
assign col_out_455 = {u0_col_out_455,u1_data_out_0[455],u1_data_out_1[455],u1_data_out_2[455],u1_data_out_3[455],partial_product_low0[455],partial_product_low1[455],96'b0};
assign col_out_456 = {u0_col_out_456,u1_data_out_0[456],u1_data_out_1[456],u1_data_out_2[456],u1_data_out_3[456],partial_product_low0[456],partial_product_low1[456],96'b0};
assign col_out_457 = {u0_col_out_457,u1_data_out_0[457],u1_data_out_1[457],u1_data_out_2[457],u1_data_out_3[457],partial_product_low0[457],partial_product_low1[457],96'b0};
assign col_out_458 = {u0_col_out_458,u1_data_out_0[458],u1_data_out_1[458],u1_data_out_2[458],u1_data_out_3[458],partial_product_low0[458],partial_product_low1[458],96'b0};
assign col_out_459 = {u0_col_out_459,u1_data_out_0[459],u1_data_out_1[459],u1_data_out_2[459],u1_data_out_3[459],partial_product_low0[459],partial_product_low1[459],96'b0};
assign col_out_460 = {u0_col_out_460,u1_data_out_0[460],u1_data_out_1[460],u1_data_out_2[460],u1_data_out_3[460],partial_product_low0[460],partial_product_low1[460],96'b0};
assign col_out_461 = {u0_col_out_461,u1_data_out_0[461],u1_data_out_1[461],u1_data_out_2[461],u1_data_out_3[461],partial_product_low0[461],partial_product_low1[461],96'b0};
assign col_out_462 = {u0_col_out_462,u1_data_out_0[462],u1_data_out_1[462],u1_data_out_2[462],u1_data_out_3[462],partial_product_low0[462],partial_product_low1[462],96'b0};
assign col_out_463 = {u0_col_out_463,u1_data_out_0[463],u1_data_out_1[463],u1_data_out_2[463],u1_data_out_3[463],partial_product_low0[463],partial_product_low1[463],96'b0};
assign col_out_464 = {u0_col_out_464,u1_data_out_0[464],u1_data_out_1[464],u1_data_out_2[464],u1_data_out_3[464],partial_product_low0[464],partial_product_low1[464],96'b0};
assign col_out_465 = {u0_col_out_465,u1_data_out_0[465],u1_data_out_1[465],u1_data_out_2[465],u1_data_out_3[465],partial_product_low0[465],partial_product_low1[465],96'b0};
assign col_out_466 = {u0_col_out_466,u1_data_out_0[466],u1_data_out_1[466],u1_data_out_2[466],u1_data_out_3[466],partial_product_low0[466],partial_product_low1[466],96'b0};
assign col_out_467 = {u0_col_out_467,u1_data_out_0[467],u1_data_out_1[467],u1_data_out_2[467],u1_data_out_3[467],partial_product_low0[467],partial_product_low1[467],96'b0};
assign col_out_468 = {u0_col_out_468,u1_data_out_0[468],u1_data_out_1[468],u1_data_out_2[468],u1_data_out_3[468],partial_product_low0[468],partial_product_low1[468],96'b0};
assign col_out_469 = {u0_col_out_469,u1_data_out_0[469],u1_data_out_1[469],u1_data_out_2[469],u1_data_out_3[469],partial_product_low0[469],partial_product_low1[469],96'b0};
assign col_out_470 = {u0_col_out_470,u1_data_out_0[470],u1_data_out_1[470],u1_data_out_2[470],u1_data_out_3[470],partial_product_low0[470],partial_product_low1[470],96'b0};
assign col_out_471 = {u0_col_out_471,u1_data_out_0[471],u1_data_out_1[471],u1_data_out_2[471],u1_data_out_3[471],partial_product_low0[471],partial_product_low1[471],96'b0};
assign col_out_472 = {u0_col_out_472,u1_data_out_0[472],u1_data_out_1[472],u1_data_out_2[472],u1_data_out_3[472],partial_product_low0[472],partial_product_low1[472],96'b0};
assign col_out_473 = {u0_col_out_473,u1_data_out_0[473],u1_data_out_1[473],u1_data_out_2[473],u1_data_out_3[473],partial_product_low0[473],partial_product_low1[473],96'b0};
assign col_out_474 = {u0_col_out_474,u1_data_out_0[474],u1_data_out_1[474],u1_data_out_2[474],u1_data_out_3[474],partial_product_low0[474],partial_product_low1[474],96'b0};
assign col_out_475 = {u0_col_out_475,u1_data_out_0[475],u1_data_out_1[475],u1_data_out_2[475],u1_data_out_3[475],partial_product_low0[475],partial_product_low1[475],96'b0};
assign col_out_476 = {u0_col_out_476,u1_data_out_0[476],u1_data_out_1[476],u1_data_out_2[476],u1_data_out_3[476],partial_product_low0[476],partial_product_low1[476],96'b0};
assign col_out_477 = {u0_col_out_477,u1_data_out_0[477],u1_data_out_1[477],u1_data_out_2[477],u1_data_out_3[477],partial_product_low0[477],partial_product_low1[477],96'b0};
assign col_out_478 = {u0_col_out_478,u1_data_out_0[478],u1_data_out_1[478],u1_data_out_2[478],u1_data_out_3[478],partial_product_low0[478],partial_product_low1[478],96'b0};
assign col_out_479 = {u0_col_out_479,u1_data_out_0[479],u1_data_out_1[479],u1_data_out_2[479],u1_data_out_3[479],partial_product_low0[479],partial_product_low1[479],96'b0};
assign col_out_480 = {u0_col_out_480,u1_data_out_0[480],u1_data_out_1[480],u1_data_out_2[480],u1_data_out_3[480],partial_product_low0[480],partial_product_low1[480],96'b0};
assign col_out_481 = {u0_col_out_481,u1_data_out_0[481],u1_data_out_1[481],u1_data_out_2[481],u1_data_out_3[481],partial_product_low0[481],partial_product_low1[481],96'b0};
assign col_out_482 = {u0_col_out_482,u1_data_out_0[482],u1_data_out_1[482],u1_data_out_2[482],u1_data_out_3[482],partial_product_low0[482],partial_product_low1[482],96'b0};
assign col_out_483 = {u0_col_out_483,u1_data_out_0[483],u1_data_out_1[483],u1_data_out_2[483],u1_data_out_3[483],partial_product_low0[483],partial_product_low1[483],96'b0};
assign col_out_484 = {u0_col_out_484,u1_data_out_0[484],u1_data_out_1[484],u1_data_out_2[484],u1_data_out_3[484],partial_product_low0[484],partial_product_low1[484],96'b0};
assign col_out_485 = {u0_col_out_485,u1_data_out_0[485],u1_data_out_1[485],u1_data_out_2[485],u1_data_out_3[485],partial_product_low0[485],partial_product_low1[485],96'b0};
assign col_out_486 = {u0_col_out_486,u1_data_out_0[486],u1_data_out_1[486],u1_data_out_2[486],u1_data_out_3[486],partial_product_low0[486],partial_product_low1[486],96'b0};
assign col_out_487 = {u0_col_out_487,u1_data_out_0[487],u1_data_out_1[487],u1_data_out_2[487],u1_data_out_3[487],partial_product_low0[487],partial_product_low1[487],96'b0};
assign col_out_488 = {u0_col_out_488,u1_data_out_0[488],u1_data_out_1[488],u1_data_out_2[488],u1_data_out_3[488],partial_product_low0[488],partial_product_low1[488],96'b0};
assign col_out_489 = {u0_col_out_489,u1_data_out_0[489],u1_data_out_1[489],u1_data_out_2[489],u1_data_out_3[489],partial_product_low0[489],partial_product_low1[489],96'b0};
assign col_out_490 = {u0_col_out_490,u1_data_out_0[490],u1_data_out_1[490],u1_data_out_2[490],u1_data_out_3[490],partial_product_low0[490],partial_product_low1[490],96'b0};
assign col_out_491 = {u0_col_out_491,u1_data_out_0[491],u1_data_out_1[491],u1_data_out_2[491],u1_data_out_3[491],partial_product_low0[491],partial_product_low1[491],96'b0};
assign col_out_492 = {u0_col_out_492,u1_data_out_0[492],u1_data_out_1[492],u1_data_out_2[492],u1_data_out_3[492],partial_product_low0[492],partial_product_low1[492],96'b0};
assign col_out_493 = {u0_col_out_493,u1_data_out_0[493],u1_data_out_1[493],u1_data_out_2[493],u1_data_out_3[493],partial_product_low0[493],partial_product_low1[493],96'b0};
assign col_out_494 = {u0_col_out_494,u1_data_out_0[494],u1_data_out_1[494],u1_data_out_2[494],u1_data_out_3[494],partial_product_low0[494],partial_product_low1[494],96'b0};
assign col_out_495 = {u0_col_out_495,u1_data_out_0[495],u1_data_out_1[495],u1_data_out_2[495],u1_data_out_3[495],partial_product_low0[495],partial_product_low1[495],96'b0};
assign col_out_496 = {u0_col_out_496,u1_data_out_0[496],u1_data_out_1[496],u1_data_out_2[496],u1_data_out_3[496],partial_product_low0[496],partial_product_low1[496],96'b0};
assign col_out_497 = {u0_col_out_497,u1_data_out_0[497],u1_data_out_1[497],u1_data_out_2[497],u1_data_out_3[497],partial_product_low0[497],partial_product_low1[497],96'b0};
assign col_out_498 = {u0_col_out_498,u1_data_out_0[498],u1_data_out_1[498],u1_data_out_2[498],u1_data_out_3[498],partial_product_low0[498],partial_product_low1[498],96'b0};
assign col_out_499 = {u0_col_out_499,u1_data_out_0[499],u1_data_out_1[499],u1_data_out_2[499],u1_data_out_3[499],partial_product_low0[499],partial_product_low1[499],96'b0};
assign col_out_500 = {u0_col_out_500,u1_data_out_0[500],u1_data_out_1[500],u1_data_out_2[500],u1_data_out_3[500],partial_product_low0[500],partial_product_low1[500],96'b0};
assign col_out_501 = {u0_col_out_501,u1_data_out_0[501],u1_data_out_1[501],u1_data_out_2[501],u1_data_out_3[501],partial_product_low0[501],partial_product_low1[501],96'b0};
assign col_out_502 = {u0_col_out_502,u1_data_out_0[502],u1_data_out_1[502],u1_data_out_2[502],u1_data_out_3[502],partial_product_low0[502],partial_product_low1[502],96'b0};
assign col_out_503 = {u0_col_out_503,u1_data_out_0[503],u1_data_out_1[503],u1_data_out_2[503],u1_data_out_3[503],partial_product_low0[503],partial_product_low1[503],96'b0};
assign col_out_504 = {u0_col_out_504,u1_data_out_0[504],u1_data_out_1[504],u1_data_out_2[504],u1_data_out_3[504],partial_product_low0[504],partial_product_low1[504],96'b0};
assign col_out_505 = {u0_col_out_505,u1_data_out_0[505],u1_data_out_1[505],u1_data_out_2[505],u1_data_out_3[505],partial_product_low0[505],partial_product_low1[505],96'b0};
assign col_out_506 = {u0_col_out_506,u1_data_out_0[506],u1_data_out_1[506],u1_data_out_2[506],u1_data_out_3[506],partial_product_low0[506],partial_product_low1[506],96'b0};
assign col_out_507 = {u0_col_out_507,u1_data_out_0[507],u1_data_out_1[507],u1_data_out_2[507],u1_data_out_3[507],partial_product_low0[507],partial_product_low1[507],96'b0};
assign col_out_508 = {u0_col_out_508,u1_data_out_0[508],u1_data_out_1[508],u1_data_out_2[508],u1_data_out_3[508],partial_product_low0[508],partial_product_low1[508],96'b0};
assign col_out_509 = {u0_col_out_509,u1_data_out_0[509],u1_data_out_1[509],u1_data_out_2[509],u1_data_out_3[509],partial_product_low0[509],partial_product_low1[509],96'b0};
assign col_out_510 = {u0_col_out_510,u1_data_out_0[510],u1_data_out_1[510],u1_data_out_2[510],u1_data_out_3[510],partial_product_low0[510],partial_product_low1[510],96'b0};
assign col_out_511 = {u0_col_out_511,u1_data_out_0[511],u1_data_out_1[511],u1_data_out_2[511],u1_data_out_3[511],partial_product_low0[511],partial_product_low1[511],96'b0};
assign col_out_512 = {u0_col_out_512,u1_data_out_0[512],u1_data_out_1[512],u1_data_out_2[512],u1_data_out_3[512],partial_product_low0[512],partial_product_low1[512],96'b0};
assign col_out_513 = {u0_col_out_513,u1_data_out_0[513],u1_data_out_1[513],u1_data_out_2[513],u1_data_out_3[513],partial_product_low0[513],partial_product_low1[513],96'b0};
assign col_out_514 = {u0_col_out_514,u1_data_out_0[514],u1_data_out_1[514],u1_data_out_2[514],u1_data_out_3[514],partial_product_low0[514],partial_product_low1[514],96'b0};
assign col_out_515 = {u0_col_out_515,u1_data_out_0[515],u1_data_out_1[515],u1_data_out_2[515],u1_data_out_3[515],partial_product_low0[515],partial_product_low1[515],96'b0};
assign col_out_516 = {u0_col_out_516,u1_data_out_0[516],u1_data_out_1[516],u1_data_out_2[516],u1_data_out_3[516],partial_product_low0[516],partial_product_low1[516],96'b0};
assign col_out_517 = {u0_col_out_517,u1_data_out_0[517],u1_data_out_1[517],u1_data_out_2[517],u1_data_out_3[517],partial_product_low0[517],partial_product_low1[517],96'b0};
assign col_out_518 = {u0_col_out_518,u1_data_out_0[518],u1_data_out_1[518],u1_data_out_2[518],u1_data_out_3[518],partial_product_low0[518],partial_product_low1[518],96'b0};
assign col_out_519 = {u0_col_out_519,u1_data_out_0[519],u1_data_out_1[519],u1_data_out_2[519],u1_data_out_3[519],partial_product_low0[519],partial_product_low1[519],96'b0};
assign col_out_520 = {u0_col_out_520,u1_data_out_0[520],u1_data_out_1[520],u1_data_out_2[520],u1_data_out_3[520],partial_product_low0[520],partial_product_low1[520],96'b0};
assign col_out_521 = {u0_col_out_521,u1_data_out_0[521],u1_data_out_1[521],u1_data_out_2[521],u1_data_out_3[521],partial_product_low0[521],partial_product_low1[521],96'b0};
assign col_out_522 = {u0_col_out_522,u1_data_out_0[522],u1_data_out_1[522],u1_data_out_2[522],u1_data_out_3[522],partial_product_low0[522],partial_product_low1[522],96'b0};
assign col_out_523 = {u0_col_out_523,u1_data_out_0[523],u1_data_out_1[523],u1_data_out_2[523],u1_data_out_3[523],partial_product_low0[523],partial_product_low1[523],96'b0};
assign col_out_524 = {u0_col_out_524,u1_data_out_0[524],u1_data_out_1[524],u1_data_out_2[524],u1_data_out_3[524],partial_product_low0[524],partial_product_low1[524],96'b0};
assign col_out_525 = {u0_col_out_525,u1_data_out_0[525],u1_data_out_1[525],u1_data_out_2[525],u1_data_out_3[525],partial_product_low0[525],partial_product_low1[525],96'b0};
assign col_out_526 = {u0_col_out_526,u1_data_out_0[526],u1_data_out_1[526],u1_data_out_2[526],u1_data_out_3[526],partial_product_low0[526],partial_product_low1[526],96'b0};
assign col_out_527 = {u0_col_out_527,u1_data_out_0[527],u1_data_out_1[527],u1_data_out_2[527],u1_data_out_3[527],partial_product_low0[527],partial_product_low1[527],96'b0};
assign col_out_528 = {u0_col_out_528,u1_data_out_0[528],u1_data_out_1[528],u1_data_out_2[528],u1_data_out_3[528],partial_product_low0[528],partial_product_low1[528],96'b0};
assign col_out_529 = {u0_col_out_529,u1_data_out_0[529],u1_data_out_1[529],u1_data_out_2[529],u1_data_out_3[529],partial_product_low0[529],partial_product_low1[529],96'b0};
assign col_out_530 = {u0_col_out_530,u1_data_out_0[530],u1_data_out_1[530],u1_data_out_2[530],u1_data_out_3[530],partial_product_low0[530],partial_product_low1[530],96'b0};
assign col_out_531 = {u0_col_out_531,u1_data_out_0[531],u1_data_out_1[531],u1_data_out_2[531],u1_data_out_3[531],partial_product_low0[531],partial_product_low1[531],96'b0};
assign col_out_532 = {u0_col_out_532,u1_data_out_0[532],u1_data_out_1[532],u1_data_out_2[532],u1_data_out_3[532],partial_product_low0[532],partial_product_low1[532],96'b0};
assign col_out_533 = {u0_col_out_533,u1_data_out_0[533],u1_data_out_1[533],u1_data_out_2[533],u1_data_out_3[533],partial_product_low0[533],partial_product_low1[533],96'b0};
assign col_out_534 = {u0_col_out_534,u1_data_out_0[534],u1_data_out_1[534],u1_data_out_2[534],u1_data_out_3[534],partial_product_low0[534],partial_product_low1[534],96'b0};
assign col_out_535 = {u0_col_out_535,u1_data_out_0[535],u1_data_out_1[535],u1_data_out_2[535],u1_data_out_3[535],partial_product_low0[535],partial_product_low1[535],96'b0};
assign col_out_536 = {u0_col_out_536,u1_data_out_0[536],u1_data_out_1[536],u1_data_out_2[536],u1_data_out_3[536],partial_product_low0[536],partial_product_low1[536],96'b0};
assign col_out_537 = {u0_col_out_537,u1_data_out_0[537],u1_data_out_1[537],u1_data_out_2[537],u1_data_out_3[537],partial_product_low0[537],partial_product_low1[537],96'b0};
assign col_out_538 = {u0_col_out_538,u1_data_out_0[538],u1_data_out_1[538],u1_data_out_2[538],u1_data_out_3[538],partial_product_low0[538],partial_product_low1[538],96'b0};
assign col_out_539 = {u0_col_out_539,u1_data_out_0[539],u1_data_out_1[539],u1_data_out_2[539],u1_data_out_3[539],partial_product_low0[539],partial_product_low1[539],96'b0};
assign col_out_540 = {u0_col_out_540,u1_data_out_0[540],u1_data_out_1[540],u1_data_out_2[540],u1_data_out_3[540],partial_product_low0[540],partial_product_low1[540],96'b0};
assign col_out_541 = {u0_col_out_541,u1_data_out_0[541],u1_data_out_1[541],u1_data_out_2[541],u1_data_out_3[541],partial_product_low0[541],partial_product_low1[541],96'b0};
assign col_out_542 = {u0_col_out_542,u1_data_out_0[542],u1_data_out_1[542],u1_data_out_2[542],u1_data_out_3[542],partial_product_low0[542],partial_product_low1[542],96'b0};
assign col_out_543 = {u0_col_out_543,u1_data_out_0[543],u1_data_out_1[543],u1_data_out_2[543],u1_data_out_3[543],partial_product_low0[543],partial_product_low1[543],96'b0};
assign col_out_544 = {u0_col_out_544,u1_data_out_0[544],u1_data_out_1[544],u1_data_out_2[544],u1_data_out_3[544],partial_product_low0[544],partial_product_low1[544],96'b0};
assign col_out_545 = {u0_col_out_545,u1_data_out_0[545],u1_data_out_1[545],u1_data_out_2[545],u1_data_out_3[545],partial_product_low0[545],partial_product_low1[545],96'b0};
assign col_out_546 = {u0_col_out_546,u1_data_out_0[546],u1_data_out_1[546],u1_data_out_2[546],u1_data_out_3[546],partial_product_low0[546],partial_product_low1[546],96'b0};
assign col_out_547 = {u0_col_out_547,u1_data_out_0[547],u1_data_out_1[547],u1_data_out_2[547],u1_data_out_3[547],partial_product_low0[547],partial_product_low1[547],96'b0};
assign col_out_548 = {u0_col_out_548,u1_data_out_0[548],u1_data_out_1[548],u1_data_out_2[548],u1_data_out_3[548],partial_product_low0[548],partial_product_low1[548],96'b0};
assign col_out_549 = {u0_col_out_549,u1_data_out_0[549],u1_data_out_1[549],u1_data_out_2[549],u1_data_out_3[549],partial_product_low0[549],partial_product_low1[549],96'b0};
assign col_out_550 = {u0_col_out_550,u1_data_out_0[550],u1_data_out_1[550],u1_data_out_2[550],u1_data_out_3[550],partial_product_low0[550],partial_product_low1[550],96'b0};
assign col_out_551 = {u0_col_out_551,u1_data_out_0[551],u1_data_out_1[551],u1_data_out_2[551],u1_data_out_3[551],partial_product_low0[551],partial_product_low1[551],96'b0};
assign col_out_552 = {u0_col_out_552,u1_data_out_0[552],u1_data_out_1[552],u1_data_out_2[552],u1_data_out_3[552],partial_product_low0[552],partial_product_low1[552],96'b0};
assign col_out_553 = {u0_col_out_553,u1_data_out_0[553],u1_data_out_1[553],u1_data_out_2[553],u1_data_out_3[553],partial_product_low0[553],partial_product_low1[553],96'b0};
assign col_out_554 = {u0_col_out_554,u1_data_out_0[554],u1_data_out_1[554],u1_data_out_2[554],u1_data_out_3[554],partial_product_low0[554],partial_product_low1[554],96'b0};
assign col_out_555 = {u0_col_out_555,u1_data_out_0[555],u1_data_out_1[555],u1_data_out_2[555],u1_data_out_3[555],partial_product_low0[555],partial_product_low1[555],96'b0};
assign col_out_556 = {u0_col_out_556,u1_data_out_0[556],u1_data_out_1[556],u1_data_out_2[556],u1_data_out_3[556],partial_product_low0[556],partial_product_low1[556],96'b0};
assign col_out_557 = {u0_col_out_557,u1_data_out_0[557],u1_data_out_1[557],u1_data_out_2[557],u1_data_out_3[557],partial_product_low0[557],partial_product_low1[557],96'b0};
assign col_out_558 = {u0_col_out_558,u1_data_out_0[558],u1_data_out_1[558],u1_data_out_2[558],u1_data_out_3[558],partial_product_low0[558],partial_product_low1[558],96'b0};
assign col_out_559 = {u0_col_out_559,u1_data_out_0[559],u1_data_out_1[559],u1_data_out_2[559],u1_data_out_3[559],partial_product_low0[559],partial_product_low1[559],96'b0};
assign col_out_560 = {u0_col_out_560,u1_data_out_0[560],u1_data_out_1[560],u1_data_out_2[560],u1_data_out_3[560],partial_product_low0[560],partial_product_low1[560],96'b0};
assign col_out_561 = {u0_col_out_561,u1_data_out_0[561],u1_data_out_1[561],u1_data_out_2[561],u1_data_out_3[561],partial_product_low0[561],partial_product_low1[561],96'b0};
assign col_out_562 = {u0_col_out_562,u1_data_out_0[562],u1_data_out_1[562],u1_data_out_2[562],u1_data_out_3[562],partial_product_low0[562],partial_product_low1[562],96'b0};
assign col_out_563 = {u0_col_out_563,u1_data_out_0[563],u1_data_out_1[563],u1_data_out_2[563],u1_data_out_3[563],partial_product_low0[563],partial_product_low1[563],96'b0};
assign col_out_564 = {u0_col_out_564,u1_data_out_0[564],u1_data_out_1[564],u1_data_out_2[564],u1_data_out_3[564],partial_product_low0[564],partial_product_low1[564],96'b0};
assign col_out_565 = {u0_col_out_565,u1_data_out_0[565],u1_data_out_1[565],u1_data_out_2[565],u1_data_out_3[565],partial_product_low0[565],partial_product_low1[565],96'b0};
assign col_out_566 = {u0_col_out_566,u1_data_out_0[566],u1_data_out_1[566],u1_data_out_2[566],u1_data_out_3[566],partial_product_low0[566],partial_product_low1[566],96'b0};
assign col_out_567 = {u0_col_out_567,u1_data_out_0[567],u1_data_out_1[567],u1_data_out_2[567],u1_data_out_3[567],partial_product_low0[567],partial_product_low1[567],96'b0};
assign col_out_568 = {u0_col_out_568,u1_data_out_0[568],u1_data_out_1[568],u1_data_out_2[568],u1_data_out_3[568],partial_product_low0[568],partial_product_low1[568],96'b0};
assign col_out_569 = {u0_col_out_569,u1_data_out_0[569],u1_data_out_1[569],u1_data_out_2[569],u1_data_out_3[569],partial_product_low0[569],partial_product_low1[569],96'b0};
assign col_out_570 = {u0_col_out_570,u1_data_out_0[570],u1_data_out_1[570],u1_data_out_2[570],u1_data_out_3[570],partial_product_low0[570],partial_product_low1[570],96'b0};
assign col_out_571 = {u0_col_out_571,u1_data_out_0[571],u1_data_out_1[571],u1_data_out_2[571],u1_data_out_3[571],partial_product_low0[571],partial_product_low1[571],96'b0};
assign col_out_572 = {u0_col_out_572,u1_data_out_0[572],u1_data_out_1[572],u1_data_out_2[572],u1_data_out_3[572],partial_product_low0[572],partial_product_low1[572],96'b0};
assign col_out_573 = {u0_col_out_573,u1_data_out_0[573],u1_data_out_1[573],u1_data_out_2[573],u1_data_out_3[573],partial_product_low0[573],partial_product_low1[573],96'b0};
assign col_out_574 = {u0_col_out_574,u1_data_out_0[574],u1_data_out_1[574],u1_data_out_2[574],u1_data_out_3[574],partial_product_low0[574],partial_product_low1[574],96'b0};
assign col_out_575 = {u0_col_out_575,u1_data_out_0[575],u1_data_out_1[575],u1_data_out_2[575],u1_data_out_3[575],partial_product_low0[575],partial_product_low1[575],96'b0};
assign col_out_576 = {u0_col_out_576,u1_data_out_0[576],u1_data_out_1[576],u1_data_out_2[576],u1_data_out_3[576],partial_product_low0[576],partial_product_low1[576],96'b0};
assign col_out_577 = {u0_col_out_577,u1_data_out_0[577],u1_data_out_1[577],u1_data_out_2[577],u1_data_out_3[577],partial_product_low0[577],partial_product_low1[577],96'b0};
assign col_out_578 = {u0_col_out_578,u1_data_out_0[578],u1_data_out_1[578],u1_data_out_2[578],u1_data_out_3[578],partial_product_low0[578],partial_product_low1[578],96'b0};
assign col_out_579 = {u0_col_out_579,u1_data_out_0[579],u1_data_out_1[579],u1_data_out_2[579],u1_data_out_3[579],partial_product_low0[579],partial_product_low1[579],96'b0};
assign col_out_580 = {u0_col_out_580,u1_data_out_0[580],u1_data_out_1[580],u1_data_out_2[580],u1_data_out_3[580],partial_product_low0[580],partial_product_low1[580],96'b0};
assign col_out_581 = {u0_col_out_581,u1_data_out_0[581],u1_data_out_1[581],u1_data_out_2[581],u1_data_out_3[581],partial_product_low0[581],partial_product_low1[581],96'b0};
assign col_out_582 = {u0_col_out_582,u1_data_out_0[582],u1_data_out_1[582],u1_data_out_2[582],u1_data_out_3[582],partial_product_low0[582],partial_product_low1[582],96'b0};
assign col_out_583 = {u0_col_out_583,u1_data_out_0[583],u1_data_out_1[583],u1_data_out_2[583],u1_data_out_3[583],partial_product_low0[583],partial_product_low1[583],96'b0};
assign col_out_584 = {u0_col_out_584,u1_data_out_0[584],u1_data_out_1[584],u1_data_out_2[584],u1_data_out_3[584],partial_product_low0[584],partial_product_low1[584],96'b0};
assign col_out_585 = {u0_col_out_585,u1_data_out_0[585],u1_data_out_1[585],u1_data_out_2[585],u1_data_out_3[585],partial_product_low0[585],partial_product_low1[585],96'b0};
assign col_out_586 = {u0_col_out_586,u1_data_out_0[586],u1_data_out_1[586],u1_data_out_2[586],u1_data_out_3[586],partial_product_low0[586],partial_product_low1[586],96'b0};
assign col_out_587 = {u0_col_out_587,u1_data_out_0[587],u1_data_out_1[587],u1_data_out_2[587],u1_data_out_3[587],partial_product_low0[587],partial_product_low1[587],96'b0};
assign col_out_588 = {u0_col_out_588,u1_data_out_0[588],u1_data_out_1[588],u1_data_out_2[588],u1_data_out_3[588],partial_product_low0[588],partial_product_low1[588],96'b0};
assign col_out_589 = {u0_col_out_589,u1_data_out_0[589],u1_data_out_1[589],u1_data_out_2[589],u1_data_out_3[589],partial_product_low0[589],partial_product_low1[589],96'b0};
assign col_out_590 = {u0_col_out_590,u1_data_out_0[590],u1_data_out_1[590],u1_data_out_2[590],u1_data_out_3[590],partial_product_low0[590],partial_product_low1[590],96'b0};
assign col_out_591 = {u0_col_out_591,u1_data_out_0[591],u1_data_out_1[591],u1_data_out_2[591],u1_data_out_3[591],partial_product_low0[591],partial_product_low1[591],96'b0};
assign col_out_592 = {u0_col_out_592,u1_data_out_0[592],u1_data_out_1[592],u1_data_out_2[592],u1_data_out_3[592],partial_product_low0[592],partial_product_low1[592],96'b0};
assign col_out_593 = {u0_col_out_593,u1_data_out_0[593],u1_data_out_1[593],u1_data_out_2[593],u1_data_out_3[593],partial_product_low0[593],partial_product_low1[593],96'b0};
assign col_out_594 = {u0_col_out_594,u1_data_out_0[594],u1_data_out_1[594],u1_data_out_2[594],u1_data_out_3[594],partial_product_low0[594],partial_product_low1[594],96'b0};
assign col_out_595 = {u0_col_out_595,u1_data_out_0[595],u1_data_out_1[595],u1_data_out_2[595],u1_data_out_3[595],partial_product_low0[595],partial_product_low1[595],96'b0};
assign col_out_596 = {u0_col_out_596,u1_data_out_0[596],u1_data_out_1[596],u1_data_out_2[596],u1_data_out_3[596],partial_product_low0[596],partial_product_low1[596],96'b0};
assign col_out_597 = {u0_col_out_597,u1_data_out_0[597],u1_data_out_1[597],u1_data_out_2[597],u1_data_out_3[597],partial_product_low0[597],partial_product_low1[597],96'b0};
assign col_out_598 = {u0_col_out_598,u1_data_out_0[598],u1_data_out_1[598],u1_data_out_2[598],u1_data_out_3[598],partial_product_low0[598],partial_product_low1[598],96'b0};
assign col_out_599 = {u0_col_out_599,u1_data_out_0[599],u1_data_out_1[599],u1_data_out_2[599],u1_data_out_3[599],partial_product_low0[599],partial_product_low1[599],96'b0};
assign col_out_600 = {u0_col_out_600,u1_data_out_0[600],u1_data_out_1[600],u1_data_out_2[600],u1_data_out_3[600],partial_product_low0[600],partial_product_low1[600],96'b0};
assign col_out_601 = {u0_col_out_601,u1_data_out_0[601],u1_data_out_1[601],u1_data_out_2[601],u1_data_out_3[601],partial_product_low0[601],partial_product_low1[601],96'b0};
assign col_out_602 = {u0_col_out_602,u1_data_out_0[602],u1_data_out_1[602],u1_data_out_2[602],u1_data_out_3[602],partial_product_low0[602],partial_product_low1[602],96'b0};
assign col_out_603 = {u0_col_out_603,u1_data_out_0[603],u1_data_out_1[603],u1_data_out_2[603],u1_data_out_3[603],partial_product_low0[603],partial_product_low1[603],96'b0};
assign col_out_604 = {u0_col_out_604,u1_data_out_0[604],u1_data_out_1[604],u1_data_out_2[604],u1_data_out_3[604],partial_product_low0[604],partial_product_low1[604],96'b0};
assign col_out_605 = {u0_col_out_605,u1_data_out_0[605],u1_data_out_1[605],u1_data_out_2[605],u1_data_out_3[605],partial_product_low0[605],partial_product_low1[605],96'b0};
assign col_out_606 = {u0_col_out_606,u1_data_out_0[606],u1_data_out_1[606],u1_data_out_2[606],u1_data_out_3[606],partial_product_low0[606],partial_product_low1[606],96'b0};
assign col_out_607 = {u0_col_out_607,u1_data_out_0[607],u1_data_out_1[607],u1_data_out_2[607],u1_data_out_3[607],partial_product_low0[607],partial_product_low1[607],96'b0};
assign col_out_608 = {u0_col_out_608,u1_data_out_0[608],u1_data_out_1[608],u1_data_out_2[608],u1_data_out_3[608],partial_product_low0[608],partial_product_low1[608],96'b0};
assign col_out_609 = {u0_col_out_609,u1_data_out_0[609],u1_data_out_1[609],u1_data_out_2[609],u1_data_out_3[609],partial_product_low0[609],partial_product_low1[609],96'b0};
assign col_out_610 = {u0_col_out_610,u1_data_out_0[610],u1_data_out_1[610],u1_data_out_2[610],u1_data_out_3[610],partial_product_low0[610],partial_product_low1[610],96'b0};
assign col_out_611 = {u0_col_out_611,u1_data_out_0[611],u1_data_out_1[611],u1_data_out_2[611],u1_data_out_3[611],partial_product_low0[611],partial_product_low1[611],96'b0};
assign col_out_612 = {u0_col_out_612,u1_data_out_0[612],u1_data_out_1[612],u1_data_out_2[612],u1_data_out_3[612],partial_product_low0[612],partial_product_low1[612],96'b0};
assign col_out_613 = {u0_col_out_613,u1_data_out_0[613],u1_data_out_1[613],u1_data_out_2[613],u1_data_out_3[613],partial_product_low0[613],partial_product_low1[613],96'b0};
assign col_out_614 = {u0_col_out_614,u1_data_out_0[614],u1_data_out_1[614],u1_data_out_2[614],u1_data_out_3[614],partial_product_low0[614],partial_product_low1[614],96'b0};
assign col_out_615 = {u0_col_out_615,u1_data_out_0[615],u1_data_out_1[615],u1_data_out_2[615],u1_data_out_3[615],partial_product_low0[615],partial_product_low1[615],96'b0};
assign col_out_616 = {u0_col_out_616,u1_data_out_0[616],u1_data_out_1[616],u1_data_out_2[616],u1_data_out_3[616],partial_product_low0[616],partial_product_low1[616],96'b0};
assign col_out_617 = {u0_col_out_617,u1_data_out_0[617],u1_data_out_1[617],u1_data_out_2[617],u1_data_out_3[617],partial_product_low0[617],partial_product_low1[617],96'b0};
assign col_out_618 = {u0_col_out_618,u1_data_out_0[618],u1_data_out_1[618],u1_data_out_2[618],u1_data_out_3[618],partial_product_low0[618],partial_product_low1[618],96'b0};
assign col_out_619 = {u0_col_out_619,u1_data_out_0[619],u1_data_out_1[619],u1_data_out_2[619],u1_data_out_3[619],partial_product_low0[619],partial_product_low1[619],96'b0};
assign col_out_620 = {u0_col_out_620,u1_data_out_0[620],u1_data_out_1[620],u1_data_out_2[620],u1_data_out_3[620],partial_product_low0[620],partial_product_low1[620],96'b0};
assign col_out_621 = {u0_col_out_621,u1_data_out_0[621],u1_data_out_1[621],u1_data_out_2[621],u1_data_out_3[621],partial_product_low0[621],partial_product_low1[621],96'b0};
assign col_out_622 = {u0_col_out_622,u1_data_out_0[622],u1_data_out_1[622],u1_data_out_2[622],u1_data_out_3[622],partial_product_low0[622],partial_product_low1[622],96'b0};
assign col_out_623 = {u0_col_out_623,u1_data_out_0[623],u1_data_out_1[623],u1_data_out_2[623],u1_data_out_3[623],partial_product_low0[623],partial_product_low1[623],96'b0};
assign col_out_624 = {u0_col_out_624,u1_data_out_0[624],u1_data_out_1[624],u1_data_out_2[624],u1_data_out_3[624],partial_product_low0[624],partial_product_low1[624],96'b0};
assign col_out_625 = {u0_col_out_625,u1_data_out_0[625],u1_data_out_1[625],u1_data_out_2[625],u1_data_out_3[625],partial_product_low0[625],partial_product_low1[625],96'b0};
assign col_out_626 = {u0_col_out_626,u1_data_out_0[626],u1_data_out_1[626],u1_data_out_2[626],u1_data_out_3[626],partial_product_low0[626],partial_product_low1[626],96'b0};
assign col_out_627 = {u0_col_out_627,u1_data_out_0[627],u1_data_out_1[627],u1_data_out_2[627],u1_data_out_3[627],partial_product_low0[627],partial_product_low1[627],96'b0};
assign col_out_628 = {u0_col_out_628,u1_data_out_0[628],u1_data_out_1[628],u1_data_out_2[628],u1_data_out_3[628],partial_product_low0[628],partial_product_low1[628],96'b0};
assign col_out_629 = {u0_col_out_629,u1_data_out_0[629],u1_data_out_1[629],u1_data_out_2[629],u1_data_out_3[629],partial_product_low0[629],partial_product_low1[629],96'b0};
assign col_out_630 = {u0_col_out_630,u1_data_out_0[630],u1_data_out_1[630],u1_data_out_2[630],u1_data_out_3[630],partial_product_low0[630],partial_product_low1[630],96'b0};
assign col_out_631 = {u0_col_out_631,u1_data_out_0[631],u1_data_out_1[631],u1_data_out_2[631],u1_data_out_3[631],partial_product_low0[631],partial_product_low1[631],96'b0};
assign col_out_632 = {u0_col_out_632,u1_data_out_0[632],u1_data_out_1[632],u1_data_out_2[632],u1_data_out_3[632],partial_product_low0[632],partial_product_low1[632],96'b0};
assign col_out_633 = {u0_col_out_633,u1_data_out_0[633],u1_data_out_1[633],u1_data_out_2[633],u1_data_out_3[633],partial_product_low0[633],partial_product_low1[633],96'b0};
assign col_out_634 = {u0_col_out_634,u1_data_out_0[634],u1_data_out_1[634],u1_data_out_2[634],u1_data_out_3[634],partial_product_low0[634],partial_product_low1[634],96'b0};
assign col_out_635 = {u0_col_out_635,u1_data_out_0[635],u1_data_out_1[635],u1_data_out_2[635],u1_data_out_3[635],partial_product_low0[635],partial_product_low1[635],96'b0};
assign col_out_636 = {u0_col_out_636,u1_data_out_0[636],u1_data_out_1[636],u1_data_out_2[636],u1_data_out_3[636],partial_product_low0[636],partial_product_low1[636],96'b0};
assign col_out_637 = {u0_col_out_637,u1_data_out_0[637],u1_data_out_1[637],u1_data_out_2[637],u1_data_out_3[637],partial_product_low0[637],partial_product_low1[637],96'b0};
assign col_out_638 = {u0_col_out_638,u1_data_out_0[638],u1_data_out_1[638],u1_data_out_2[638],u1_data_out_3[638],partial_product_low0[638],partial_product_low1[638],96'b0};
assign col_out_639 = {u0_col_out_639,u1_data_out_0[639],u1_data_out_1[639],u1_data_out_2[639],u1_data_out_3[639],partial_product_low0[639],partial_product_low1[639],96'b0};
assign col_out_640 = {u0_col_out_640,u1_data_out_0[640],u1_data_out_1[640],u1_data_out_2[640],u1_data_out_3[640],partial_product_low0[640],partial_product_low1[640],96'b0};
assign col_out_641 = {u0_col_out_641,u1_data_out_0[641],u1_data_out_1[641],u1_data_out_2[641],u1_data_out_3[641],partial_product_low0[641],partial_product_low1[641],96'b0};
assign col_out_642 = {u0_col_out_642,u1_data_out_0[642],u1_data_out_1[642],u1_data_out_2[642],u1_data_out_3[642],partial_product_low0[642],partial_product_low1[642],96'b0};
assign col_out_643 = {u0_col_out_643,u1_data_out_0[643],u1_data_out_1[643],u1_data_out_2[643],u1_data_out_3[643],partial_product_low0[643],partial_product_low1[643],96'b0};
assign col_out_644 = {u0_col_out_644,u1_data_out_0[644],u1_data_out_1[644],u1_data_out_2[644],u1_data_out_3[644],partial_product_low0[644],partial_product_low1[644],96'b0};
assign col_out_645 = {u0_col_out_645,u1_data_out_0[645],u1_data_out_1[645],u1_data_out_2[645],u1_data_out_3[645],partial_product_low0[645],partial_product_low1[645],96'b0};
assign col_out_646 = {u0_col_out_646,u1_data_out_0[646],u1_data_out_1[646],u1_data_out_2[646],u1_data_out_3[646],partial_product_low0[646],partial_product_low1[646],96'b0};
assign col_out_647 = {u0_col_out_647,u1_data_out_0[647],u1_data_out_1[647],u1_data_out_2[647],u1_data_out_3[647],partial_product_low0[647],partial_product_low1[647],96'b0};
assign col_out_648 = {u0_col_out_648,u1_data_out_0[648],u1_data_out_1[648],u1_data_out_2[648],u1_data_out_3[648],partial_product_low0[648],partial_product_low1[648],96'b0};
assign col_out_649 = {u0_col_out_649,u1_data_out_0[649],u1_data_out_1[649],u1_data_out_2[649],u1_data_out_3[649],partial_product_low0[649],partial_product_low1[649],96'b0};
assign col_out_650 = {u0_col_out_650,u1_data_out_0[650],u1_data_out_1[650],u1_data_out_2[650],u1_data_out_3[650],partial_product_low0[650],partial_product_low1[650],96'b0};
assign col_out_651 = {u0_col_out_651,u1_data_out_0[651],u1_data_out_1[651],u1_data_out_2[651],u1_data_out_3[651],partial_product_low0[651],partial_product_low1[651],96'b0};
assign col_out_652 = {u0_col_out_652,u1_data_out_0[652],u1_data_out_1[652],u1_data_out_2[652],u1_data_out_3[652],partial_product_low0[652],partial_product_low1[652],96'b0};
assign col_out_653 = {u0_col_out_653,u1_data_out_0[653],u1_data_out_1[653],u1_data_out_2[653],u1_data_out_3[653],partial_product_low0[653],partial_product_low1[653],96'b0};
assign col_out_654 = {u0_col_out_654,u1_data_out_0[654],u1_data_out_1[654],u1_data_out_2[654],u1_data_out_3[654],partial_product_low0[654],partial_product_low1[654],96'b0};
assign col_out_655 = {u0_col_out_655,u1_data_out_0[655],u1_data_out_1[655],u1_data_out_2[655],u1_data_out_3[655],partial_product_low0[655],partial_product_low1[655],96'b0};
assign col_out_656 = {u0_col_out_656,u1_data_out_0[656],u1_data_out_1[656],u1_data_out_2[656],u1_data_out_3[656],partial_product_low0[656],partial_product_low1[656],96'b0};
assign col_out_657 = {u0_col_out_657,u1_data_out_0[657],u1_data_out_1[657],u1_data_out_2[657],u1_data_out_3[657],partial_product_low0[657],partial_product_low1[657],96'b0};
assign col_out_658 = {u0_col_out_658,u1_data_out_0[658],u1_data_out_1[658],u1_data_out_2[658],u1_data_out_3[658],partial_product_low0[658],partial_product_low1[658],96'b0};
assign col_out_659 = {u0_col_out_659,u1_data_out_0[659],u1_data_out_1[659],u1_data_out_2[659],u1_data_out_3[659],partial_product_low0[659],partial_product_low1[659],96'b0};
assign col_out_660 = {u0_col_out_660,u1_data_out_0[660],u1_data_out_1[660],u1_data_out_2[660],u1_data_out_3[660],partial_product_low0[660],partial_product_low1[660],96'b0};
assign col_out_661 = {u0_col_out_661,u1_data_out_0[661],u1_data_out_1[661],u1_data_out_2[661],u1_data_out_3[661],partial_product_low0[661],partial_product_low1[661],96'b0};
assign col_out_662 = {u0_col_out_662,u1_data_out_0[662],u1_data_out_1[662],u1_data_out_2[662],u1_data_out_3[662],partial_product_low0[662],partial_product_low1[662],96'b0};
assign col_out_663 = {u0_col_out_663,u1_data_out_0[663],u1_data_out_1[663],u1_data_out_2[663],u1_data_out_3[663],partial_product_low0[663],partial_product_low1[663],96'b0};
assign col_out_664 = {u0_col_out_664,u1_data_out_0[664],u1_data_out_1[664],u1_data_out_2[664],u1_data_out_3[664],partial_product_low0[664],partial_product_low1[664],96'b0};
assign col_out_665 = {u0_col_out_665,u1_data_out_0[665],u1_data_out_1[665],u1_data_out_2[665],u1_data_out_3[665],partial_product_low0[665],partial_product_low1[665],96'b0};
assign col_out_666 = {u0_col_out_666,u1_data_out_0[666],u1_data_out_1[666],u1_data_out_2[666],u1_data_out_3[666],partial_product_low0[666],partial_product_low1[666],96'b0};
assign col_out_667 = {u0_col_out_667,u1_data_out_0[667],u1_data_out_1[667],u1_data_out_2[667],u1_data_out_3[667],partial_product_low0[667],partial_product_low1[667],96'b0};
assign col_out_668 = {u0_col_out_668,u1_data_out_0[668],u1_data_out_1[668],u1_data_out_2[668],u1_data_out_3[668],partial_product_low0[668],partial_product_low1[668],96'b0};
assign col_out_669 = {u0_col_out_669,u1_data_out_0[669],u1_data_out_1[669],u1_data_out_2[669],u1_data_out_3[669],partial_product_low0[669],partial_product_low1[669],96'b0};
assign col_out_670 = {u0_col_out_670,u1_data_out_0[670],u1_data_out_1[670],u1_data_out_2[670],u1_data_out_3[670],partial_product_low0[670],partial_product_low1[670],96'b0};
assign col_out_671 = {u0_col_out_671,u1_data_out_0[671],u1_data_out_1[671],u1_data_out_2[671],u1_data_out_3[671],partial_product_low0[671],partial_product_low1[671],96'b0};
assign col_out_672 = {u0_col_out_672,u1_data_out_0[672],u1_data_out_1[672],u1_data_out_2[672],u1_data_out_3[672],partial_product_low0[672],partial_product_low1[672],96'b0};
assign col_out_673 = {u0_col_out_673,u1_data_out_0[673],u1_data_out_1[673],u1_data_out_2[673],u1_data_out_3[673],partial_product_low0[673],partial_product_low1[673],96'b0};
assign col_out_674 = {u0_col_out_674,u1_data_out_0[674],u1_data_out_1[674],u1_data_out_2[674],u1_data_out_3[674],partial_product_low0[674],partial_product_low1[674],96'b0};
assign col_out_675 = {u0_col_out_675,u1_data_out_0[675],u1_data_out_1[675],u1_data_out_2[675],u1_data_out_3[675],partial_product_low0[675],partial_product_low1[675],96'b0};
assign col_out_676 = {u0_col_out_676,u1_data_out_0[676],u1_data_out_1[676],u1_data_out_2[676],u1_data_out_3[676],partial_product_low0[676],partial_product_low1[676],96'b0};
assign col_out_677 = {u0_col_out_677,u1_data_out_0[677],u1_data_out_1[677],u1_data_out_2[677],u1_data_out_3[677],partial_product_low0[677],partial_product_low1[677],96'b0};
assign col_out_678 = {u0_col_out_678,u1_data_out_0[678],u1_data_out_1[678],u1_data_out_2[678],u1_data_out_3[678],partial_product_low0[678],partial_product_low1[678],96'b0};
assign col_out_679 = {u0_col_out_679,u1_data_out_0[679],u1_data_out_1[679],u1_data_out_2[679],u1_data_out_3[679],partial_product_low0[679],partial_product_low1[679],96'b0};
assign col_out_680 = {u0_col_out_680,u1_data_out_0[680],u1_data_out_1[680],u1_data_out_2[680],u1_data_out_3[680],partial_product_low0[680],partial_product_low1[680],96'b0};
assign col_out_681 = {u0_col_out_681,u1_data_out_0[681],u1_data_out_1[681],u1_data_out_2[681],u1_data_out_3[681],partial_product_low0[681],partial_product_low1[681],96'b0};
assign col_out_682 = {u0_col_out_682,u1_data_out_0[682],u1_data_out_1[682],u1_data_out_2[682],u1_data_out_3[682],partial_product_low0[682],partial_product_low1[682],96'b0};
assign col_out_683 = {u0_col_out_683,u1_data_out_0[683],u1_data_out_1[683],u1_data_out_2[683],u1_data_out_3[683],partial_product_low0[683],partial_product_low1[683],96'b0};
assign col_out_684 = {u0_col_out_684,u1_data_out_0[684],u1_data_out_1[684],u1_data_out_2[684],u1_data_out_3[684],partial_product_low0[684],partial_product_low1[684],96'b0};
assign col_out_685 = {u0_col_out_685,u1_data_out_0[685],u1_data_out_1[685],u1_data_out_2[685],u1_data_out_3[685],partial_product_low0[685],partial_product_low1[685],96'b0};
assign col_out_686 = {u0_col_out_686,u1_data_out_0[686],u1_data_out_1[686],u1_data_out_2[686],u1_data_out_3[686],partial_product_low0[686],partial_product_low1[686],96'b0};
assign col_out_687 = {u0_col_out_687,u1_data_out_0[687],u1_data_out_1[687],u1_data_out_2[687],u1_data_out_3[687],partial_product_low0[687],partial_product_low1[687],96'b0};
assign col_out_688 = {u0_col_out_688,u1_data_out_0[688],u1_data_out_1[688],u1_data_out_2[688],u1_data_out_3[688],partial_product_low0[688],partial_product_low1[688],96'b0};
assign col_out_689 = {u0_col_out_689,u1_data_out_0[689],u1_data_out_1[689],u1_data_out_2[689],u1_data_out_3[689],partial_product_low0[689],partial_product_low1[689],96'b0};
assign col_out_690 = {u0_col_out_690,u1_data_out_0[690],u1_data_out_1[690],u1_data_out_2[690],u1_data_out_3[690],partial_product_low0[690],partial_product_low1[690],96'b0};
assign col_out_691 = {u0_col_out_691,u1_data_out_0[691],u1_data_out_1[691],u1_data_out_2[691],u1_data_out_3[691],partial_product_low0[691],partial_product_low1[691],96'b0};
assign col_out_692 = {u0_col_out_692,u1_data_out_0[692],u1_data_out_1[692],u1_data_out_2[692],u1_data_out_3[692],partial_product_low0[692],partial_product_low1[692],96'b0};
assign col_out_693 = {u0_col_out_693,u1_data_out_0[693],u1_data_out_1[693],u1_data_out_2[693],u1_data_out_3[693],partial_product_low0[693],partial_product_low1[693],96'b0};
assign col_out_694 = {u0_col_out_694,u1_data_out_0[694],u1_data_out_1[694],u1_data_out_2[694],u1_data_out_3[694],partial_product_low0[694],partial_product_low1[694],96'b0};
assign col_out_695 = {u0_col_out_695,u1_data_out_0[695],u1_data_out_1[695],u1_data_out_2[695],u1_data_out_3[695],partial_product_low0[695],partial_product_low1[695],96'b0};
assign col_out_696 = {u0_col_out_696,u1_data_out_0[696],u1_data_out_1[696],u1_data_out_2[696],u1_data_out_3[696],partial_product_low0[696],partial_product_low1[696],96'b0};
assign col_out_697 = {u0_col_out_697,u1_data_out_0[697],u1_data_out_1[697],u1_data_out_2[697],u1_data_out_3[697],partial_product_low0[697],partial_product_low1[697],96'b0};
assign col_out_698 = {u0_col_out_698,u1_data_out_0[698],u1_data_out_1[698],u1_data_out_2[698],u1_data_out_3[698],partial_product_low0[698],partial_product_low1[698],96'b0};
assign col_out_699 = {u0_col_out_699,u1_data_out_0[699],u1_data_out_1[699],u1_data_out_2[699],u1_data_out_3[699],partial_product_low0[699],partial_product_low1[699],96'b0};
assign col_out_700 = {u0_col_out_700,u1_data_out_0[700],u1_data_out_1[700],u1_data_out_2[700],u1_data_out_3[700],partial_product_low0[700],partial_product_low1[700],96'b0};
assign col_out_701 = {u0_col_out_701,u1_data_out_0[701],u1_data_out_1[701],u1_data_out_2[701],u1_data_out_3[701],partial_product_low0[701],partial_product_low1[701],96'b0};
assign col_out_702 = {u0_col_out_702,u1_data_out_0[702],u1_data_out_1[702],u1_data_out_2[702],u1_data_out_3[702],partial_product_low0[702],partial_product_low1[702],96'b0};
assign col_out_703 = {u0_col_out_703,u1_data_out_0[703],u1_data_out_1[703],u1_data_out_2[703],u1_data_out_3[703],partial_product_low0[703],partial_product_low1[703],96'b0};
assign col_out_704 = {u0_col_out_704,u1_data_out_0[704],u1_data_out_1[704],u1_data_out_2[704],u1_data_out_3[704],partial_product_low0[704],partial_product_low1[704],96'b0};
assign col_out_705 = {u0_col_out_705,u1_data_out_0[705],u1_data_out_1[705],u1_data_out_2[705],u1_data_out_3[705],partial_product_low0[705],partial_product_low1[705],96'b0};
assign col_out_706 = {u0_col_out_706,u1_data_out_0[706],u1_data_out_1[706],u1_data_out_2[706],u1_data_out_3[706],partial_product_low0[706],partial_product_low1[706],96'b0};
assign col_out_707 = {u0_col_out_707,u1_data_out_0[707],u1_data_out_1[707],u1_data_out_2[707],u1_data_out_3[707],partial_product_low0[707],partial_product_low1[707],96'b0};
assign col_out_708 = {u0_col_out_708,u1_data_out_0[708],u1_data_out_1[708],u1_data_out_2[708],u1_data_out_3[708],partial_product_low0[708],partial_product_low1[708],96'b0};
assign col_out_709 = {u0_col_out_709,u1_data_out_0[709],u1_data_out_1[709],u1_data_out_2[709],u1_data_out_3[709],partial_product_low0[709],partial_product_low1[709],96'b0};
assign col_out_710 = {u0_col_out_710,u1_data_out_0[710],u1_data_out_1[710],u1_data_out_2[710],u1_data_out_3[710],partial_product_low0[710],partial_product_low1[710],96'b0};
assign col_out_711 = {u0_col_out_711,u1_data_out_0[711],u1_data_out_1[711],u1_data_out_2[711],u1_data_out_3[711],partial_product_low0[711],partial_product_low1[711],96'b0};
assign col_out_712 = {u0_col_out_712,u1_data_out_0[712],u1_data_out_1[712],u1_data_out_2[712],u1_data_out_3[712],partial_product_low0[712],partial_product_low1[712],96'b0};
assign col_out_713 = {u0_col_out_713,u1_data_out_0[713],u1_data_out_1[713],u1_data_out_2[713],u1_data_out_3[713],partial_product_low0[713],partial_product_low1[713],96'b0};
assign col_out_714 = {u0_col_out_714,u1_data_out_0[714],u1_data_out_1[714],u1_data_out_2[714],u1_data_out_3[714],partial_product_low0[714],partial_product_low1[714],96'b0};
assign col_out_715 = {u0_col_out_715,u1_data_out_0[715],u1_data_out_1[715],u1_data_out_2[715],u1_data_out_3[715],partial_product_low0[715],partial_product_low1[715],96'b0};
assign col_out_716 = {u0_col_out_716,u1_data_out_0[716],u1_data_out_1[716],u1_data_out_2[716],u1_data_out_3[716],partial_product_low0[716],partial_product_low1[716],96'b0};
assign col_out_717 = {u0_col_out_717,u1_data_out_0[717],u1_data_out_1[717],u1_data_out_2[717],u1_data_out_3[717],partial_product_low0[717],partial_product_low1[717],96'b0};
assign col_out_718 = {u0_col_out_718,u1_data_out_0[718],u1_data_out_1[718],u1_data_out_2[718],u1_data_out_3[718],partial_product_low0[718],partial_product_low1[718],96'b0};
assign col_out_719 = {u0_col_out_719,u1_data_out_0[719],u1_data_out_1[719],u1_data_out_2[719],u1_data_out_3[719],partial_product_low0[719],partial_product_low1[719],96'b0};
assign col_out_720 = {u0_col_out_720,u1_data_out_0[720],u1_data_out_1[720],u1_data_out_2[720],u1_data_out_3[720],partial_product_low0[720],partial_product_low1[720],96'b0};
assign col_out_721 = {u0_col_out_721,u1_data_out_0[721],u1_data_out_1[721],u1_data_out_2[721],u1_data_out_3[721],partial_product_low0[721],partial_product_low1[721],96'b0};
assign col_out_722 = {u0_col_out_722,u1_data_out_0[722],u1_data_out_1[722],u1_data_out_2[722],u1_data_out_3[722],partial_product_low0[722],partial_product_low1[722],96'b0};
assign col_out_723 = {u0_col_out_723,u1_data_out_0[723],u1_data_out_1[723],u1_data_out_2[723],u1_data_out_3[723],partial_product_low0[723],partial_product_low1[723],96'b0};
assign col_out_724 = {u0_col_out_724,u1_data_out_0[724],u1_data_out_1[724],u1_data_out_2[724],u1_data_out_3[724],partial_product_low0[724],partial_product_low1[724],96'b0};
assign col_out_725 = {u0_col_out_725,u1_data_out_0[725],u1_data_out_1[725],u1_data_out_2[725],u1_data_out_3[725],partial_product_low0[725],partial_product_low1[725],96'b0};
assign col_out_726 = {u0_col_out_726,u1_data_out_0[726],u1_data_out_1[726],u1_data_out_2[726],u1_data_out_3[726],partial_product_low0[726],partial_product_low1[726],96'b0};
assign col_out_727 = {u0_col_out_727,u1_data_out_0[727],u1_data_out_1[727],u1_data_out_2[727],u1_data_out_3[727],partial_product_low0[727],partial_product_low1[727],96'b0};
assign col_out_728 = {u0_col_out_728,u1_data_out_0[728],u1_data_out_1[728],u1_data_out_2[728],u1_data_out_3[728],partial_product_low0[728],partial_product_low1[728],96'b0};
assign col_out_729 = {u0_col_out_729,u1_data_out_0[729],u1_data_out_1[729],u1_data_out_2[729],u1_data_out_3[729],partial_product_low0[729],partial_product_low1[729],96'b0};
assign col_out_730 = {u0_col_out_730,u1_data_out_0[730],u1_data_out_1[730],u1_data_out_2[730],u1_data_out_3[730],partial_product_low0[730],partial_product_low1[730],96'b0};
assign col_out_731 = {u0_col_out_731,u1_data_out_0[731],u1_data_out_1[731],u1_data_out_2[731],u1_data_out_3[731],partial_product_low0[731],partial_product_low1[731],96'b0};
assign col_out_732 = {u0_col_out_732,u1_data_out_0[732],u1_data_out_1[732],u1_data_out_2[732],u1_data_out_3[732],partial_product_low0[732],partial_product_low1[732],96'b0};
assign col_out_733 = {u0_col_out_733,u1_data_out_0[733],u1_data_out_1[733],u1_data_out_2[733],u1_data_out_3[733],partial_product_low0[733],partial_product_low1[733],96'b0};
assign col_out_734 = {u0_col_out_734,u1_data_out_0[734],u1_data_out_1[734],u1_data_out_2[734],u1_data_out_3[734],partial_product_low0[734],partial_product_low1[734],96'b0};
assign col_out_735 = {u0_col_out_735,u1_data_out_0[735],u1_data_out_1[735],u1_data_out_2[735],u1_data_out_3[735],partial_product_low0[735],partial_product_low1[735],96'b0};
assign col_out_736 = {u0_col_out_736,u1_data_out_0[736],u1_data_out_1[736],u1_data_out_2[736],u1_data_out_3[736],partial_product_low0[736],partial_product_low1[736],96'b0};
assign col_out_737 = {u0_col_out_737,u1_data_out_0[737],u1_data_out_1[737],u1_data_out_2[737],u1_data_out_3[737],partial_product_low0[737],partial_product_low1[737],96'b0};
assign col_out_738 = {u0_col_out_738,u1_data_out_0[738],u1_data_out_1[738],u1_data_out_2[738],u1_data_out_3[738],partial_product_low0[738],partial_product_low1[738],96'b0};
assign col_out_739 = {u0_col_out_739,u1_data_out_0[739],u1_data_out_1[739],u1_data_out_2[739],u1_data_out_3[739],partial_product_low0[739],partial_product_low1[739],96'b0};
assign col_out_740 = {u0_col_out_740,u1_data_out_0[740],u1_data_out_1[740],u1_data_out_2[740],u1_data_out_3[740],partial_product_low0[740],partial_product_low1[740],96'b0};
assign col_out_741 = {u0_col_out_741,u1_data_out_0[741],u1_data_out_1[741],u1_data_out_2[741],u1_data_out_3[741],partial_product_low0[741],partial_product_low1[741],96'b0};
assign col_out_742 = {u0_col_out_742,u1_data_out_0[742],u1_data_out_1[742],u1_data_out_2[742],u1_data_out_3[742],partial_product_low0[742],partial_product_low1[742],96'b0};
assign col_out_743 = {u0_col_out_743,u1_data_out_0[743],u1_data_out_1[743],u1_data_out_2[743],u1_data_out_3[743],partial_product_low0[743],partial_product_low1[743],96'b0};
assign col_out_744 = {u0_col_out_744,u1_data_out_0[744],u1_data_out_1[744],u1_data_out_2[744],u1_data_out_3[744],partial_product_low0[744],partial_product_low1[744],96'b0};
assign col_out_745 = {u0_col_out_745,u1_data_out_0[745],u1_data_out_1[745],u1_data_out_2[745],u1_data_out_3[745],partial_product_low0[745],partial_product_low1[745],96'b0};
assign col_out_746 = {u0_col_out_746,u1_data_out_0[746],u1_data_out_1[746],u1_data_out_2[746],u1_data_out_3[746],partial_product_low0[746],partial_product_low1[746],96'b0};
assign col_out_747 = {u0_col_out_747,u1_data_out_0[747],u1_data_out_1[747],u1_data_out_2[747],u1_data_out_3[747],partial_product_low0[747],partial_product_low1[747],96'b0};
assign col_out_748 = {u0_col_out_748,u1_data_out_0[748],u1_data_out_1[748],u1_data_out_2[748],u1_data_out_3[748],partial_product_low0[748],partial_product_low1[748],96'b0};
assign col_out_749 = {u0_col_out_749,u1_data_out_0[749],u1_data_out_1[749],u1_data_out_2[749],u1_data_out_3[749],partial_product_low0[749],partial_product_low1[749],96'b0};
assign col_out_750 = {u0_col_out_750,u1_data_out_0[750],u1_data_out_1[750],u1_data_out_2[750],u1_data_out_3[750],partial_product_low0[750],partial_product_low1[750],96'b0};
assign col_out_751 = {u0_col_out_751,u1_data_out_0[751],u1_data_out_1[751],u1_data_out_2[751],u1_data_out_3[751],partial_product_low0[751],partial_product_low1[751],96'b0};
assign col_out_752 = {u0_col_out_752,u1_data_out_0[752],u1_data_out_1[752],u1_data_out_2[752],u1_data_out_3[752],partial_product_low0[752],partial_product_low1[752],96'b0};
assign col_out_753 = {u0_col_out_753,u1_data_out_0[753],u1_data_out_1[753],u1_data_out_2[753],u1_data_out_3[753],partial_product_low0[753],partial_product_low1[753],96'b0};
assign col_out_754 = {u0_col_out_754,u1_data_out_0[754],u1_data_out_1[754],u1_data_out_2[754],u1_data_out_3[754],partial_product_low0[754],partial_product_low1[754],96'b0};
assign col_out_755 = {u0_col_out_755,u1_data_out_0[755],u1_data_out_1[755],u1_data_out_2[755],u1_data_out_3[755],partial_product_low0[755],partial_product_low1[755],96'b0};
assign col_out_756 = {u0_col_out_756,u1_data_out_0[756],u1_data_out_1[756],u1_data_out_2[756],u1_data_out_3[756],partial_product_low0[756],partial_product_low1[756],96'b0};
assign col_out_757 = {u0_col_out_757,u1_data_out_0[757],u1_data_out_1[757],u1_data_out_2[757],u1_data_out_3[757],partial_product_low0[757],partial_product_low1[757],96'b0};
assign col_out_758 = {u0_col_out_758,u1_data_out_0[758],u1_data_out_1[758],u1_data_out_2[758],u1_data_out_3[758],partial_product_low0[758],partial_product_low1[758],96'b0};
assign col_out_759 = {u0_col_out_759,u1_data_out_0[759],u1_data_out_1[759],u1_data_out_2[759],u1_data_out_3[759],partial_product_low0[759],partial_product_low1[759],96'b0};
assign col_out_760 = {u0_col_out_760,u1_data_out_0[760],u1_data_out_1[760],u1_data_out_2[760],u1_data_out_3[760],partial_product_low0[760],partial_product_low1[760],96'b0};
assign col_out_761 = {u0_col_out_761,u1_data_out_0[761],u1_data_out_1[761],u1_data_out_2[761],u1_data_out_3[761],partial_product_low0[761],partial_product_low1[761],96'b0};
assign col_out_762 = {u0_col_out_762,u1_data_out_0[762],u1_data_out_1[762],u1_data_out_2[762],u1_data_out_3[762],partial_product_low0[762],partial_product_low1[762],96'b0};
assign col_out_763 = {u0_col_out_763,u1_data_out_0[763],u1_data_out_1[763],u1_data_out_2[763],u1_data_out_3[763],partial_product_low0[763],partial_product_low1[763],96'b0};
assign col_out_764 = {u0_col_out_764,u1_data_out_0[764],u1_data_out_1[764],u1_data_out_2[764],u1_data_out_3[764],partial_product_low0[764],partial_product_low1[764],96'b0};
assign col_out_765 = {u0_col_out_765,u1_data_out_0[765],u1_data_out_1[765],u1_data_out_2[765],u1_data_out_3[765],partial_product_low0[765],partial_product_low1[765],96'b0};
assign col_out_766 = {u0_col_out_766,u1_data_out_0[766],u1_data_out_1[766],u1_data_out_2[766],u1_data_out_3[766],partial_product_low0[766],partial_product_low1[766],96'b0};
assign col_out_767 = {u0_col_out_767,u1_data_out_0[767],u1_data_out_1[767],u1_data_out_2[767],u1_data_out_3[767],partial_product_low0[767],partial_product_low1[767],96'b0};
assign col_out_768 = {u0_col_out_768,u1_data_out_0[768],u1_data_out_1[768],u1_data_out_2[768],u1_data_out_3[768],partial_product_low0[768],partial_product_low1[768],96'b0};
assign col_out_769 = {u0_col_out_769,u1_data_out_0[769],u1_data_out_1[769],u1_data_out_2[769],u1_data_out_3[769],partial_product_low0[769],partial_product_low1[769],96'b0};
assign col_out_770 = {u0_col_out_770,u1_data_out_0[770],u1_data_out_1[770],u1_data_out_2[770],u1_data_out_3[770],partial_product_low0[770],partial_product_low1[770],96'b0};
assign col_out_771 = {u0_col_out_771,u1_data_out_0[771],u1_data_out_1[771],u1_data_out_2[771],u1_data_out_3[771],partial_product_low0[771],partial_product_low1[771],96'b0};
assign col_out_772 = {u0_col_out_772,u1_data_out_0[772],u1_data_out_1[772],u1_data_out_2[772],u1_data_out_3[772],partial_product_low0[772],partial_product_low1[772],96'b0};
assign col_out_773 = {u0_col_out_773,u1_data_out_0[773],u1_data_out_1[773],u1_data_out_2[773],u1_data_out_3[773],partial_product_low0[773],partial_product_low1[773],96'b0};
assign col_out_774 = {u0_col_out_774,u1_data_out_0[774],u1_data_out_1[774],u1_data_out_2[774],u1_data_out_3[774],partial_product_low0[774],partial_product_low1[774],96'b0};
assign col_out_775 = {u0_col_out_775,u1_data_out_0[775],u1_data_out_1[775],u1_data_out_2[775],u1_data_out_3[775],partial_product_low0[775],partial_product_low1[775],96'b0};
assign col_out_776 = {u0_col_out_776,u1_data_out_0[776],u1_data_out_1[776],u1_data_out_2[776],u1_data_out_3[776],partial_product_low0[776],partial_product_low1[776],96'b0};
assign col_out_777 = {u0_col_out_777,u1_data_out_0[777],u1_data_out_1[777],u1_data_out_2[777],u1_data_out_3[777],partial_product_low0[777],partial_product_low1[777],96'b0};
assign col_out_778 = {u0_col_out_778,u1_data_out_0[778],u1_data_out_1[778],u1_data_out_2[778],u1_data_out_3[778],partial_product_low0[778],partial_product_low1[778],96'b0};
assign col_out_779 = {u0_col_out_779,u1_data_out_0[779],u1_data_out_1[779],u1_data_out_2[779],u1_data_out_3[779],partial_product_low0[779],partial_product_low1[779],96'b0};
assign col_out_780 = {u0_col_out_780,u1_data_out_0[780],u1_data_out_1[780],u1_data_out_2[780],u1_data_out_3[780],partial_product_low0[780],partial_product_low1[780],96'b0};
assign col_out_781 = {u0_col_out_781,u1_data_out_0[781],u1_data_out_1[781],u1_data_out_2[781],u1_data_out_3[781],partial_product_low0[781],partial_product_low1[781],96'b0};
assign col_out_782 = {u0_col_out_782,u1_data_out_0[782],u1_data_out_1[782],u1_data_out_2[782],u1_data_out_3[782],partial_product_low0[782],partial_product_low1[782],96'b0};
assign col_out_783 = {u0_col_out_783,u1_data_out_0[783],u1_data_out_1[783],u1_data_out_2[783],u1_data_out_3[783],partial_product_low0[783],partial_product_low1[783],96'b0};
assign col_out_784 = {u0_col_out_784,u1_data_out_0[784],u1_data_out_1[784],u1_data_out_2[784],u1_data_out_3[784],partial_product_low0[784],partial_product_low1[784],96'b0};
assign col_out_785 = {u0_col_out_785,u1_data_out_0[785],u1_data_out_1[785],u1_data_out_2[785],u1_data_out_3[785],partial_product_low0[785],partial_product_low1[785],96'b0};
assign col_out_786 = {u0_col_out_786,u1_data_out_0[786],u1_data_out_1[786],u1_data_out_2[786],u1_data_out_3[786],partial_product_low0[786],partial_product_low1[786],96'b0};
assign col_out_787 = {u0_col_out_787,u1_data_out_0[787],u1_data_out_1[787],u1_data_out_2[787],u1_data_out_3[787],partial_product_low0[787],partial_product_low1[787],96'b0};
assign col_out_788 = {u0_col_out_788,u1_data_out_0[788],u1_data_out_1[788],u1_data_out_2[788],u1_data_out_3[788],partial_product_low0[788],partial_product_low1[788],96'b0};
assign col_out_789 = {u0_col_out_789,u1_data_out_0[789],u1_data_out_1[789],u1_data_out_2[789],u1_data_out_3[789],partial_product_low0[789],partial_product_low1[789],96'b0};
assign col_out_790 = {u0_col_out_790,u1_data_out_0[790],u1_data_out_1[790],u1_data_out_2[790],u1_data_out_3[790],partial_product_low0[790],partial_product_low1[790],96'b0};
assign col_out_791 = {u0_col_out_791,u1_data_out_0[791],u1_data_out_1[791],u1_data_out_2[791],u1_data_out_3[791],partial_product_low0[791],partial_product_low1[791],96'b0};
assign col_out_792 = {u0_col_out_792,u1_data_out_0[792],u1_data_out_1[792],u1_data_out_2[792],u1_data_out_3[792],partial_product_low0[792],partial_product_low1[792],96'b0};
assign col_out_793 = {u0_col_out_793,u1_data_out_0[793],u1_data_out_1[793],u1_data_out_2[793],u1_data_out_3[793],partial_product_low0[793],partial_product_low1[793],96'b0};
assign col_out_794 = {u0_col_out_794,u1_data_out_0[794],u1_data_out_1[794],u1_data_out_2[794],u1_data_out_3[794],partial_product_low0[794],partial_product_low1[794],96'b0};
assign col_out_795 = {u0_col_out_795,u1_data_out_0[795],u1_data_out_1[795],u1_data_out_2[795],u1_data_out_3[795],partial_product_low0[795],partial_product_low1[795],96'b0};
assign col_out_796 = {u0_col_out_796,u1_data_out_0[796],u1_data_out_1[796],u1_data_out_2[796],u1_data_out_3[796],partial_product_low0[796],partial_product_low1[796],96'b0};
assign col_out_797 = {u0_col_out_797,u1_data_out_0[797],u1_data_out_1[797],u1_data_out_2[797],u1_data_out_3[797],partial_product_low0[797],partial_product_low1[797],96'b0};
assign col_out_798 = {u0_col_out_798,u1_data_out_0[798],u1_data_out_1[798],u1_data_out_2[798],u1_data_out_3[798],partial_product_low0[798],partial_product_low1[798],96'b0};
assign col_out_799 = {u0_col_out_799,u1_data_out_0[799],u1_data_out_1[799],u1_data_out_2[799],u1_data_out_3[799],partial_product_low0[799],partial_product_low1[799],96'b0};
assign col_out_800 = {u0_col_out_800,u1_data_out_0[800],u1_data_out_1[800],u1_data_out_2[800],u1_data_out_3[800],partial_product_low0[800],partial_product_low1[800],96'b0};
assign col_out_801 = {u0_col_out_801,u1_data_out_0[801],u1_data_out_1[801],u1_data_out_2[801],u1_data_out_3[801],partial_product_low0[801],partial_product_low1[801],96'b0};
assign col_out_802 = {u0_col_out_802,u1_data_out_0[802],u1_data_out_1[802],u1_data_out_2[802],u1_data_out_3[802],partial_product_low0[802],partial_product_low1[802],96'b0};
assign col_out_803 = {u0_col_out_803,u1_data_out_0[803],u1_data_out_1[803],u1_data_out_2[803],u1_data_out_3[803],partial_product_low0[803],partial_product_low1[803],96'b0};
assign col_out_804 = {u0_col_out_804,u1_data_out_0[804],u1_data_out_1[804],u1_data_out_2[804],u1_data_out_3[804],partial_product_low0[804],partial_product_low1[804],96'b0};
assign col_out_805 = {u0_col_out_805,u1_data_out_0[805],u1_data_out_1[805],u1_data_out_2[805],u1_data_out_3[805],partial_product_low0[805],partial_product_low1[805],96'b0};
assign col_out_806 = {u0_col_out_806,u1_data_out_0[806],u1_data_out_1[806],u1_data_out_2[806],u1_data_out_3[806],partial_product_low0[806],partial_product_low1[806],96'b0};
assign col_out_807 = {u0_col_out_807,u1_data_out_0[807],u1_data_out_1[807],u1_data_out_2[807],u1_data_out_3[807],partial_product_low0[807],partial_product_low1[807],96'b0};
assign col_out_808 = {u0_col_out_808,u1_data_out_0[808],u1_data_out_1[808],u1_data_out_2[808],u1_data_out_3[808],partial_product_low0[808],partial_product_low1[808],96'b0};
assign col_out_809 = {u0_col_out_809,u1_data_out_0[809],u1_data_out_1[809],u1_data_out_2[809],u1_data_out_3[809],partial_product_low0[809],partial_product_low1[809],96'b0};
assign col_out_810 = {u0_col_out_810,u1_data_out_0[810],u1_data_out_1[810],u1_data_out_2[810],u1_data_out_3[810],partial_product_low0[810],partial_product_low1[810],96'b0};
assign col_out_811 = {u0_col_out_811,u1_data_out_0[811],u1_data_out_1[811],u1_data_out_2[811],u1_data_out_3[811],partial_product_low0[811],partial_product_low1[811],96'b0};
assign col_out_812 = {u0_col_out_812,u1_data_out_0[812],u1_data_out_1[812],u1_data_out_2[812],u1_data_out_3[812],partial_product_low0[812],partial_product_low1[812],96'b0};
assign col_out_813 = {u0_col_out_813,u1_data_out_0[813],u1_data_out_1[813],u1_data_out_2[813],u1_data_out_3[813],partial_product_low0[813],partial_product_low1[813],96'b0};
assign col_out_814 = {u0_col_out_814,u1_data_out_0[814],u1_data_out_1[814],u1_data_out_2[814],u1_data_out_3[814],partial_product_low0[814],partial_product_low1[814],96'b0};
assign col_out_815 = {u0_col_out_815,u1_data_out_0[815],u1_data_out_1[815],u1_data_out_2[815],u1_data_out_3[815],partial_product_low0[815],partial_product_low1[815],96'b0};
assign col_out_816 = {u0_col_out_816,u1_data_out_0[816],u1_data_out_1[816],u1_data_out_2[816],u1_data_out_3[816],partial_product_low0[816],partial_product_low1[816],96'b0};
assign col_out_817 = {u0_col_out_817,u1_data_out_0[817],u1_data_out_1[817],u1_data_out_2[817],u1_data_out_3[817],partial_product_low0[817],partial_product_low1[817],96'b0};
assign col_out_818 = {u0_col_out_818,u1_data_out_0[818],u1_data_out_1[818],u1_data_out_2[818],u1_data_out_3[818],partial_product_low0[818],partial_product_low1[818],96'b0};
assign col_out_819 = {u0_col_out_819,u1_data_out_0[819],u1_data_out_1[819],u1_data_out_2[819],u1_data_out_3[819],partial_product_low0[819],partial_product_low1[819],96'b0};
assign col_out_820 = {u0_col_out_820,u1_data_out_0[820],u1_data_out_1[820],u1_data_out_2[820],u1_data_out_3[820],partial_product_low0[820],partial_product_low1[820],96'b0};
assign col_out_821 = {u0_col_out_821,u1_data_out_0[821],u1_data_out_1[821],u1_data_out_2[821],u1_data_out_3[821],partial_product_low0[821],partial_product_low1[821],96'b0};
assign col_out_822 = {u0_col_out_822,u1_data_out_0[822],u1_data_out_1[822],u1_data_out_2[822],u1_data_out_3[822],partial_product_low0[822],partial_product_low1[822],96'b0};
assign col_out_823 = {u0_col_out_823,u1_data_out_0[823],u1_data_out_1[823],u1_data_out_2[823],u1_data_out_3[823],partial_product_low0[823],partial_product_low1[823],96'b0};
assign col_out_824 = {u0_col_out_824,u1_data_out_0[824],u1_data_out_1[824],u1_data_out_2[824],u1_data_out_3[824],partial_product_low0[824],partial_product_low1[824],96'b0};
assign col_out_825 = {u0_col_out_825,u1_data_out_0[825],u1_data_out_1[825],u1_data_out_2[825],u1_data_out_3[825],partial_product_low0[825],partial_product_low1[825],96'b0};
assign col_out_826 = {u0_col_out_826,u1_data_out_0[826],u1_data_out_1[826],u1_data_out_2[826],u1_data_out_3[826],partial_product_low0[826],partial_product_low1[826],96'b0};
assign col_out_827 = {u0_col_out_827,u1_data_out_0[827],u1_data_out_1[827],u1_data_out_2[827],u1_data_out_3[827],partial_product_low0[827],partial_product_low1[827],96'b0};
assign col_out_828 = {u0_col_out_828,u1_data_out_0[828],u1_data_out_1[828],u1_data_out_2[828],u1_data_out_3[828],partial_product_low0[828],partial_product_low1[828],96'b0};
assign col_out_829 = {u0_col_out_829,u1_data_out_0[829],u1_data_out_1[829],u1_data_out_2[829],u1_data_out_3[829],partial_product_low0[829],partial_product_low1[829],96'b0};
assign col_out_830 = {u0_col_out_830,u1_data_out_0[830],u1_data_out_1[830],u1_data_out_2[830],u1_data_out_3[830],partial_product_low0[830],partial_product_low1[830],96'b0};
assign col_out_831 = {u0_col_out_831,u1_data_out_0[831],u1_data_out_1[831],u1_data_out_2[831],u1_data_out_3[831],partial_product_low0[831],partial_product_low1[831],96'b0};
assign col_out_832 = {u0_col_out_832,u1_data_out_0[832],u1_data_out_1[832],u1_data_out_2[832],u1_data_out_3[832],partial_product_low0[832],partial_product_low1[832],96'b0};
assign col_out_833 = {u0_col_out_833,u1_data_out_0[833],u1_data_out_1[833],u1_data_out_2[833],u1_data_out_3[833],partial_product_low0[833],partial_product_low1[833],96'b0};
assign col_out_834 = {u0_col_out_834,u1_data_out_0[834],u1_data_out_1[834],u1_data_out_2[834],u1_data_out_3[834],partial_product_low0[834],partial_product_low1[834],96'b0};
assign col_out_835 = {u0_col_out_835,u1_data_out_0[835],u1_data_out_1[835],u1_data_out_2[835],u1_data_out_3[835],partial_product_low0[835],partial_product_low1[835],96'b0};
assign col_out_836 = {u0_col_out_836,u1_data_out_0[836],u1_data_out_1[836],u1_data_out_2[836],u1_data_out_3[836],partial_product_low0[836],partial_product_low1[836],96'b0};
assign col_out_837 = {u0_col_out_837,u1_data_out_0[837],u1_data_out_1[837],u1_data_out_2[837],u1_data_out_3[837],partial_product_low0[837],partial_product_low1[837],96'b0};
assign col_out_838 = {u0_col_out_838,u1_data_out_0[838],u1_data_out_1[838],u1_data_out_2[838],u1_data_out_3[838],partial_product_low0[838],partial_product_low1[838],96'b0};
assign col_out_839 = {u0_col_out_839,u1_data_out_0[839],u1_data_out_1[839],u1_data_out_2[839],u1_data_out_3[839],partial_product_low0[839],partial_product_low1[839],96'b0};
assign col_out_840 = {u0_col_out_840,u1_data_out_0[840],u1_data_out_1[840],u1_data_out_2[840],u1_data_out_3[840],partial_product_low0[840],partial_product_low1[840],96'b0};
assign col_out_841 = {u0_col_out_841,u1_data_out_0[841],u1_data_out_1[841],u1_data_out_2[841],u1_data_out_3[841],partial_product_low0[841],partial_product_low1[841],96'b0};
assign col_out_842 = {u0_col_out_842,u1_data_out_0[842],u1_data_out_1[842],u1_data_out_2[842],u1_data_out_3[842],partial_product_low0[842],partial_product_low1[842],96'b0};
assign col_out_843 = {u0_col_out_843,u1_data_out_0[843],u1_data_out_1[843],u1_data_out_2[843],u1_data_out_3[843],partial_product_low0[843],partial_product_low1[843],96'b0};
assign col_out_844 = {u0_col_out_844,u1_data_out_0[844],u1_data_out_1[844],u1_data_out_2[844],u1_data_out_3[844],partial_product_low0[844],partial_product_low1[844],96'b0};
assign col_out_845 = {u0_col_out_845,u1_data_out_0[845],u1_data_out_1[845],u1_data_out_2[845],u1_data_out_3[845],partial_product_low0[845],partial_product_low1[845],96'b0};
assign col_out_846 = {u0_col_out_846,u1_data_out_0[846],u1_data_out_1[846],u1_data_out_2[846],u1_data_out_3[846],partial_product_low0[846],partial_product_low1[846],96'b0};
assign col_out_847 = {u0_col_out_847,u1_data_out_0[847],u1_data_out_1[847],u1_data_out_2[847],u1_data_out_3[847],partial_product_low0[847],partial_product_low1[847],96'b0};
assign col_out_848 = {u0_col_out_848,u1_data_out_0[848],u1_data_out_1[848],u1_data_out_2[848],u1_data_out_3[848],partial_product_low0[848],partial_product_low1[848],96'b0};
assign col_out_849 = {u0_col_out_849,u1_data_out_0[849],u1_data_out_1[849],u1_data_out_2[849],u1_data_out_3[849],partial_product_low0[849],partial_product_low1[849],96'b0};
assign col_out_850 = {u0_col_out_850,u1_data_out_0[850],u1_data_out_1[850],u1_data_out_2[850],u1_data_out_3[850],partial_product_low0[850],partial_product_low1[850],96'b0};
assign col_out_851 = {u0_col_out_851,u1_data_out_0[851],u1_data_out_1[851],u1_data_out_2[851],u1_data_out_3[851],partial_product_low0[851],partial_product_low1[851],96'b0};
assign col_out_852 = {u0_col_out_852,u1_data_out_0[852],u1_data_out_1[852],u1_data_out_2[852],u1_data_out_3[852],partial_product_low0[852],partial_product_low1[852],96'b0};
assign col_out_853 = {u0_col_out_853,u1_data_out_0[853],u1_data_out_1[853],u1_data_out_2[853],u1_data_out_3[853],partial_product_low0[853],partial_product_low1[853],96'b0};
assign col_out_854 = {u0_col_out_854,u1_data_out_0[854],u1_data_out_1[854],u1_data_out_2[854],u1_data_out_3[854],partial_product_low0[854],partial_product_low1[854],96'b0};
assign col_out_855 = {u0_col_out_855,u1_data_out_0[855],u1_data_out_1[855],u1_data_out_2[855],u1_data_out_3[855],partial_product_low0[855],partial_product_low1[855],96'b0};
assign col_out_856 = {u0_col_out_856,u1_data_out_0[856],u1_data_out_1[856],u1_data_out_2[856],u1_data_out_3[856],partial_product_low0[856],partial_product_low1[856],96'b0};
assign col_out_857 = {u0_col_out_857,u1_data_out_0[857],u1_data_out_1[857],u1_data_out_2[857],u1_data_out_3[857],partial_product_low0[857],partial_product_low1[857],96'b0};
assign col_out_858 = {u0_col_out_858,u1_data_out_0[858],u1_data_out_1[858],u1_data_out_2[858],u1_data_out_3[858],partial_product_low0[858],partial_product_low1[858],96'b0};
assign col_out_859 = {u0_col_out_859,u1_data_out_0[859],u1_data_out_1[859],u1_data_out_2[859],u1_data_out_3[859],partial_product_low0[859],partial_product_low1[859],96'b0};
assign col_out_860 = {u0_col_out_860,u1_data_out_0[860],u1_data_out_1[860],u1_data_out_2[860],u1_data_out_3[860],partial_product_low0[860],partial_product_low1[860],96'b0};
assign col_out_861 = {u0_col_out_861,u1_data_out_0[861],u1_data_out_1[861],u1_data_out_2[861],u1_data_out_3[861],partial_product_low0[861],partial_product_low1[861],96'b0};
assign col_out_862 = {u0_col_out_862,u1_data_out_0[862],u1_data_out_1[862],u1_data_out_2[862],u1_data_out_3[862],partial_product_low0[862],partial_product_low1[862],96'b0};
assign col_out_863 = {u0_col_out_863,u1_data_out_0[863],u1_data_out_1[863],u1_data_out_2[863],u1_data_out_3[863],partial_product_low0[863],partial_product_low1[863],96'b0};
assign col_out_864 = {u0_col_out_864,u1_data_out_0[864],u1_data_out_1[864],u1_data_out_2[864],u1_data_out_3[864],partial_product_low0[864],partial_product_low1[864],96'b0};
assign col_out_865 = {u0_col_out_865,u1_data_out_0[865],u1_data_out_1[865],u1_data_out_2[865],u1_data_out_3[865],partial_product_low0[865],partial_product_low1[865],96'b0};
assign col_out_866 = {u0_col_out_866,u1_data_out_0[866],u1_data_out_1[866],u1_data_out_2[866],u1_data_out_3[866],partial_product_low0[866],partial_product_low1[866],96'b0};
assign col_out_867 = {u0_col_out_867,u1_data_out_0[867],u1_data_out_1[867],u1_data_out_2[867],u1_data_out_3[867],partial_product_low0[867],partial_product_low1[867],96'b0};
assign col_out_868 = {u0_col_out_868,u1_data_out_0[868],u1_data_out_1[868],u1_data_out_2[868],u1_data_out_3[868],partial_product_low0[868],partial_product_low1[868],96'b0};
assign col_out_869 = {u0_col_out_869,u1_data_out_0[869],u1_data_out_1[869],u1_data_out_2[869],u1_data_out_3[869],partial_product_low0[869],partial_product_low1[869],96'b0};
assign col_out_870 = {u0_col_out_870,u1_data_out_0[870],u1_data_out_1[870],u1_data_out_2[870],u1_data_out_3[870],partial_product_low0[870],partial_product_low1[870],96'b0};
assign col_out_871 = {u0_col_out_871,u1_data_out_0[871],u1_data_out_1[871],u1_data_out_2[871],u1_data_out_3[871],partial_product_low0[871],partial_product_low1[871],96'b0};
assign col_out_872 = {u0_col_out_872,u1_data_out_0[872],u1_data_out_1[872],u1_data_out_2[872],u1_data_out_3[872],partial_product_low0[872],partial_product_low1[872],96'b0};
assign col_out_873 = {u0_col_out_873,u1_data_out_0[873],u1_data_out_1[873],u1_data_out_2[873],u1_data_out_3[873],partial_product_low0[873],partial_product_low1[873],96'b0};
assign col_out_874 = {u0_col_out_874,u1_data_out_0[874],u1_data_out_1[874],u1_data_out_2[874],u1_data_out_3[874],partial_product_low0[874],partial_product_low1[874],96'b0};
assign col_out_875 = {u0_col_out_875,u1_data_out_0[875],u1_data_out_1[875],u1_data_out_2[875],u1_data_out_3[875],partial_product_low0[875],partial_product_low1[875],96'b0};
assign col_out_876 = {u0_col_out_876,u1_data_out_0[876],u1_data_out_1[876],u1_data_out_2[876],u1_data_out_3[876],partial_product_low0[876],partial_product_low1[876],96'b0};
assign col_out_877 = {u0_col_out_877,u1_data_out_0[877],u1_data_out_1[877],u1_data_out_2[877],u1_data_out_3[877],partial_product_low0[877],partial_product_low1[877],96'b0};
assign col_out_878 = {u0_col_out_878,u1_data_out_0[878],u1_data_out_1[878],u1_data_out_2[878],u1_data_out_3[878],partial_product_low0[878],partial_product_low1[878],96'b0};
assign col_out_879 = {u0_col_out_879,u1_data_out_0[879],u1_data_out_1[879],u1_data_out_2[879],u1_data_out_3[879],partial_product_low0[879],partial_product_low1[879],96'b0};
assign col_out_880 = {u0_col_out_880,u1_data_out_0[880],u1_data_out_1[880],u1_data_out_2[880],u1_data_out_3[880],partial_product_low0[880],partial_product_low1[880],96'b0};
assign col_out_881 = {u0_col_out_881,u1_data_out_0[881],u1_data_out_1[881],u1_data_out_2[881],u1_data_out_3[881],partial_product_low0[881],partial_product_low1[881],96'b0};
assign col_out_882 = {u0_col_out_882,u1_data_out_0[882],u1_data_out_1[882],u1_data_out_2[882],u1_data_out_3[882],partial_product_low0[882],partial_product_low1[882],96'b0};
assign col_out_883 = {u0_col_out_883,u1_data_out_0[883],u1_data_out_1[883],u1_data_out_2[883],u1_data_out_3[883],partial_product_low0[883],partial_product_low1[883],96'b0};
assign col_out_884 = {u0_col_out_884,u1_data_out_0[884],u1_data_out_1[884],u1_data_out_2[884],u1_data_out_3[884],partial_product_low0[884],partial_product_low1[884],96'b0};
assign col_out_885 = {u0_col_out_885,u1_data_out_0[885],u1_data_out_1[885],u1_data_out_2[885],u1_data_out_3[885],partial_product_low0[885],partial_product_low1[885],96'b0};
assign col_out_886 = {u0_col_out_886,u1_data_out_0[886],u1_data_out_1[886],u1_data_out_2[886],u1_data_out_3[886],partial_product_low0[886],partial_product_low1[886],96'b0};
assign col_out_887 = {u0_col_out_887,u1_data_out_0[887],u1_data_out_1[887],u1_data_out_2[887],u1_data_out_3[887],partial_product_low0[887],partial_product_low1[887],96'b0};
assign col_out_888 = {u0_col_out_888,u1_data_out_0[888],u1_data_out_1[888],u1_data_out_2[888],u1_data_out_3[888],partial_product_low0[888],partial_product_low1[888],96'b0};
assign col_out_889 = {u0_col_out_889,u1_data_out_0[889],u1_data_out_1[889],u1_data_out_2[889],u1_data_out_3[889],partial_product_low0[889],partial_product_low1[889],96'b0};
assign col_out_890 = {u0_col_out_890,u1_data_out_0[890],u1_data_out_1[890],u1_data_out_2[890],u1_data_out_3[890],partial_product_low0[890],partial_product_low1[890],96'b0};
assign col_out_891 = {u0_col_out_891,u1_data_out_0[891],u1_data_out_1[891],u1_data_out_2[891],u1_data_out_3[891],partial_product_low0[891],partial_product_low1[891],96'b0};
assign col_out_892 = {u0_col_out_892,u1_data_out_0[892],u1_data_out_1[892],u1_data_out_2[892],u1_data_out_3[892],partial_product_low0[892],partial_product_low1[892],96'b0};
assign col_out_893 = {u0_col_out_893,u1_data_out_0[893],u1_data_out_1[893],u1_data_out_2[893],u1_data_out_3[893],partial_product_low0[893],partial_product_low1[893],96'b0};
assign col_out_894 = {u0_col_out_894,u1_data_out_0[894],u1_data_out_1[894],u1_data_out_2[894],u1_data_out_3[894],partial_product_low0[894],partial_product_low1[894],96'b0};
assign col_out_895 = {u0_col_out_895,u1_data_out_0[895],u1_data_out_1[895],u1_data_out_2[895],u1_data_out_3[895],partial_product_low0[895],partial_product_low1[895],96'b0};
assign col_out_896 = {u0_col_out_896,u1_data_out_0[896],u1_data_out_1[896],u1_data_out_2[896],u1_data_out_3[896],partial_product_low0[896],partial_product_low1[896],96'b0};
assign col_out_897 = {u0_col_out_897,u1_data_out_0[897],u1_data_out_1[897],u1_data_out_2[897],u1_data_out_3[897],partial_product_low0[897],partial_product_low1[897],96'b0};
assign col_out_898 = {u0_col_out_898,u1_data_out_0[898],u1_data_out_1[898],u1_data_out_2[898],u1_data_out_3[898],partial_product_low0[898],partial_product_low1[898],96'b0};
assign col_out_899 = {u0_col_out_899,u1_data_out_0[899],u1_data_out_1[899],u1_data_out_2[899],u1_data_out_3[899],partial_product_low0[899],partial_product_low1[899],96'b0};
assign col_out_900 = {u0_col_out_900,u1_data_out_0[900],u1_data_out_1[900],u1_data_out_2[900],u1_data_out_3[900],partial_product_low0[900],partial_product_low1[900],96'b0};
assign col_out_901 = {u0_col_out_901,u1_data_out_0[901],u1_data_out_1[901],u1_data_out_2[901],u1_data_out_3[901],partial_product_low0[901],partial_product_low1[901],96'b0};
assign col_out_902 = {u0_col_out_902,u1_data_out_0[902],u1_data_out_1[902],u1_data_out_2[902],u1_data_out_3[902],partial_product_low0[902],partial_product_low1[902],96'b0};
assign col_out_903 = {u0_col_out_903,u1_data_out_0[903],u1_data_out_1[903],u1_data_out_2[903],u1_data_out_3[903],partial_product_low0[903],partial_product_low1[903],96'b0};
assign col_out_904 = {u0_col_out_904,u1_data_out_0[904],u1_data_out_1[904],u1_data_out_2[904],u1_data_out_3[904],partial_product_low0[904],partial_product_low1[904],96'b0};
assign col_out_905 = {u0_col_out_905,u1_data_out_0[905],u1_data_out_1[905],u1_data_out_2[905],u1_data_out_3[905],partial_product_low0[905],partial_product_low1[905],96'b0};
assign col_out_906 = {u0_col_out_906,u1_data_out_0[906],u1_data_out_1[906],u1_data_out_2[906],u1_data_out_3[906],partial_product_low0[906],partial_product_low1[906],96'b0};
assign col_out_907 = {u0_col_out_907,u1_data_out_0[907],u1_data_out_1[907],u1_data_out_2[907],u1_data_out_3[907],partial_product_low0[907],partial_product_low1[907],96'b0};
assign col_out_908 = {u0_col_out_908,u1_data_out_0[908],u1_data_out_1[908],u1_data_out_2[908],u1_data_out_3[908],partial_product_low0[908],partial_product_low1[908],96'b0};
assign col_out_909 = {u0_col_out_909,u1_data_out_0[909],u1_data_out_1[909],u1_data_out_2[909],u1_data_out_3[909],partial_product_low0[909],partial_product_low1[909],96'b0};
assign col_out_910 = {u0_col_out_910,u1_data_out_0[910],u1_data_out_1[910],u1_data_out_2[910],u1_data_out_3[910],partial_product_low0[910],partial_product_low1[910],96'b0};
assign col_out_911 = {u0_col_out_911,u1_data_out_0[911],u1_data_out_1[911],u1_data_out_2[911],u1_data_out_3[911],partial_product_low0[911],partial_product_low1[911],96'b0};
assign col_out_912 = {u0_col_out_912,u1_data_out_0[912],u1_data_out_1[912],u1_data_out_2[912],u1_data_out_3[912],partial_product_low0[912],partial_product_low1[912],96'b0};
assign col_out_913 = {u0_col_out_913,u1_data_out_0[913],u1_data_out_1[913],u1_data_out_2[913],u1_data_out_3[913],partial_product_low0[913],partial_product_low1[913],96'b0};
assign col_out_914 = {u0_col_out_914,u1_data_out_0[914],u1_data_out_1[914],u1_data_out_2[914],u1_data_out_3[914],partial_product_low0[914],partial_product_low1[914],96'b0};
assign col_out_915 = {u0_col_out_915,u1_data_out_0[915],u1_data_out_1[915],u1_data_out_2[915],u1_data_out_3[915],partial_product_low0[915],partial_product_low1[915],96'b0};
assign col_out_916 = {u0_col_out_916,u1_data_out_0[916],u1_data_out_1[916],u1_data_out_2[916],u1_data_out_3[916],partial_product_low0[916],partial_product_low1[916],96'b0};
assign col_out_917 = {u0_col_out_917,u1_data_out_0[917],u1_data_out_1[917],u1_data_out_2[917],u1_data_out_3[917],partial_product_low0[917],partial_product_low1[917],96'b0};
assign col_out_918 = {u0_col_out_918,u1_data_out_0[918],u1_data_out_1[918],u1_data_out_2[918],u1_data_out_3[918],partial_product_low0[918],partial_product_low1[918],96'b0};
assign col_out_919 = {u0_col_out_919,u1_data_out_0[919],u1_data_out_1[919],u1_data_out_2[919],u1_data_out_3[919],partial_product_low0[919],partial_product_low1[919],96'b0};
assign col_out_920 = {u0_col_out_920,u1_data_out_0[920],u1_data_out_1[920],u1_data_out_2[920],u1_data_out_3[920],partial_product_low0[920],partial_product_low1[920],96'b0};
assign col_out_921 = {u0_col_out_921,u1_data_out_0[921],u1_data_out_1[921],u1_data_out_2[921],u1_data_out_3[921],partial_product_low0[921],partial_product_low1[921],96'b0};
assign col_out_922 = {u0_col_out_922,u1_data_out_0[922],u1_data_out_1[922],u1_data_out_2[922],u1_data_out_3[922],partial_product_low0[922],partial_product_low1[922],96'b0};
assign col_out_923 = {u0_col_out_923,u1_data_out_0[923],u1_data_out_1[923],u1_data_out_2[923],u1_data_out_3[923],partial_product_low0[923],partial_product_low1[923],96'b0};
assign col_out_924 = {u0_col_out_924,u1_data_out_0[924],u1_data_out_1[924],u1_data_out_2[924],u1_data_out_3[924],partial_product_low0[924],partial_product_low1[924],96'b0};
assign col_out_925 = {u0_col_out_925,u1_data_out_0[925],u1_data_out_1[925],u1_data_out_2[925],u1_data_out_3[925],partial_product_low0[925],partial_product_low1[925],96'b0};
assign col_out_926 = {u0_col_out_926,u1_data_out_0[926],u1_data_out_1[926],u1_data_out_2[926],u1_data_out_3[926],partial_product_low0[926],partial_product_low1[926],96'b0};
assign col_out_927 = {u0_col_out_927,u1_data_out_0[927],u1_data_out_1[927],u1_data_out_2[927],u1_data_out_3[927],partial_product_low0[927],partial_product_low1[927],96'b0};
assign col_out_928 = {u0_col_out_928,u1_data_out_0[928],u1_data_out_1[928],u1_data_out_2[928],u1_data_out_3[928],partial_product_low0[928],partial_product_low1[928],96'b0};
assign col_out_929 = {u0_col_out_929,u1_data_out_0[929],u1_data_out_1[929],u1_data_out_2[929],u1_data_out_3[929],partial_product_low0[929],partial_product_low1[929],96'b0};
assign col_out_930 = {u0_col_out_930,u1_data_out_0[930],u1_data_out_1[930],u1_data_out_2[930],u1_data_out_3[930],partial_product_low0[930],partial_product_low1[930],96'b0};
assign col_out_931 = {u0_col_out_931,u1_data_out_0[931],u1_data_out_1[931],u1_data_out_2[931],u1_data_out_3[931],partial_product_low0[931],partial_product_low1[931],96'b0};
assign col_out_932 = {u0_col_out_932,u1_data_out_0[932],u1_data_out_1[932],u1_data_out_2[932],u1_data_out_3[932],partial_product_low0[932],partial_product_low1[932],96'b0};
assign col_out_933 = {u0_col_out_933,u1_data_out_0[933],u1_data_out_1[933],u1_data_out_2[933],u1_data_out_3[933],partial_product_low0[933],partial_product_low1[933],96'b0};
assign col_out_934 = {u0_col_out_934,u1_data_out_0[934],u1_data_out_1[934],u1_data_out_2[934],u1_data_out_3[934],partial_product_low0[934],partial_product_low1[934],96'b0};
assign col_out_935 = {u0_col_out_935,u1_data_out_0[935],u1_data_out_1[935],u1_data_out_2[935],u1_data_out_3[935],partial_product_low0[935],partial_product_low1[935],96'b0};
assign col_out_936 = {u0_col_out_936,u1_data_out_0[936],u1_data_out_1[936],u1_data_out_2[936],u1_data_out_3[936],partial_product_low0[936],partial_product_low1[936],96'b0};
assign col_out_937 = {u0_col_out_937,u1_data_out_0[937],u1_data_out_1[937],u1_data_out_2[937],u1_data_out_3[937],partial_product_low0[937],partial_product_low1[937],96'b0};
assign col_out_938 = {u0_col_out_938,u1_data_out_0[938],u1_data_out_1[938],u1_data_out_2[938],u1_data_out_3[938],partial_product_low0[938],partial_product_low1[938],96'b0};
assign col_out_939 = {u0_col_out_939,u1_data_out_0[939],u1_data_out_1[939],u1_data_out_2[939],u1_data_out_3[939],partial_product_low0[939],partial_product_low1[939],96'b0};
assign col_out_940 = {u0_col_out_940,u1_data_out_0[940],u1_data_out_1[940],u1_data_out_2[940],u1_data_out_3[940],partial_product_low0[940],partial_product_low1[940],96'b0};
assign col_out_941 = {u0_col_out_941,u1_data_out_0[941],u1_data_out_1[941],u1_data_out_2[941],u1_data_out_3[941],partial_product_low0[941],partial_product_low1[941],96'b0};
assign col_out_942 = {u0_col_out_942,u1_data_out_0[942],u1_data_out_1[942],u1_data_out_2[942],u1_data_out_3[942],partial_product_low0[942],partial_product_low1[942],96'b0};
assign col_out_943 = {u0_col_out_943,u1_data_out_0[943],u1_data_out_1[943],u1_data_out_2[943],u1_data_out_3[943],partial_product_low0[943],partial_product_low1[943],96'b0};
assign col_out_944 = {u0_col_out_944,u1_data_out_0[944],u1_data_out_1[944],u1_data_out_2[944],u1_data_out_3[944],partial_product_low0[944],partial_product_low1[944],96'b0};
assign col_out_945 = {u0_col_out_945,u1_data_out_0[945],u1_data_out_1[945],u1_data_out_2[945],u1_data_out_3[945],partial_product_low0[945],partial_product_low1[945],96'b0};
assign col_out_946 = {u0_col_out_946,u1_data_out_0[946],u1_data_out_1[946],u1_data_out_2[946],u1_data_out_3[946],partial_product_low0[946],partial_product_low1[946],96'b0};
assign col_out_947 = {u0_col_out_947,u1_data_out_0[947],u1_data_out_1[947],u1_data_out_2[947],u1_data_out_3[947],partial_product_low0[947],partial_product_low1[947],96'b0};
assign col_out_948 = {u0_col_out_948,u1_data_out_0[948],u1_data_out_1[948],u1_data_out_2[948],u1_data_out_3[948],partial_product_low0[948],partial_product_low1[948],96'b0};
assign col_out_949 = {u0_col_out_949,u1_data_out_0[949],u1_data_out_1[949],u1_data_out_2[949],u1_data_out_3[949],partial_product_low0[949],partial_product_low1[949],96'b0};
assign col_out_950 = {u0_col_out_950,u1_data_out_0[950],u1_data_out_1[950],u1_data_out_2[950],u1_data_out_3[950],partial_product_low0[950],partial_product_low1[950],96'b0};
assign col_out_951 = {u0_col_out_951,u1_data_out_0[951],u1_data_out_1[951],u1_data_out_2[951],u1_data_out_3[951],partial_product_low0[951],partial_product_low1[951],96'b0};
assign col_out_952 = {u0_col_out_952,u1_data_out_0[952],u1_data_out_1[952],u1_data_out_2[952],u1_data_out_3[952],partial_product_low0[952],partial_product_low1[952],96'b0};
assign col_out_953 = {u0_col_out_953,u1_data_out_0[953],u1_data_out_1[953],u1_data_out_2[953],u1_data_out_3[953],partial_product_low0[953],partial_product_low1[953],96'b0};
assign col_out_954 = {u0_col_out_954,u1_data_out_0[954],u1_data_out_1[954],u1_data_out_2[954],u1_data_out_3[954],partial_product_low0[954],partial_product_low1[954],96'b0};
assign col_out_955 = {u0_col_out_955,u1_data_out_0[955],u1_data_out_1[955],u1_data_out_2[955],u1_data_out_3[955],partial_product_low0[955],partial_product_low1[955],96'b0};
assign col_out_956 = {u0_col_out_956,u1_data_out_0[956],u1_data_out_1[956],u1_data_out_2[956],u1_data_out_3[956],partial_product_low0[956],partial_product_low1[956],96'b0};
assign col_out_957 = {u0_col_out_957,u1_data_out_0[957],u1_data_out_1[957],u1_data_out_2[957],u1_data_out_3[957],partial_product_low0[957],partial_product_low1[957],96'b0};
assign col_out_958 = {u0_col_out_958,u1_data_out_0[958],u1_data_out_1[958],u1_data_out_2[958],u1_data_out_3[958],partial_product_low0[958],partial_product_low1[958],96'b0};
assign col_out_959 = {u0_col_out_959,u1_data_out_0[959],u1_data_out_1[959],u1_data_out_2[959],u1_data_out_3[959],partial_product_low0[959],partial_product_low1[959],96'b0};
assign col_out_960 = {u0_col_out_960,u1_data_out_0[960],u1_data_out_1[960],u1_data_out_2[960],u1_data_out_3[960],partial_product_low0[960],partial_product_low1[960],96'b0};
assign col_out_961 = {u0_col_out_961,u1_data_out_0[961],u1_data_out_1[961],u1_data_out_2[961],u1_data_out_3[961],partial_product_low0[961],partial_product_low1[961],96'b0};
assign col_out_962 = {u0_col_out_962,u1_data_out_0[962],u1_data_out_1[962],u1_data_out_2[962],u1_data_out_3[962],partial_product_low0[962],partial_product_low1[962],96'b0};
assign col_out_963 = {u0_col_out_963,u1_data_out_0[963],u1_data_out_1[963],u1_data_out_2[963],u1_data_out_3[963],partial_product_low0[963],partial_product_low1[963],96'b0};
assign col_out_964 = {u0_col_out_964,u1_data_out_0[964],u1_data_out_1[964],u1_data_out_2[964],u1_data_out_3[964],partial_product_low0[964],partial_product_low1[964],96'b0};
assign col_out_965 = {u0_col_out_965,u1_data_out_0[965],u1_data_out_1[965],u1_data_out_2[965],u1_data_out_3[965],partial_product_low0[965],partial_product_low1[965],96'b0};
assign col_out_966 = {u0_col_out_966,u1_data_out_0[966],u1_data_out_1[966],u1_data_out_2[966],u1_data_out_3[966],partial_product_low0[966],partial_product_low1[966],96'b0};
assign col_out_967 = {u0_col_out_967,u1_data_out_0[967],u1_data_out_1[967],u1_data_out_2[967],u1_data_out_3[967],partial_product_low0[967],partial_product_low1[967],96'b0};
assign col_out_968 = {u0_col_out_968,u1_data_out_0[968],u1_data_out_1[968],u1_data_out_2[968],u1_data_out_3[968],partial_product_low0[968],partial_product_low1[968],96'b0};
assign col_out_969 = {u0_col_out_969,u1_data_out_0[969],u1_data_out_1[969],u1_data_out_2[969],u1_data_out_3[969],partial_product_low0[969],partial_product_low1[969],96'b0};
assign col_out_970 = {u0_col_out_970,u1_data_out_0[970],u1_data_out_1[970],u1_data_out_2[970],u1_data_out_3[970],partial_product_low0[970],partial_product_low1[970],96'b0};
assign col_out_971 = {u0_col_out_971,u1_data_out_0[971],u1_data_out_1[971],u1_data_out_2[971],u1_data_out_3[971],partial_product_low0[971],partial_product_low1[971],96'b0};
assign col_out_972 = {u0_col_out_972,u1_data_out_0[972],u1_data_out_1[972],u1_data_out_2[972],u1_data_out_3[972],partial_product_low0[972],partial_product_low1[972],96'b0};
assign col_out_973 = {u0_col_out_973,u1_data_out_0[973],u1_data_out_1[973],u1_data_out_2[973],u1_data_out_3[973],partial_product_low0[973],partial_product_low1[973],96'b0};
assign col_out_974 = {u0_col_out_974,u1_data_out_0[974],u1_data_out_1[974],u1_data_out_2[974],u1_data_out_3[974],partial_product_low0[974],partial_product_low1[974],96'b0};
assign col_out_975 = {u0_col_out_975,u1_data_out_0[975],u1_data_out_1[975],u1_data_out_2[975],u1_data_out_3[975],partial_product_low0[975],partial_product_low1[975],96'b0};
assign col_out_976 = {u0_col_out_976,u1_data_out_0[976],u1_data_out_1[976],u1_data_out_2[976],u1_data_out_3[976],partial_product_low0[976],partial_product_low1[976],96'b0};
assign col_out_977 = {u0_col_out_977,u1_data_out_0[977],u1_data_out_1[977],u1_data_out_2[977],u1_data_out_3[977],partial_product_low0[977],partial_product_low1[977],96'b0};
assign col_out_978 = {u0_col_out_978,u1_data_out_0[978],u1_data_out_1[978],u1_data_out_2[978],u1_data_out_3[978],partial_product_low0[978],partial_product_low1[978],96'b0};
assign col_out_979 = {u0_col_out_979,u1_data_out_0[979],u1_data_out_1[979],u1_data_out_2[979],u1_data_out_3[979],partial_product_low0[979],partial_product_low1[979],96'b0};
assign col_out_980 = {u0_col_out_980,u1_data_out_0[980],u1_data_out_1[980],u1_data_out_2[980],u1_data_out_3[980],partial_product_low0[980],partial_product_low1[980],96'b0};
assign col_out_981 = {u0_col_out_981,u1_data_out_0[981],u1_data_out_1[981],u1_data_out_2[981],u1_data_out_3[981],partial_product_low0[981],partial_product_low1[981],96'b0};
assign col_out_982 = {u0_col_out_982,u1_data_out_0[982],u1_data_out_1[982],u1_data_out_2[982],u1_data_out_3[982],partial_product_low0[982],partial_product_low1[982],96'b0};
assign col_out_983 = {u0_col_out_983,u1_data_out_0[983],u1_data_out_1[983],u1_data_out_2[983],u1_data_out_3[983],partial_product_low0[983],partial_product_low1[983],96'b0};
assign col_out_984 = {u0_col_out_984,u1_data_out_0[984],u1_data_out_1[984],u1_data_out_2[984],u1_data_out_3[984],partial_product_low0[984],partial_product_low1[984],96'b0};
assign col_out_985 = {u0_col_out_985,u1_data_out_0[985],u1_data_out_1[985],u1_data_out_2[985],u1_data_out_3[985],partial_product_low0[985],partial_product_low1[985],96'b0};
assign col_out_986 = {u0_col_out_986,u1_data_out_0[986],u1_data_out_1[986],u1_data_out_2[986],u1_data_out_3[986],partial_product_low0[986],partial_product_low1[986],96'b0};
assign col_out_987 = {u0_col_out_987,u1_data_out_0[987],u1_data_out_1[987],u1_data_out_2[987],u1_data_out_3[987],partial_product_low0[987],partial_product_low1[987],96'b0};
assign col_out_988 = {u0_col_out_988,u1_data_out_0[988],u1_data_out_1[988],u1_data_out_2[988],u1_data_out_3[988],partial_product_low0[988],partial_product_low1[988],96'b0};
assign col_out_989 = {u0_col_out_989,u1_data_out_0[989],u1_data_out_1[989],u1_data_out_2[989],u1_data_out_3[989],partial_product_low0[989],partial_product_low1[989],96'b0};
assign col_out_990 = {u0_col_out_990,u1_data_out_0[990],u1_data_out_1[990],u1_data_out_2[990],u1_data_out_3[990],partial_product_low0[990],partial_product_low1[990],96'b0};
assign col_out_991 = {u0_col_out_991,u1_data_out_0[991],u1_data_out_1[991],u1_data_out_2[991],u1_data_out_3[991],partial_product_low0[991],partial_product_low1[991],96'b0};
assign col_out_992 = {u0_col_out_992,u1_data_out_0[992],u1_data_out_1[992],u1_data_out_2[992],u1_data_out_3[992],partial_product_low0[992],partial_product_low1[992],96'b0};
assign col_out_993 = {u0_col_out_993,u1_data_out_0[993],u1_data_out_1[993],u1_data_out_2[993],u1_data_out_3[993],partial_product_low0[993],partial_product_low1[993],96'b0};
assign col_out_994 = {u0_col_out_994,u1_data_out_0[994],u1_data_out_1[994],u1_data_out_2[994],u1_data_out_3[994],partial_product_low0[994],partial_product_low1[994],96'b0};
assign col_out_995 = {u0_col_out_995,u1_data_out_0[995],u1_data_out_1[995],u1_data_out_2[995],u1_data_out_3[995],partial_product_low0[995],partial_product_low1[995],96'b0};
assign col_out_996 = {u0_col_out_996,u1_data_out_0[996],u1_data_out_1[996],u1_data_out_2[996],u1_data_out_3[996],partial_product_low0[996],partial_product_low1[996],96'b0};
assign col_out_997 = {u0_col_out_997,u1_data_out_0[997],u1_data_out_1[997],u1_data_out_2[997],u1_data_out_3[997],partial_product_low0[997],partial_product_low1[997],96'b0};
assign col_out_998 = {u0_col_out_998,u1_data_out_0[998],u1_data_out_1[998],u1_data_out_2[998],u1_data_out_3[998],partial_product_low0[998],partial_product_low1[998],96'b0};
assign col_out_999 = {u0_col_out_999,u1_data_out_0[999],u1_data_out_1[999],u1_data_out_2[999],u1_data_out_3[999],partial_product_low0[999],partial_product_low1[999],96'b0};
assign col_out_1000 = {u0_col_out_1000,u1_data_out_0[1000],u1_data_out_1[1000],u1_data_out_2[1000],u1_data_out_3[1000],partial_product_low0[1000],partial_product_low1[1000],96'b0};
assign col_out_1001 = {u0_col_out_1001,u1_data_out_0[1001],u1_data_out_1[1001],u1_data_out_2[1001],u1_data_out_3[1001],partial_product_low0[1001],partial_product_low1[1001],96'b0};
assign col_out_1002 = {u0_col_out_1002,u1_data_out_0[1002],u1_data_out_1[1002],u1_data_out_2[1002],u1_data_out_3[1002],partial_product_low0[1002],partial_product_low1[1002],96'b0};
assign col_out_1003 = {u0_col_out_1003,u1_data_out_0[1003],u1_data_out_1[1003],u1_data_out_2[1003],u1_data_out_3[1003],partial_product_low0[1003],partial_product_low1[1003],96'b0};
assign col_out_1004 = {u0_col_out_1004,u1_data_out_0[1004],u1_data_out_1[1004],u1_data_out_2[1004],u1_data_out_3[1004],partial_product_low0[1004],partial_product_low1[1004],96'b0};
assign col_out_1005 = {u0_col_out_1005,u1_data_out_0[1005],u1_data_out_1[1005],u1_data_out_2[1005],u1_data_out_3[1005],partial_product_low0[1005],partial_product_low1[1005],96'b0};
assign col_out_1006 = {u0_col_out_1006,u1_data_out_0[1006],u1_data_out_1[1006],u1_data_out_2[1006],u1_data_out_3[1006],partial_product_low0[1006],partial_product_low1[1006],96'b0};
assign col_out_1007 = {u0_col_out_1007,u1_data_out_0[1007],u1_data_out_1[1007],u1_data_out_2[1007],u1_data_out_3[1007],partial_product_low0[1007],partial_product_low1[1007],96'b0};
assign col_out_1008 = {u0_col_out_1008,u1_data_out_0[1008],u1_data_out_1[1008],u1_data_out_2[1008],u1_data_out_3[1008],partial_product_low0[1008],partial_product_low1[1008],96'b0};
assign col_out_1009 = {u0_col_out_1009,u1_data_out_0[1009],u1_data_out_1[1009],u1_data_out_2[1009],u1_data_out_3[1009],partial_product_low0[1009],partial_product_low1[1009],96'b0};
assign col_out_1010 = {u0_col_out_1010,u1_data_out_0[1010],u1_data_out_1[1010],u1_data_out_2[1010],u1_data_out_3[1010],partial_product_low0[1010],partial_product_low1[1010],96'b0};
assign col_out_1011 = {u0_col_out_1011,u1_data_out_0[1011],u1_data_out_1[1011],u1_data_out_2[1011],u1_data_out_3[1011],partial_product_low0[1011],partial_product_low1[1011],96'b0};
assign col_out_1012 = {u0_col_out_1012,u1_data_out_0[1012],u1_data_out_1[1012],u1_data_out_2[1012],u1_data_out_3[1012],partial_product_low0[1012],partial_product_low1[1012],96'b0};
assign col_out_1013 = {u0_col_out_1013,u1_data_out_0[1013],u1_data_out_1[1013],u1_data_out_2[1013],u1_data_out_3[1013],partial_product_low0[1013],partial_product_low1[1013],96'b0};
assign col_out_1014 = {u0_col_out_1014,u1_data_out_0[1014],u1_data_out_1[1014],u1_data_out_2[1014],u1_data_out_3[1014],partial_product_low0[1014],partial_product_low1[1014],96'b0};
assign col_out_1015 = {u0_col_out_1015,u1_data_out_0[1015],u1_data_out_1[1015],u1_data_out_2[1015],u1_data_out_3[1015],partial_product_low0[1015],partial_product_low1[1015],96'b0};
assign col_out_1016 = {u0_col_out_1016,u1_data_out_0[1016],u1_data_out_1[1016],u1_data_out_2[1016],u1_data_out_3[1016],partial_product_low0[1016],partial_product_low1[1016],96'b0};
assign col_out_1017 = {u0_col_out_1017,u1_data_out_0[1017],u1_data_out_1[1017],u1_data_out_2[1017],u1_data_out_3[1017],partial_product_low0[1017],partial_product_low1[1017],96'b0};
assign col_out_1018 = {u0_col_out_1018,u1_data_out_0[1018],u1_data_out_1[1018],u1_data_out_2[1018],u1_data_out_3[1018],partial_product_low0[1018],partial_product_low1[1018],96'b0};
assign col_out_1019 = {u0_col_out_1019,u1_data_out_0[1019],u1_data_out_1[1019],u1_data_out_2[1019],u1_data_out_3[1019],partial_product_low0[1019],partial_product_low1[1019],96'b0};
assign col_out_1020 = {u0_col_out_1020,u1_data_out_0[1020],u1_data_out_1[1020],u1_data_out_2[1020],u1_data_out_3[1020],partial_product_low0[1020],partial_product_low1[1020],96'b0};
assign col_out_1021 = {u0_col_out_1021,u1_data_out_0[1021],u1_data_out_1[1021],u1_data_out_2[1021],u1_data_out_3[1021],partial_product_low0[1021],partial_product_low1[1021],96'b0};
assign col_out_1022 = {u0_col_out_1022,u1_data_out_0[1022],u1_data_out_1[1022],u1_data_out_2[1022],u1_data_out_3[1022],partial_product_low0[1022],partial_product_low1[1022],96'b0};
assign col_out_1023 = {u0_col_out_1023,u1_data_out_0[1023],u1_data_out_1[1023],u1_data_out_2[1023],u1_data_out_3[1023],partial_product_low0[1023],partial_product_low1[1023],96'b0};




















endmodule
module xpb_5_880
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h878e88032bc2f32fe65fdb211e53d13e3735dafd4017050edc2d6518cbaaedfd56e6850da4221acc69acb8636d1b571716f84dc4cc4b63eeaf4ed568099a4db8a25dcd8b794cff37e937379c53540d84b6164b1bb06bef2178218604ba94c5d8b47636bb4af4b17cb3081da61d3bcdf9a45a0f5f8c8fa9e6c6b2374e3c75335d;
    5'b00010 : xpb = 1024'h5e6fcab09597b19701ba3e6b2c4d5b2afcf5b2c9aab669a63a7e10dbe4532ef2aa848ca27e1db70a33fb317ff6d89d63c9d673a375e3f791adfe6b71d86226bfd06c66684309012abfd46c960dcc56d878279c9ed451b1323ab67a0ebafee91f39e4db4ce5206a6bdf50546d42a775c9f9da3fdcc8d3f69d46f4f397f008004f;
    5'b00011 : xpb = 1024'h35510d5dff6c6ffe1d14a1b53a46e517c2b58a961555ce3d98cebc9efcfb6fe7fe22943758195347fe49aa9c8095e3b07cb499821f7c8b34acae017ba729ffc6fe7aff450cc5031d9671a18fc844a02c3a38ee21f8377342fd4b6e18bb690c65bf537fde7f4c235b0b988b3468131d9a4f5a705a05184353c737afe1a39acd41;
    5'b00100 : xpb = 1024'hc32500b69412e65386f04ff48406f04887562627ff532d4f71f686215a3b0dd51c09bcc3214ef85c89823b90a5329fd2f92bf60c9151ed7ab5d978575f1d8ce2c899821d68105106d0ed68982bce97ffc4a3fa51c1d3553bfe06222bbd32fac44c224701977dc4a37e0c1fb8d7ec56aa4daa0d7415c900a477a6c2b572d9a33;
    5'b00101 : xpb = 1024'h93c0d80e950421951ecee02066944042bfab3d5fc00c37e3d34ccd7ae14e9edaa8a720d9d6370a523244dc1c776e8114468b0d25956082c65aac6ced7f8c2686cee765ad4fce044856460e25d610f704b2608ac0cc8924753801e8277667f584f9385b2b646c8dc6eae8dfa1aaba93644934b036cdec39f10e2ca37993a2cd90;
    5'b00110 : xpb = 1024'h6aa21abbfed8dffc3a29436a748dca2f856b152c2aab9c7b319d793df9f6dfcffc45286eb032a68ffc935539012bc760f96933043ef91669595c02f74e53ff8dfcf5fe8a198a063b2ce3431f908940587471dc43f06ee685fa96dc3176d218cb7ea6ffbcfe9846b617311668d0263b349eb4e0b40a3086a78e6f5fc347359a82;
    5'b00111 : xpb = 1024'h41835d6968ad9e635583a6b48287541c4b2aecf8954b01128fee2501129f20c54fe330038a2e42cdc6e1ce558ae90dadac4758e2e891aa0c580b99011d1bd8952b049766e346082e038078194b0189ac36832dc71454a896bd2bd03b773c3c120415a44e98c3ffa543794d2ff591e304f43511314674d35e0eb21c0cfac86774;
    5'b01000 : xpb = 1024'h1864a016d2825cca70de09fe9080de0910eac4c4ffea65a9ee3ed0c42b4761baa38137986429df0b9130477214a653fa5f257ec1922a3daf56bb2f0aebe3b19c59133043ad020a20da1dad130579d2fff8947f4a383a6aa77fc0c44577a65f58898448e032efb8946fc183f71afd8ad549b541ae82b920148ef4d856ae5b3466;
    5'b01001 : xpb = 1024'h9ff32819fe454ffa573de51faed4af4748209fc240016ab8ca6c35dcf6f24fb7fa67bca6084bf9d7fadcffd581c1ab11761dcc865e75a19e060a0472f57dff54fb70fdcf264f0958c354e4af58cde084aeaaca65e8a659c8f7e24a4a323b25313dfa7f9b7de46a1122c9a19d383958ceee0f510e0f48c9fb55a70fa4ead067c3;
    5'b01010 : xpb = 1024'h76d46ac7681a0e6172984869bcce39340de0778eaaa0cf5028bce1a00f9a90ad4e05c43ae2479615c52b78f20b7ef15e28fbf265080e354104b99a7cc445d85c297f96abf00b0b4b99f219a9134629d870bc1be90c8c1bd9ba773e5432a54877c369242d181023004f11d8645da5009f438f818b4b8d16b1d5e9cbee9e6334b5;
    5'b01011 : xpb = 1024'h4db5ad74d1eeccc88df2abb3cac7c320d3a04f5b154033e7870d8d632842d1a2a1a3cbcfbc4332538f79f20e953c37aadbda1843b1a6c8e403693086930db163578e2f88b9c70d3e708f4ea2cdbe732c32cd6d6c3071ddea7d0c325e330f6bbe48d7c8beb23bdbef7b5a0f2b8310a86f990fb20887d16368562c883851f601a7;
    5'b01100 : xpb = 1024'h2496f0223bc38b2fa94d0efdd8c14d0d996027277fdf987ee55e392640eb1297f541d364963ece9159c86b2b1ef97df78eb83e225b3f5c870218c69061d58a6a859cc86583830f31472c839c8836bc7ff4debeef54579ffb3fa1266833798f04ce466d504c6794dea7a245f2a87c503fee8fe285c415b01ed66f44820588ce99;
    5'b01101 : xpb = 1024'hac25782567867e5f8facea1ef7151e4bd0960224bff69d8dc18b9e3f0c9600954c2858723a60e95dc375238e8c14d50ea5b08be7278ac075b1679bf86b6fd82327fa95f0fcd00e693063bb38db8aca04aaf50a0b04c38f1cb7c2ac6cee0e54dd82bca40b975c465b5aaa6398c5b81e3992e9f1e550a55a059d217bd041fe01f6;
    5'b01110 : xpb = 1024'h8306bad2d15b3cc6ab074d69050ea8389655d9f12a9602251fdc4a02253e418a9fc66007145c859b8dc39cab15d21b5b588eb1c5d1235418b01732023a37b12a56092ecdc68c105c0700f032960313586d065b8e28a9512d7a57a076ee787824082b489d3187ff4a86f29a5feb23c609e86a22628ce9a6bc1d643819f590cee8;
    5'b01111 : xpb = 1024'h59e7fd803b2ffb2dc661b0b3130832255c15b1bd953566bc7e2cf5c53de6827ff364679bee5821d9581215c79f8f61a80b6cd7a47abbe7bbaec6c80c08ff8a318417c7aa9048124edd9e252c507b5cac2f17ad114c8f133e3cec9480eee29b6a8d99ed2ecbb3b839b33ad127108f6dda3dea52dfc92df3729da6f463a9239bda;
    5'b10000 : xpb = 1024'h30c9402da504b994e1bc13fd2101bc1221d58989ffd4cb53dc7da188568ec37547026f30c853be1722608ee4294ca7f4be4afd8324547b5ead765e15d7c76338b22660875a041441b43b5a260af3a5fff128fe947074d54eff81888aef4cbeb1130891c065df7128df8307ee35fb15aa936a835d057240291de9b0ad5cb668cc;
    5'b10001 : xpb = 1024'h7aa82db0ed977fbfd1677472efb45fee79561566a742feb3ace4d4b6f37046a9aa076c5a24f5a54ecaf0800b309ee4171292361cded0f01ac25f41fa68f3c3fe034f96423c016348ad88f1fc56bef53b33a5017945a975fc2167c94efb6e1f798773652000b2a180bcb3eb55b66bd7ae8eab3da41b68cdf9e2c6cf7104935be;
    5'b10010 : xpb = 1024'h8f390ade3a9c6b2be37652684d4f173d1ecb3c53aa8b34fa16fbb2643ae1f267f186fbd346717521565bc06420254558882171269a3872f05b74c987b02989f88292c6ef9d0d156c740fc6bc18bffcd869509b3344c686813a380299aa4ba7d04ced6d0d4affdb94bed35c5b78a28b748d44c339ce4636c664dea4454cbe691b;
    5'b10011 : xpb = 1024'h661a4d8ba4712992fed0b5b25b48a129e48b1420152a9991754c5e27538a335d45250368206d115f20aa3980a9e28ba53aff970543d106935a245f917ef162ffb0a15fcc66c9175f4aacfbb5d338462c2b61ecb668ac4891fcccf6a3aab5cb16d25c119ee52b9483eb1b93229e0e3344e2c4f3b70a8a837ce521608f0051360d;
    5'b10100 : xpb = 1024'h3cfb90390e45e7fa1a2b18fc69422b16aa4aebec7fc9fe28d39d09ea6c32745298c30afcfa68ad9ceaf8b29d339fd1f1edddbce3ed699a3658d3f59b4db93c06deaff8a930851952214a30af8db08f7fed733e398c920aa2bf61eaadab1fee5d57cab6307f574d731763c9e9c379db153845243446ced03365641cd8b3e402ff;
    5'b10101 : xpb = 1024'h13dcd2e6781aa66135857c46773bb503700ac3b8ea6962c031edb5ad84dab547ec611291d46449dab5472bb9bd5d183ea0bbe2c297022dd957838ba51c81150e0cbe9185fa411b44f7e765a94828d8d3af848fbcb077ccb381f6deb7ab8a11a3dd395ac21983066243ac00b0e8e582e58dc554b183131ce9e5a6d9226776cff1;
    5'b10110 : xpb = 1024'h9b6b5ae9a3dd99911be55767958f8641a7409eb62a8067cf0e1b1ac65085a3454347979f788664a71ef3e41d2a786f55b7b43087634d91c806d2610d261b62c6af1c5f11738e1a7ce11e9d459b7ce658659adad860e3bbd4fa1864bc661ed77c91af917d6477b7def6b41e57062150df321f64110fa2c6d0ac591070a3ec034e;
    5'b10111 : xpb = 1024'h724c9d970db257f8373fbab1a389102e6d007682951fcc666c6bc689692de43a96e59f34528200e4e9425d39b435b5a26a9256660ce6256b0581f716f4e33bcddd2af7ee3d4a1c6fb7bbd23f55f52fac27ac2c5b84c97de5bcad58c66688fac3171e360efea370ce22fc551e2b8cf8af879f948e4be713872c9bccba577ed040;
    5'b11000 : xpb = 1024'h492de0447787165f529a1dfbb1829a1b32c04e4effbf30fdcabc724c81d6252fea83a6c92c7d9d22b390d6563df2fbef1d707c44b67eb90e04318d20c3ab14d50b3990cb07061e628e590739106d78ffe9bd7ddea8af3ff67f424cd066f31e099c8cdaa098cf29bd4f448be550f8a07fdd1fc50b882b603dacde89040b119d32;
    5'b11001 : xpb = 1024'h200f22f1e15bd4c66df48145bf7c2407f880261b6a5e9595290d1e0f9a7e66253e21ae5e067939607ddf4f72c7b0423bd04ea22360174cb102e1232a9272eddc394829a7d0c2205564f63c32cae5c253abcecf61cc95020741d740da675d415021fb7f3232fae2ac7b8cc2ac76644850329ff588c46facf42d21454dbea46a24;
    5'b11010 : xpb = 1024'ha79daaf50d1ec7f654545c66ddcff5462fb60118aa759aa4053a8328662954229508336baa9b542ce78c07d634cb9952e746efe82c62b09fb22ff8929c0d3b94dba5f7334a0f1f8d4e2d73cf1e39cfd861e51a7d7d00f128b9f8c6df21f20728d671b5ed7def94292e94e05293a01649d6fa04e850ff56daf3d37c9bfb199d81;
    5'b11011 : xpb = 1024'h7e7eeda276f3865d6faebfb0ebc97f32f575d8e51514ff3b638b2eeb7ed19517e8a63b008496f06ab1da80f2be88df9f9a2515c6d5fb4442b0df8e9c6ad5149c09b4901013cb218024caa8c8d8b2192c23f66c00a0e6b3397c8dbae9225c2a6f5be05a7f181b4d185add1719b90bbe1a2c7a35658d43a391741638e5aeac6a73;
    5'b11100 : xpb = 1024'h5560304fe0c844c48b0922faf9c3091fbb35b0b17fb463d2c1dbdaae9779d60d3c4442955e928ca87c28fa0f484625ec4d033ba57f93d7e5af8f24a6399ceda337c328ecdd872372fb67ddc2932a627fe607bd83c4cc754a3f22aef322c64db5e14eff10b247060787254de0de7765ea81fa65e2c987f047f458f52f623f3765;
    5'b11101 : xpb = 1024'h2c4172fd4a9d032ba663864507bc930c80f5887dea53c86a202c8671b02217028fe24a2a388e28e64677732bd2036c38ffe16184292c6b88ae3ebab00864c6aa65d1c1c9a7432565d20512bc4da2abd3a8190f06e8b2375b01b7a2fd233070fc66bda3a24c72bef6b36d84a803e30dbad77a966005cc3cfe749bb17915d20457;
    5'b11110 : xpb = 1024'h322b5aab471c192c1bde98f15b61cf946b5604a54f32d017e7d3234c8ca57f7e38051bf1289c52410c5ec485bc0b285b2bf8762d2c4ff2bacee50b9d72c9fb193e05aa670ff2758a8a247b6081af5276a2a608a0c97f96bc44c9707239a9442ec2c4833e69e77e5dfb5bb6f294eb58b2cfac6dd421089b4f4de6dc2c964d149;
    5'b11111 : xpb = 1024'h8ab13dade034b4c2a81dc4b03409ee377deb3b47950a32105aaa974d947545f53a66d6ccb6abdff07a72a4abc8dc099cc9b7d5279f10631a5c3d2621e0c6ed6a363e2831ea4c269091d97f525b6f02ac2040aba5bd03e88d3c6e1d0bde2f5a1ba0a27eef3193296292bdd915468a8384d154d63ccea0339bbb90a51105da04a6;
    endcase
end

endmodule

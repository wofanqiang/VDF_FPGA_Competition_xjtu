module xpb_5_70
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'habdc29827794f14340fe07dfefd539c6d34cfcc7faaa4199747d85a63407c9a69924b2bc6981df24c3379c4dbaa771f05315d03e7f641fd483e359c9f089b0cf194b9aecb25b3770cafbfbdcb5ca3c899b26e333e9a664799a8e2fbd7c4be896846de0a78e70854dbc9371701ab1d23eea1d642704797b64a7a4370e214e8adb;
    5'b00010 : xpb = 1024'ha70b0daf2d3badbdb6f697e8cf502c3c3523f65f1fdce2bb6b1e51f6b50ce6452f00e80008dd3fbae710f95491f0d31642117896dc156f5d57277435a640ececbe48012ab525719c835df516d2b8b4e24248cccf46c69be27f8fcd803e6d2e9ad9d42f256c18120df266fc013d937e548560e96bb8a7999908d8f317b9baaf4b;
    5'b00011 : xpb = 1024'ha239f1dbe2e26a382cef27f1aecb1eb196faeff6450f83dd61bf1e47361202e3c4dd1d43a838a0510aea565b693a343c310d20ef38c6bee62a6b8ea15bf8290a63446768b7efabc83bbfee50efa72d3ae96ab66aa3e6d34b64916b43008e749f2f3a7da349bf9ece283a869260752a6a20a46eb06cd5b7cd6a0daf215226d3bb;
    5'b00100 : xpb = 1024'h9d68d608988926b2a2e7b7fa8e461126f8d1e98d6a4224ff585fea97b7171f825ab95287479400e72ec3b362408395622008c94795780e6efdafa90d11af65280840cda6bab9e5f3f421e78b0c95a593908ca00601070ab449930905c2afbaa384a0cc2127672b8e5e0e11238356d67fbbe7f3f52103d601cb426b2aea92f82b;
    5'b00101 : xpb = 1024'h9897ba354e2fe32d18e048036dc1039c5aa8e3248f74c6214f00b6e8381c3c20f09587cae6ef617d529d106917ccf6880f04719ff2295df7d0f3c378c766a145ad3d33e4bd84201fac83e0c529841dec37ae89a15e27421d2e94a6c884d100a7da071a9f050eb84e93e19bb4a6388295572b7939d531f4362c77273482ff1c9b;
    5'b00110 : xpb = 1024'h93c69e6203d69fa78ed8d80c4d3bf611bc7fdcbbb4a7674345a18338b92158bf8671bd0e864ac21376766d6fef1657adfe0019f84edaad80a437dde47d1ddd6352399a22c04e5a4b64e5d9ff46729644ded0733cbb4779861396448b46f246ac2f6d691ce2b6450ec9b52645c91a2eaaf26efe7e8960126a8dabe33e1b6b410b;
    5'b00111 : xpb = 1024'h8ef5828eb97d5c2204d168152cb6e8871e56d652d9da08653c424f893a26755e1c4df25225a622a99a4fca76c65fb8d3ecfbc250ab8bfd09777bf85032d51980f7360060c31894771d47d33963610e9d85f25cd81867b0eef897e24e09138cb084d3b79ac05dd1ceff88b0d6ebfbdac08db283c33d8e309eeee09f47b3d7657b;
    5'b01000 : xpb = 1024'h8a2466bb6f24189c7ac9f81e0c31dafc802dcfe9ff0ca98732e31bd9bb2b91fcb22a2795c501833fbe29277d9da919f9dbf76aa9083d4c924ac012bbe88c559e9c32669ec5e2cea2d5a9cc73804f86f62d1446737587e857dd998010cb34d2b4da3a06189e055e8f355c3b680edd86d628f60907f1bc4ed350155b514c4389eb;
    5'b01001 : xpb = 1024'h85534ae824cad516f0c28826ebaccd71e204c981243f4aa92983e82a3c30ae9b48065cd9645ce3d5e202848474f27b1fcaf3130164ee9c1b1e042d279e4391bc412eccdcc8ad08ce8e0bc5ad9d3dff4ed436300ed2a81fc0c29b1dd38d5618b92fa054967baceb4f6b2fc5f931bf32ebc4398e4ca5ea6d07b14a175ae4afae5b;
    5'b01010 : xpb = 1024'h80822f14da71919166bb182fcb27bfe743dbc3184971ebcb2024b47abd35cb39dde2921d03b8446c05dbe18b4c3bdc45b9eebb59c19feba3f148479353facdd9e62b331acb7742fa466dbee7ba2c77a77b5819aa2fc85729a79cbb964f775ebd8506a3145954780fa103508a54a0df015f7d13915a188b3c127ed3647d1bd2cb;
    5'b01011 : xpb = 1024'h7bb1134190184e0bdcb3a838aaa2b25ca5b2bcaf6ea48ced16c580cb3e3ae7d873bec760a313a50229b53e9223853d6ba8ea63b21e513b2cc48c61ff09b209f78b279958ce417d25fecfb821d71af000227a03458ce88e928c9e59591198a4c1da6cf19236fc04cfd6d6db1b77828b16fac098d60e46a97073b38f6e1587f73b;
    5'b01100 : xpb = 1024'h76dff76e45bf0a8652ac38418a1da4d20789b64693d72e0f0d664d1bbf400477099afca4426f05984d8e9b98face9e9197e60c0a7b028ab597d07c6abf6946153023ff96d10bb751b731b15bf4096858c99bece0ea08c5fb719ff71bd3b9eac62fd3401014a391900caa65ac9a64372c96041e1ac274c7a4d4e84b77adf41bab;
    5'b01101 : xpb = 1024'h720edb9afb65c700c8a4c84a699897476960afddb909cf310407196c404521159f7731e7e1ca662e7167f89fd217ffb786e1b462d7b3da3e6b1496d675208232d52065d4d3d5f17d6f93aa9610f7e0b170bdd67c4728fd6456a194de95db30ca85398e8df24b1e50427df03dbd45e3423147a35f76a2e5d9361d07814660401b;
    5'b01110 : xpb = 1024'h6d3dbfc7b10c837b3e9d5853491389bccb37a974de3c7052faa7e5bcc14a3db43553672b8125c6c4954155a6a96160dd75dd5cbb346529c73e58b1422ad7be507a1ccc12d6a02ba927f5a3d02de6590a17dfc017a44934cd3ba332a157fc76ceda9fdd0bcff2ab1078517acee0278f57cc8b28a42ad1040d9751c38adecc648b;
    5'b01111 : xpb = 1024'h686ca3f466b33ff5b495e85c288e7c322d0ea30c036f1174f148b20d424f5a52cb2f9c6f2081275ab91ab2ad80aac20364d9051391167950119ccbade08efa6e1f193250d96a65d4e0579d0a4ad4d162bf01a9b301696c3620a4d0641a1dbcd330062b89ad9a37d0ae25056003093b6d67ceade8deff2241f8867f94773888fb;
    5'b10000 : xpb = 1024'h639b88211c59fc702a8e786508096ea78ee59ca328a1b296e7e97e5dc35476f1610bd1b2bfdc87f0dcf40fb457f4232953d4ad6bedc7c8d8e4e0e6199646368bc415988edc34a00098b9964467c349bb6623934e5e89a39f05a66e26dc3f02d7856c7a078b41c490e3f88ff125eae7830312332d932d407659bb3b9e0fa4ad6b;
    5'b10001 : xpb = 1024'h5eca6c4dd200b8eaa087086de784611cf0bc963a4dd453b8de8a4aae4459938ff6e806f65f37e88700cd6cbb2f3d844f42d055c44a791861b82500854bfd72a96911feccdefeda2c511b8f7e84b1c2140d457ce9bba9db07eaa80be99e6048dbdad2c88568e9515119cc1a8248cc93989e55b872475b5eaabaeff7a7a810d1db;
    5'b10010 : xpb = 1024'h59f9507a87a77565167f9876c6ff539252938fd17306f4dad52b16fec55eb02e8cc43c39fe93491d24a6c9c20686e57531cbfe1ca72a67ea8b691af101b4aec70e0e650ae1c91458097d88b8a1a03a6cb467668518ca1270cfa9a9ac60818ee0303917034690de114f9fa5136bae3fae39993db6fb897cdf1c24b3b1407cf64b;
    5'b10011 : xpb = 1024'h552834a73d4e31df8c78287fa67a4607b46a8968983995fccbcbe34f4663cccd22a0717d9deea9b3488026c8ddd0469b20c7a67503dbb7735ead355cb76beae4b30acb48e4934e83c1df81f2be8eb2c55b89502075ea49d9b4ab476f22a2d4e4859f658124386ad185732fa48e8febc3d4dcc2fbafb79b137d596fbad8e91abb;
    5'b10100 : xpb = 1024'h505718d3f2f4ee5a0270b88885f5387d164182ffbd6c371ec26caf9fc768e96bb87ca6c13d4a0a496c5983cfb519a7c10fc34ecd608d06fc31f14fc86d23270258073186e75d88af7a417b2cdb7d2b1e02ab39bbd30a814299ace531e4c41ae8db05b3ff01dff791bb46ba35b17197d97020484063e5b947de8e2bc471553f2b;
    5'b10101 : xpb = 1024'h4b85fd00a89baad47869489165702af278187c96e29ed840b90d7bf0486e060a4e58dc04dca56adf9032e0d68c6308e6febef725bd3e568505356a3422da631ffd0397c4ea27c2db32a37466f86ba376a9cd2357302ab8ab7eae82f4a6e560ed306c027cdf878451f11a44c6d45343ef0b63cd851813d77c3fc2e7ce09c1639b;
    5'b10110 : xpb = 1024'h46b4e12d5e42674eee61d89a44eb1d67d9ef762e07d17962afae4840c97322a8e43511487c00cb75b40c3ddd63ac6a0cedba9f7e19efa60dd879849fd8919f3da1fffe02ecf1fd06eb056da1155a1bcf50ef0cf28d4af01463b020b76906a6f185d250fabd2f111226edcf57f734f004a6a752c9cc41f5b0a0f7a3d7a22d880b;
    5'b10111 : xpb = 1024'h41e3c55a13e923c9645a68a324660fdd3bc66fc52d041a84a64f14914a783f477a11468c1b5c2c0bd7e59ae43af5cb32dcb647d676a0f596abbd9f0b8e48db5b46fc6440efbc3732a36766db32489427f810f68dea6b277d48b1be7a2b27ecf5db389f789ad69dd25cc159e91a169c1a41ead80e807013e5022c5fe13a99ac7b;
    5'b11000 : xpb = 1024'h3d12a986c98fe043da52f8ac03e102529d9d695c5236bba69cefe0e1cb7d5be60fed7bcfbab78ca1fbbef7eb123f2c58cbb1f02ed352451f7f01b97744001778ebf8ca7ef286715e5bc960154f370c809f32e029478b5ee62db35c3ced4932fa309eedf6787e2a929294e47a3cf8482fdd2e5d53349e321963611bead305d0eb;
    5'b11001 : xpb = 1024'h38418db37f369cbe504b88b4e35bf4c7ff7462f377695cc89390ad324c827884a5c9b1135a12ed381f9854f1e9888d7ebaad9887300394a85245d3e2f9b7539690f530bcf550ab8a142b594f6c2584d94654c9c4a4ab964f12b4f9ffaf6a78fe86053c745625b752c8686f0b5fd9f4457871e297e8cc504dc495d7f46b71f55b;
    5'b11010 : xpb = 1024'h337071e034dd5938c64418bdc2d6e73d614b5c8a9c9bfdea8a317982cd8795233ba5e656f96e4dce4371b1f8c0d1eea4a9a940df8cb4e4312589ee4eaf6e8fb435f196faf81ae5b5cc8d52898913fd31ed76b36001cbcdb7f7b697c2718bbf02db6b8af233cd4412fe3bf99c82bba05b13b567dc9cfa6e8225ca93fe03de19cb;
    5'b11011 : xpb = 1024'h2e9f560cea8415b33c3ca8c6a251d9b2c3225621c1ce9f0c80d245d34e8cb1c1d1821b9a98c9ae64674b0eff981b4fca98a4e937e96633b9f8ce08ba6525cbd1daedfd38fae51fe184ef4bc3a602758a94989cfb5eec0520dcb8358533ad050730d1d9701174d0d3340f842da59d4c70aef8ed2151288cb686ff50079c4a3e3b;
    5'b11100 : xpb = 1024'h29ce3a39a02ad22db23538cf81cccc2824f94fb8e701402e77731223cf91ce60675e50de38250efa8b246c066f64b0f087a0919046178342cc1223261add07ef7fea6376fdaf5a0d3d5144fdc2f0ede33bba8696bc0c3c89c1b9d347f5ce4b0b863827edef1c5d9369e30ebec87ef8864a3c72660556aaeae8340c1134b662ab;
    5'b11101 : xpb = 1024'h24fd1e6655d18ea8282dc8d86147be9d86d049500c33e1506e13de745096eafefd3a8621d7806f90aefdc90d46ae1216769c39e8a2c8d2cb9f563d91d094440d24e6c9b500799438f5b33e37dfdf663be2dc7032192c73f2a6bb710ab7ef910fdb9e766bccc3ea539fb6994feb60a49be57ff7aab984c91f4968c81acd22871b;
    5'b11110 : xpb = 1024'h202c02930b784b229e2658e140c2b112e8a742e73166827264b4aac4d19c079d9316bb6576dbd026d2d726141df7733c6597e240ff7a2254729a57fd864b802ac9e32ff30343ce64ae153771fccdde9489fe59cd764cab5b8bbd0ecd7a10d7143104c4e9aa6b7713d58a23e10e4250b180c37cef6db2e753aa9d8424658eab8b;
    5'b11111 : xpb = 1024'h1b5ae6bfc11f079d141ee8ea203da3884a7e3c7e569923945b55771552a1243c28f2f0a9163730bcf6b0831af540d46254938a995c2b71dd45de72693c02bc486edf9631060e0890667730ac19bc56ed31204368d36ce2c470beac903c321d18866b1367881303d40b5dae723123fcc71c07023421e105880bd2402dfdfacffb;
    endcase
end

endmodule

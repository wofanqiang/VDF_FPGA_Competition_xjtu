module xpb_5_280
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h63350e0debf7ca1cf0735dd8be6a1f619cc73fd3d4d62853e7ef12cbd23e7391e77864b9e26d3c167ba851682e16c1c673c1a4c68ad8ed63868b91a2326e5586c4f7d392adeea583014eda2198cfc6ded9c59962f260d6abf5c3b2a87aa6267f9a9d9e02784f9e2beb54e0aa53c89056d01f97752c1437823bb0f241e70d838f;
    5'b00010 : xpb = 1024'h15bcd6c616015f7115e143da6c79f771c8187c76d434b03052016c41f17a3a1bcba84bfafab3f99e57f2638978cf72c2836921a6f2ff0a7b5c77e3e62a0a365c15a07276ac4c4dc0f003b1a098c3c98cbf86392d583b804735fad3563b21aa6d0633a9db3fd643ca4fe9da75afc0fa845165500807dd11d430f2697f4538a0b3;
    5'b00011 : xpb = 1024'h78f1e4d401f9298e0654a1b32ae416d364dfbc4aa90ad88439f07f0dc3b8adadb320b0b4dd2135b4d39ab4f1a6e63488f72ac66d7dd7f7dee30375885c788be2da9846095a3af343f1528bc23193906b994bd2904a9c56f32bbe85feb5c7d0eca0d147ddb825e1f63b3ebb2003898adb2184e77d33f149566ca35bc12c462442;
    5'b00100 : xpb = 1024'h2b79ad8c2c02bee22bc287b4d8f3eee39030f8eda8696060a402d883e2f47437975097f5f567f33cafe4c712f19ee58506d2434de5fe14f6b8efc7cc54146cb82b40e4ed58989b81e0076341318793197f0c725ab077008e6bf5a6ac764354da0c6753b67fac87949fd3b4eb5f81f508a2caa0100fba23a861e4d2fe8a714166;
    5'b00101 : xpb = 1024'h8eaebb9a17fa88ff1c35e58d975e0e452cf838c17d3f88b48bf1eb4fb532e7c97ec8fcafd7d52f532b8d187b1fb5a74b7a93e81470d7025a3f7b596e8682c23ef038b88006874104e1563d62ca5759f858d20bbda2d7d73a61b95954f0e97b59a704f1b8f7fc25c08b289595b34a855f72ea37853bce5b2a9d95c540717ec4f5;
    5'b00110 : xpb = 1024'h4136845242041e5341a3cb8f456de655584975647c9e1090f60444c5d46eae5362f8e3f0f01becdb07d72a9c6a6e58478a3b64f4d8fd1f721567abb27e1ea31440e1576404e4e942d00b14e1ca4b5ca63e92ab8808b280d5a1f07a02b164ff47129afd91bf82cb5eefbd8f610f42ef8cf42ff0181797357c92d73c7dcfa9e219;
    5'b00111 : xpb = 1024'ha46b92602dfbe8703217296803d805b6f510b538517438e4ddf35791a6ad21e54a7148aad28928f1837f7c0498851a0dfdfd09bb63d60cd59bf33d54b08cf89b05d92af6b2d38ec5d159ef03631b2385185844eafb13578197b42cab2c0b25c6ad389b9437d2698adb12700b630b7fe3c44f878d43ab6cfece882ebfb6b765a8;
    5'b01000 : xpb = 1024'h56f35b1858057dc457850f69b1e7ddc72061f1db50d2c0c14805b107c5e8e86f2ea12febeacfe6795fc98e25e33dcb0a0da4869bcbfc29ed71df8f98a828d9705681c9dab1313703c00ec682630f2632fe18e4b560ee011cd7eb4d58ec86a9b418cea76cff590f293fa769d6bf03ea11459540201f744750c3c9a5fd14e282cc;
    5'b01001 : xpb = 1024'h97b23d0820f13187cf2f56b5ff7b5d74bb32e7e5031489db2180a7de524aef912d1172d0316a4013c13a0472df67c061d4c037c3422470547cbe1dc9fc4ba45a72a68beaf8edf41aec39e01630328e0e3d9847fc6c8aab818226e06ad022da18464b345c6dfb4c7a43c63a21afc543ec6daf8b2fb3d21a2b90b1d3a730d9ff0;
    5'b01010 : xpb = 1024'h6cb031de6e06dd356d6653441e61d538e87a6e52250770f19a071d49b763228afa497be6e583e017b7bbf1af5c0d3dcc910da842befb3468ce57737ed2330fcc6c223c515d7d84c4b0127822fbd2efbfbd9f1de2b92981640de620af27a854211f0251483f2f52f38f91444c6ec4e49596fa902827515924f4bc0f7c5a1b237f;
    5'b01011 : xpb = 1024'h1f37fa969810728992d43945cc71ad4913cbaaf52465f8ce041976bfd69ee914de796327fdca9d9f940603d0a6c5eec8a0b5252327215180a443c5c2c9cef0a1bccadb355bdb2d029ec74fa1fbc6f26da35fbdad1f042aff4e1d415ce823d80e8a985d2106b5f891f4263e17cabd4ec3184048bb031a3376e9fd86b9b84640a3;
    5'b01100 : xpb = 1024'h826d08a484083ca68347971e8adbccaab092eac8f93c2121ec08898ba8dd5ca6c5f1c7e1e037d9b60fae5538d4dcb08f1476c9e9b1fa3ee42acf5764fc3d462881c2aec809c9d285a01629c39496b94c7d255710116501ab43e0f40562c9fe8e2535fb237f0596bddf7b1ec21e85df19e85fe0302f2e6af925ae78fb9f53c432;
    5'b01101 : xpb = 1024'h34f4d15cae11d1faa8b57d2038eba4badbe4276bf89aa8fe561ae301c8192330aa21af22f87e973debf8675a1f95618b241e46ca1a205bfc00bba9a8f3d926fdd26b4dac08277ac38ecb0142948abbfa62e5f6da773fab46841814b32345827b90cc06fc468c3c5c4410188d7a7e494769a598c30af7454b1aeff038fd7ee156;
    5'b01110 : xpb = 1024'h9829df6a9a099c179928daf8f755c41c78ab673fcd70d1523e09f5cd9a5796c2919a13dcdaebd35467a0b8c24dac235197dfeb90a4f9495f87473b4b26477c849763213eb61620469019db642d5a82d93cab903d69a081f279dbc75b9deba8fb2b69a4febedbda882f64f937ce46d99e39c53038370b7ccd56a0e27ae48c64e5;
    5'b01111 : xpb = 1024'h4ab1a822c413316bbe96c0faa5659c2ca3fca3e2cccf592ea81c4f43b9935d4c75c9fb1df33290dc43eacae39864d44da78768710d1f66775d338d8f1de35d59e80bc022b473c8847eceb2e32d4e8587226c3007cf7b2b8dba12e8095e672ce896ffb0d78662802693f9f3032a3f43cbbb0ae8cb12d4571f4be259b842b78209;
    5'b10000 : xpb = 1024'hade6b630b00afb88af0a1ed363cfbb8e40c3e3b6a1a58182900b620f8bd1d0de5d425fd7d59fccf2bf931c4bc67b96141b490d3797f853dae3bf1f315051b2e0ad0393b562626e07801d8d04c61e4c65fc31c96ac1dc0239afd69ab1d90d5368319d4ed9feb21e527f4ed3ad7e07d4228b2a80403ee88ea187934bfa29c50598;
    5'b10001 : xpb = 1024'h606e7ee8da1490dcd47804d511df939e6c152059a104095efa1dbb85ab0d976841724718ede68a7a9bdd2e6d113447102af08a18001e70f2b9ab717547ed93b5fdac329960c016456ed26483c6124f13e1f2693527b6abd4f00dbb5f9988d7559d335ab2c638c3f0e3e3cd78da003e500c7038d31ab168f37cd4c33787f022bc;
    5'b10010 : xpb = 1024'h12f647a1041e2630f9e5ead6bfef6bae97665cfca062913b643014fbca495df225a22e5a062d48027827408e5becf80c3a9806f868448e0a8f97c3b93f89748b4e54d17d5f1dbe835d873c02c60651c1c7b308ff8d9155703044dc0d5a045b4308c9668b8dbf698f4878c74435f8a87d8db5f165f67a434572163a74e61b3fe0;
    5'b10011 : xpb = 1024'h762b55aef015f04dea5948af7e598b10342d9cd07538b98f4c1f27c79c87d1840d1a9313e89a8418f3cf91f68a03b9d2ae59abbef31d7b6e1623555b71f7ca12134ca5100d0c64065ed616245ed618a0a178a2627ff22c1c26088eb5d4aa81c2a367048e060f07bb33cda7ee89c138d45dd588db228e7ac7adc72cb6cd28c36f;
    5'b10100 : xpb = 1024'h28b31e671a1f85a20fc72eb12c6963205f7ed9737497416bb631813dbbc3980df14a7a5500e141a0d019a417d4bc6acebe01289f5b439885ec0fa79f6993aae763f543f40b6a0c444d8aeda35eca1b4e8739422ce5ccd5b7663faf63952605b00efd1066cd95ad599862a1b9e5b9a301df1b416dfe575519a308a3f42b53e093;
    5'b10101 : xpb = 1024'h8be82c7506174fbf003a8c89ead38281fc461947496d69bf9e2094098e020b9fd8c2df0ee34e7db74bc1f58002d32c9531c2cd65e61c85e9729b39419c02006e28ed1786b958b1c74ed9c7c4f799e22d60fedb8fd82dac635c03620c0fcc2c2fa99aae6945e54b8583b7826439823358af3ad8e32a6b8c9bdeb9963612616422;
    5'b10110 : xpb = 1024'h3e6ff52d3020e51325a8728b98e35a92279755ea48cbf19c0832ed7fad3dd229bcf2c64ffb953b3f280c07a14d8bdd91416a4a464e42a30148878b85939de1437995b66ab7b65a053d8e9f43f78de4db46bf7b5a3e0855fe9c3a82b9d047b01d1530ba420d6bf123e84c7c2f957a9d8630809176063466edd3fb0d73708c8146;
    5'b10111 : xpb = 1024'ha1a5033b1c18af30161bd064574d79f3c45e95be1da219eff022004b7f7c45bba46b2b09de027755a3b459097ba29f57b52bef0cd91b9064cf131d27c60c36ca3e8d89fd65a4ff883edd7965905dabba208514bd30692caa91fe35624aedd69cafce584485bb8f4fd3a15cd9e9432ddd00a028eb32489e700fabffb5579a04d5;
    5'b11000 : xpb = 1024'h542ccbf3462244843b89b666055d5203efafd2611d00a1cc5a3459c19eb80c45889b124af64934dd7ffe6b2ac65b5053c4d36bed4141ad7ca4ff6f6bbda8179f8f3628e16402a7c62d9250e49051ae680645b4879643d645d23556100b695a8a1b64641d4d4234ee383656a5453b980a81e5e17e0e1178c204ed76f2b5c521f9;
    5'b11001 : xpb = 1024'h6b494ab702bd9d860f79c67b36d2a141b010f041c5f29a8c446b337bdf3d2cf6ccaf98c0e8ff2655c487d4c1114014fd47ae8cda967ca947aebc1afb543f874dfdec7c5626050041c4728639045b115ec065451fc1e7fe1126c76bdcbe4de7786fa6ff614c8da8c9ccb5070a1340238032b9a10e9da5313fa2eee3013f03f1d;
    5'b11010 : xpb = 1024'h69e9a2b95c23a3f5516afa4071d74975b7c84ed7f13551fcac35c6039032466154435e45f0fd2e7bd7f0ceb43f2ac316483c8d943440b7f801775351e7b24dfba4d69b58104ef5871d960285291577f4c5cbedb4ee7f568d08302966468b04f721980df88d1878b88820311af4fc928ed34b318615ee8a9635dfe071fafdc2ac;
    5'b11011 : xpb = 1024'h1c716b71862d394976d8e0421fe72185e3198b7af093d9d916481f79af6e0ceb387345870943ec03b43ae0d589e3741257e40a749c66d50fd763a595df4e2ed0f57f3a3c0eac9dc50c4ada0429097aa2ab8c8d7f545a002848674a14070688e48d2e19d1549f1e56ecb52ae650f4fcbc5490ea18f1b764e82b2157af5928dfd0;
    5'b11100 : xpb = 1024'h7fa6797f72250366674c3e1ade5140e77fe0cb4ec56a022cfe37324581ac807d1febaa40ebb1281a2fe3323db7fa35d8cba5af3b273fc2735def373811bc8457ba770dcebc9b43480d99b425c1d94181855226e246bad6d43e2afcbc81acaf6427cbb7d3cceebc82d80a0b90a4bd8d1324b0818e1dcb9c6a66d249f14036635f;
    5'b11101 : xpb = 1024'h322e42379c2e98ba8cba241c8c6118f7ab3207f1c4c88a0968498bbba0e84707041b918203f7e5a20c2d445f02b2e6d4db4d2c1b8f65df8b33db897c0958652d0b1facb2baf8eb85fc4e8ba4c1cd442f6b12c6acac95806f7e621d6a422833519361c3ac947562213c9f055c00b5f740a5f63a20f99476bc5c13c12e9e618083;
    5'b11110 : xpb = 1024'h95635045882662d77d2d81f54acb385947f947c5999eb25d50389e877326ba98eb93f63be66521b887d595c730c9a89b4f0ed0e21a3ecceeba671b1e3bc6bab3d017804568e79108fd9d65c65a9d0b0e44d8600f9ef6571b7425d012bcce59d12dff61af0cc5004d27f3e606547e87977615d19625a8ae3e97c4b370856f0412;
    5'b11111 : xpb = 1024'h47eb18fdb22ff82ba29b67f6f8db1069734a846898fd3a39ba4af7fd92628122cfc3dd7cfeabdf40641fa7e87b8259975eb64dc28264ea0690536d6233629b8920c01f2967453946ec523d455a910dbc2a98ffda04d100b6b45cf0c07d49ddbe99956d87d44ba5eb8c88dfd1b076f1c4f75b8a29017188908d062aade39a2136;
    endcase
end

endmodule

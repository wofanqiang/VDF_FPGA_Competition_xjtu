module reduction
#(
    parameter BIT_LEN_FLAG  = 18,
    parameter BIT_LEN_XPB   = 27,
    parameter NUM_XPB       = 38,
    parameter NUM_FLAG      = 64,
    localparam NUM_ELEMENTS_OUT = 62*17
)
(
    input logic [NUM_XPB-1:0][BIT_LEN_XPB-1:0] rest0,
    input logic [NUM_XPB-1:0][BIT_LEN_XPB-1:0] rest1,
    input logic [NUM_FLAG-1:0][BIT_LEN_FLAG-1:0] xpb_flag,

    output logic [NUM_ELEMENTS_OUT-1:0] C,
    output logic [NUM_ELEMENTS_OUT-1:0] S
);

    logic [NUM_XPB-1:0][BIT_LEN_XPB-1:0] xpb_primes[NUM_FLAG];
    //initial begin
    //    $readmemh("reduction_lut.mem", xpb_primes);
    //end

    assign xpb_primes[0] = 1026'h4f52baaa3e11cb3734fa8828efa5b8ae8e89fccf2a885f88822346aa4cfd52f7fcb7828735d9817160a1c0b91ca1ef359be5d819dd4d2fb44f60c0a1c52d8b4e8bb0cb51506f02baed65fd5d67243bcf0bfb06677379d2ef4a736e0545d55d6dd0f86dd64f37077279401921082fd9d6b126211dafb4a2cfb99084fb771d9995;
assign xpb_primes[1] = 1026'h8f5f5ff592b6d170525b195370ed22a392f6de92c951589978457f3251d3148450ac12a67c24ee775fbeb120aa758bf317ba1c18315177d432dc0ca796e6b3c26b8379a6639a71fd02370fe8b9ae67090934055d36ad60f1f80219ba6c4b40881e5500f9497dd5ae27928078a33930c7ae11c671e99d1711f5cfb6d5705511cb;
assign xpb_primes[2] = 1026'h48978a828bed9255febb322bffef938c78cfdcee5e1f81a13708f0f21d3cd4240ac962138b203e0e6806c3ff791df52554d6fcea4160cdbc6472bacdbe68a586368813fbcf2c5dd172f296ce8093af1dc7b33ba92dd8059d62b8af5936de839df45631343f167d26a4b9feb7eadfe94e2b0afd711d91860e973ef090d1e4ef2c;
assign xpb_primes[3] = 1026'h1285494887e7e5315c07937d1771f2a541e981347fb37cf29acfe029bb5bf9f0189bee12ae2958f3b37b8fb143fa793fc37f13ca2ef23637f926ebf70e0c027e79aafa2f54a33d4602e6a80ef6995d40c8bf926660fe8461655526f5b2384c6ae7ba9fd9349decf31796289814e0703c4e0cbe2bbdff5cfc9148bfd5e3329eb6;
assign xpb_primes[4] = 1026'haf78fe60ef57e3e768839bd9483903eec9ebc1969ec448bffb84ec69d343f42fa8bf8ac9b1fd56b42854968899306913dfd911fc39df242de57045f9284043b8dd8e4e3e30438bd000b280f1201762471dcd73ff63ce3aeaeeccf96b6ab2f413446125c92832dbbd9434c9834088912eb5aac0337d56e4bd5ebcaa06eefd6f87;
assign xpb_primes[5] = 1026'h6f2e7c4e9c199031451cf0c8947fbf55b6eab722c8535c99eef779c9b1a78ce991c7fb7fa2b907fd39a46532b3119a4767838405d437d1f4d95525ed090256325fb8fb6e396a5367f27242490ba376851e2d514ad845d2dacfc72aa6c3e5e53363af5c6b243419265770d0163ef011e31f7ab46b76499f305754660c18d9a9aa;
assign xpb_primes[6] = 1026'h858fcf85a177aba559c33e6cbf550f36d535849c90003a48bd596568c5a943de2504d596294656f91e65e04e7b10f59694c065d7f2fdcfb97f0b2ba07882c07d9f206fe1fded8c012b2d0f40a55857dcb7ab0fff6ed1cdf0103ba6a9cd9727aa03834be6e26a1fbfee4cf29fed1ed5b5f7f0bb60c471c2a2d19676a3d249691a;
assign xpb_primes[7] = 1026'h5c0d413a27845a21e62d32ebfada5716df220a0f07210e53c92db05b203b6a2e787dc596e85b6138fcd568a48a6491bc7f0d0f168c92df1f1c006f2231099b8c6cb06e54f351174481958b81a1eb3c542679add16696719def59809ad3c25ef936ec04cc4c452286cbe296c7459676bcae739213346900e8c370f6514fea526;
assign xpb_primes[8] = 1026'h1f6753335bec392ce73389d6a9c5da14a5c4aebd3b6330ff5a298342fca90d78fc27034132612dd1b5cd9f75edf7a1a4bdd1a0c7debb359b6eefcf2486c00f16f5484e131daa14a091cc4570f79fa4aaf2c8f18c013c6b586c819a608d10c9b56e60ba794dc101f9cb7bdb674c9b5d1fd9f2817a77a77797d4333a632bc8801c;
assign xpb_primes[9] = 1026'h5e13f69303a83973570e68e48c7510e2f8e217b4067c9a1e12c7c95a746d721b3e9ff76de2803a661f0f69d5eff379439146c73ab87925cb52234f3913e06187001cee3cefa898b6b958204691bcbaa32a59ceec9825bb69875067f9b176437794f63780e2d04f83f8fd7040c4dedeb441e09de1d4c4222c8d9c3fe3fced9095;
assign xpb_primes[10] = 1026'h5d508fea213ef5688fec171dcde47acff5625430409a437681c926cc4ac7ab0d5ac07c7a1f89e89d6cc83771f29781e6b83ac72591e68b7a657ef9fede39c5a1a60ee3c0a93c936d84ab62b39c02a73e9812873fa08c92891e49c756b38f772a0eafb6937c4493fb5c48957c32479d5d914290161a4d7d57a874f8bf513804a;
assign xpb_primes[11] = 1026'h81fb9cfcbf5d18e6c47c9d7e39c8d468fa4c1cdc04ed2d0044f5ab29f629b5f09496fcc936950f7ff44cf66cc8ad1aefc6e6774e77c36da53c3709713854460e6a03d53cc655d35d15cdebdd43327fc6c4d62c3aeef39b6d5380038c026e0f8f3ce283072e6743f603d82a794c46d41ddc565ef0d62237485f3f1b85dec54bde;
assign xpb_primes[12] = 1026'ha65e699a845ebe4f35411f5ff2b5dc97c6d225218f01f7d79a181527d1ebc8e94603bc282ef469972dda71398346e1367a3bce24a3d1b9922192f83775ace09647432c135e309356ff2deb5e520649ff2e7c29d2a1777afe2b248b02f75d4555f03bc8d132433994e36c310780b51cc9266fc8832a78803a9a977769076d3b46;
assign xpb_primes[13] = 1026'h8100e6e2bf75c328926dfdbfb39f4bd5e980c5fe049a2a46d9c51e1627b3d4d893034233141601d18387a59a3b0dcab1d9e4fd8a709bb724073794d22727db5aad0f3ffc37b248b38a862bebb121ab687514d748c45d3e5fb9999cdeff4051a56f7da075f6103d72396256f557b3c13f80245d791194aa883b44248f1569bca0;
assign xpb_primes[14] = 1026'h458d0affd26c0ba1b745eef54195fbf8ddc330f8ead034556fe61145b9527a7b206b4bb75cc27084817cc903af8ea52b68e0e67b9dea063a1bf28b19711c55ecf56176322e0bbeaa400e405a28880d508ab3ab446be014943a7081b37072b51d8a91da5e7f2c8605609d043423449d8ac15e5537c6b27f2c6cd0c38e1affaeb8;
assign xpb_primes[15] = 1026'ha72da027db07fc3f5ca2e0a03df3a43c9fab8ef13520bb204985b8e8f9efbd0dab549cc8650d4bc2c119d4650fa98e5bd2168ee67b9403c151cbfc4cd7ddc023817fb59440cc831433530dac3afd2a813cd9eccdd595710f0d00ba6acf02120acc72f6b3169c3ec9db1264957a9e8e9dd963ad14860418cedaf6a01ad712da6;
assign xpb_primes[16] = 1026'h65d6b3de4c47c0196984972e5722411325c38b14de68874cf12dad7f019cc7cf2bca187115f687e7fbfec6a71cbd1a65fdeec68dec778688d9f1fcf4bdf947576c8e7313e17e30142cafbe5d7f5f016efaf8a0ebfba36cb744357b85a1612180709bf68bf2fbb657704b8672b2a04e7a0f173a9369475aba3aadb495dc810e53;
assign xpb_primes[17] = 1026'h57db60b385870cc54b9a57617f08ceeb5b3213ea5b33c1d9c3b1d090cce727d34284c95a39504b12a5f9dfe3470eba0149f6d214cb634232149b39c0eaba3a988adb158509bf1592c30b4ee8412ccad1f99ef3df3740d22ffecda8de9680bd5281bf28336dedb12c989d80afbec5e550d8ee0aa023f18b586ae999b8a5364c0b;
assign xpb_primes[18] = 1026'h8e603f0d17df9cfb2091847834c500d2cfac573a688670a0ea7714a3f85c7af5ac9b1f64c96ba8085e4c27e158c3aadb78d73fe83a27c27032d6386842ced18f9d1f1036b2a2a2149e8d98df94c75bae2d1aed4ffaf24d6ca25697772fb22ce482d3915fa2d740658add618a318dc0c67b0ba81402e4e0e63852c9e19e4639a2;
assign xpb_primes[19] = 1026'haf5bb62f5a58e64e5cdabaff0e9ed11f1ca5150c6829ef4b6174068aad90a239e8830508b6190df6298ca3e0f792f9e93f83bed00c8182f97a7ffa1c789e500244dc650fee6b4e33775e85fac45503c01f54790ae21718272fb9cee78aa9898d7fdd24068aac44862d4910668bbac808d3d974e7ac80d7011276a8a4720960d;
assign xpb_primes[20] = 1026'h9811fdd24de17adbd3b805de8716fb1f5cd03829fcd35963651b8213194c24981c8060bf473f97d0656695b1adebec717132e6f63da42b90dde9208bba625d0bd13aea29cf3b235311b7a8d02d2b69450922bda425e1b9519fa8f4c8f332c982161101553a2b4717c7aadc7d58a52ea10b84a656217aab31f4b3c83e06216dea;
assign xpb_primes[21] = 1026'h4ac4626754c0baa46fb8e607d3f6f4e283fd5fd7f4377459ffec2aaeaf0d0d1e4b83289417e2846fe77c50af7fd6a69a3435987037d9feb6e12af845603f3dc4703f3edb0184eb4c09d11316963490436d987c3ac695ebac87a0811941e843a7b36bda9e80875e1b97cd73344c0b4f350f42e7a4a1d81f741f832db17434805;
assign xpb_primes[22] = 1026'h82602f84743de76a64b874bb7852bbd58433cb5cc8e8ae2f76f09397ff691af3f19fbd9b636085f5d8113a387d43f25768edd52976debb6012f8ba3f8258a3772f7c1b1b9c64780c493b255d029a2eeb442c0d742cd76cba0ef2bba08337e73cbed2e79d6ace46d74c3ac2ba41c1f6a2cb30f027e792d456c45ea32146cb5b52;
assign xpb_primes[23] = 1026'h45cabd8aedb1c9bf517eeb251a959781b938096514ed5381db30c1e66ce525d708f8f7f887f7d671edf1ad8bdacafe6b081c49dbab51d0c00d8b44c51871511e28a8c0f0662e17683a8268b755a380d49b41f399fb058ad486f70a9a4e16da7914c58a1192ca48ec610ac5ab1c537360585bb140ce9eff6952a5f6490418693a;
assign xpb_primes[24] = 1026'h970edaed224b0098c45c8c7fdc2b5a8c96c4d534e47d4f31e260e51d6e7a7d59ead0623ac367ae7b2599f474ec122aa2e9b1c5b9dc704eccb9b9fee9dd8b1f2dee81ca27e2b8a312a4d9b60361e989baf9033106148e9a7fc6e0469986022be358e9b5a9cb7af2606f30915eb49a8e2bc22b514e747341a659a1b30bf509f740;
assign xpb_primes[25] = 1026'hb30558d6a92c5fee948c87234f11b233b890193a4d0305aa0971f6fc14e07f38957403275c0ed134179e24c75539d230985a33f148665984df9db4469ac82fe3b5ba75db9ee729a6cd135ac1703b460f8359ba1ac63e12e037b6c387bf3f4c3db15a896dc2aec1b7035d736ff76156ef809ae55041cac71b89df2f9ba19bbea;
assign xpb_primes[26] = 1026'h7956dcb9f4e6747b3b9af91c0746328764f7d6575e2e9f098e969c14352512e40e20e347c2174adcc0ed5c538c7db125c6788f9fcdb745f14b6e503de69d0d5056bb6438b4615e2b520abe5373850d43a5f6fadbb41eed38aee40adc0b38da9e87b6d8a6245c53ded89cb9e19a48accadce3b6b60d7218103f8afd2d6b836adc;
assign xpb_primes[27] = 1026'h59bd74a295d9c1c8f97259084424fdd511a0c2c7235bbbfdf05ea19e32d8a0af4ea78093e1d7df17a640dc6187bf6d9de9fdd2396b22ffcc83d380f2537386b295168f7fd754a9de8d944c900d760660b8594d08f5bef049769cf087715bc0708d1aa0f33bc65be910c765b2238af086cef4c3960baa55f68e23c679cc067b4a;
assign xpb_primes[28] = 1026'h94b302b73900ecef3f08161455f13e4004667e0d77001de8b7127fdd0c7a56813079bc4ccd65084aa9f95b6bffab4a753664c48c5b91f3d5ec343ca3dc8c19a6dcda2e1dc9041d38176cd025e49f39ff40485cd55ef150dc798faff34b451be0d0028f8f3f9bd468ffab4c55f5196d68a20a2e856cdd9eea337ac7c3014b53bb;
assign xpb_primes[29] = 1026'h1b3c7b34f59c8ff1d3d2f427c57b7d2429f3f66c8200ca9438f14b4527e7680caf050be30c8518c77dac9814f9fefe1151f760b390f4aff62a09076c794814c018b99618d75cadedc9e43e9865db698f69d66937b65556c5e51cdeb2fb6236430ca1b9d71e0f248809f89066c6d4b38db7d13e3aa1d36825601efc7c2eb7db5c;
assign xpb_primes[30] = 1026'h9ae099be02479be649bc11e154f97cefed9f2ec182847ae9d0ba9eed45e6bc9ef76f229f515c5cc0eea1c616d4ef6e101d081348c4ea6e2f061c9267951c17ba5cd0af82a5760f2b57ced09c59e3480165c7df9fb398fa70d5c86ced15850d999b2337a86346d9dce8cce1bc8fc7855e1ad8f7ab8420c516cc48188801ea94f1;
assign xpb_primes[31] = 1026'h5b55cb7f8417aeaf3c88871282a88c8f53a8ee37ab6942b63c97d0e63f3b4b84b4ebd666be4df6d142c3748cd8363411df2fea6d5677e8bfe2a9089d67c7ffd3e58b2bb3ae9d0f21c7abfc41fb8a6c2dea5ab88b536d4915378713980d8f657c6c4a58d14b1d4923df47a41c876477a8abb8473578fb4e830be5af8c240c55cf;
assign xpb_primes[32] = 1026'h210c329225195270a1d2506fd1dbe9a39978cc4d3b2a8db4f8c96c4675c4ddfaacdb26920aceedaec66b547df9858cca6dd412d5b27553701b05517cc17305d626ee34c294f731f16e847c4bb7ce3b99804ab6a823f86569158dc0bd902cf626bcbaad6b7893e2da44f44ccee0aca7e2f9a2327401679b28420682d59f3ba4db;
assign xpb_primes[33] = 1026'h23131c3d02fc21c95e319c26bd57182a7d9ae28971cf1dea14eb7f28fcb03953dfcbb4a602c73bf20bf9f31e39f6d4c368bc49f197f9d5409fe9c78eae6aa7248404cc5a7b5354fa811911c34846dc5bccdc9966dcd849e0a222bf52d72a1f835ac5fe7826d0bffeb14459ce5e6f4137dd8982db74bce3c3733ae52def7b7aa9;
assign xpb_primes[34] = 1026'had1ec5850c25b3a80084db74185c29458636941d48e238a247cc6ed9b6acbd29b55afc6bc74cbfb59ee4f2cfe4a436522163d4d4e3c5f2a795189742976c4377d62e4b79fd26819b75d2ba1517869a16e924a4859e04cdf0bb003e422992e357df6c382cf52e51b4aa96de42a208fc808d34d6d09b7b27beaf68460df1e02c74;
assign xpb_primes[35] = 1026'h4a8c537924508ce3a4987205568d5a11c163cb3dbc84c3a9e16291c478d919bed62b6a7865209f4a43a04e4e21be90f1437ecf85f60905346966f593fd0db50c2a16afeee04fa17c3086277b6d475ee2d5231e8ddcea9a26dca3b6759f0d41bc1b1244901a08829e030448ee4767e089c7cd35594e027697ad47f5baa1efc905;
assign xpb_primes[36] = 1026'h3e5a7cfc4bde02d523bc00bef4ca492f06a4283516ba4c5f7a661ea4a666d4498d867671a871bdc57ce83a27c5692b6a087657b3f25fa31e58173e29c63c7fcd74a18258c12d31ecb55391ddf08276a976563ce70d900a826fce8f35fecd27527e88e3703c73df5cea514fe16a8f5d9ed0fad25083e8586f61be1d37bbaa1e3d;
assign xpb_primes[37] = 1026'h4cbe15bfb0ec651aff6d5e8bb97332e0721d9f680ebd5d3787802d594f0d292bac4324c3dbcab2976049b3aa1b9e15d0b12a56556b72a35db50b3b981f39001874940d725ef4bf8beacbb87c1e92170f4ed94c400809ca580c0a325ee2b12a5bc0d7879d84397f7bffff87d811ae0dcba06cedffdef20664de6cbdeddf0b8d9a;
assign xpb_primes[38] = 1026'h3502a8d6b5750b93e602aadea84a20b5247c8218c51520b649e52e0e603c2184211f77a0423f241acc45c718e4f53fac7fbf8702858d990faf68874249f6fc4887f578be7f4203358bec326f4b47c2c602174d07c8abd30cddb0c005e8ea9939f07e36b1f823354e7bc4b27dd560602cd0c28cf9043e1bb905324698c510cdc9;
assign xpb_primes[39] = 1026'h79f19bf46a901f8f8b8593b24b8509403fd5f412d387f5a45416c417af5004e923d65a7b8a9c0b73ed71f000fe39bf73fedb86ec692c33f2ebce73fa81c87305dcedf1753ff81d3cba3c6373ccbe7f011cc5f9c2dd4c17fba7e4dd816cf8a15b1553db9813e021a02d004296f433dbcea6b57ef4df14f502d6e6c8147be708b;
assign xpb_primes[40] = 1026'h20a53948e0f026bcc7b1818d7744e73ada17e1e65ea27b6d0f9dab2a63839582484c4792d33f5bba727698259867a9dc973058632d39f5caf15dc511ea43745ef0d91de5776de3beb6f8467bca21126b5957cc79e79825f2ed1016136a88da0fca3cddb58d927fe1f5fdde114c4f00832ffe01893e2432a936db9955a8d400ce;
assign xpb_primes[41] = 1026'h8ae08f142ccc140cdfcfdf28d1f6e5882da2e3829ff7b722937fd1be7fdf8891f777d19af9d4649cb65d18ae02f8c3dede63d9456388ca58d1131c3e3f4a863d2ecd194eed45b58ecf5a4a517e98b3a2fa4fa5d27ea29b6957fcf3e20ec81b44a931df26db9a6f5e35ebd77e7fcc402e942b4ea86bc4a4cfe46fa6aa87cf19a2;
assign xpb_primes[42] = 1026'h4816fede7758510c5ea226f58dcfdee19b131b68049d2cbe8293b87a0d34451e4e0cee03f2e59f495bebc981e7623f16dfef2866ede194346e329025af0c5fdba9b07703802366ed3c1c74d870c06b0ff56d5de24abbda403149ada22dc377ba5c52728b7c94958fc0be5a8c624ed9a373be98043ed863340d34b7981ef72b19;
assign xpb_primes[43] = 1026'h67b3261195678d8f14924b9881a620d60fcf7456dd3ae2228c79c9f670369d23f91b8e9bfab5a68bf2d29e831fec0653f4948f1c4a6bc7fffbde218a375aef5db7221ea3351bd53dd9605f5126b2940898717772c9c3cadbe7b7c710da8ffb61f0711193fa424b3124da7a5507d29bd366a4c0787619103ebfc59795ccebd89d;
assign xpb_primes[44] = 1026'h258aeb53f66fa3b17fef313e078be8aa1c16db1f828a53d804ece275ca21563c78cdb63df4ef81589e468cd8947a137ed9fa51841fb3ddba92b55530e9774e7772b28a673aec2956ac22666cccd6a9af47d61c31e3b8fe1136949dae0244be6503f7bbd9eb7c46d29729ba45839ab7958768c968686ce01c3986db17cc77ccd4;
assign xpb_primes[45] = 1026'ha401c40e013a6eff16974ca7c3a74ebaf451e34cea2161ffd8b475c8985a5ade3d1175ce78c6b638f74313d22c51013c39758546c7ca0ae26d5ed2652ed17f9c6fc5fd41efdb5ea6139cea41665555e89f258031f2b9a451f74e7c2de065722cfb095954956c6140a4f8e3db1d035ecc220599844925300ed3e322978aeba527;
assign xpb_primes[46] = 1026'h57ba6381570ec4025a69c77a81bdbc35e57d5271c39cd944f99b0d7465edf1ca7e6a887f24cbb4b575ba04d286dc32425b2a54788afdd4bc7d6cb3fdf582cad44d7ceed35695c248d64e5d4fe8fb3bc123dfa5cecd49410e15f67ad96cb6ffb26c54b41a24ccc91dd05d9581d43ee31ec533f7a7f502df819c931294b698a8e8;
assign xpb_primes[47] = 1026'h24489cef7dbf511d57cb02b120da8ca26786572bcec168cb19270d7efa4928ba62cb862ea0fa3e75cc2422caa92e085da3538d843f97e029b268d1f1375fa4ad792036b732dcc53ca283e2d330337e5a1ed2b8fcfe7934f1a5766feeca44564f0e703c966d4dec6ab5b8393a2367c2a697f50032772ed9234d69935524043b57;
assign xpb_primes[48] = 1026'h9f63c98ee726b34b6f70b9eab4f818bde0fa1fe5e67afe69621304c359197a15d76c94957b72ce4d950219db9f3fd657e8e356b1650c3e6fcbe0a00077134be621602277b2a3556aea4f4e34c178ce7c22e258431202ed0bfaaca4f047c6a8759221a112ddd772b7430674f15490ba9a3e7ce4b92e2955f53f18a43bd1f34f89;
assign xpb_primes[49] = 1026'h20e8cfb17397a8196917fe6ddd97be255a8ffb7cf1e9caacfd9c22829b2a1eb4a8cf3adfe1f82255adb97e181e9234e33fef5cf32c6d56661b32103287c1682daf98497e26ebe8cb7cb254f5ee5e162b8a9136516dde3457552855108db133aa301bc4b6787f62b0bff9d1ae03a9aab54c7cb384811978caf958784f6858e673;
assign xpb_primes[50] = 1026'h73089ebab524ed1e6960eb25faad4c1d827598adcee0b7a325325b6e8437cf755a91de91c191f5f07e19b2bd05013a68437d4b7993d7a40e2d67d3151dc6abde795a228c8c5d5820ae648e4e7dd6e09afa2f999304b0eaced657763c39586f167567cd154759b6faf238837e18d3418b99532f4d7e54d0d3b508f63b85c2afb6;
assign xpb_primes[51] = 1026'h5bfff2354df8aa82c37223cb4904730fe8cbf2881c8d30bb5e75f3c8cee119fd43e04cc7336bfba4874c16c7632b3a0897a675d836e70add0781e32c72502ea3711aef93feb37ec417d68868f407c55d08b0e7c4ccc6be85d410d86c81625719da51ccc27a6c794cfab5312bb2a5c03ca16280e2be5a21199961efd5aed6028c;
assign xpb_primes[52] = 1026'h30c9402da504b994e1bc13fd2101bc1221d58989ffd4cb53dc7da188568ec37547026f30c853be1722608ee4294ca7f4be4afd8324547b5ead765e15d7c76338b22660875a041441b43b5a260af3a5fff128fe947074d54eff81888aef4cbeb1130891c065df7128df8307ee35fb15aa936a835d057240291de9b0ad5cb668cc;
assign xpb_primes[53] = 1026'h1f83c8bac4d52b9137e665848ca76251159ae495d0f21b62005a400c3999942cb2ce7e8bafe3c2efd2384d825a05a6c3a52369595442bdf719edc674926d70000f078724c714660bd47d881a55ab955ec9cd48b684f4b7afda6b760f77b008c62621739435459e2e4efd22fca071f0c02669f0ea917055bd4a5b9d5041664275;
assign xpb_primes[54] = 1026'hf54d970835bdbf3ba453ed4fa8d1279b5039fca578dfc1bdca2c7277f6c5d124b4444982416afdcf99bdf642b1d648adeec2ac8936f33cfd21db06c376bf7cbc922c6ea67d00b436bc01a6e3e3ccccbb11e9e7a153fad2621ae8edd3c4fd93c7b7a305ca10c0a3d7f03da393a3183e901d8e13889fd7d67d5188a720385be4;
assign xpb_primes[55] = 1026'h9a9fc493a0d8126596b040da47ed6abfc6ac7181b5bc702d46baec3f1236652f6d8707822f389fa57c8906c915aeca8be4ce6a29aa8c4857dc63c7965b49d4fbc531307f1549ffe66c2a78d3a817565f0e0305923983c7de4dfeca29a8e8ae00d70c348133e6575cc30cd8e2e53349aa6be6e994fea886bfb81f11dd13dff33e;
assign xpb_primes[56] = 1026'h703ff39adc050c0cb27e6eea60949e792bd3ac8459ca06774553847506534996e7edb6d3b85c035ccd5e6e1a8a421840102702b2861a8ce401f91e2c14d882e651aebba47e8d3692c134881259a9d09769e7106820d151c7453b6e8005ad40a8ef8b50ae19b38592c281dab20cd9201a778aea77f3a595a4b86e2acb66e98c63;
assign xpb_primes[57] = 1026'h2b6c88b6de4d046b72169d64d5f50dc04968c544a42ad4dbf1f5f448bbb9f257702055b1eec776a185438c1928a043ed7d1431bbecf4e68b523df8689bff2ab7d632c909ec229e8f17ad81a1d8ba33ac527c778b21092016377df88dd670a88e3d9573c11cb9077b9b1265c465c74fe123264b0df7e6da4c2bc101b7926c27a7;
assign xpb_primes[58] = 1026'h150da1e2da0284690dae034f4adbe904a0ddc216f8e5c71c6db2f8123ef2a4eb843e82685b231cee3b258fb2a5a80d4d8c04f8b15934bfacd921fd222bb5059236d54dd5feaec04330a21642b7faf8b591092656b77b6d4dd4c5a66825ec916eb5c81d1c74d15c7ceca3074bdd500e1afb4d3e8778cc81926cbd9d32cd27bd23;
assign xpb_primes[59] = 1026'h98e5ba23c261d96a230567242e564b0f827f488c620d21795c419f924096c5a4b859f32979677d346b94e894e9debc9aedac8c589e520896a6ec64a96fb13b90d37ff42a950af14b54b0ac4461f3ef8b352a2249c8d2542762ee698785cb51370e55d62f742e2f0f4714cbd5937dd27df53f46b26d599e521d368fa87619b42a;
assign xpb_primes[60] = 1026'h6e6828cdd3044576e56ee6e4f4f2f4a7996efc81e7fc27717975470a87a1b4552cf8249cfe1929200790b83228122ebb3b6690d1a75c6cb408fb5d7f391c8b7ad95c5942e5da5e413cbd2b6a6fb2d7dab03b235c64cafc42f85d9fe2db712cb987ca33db66bc49d1eea978fd270f277ec1fa124debe7ae6427db80efdda409ce;
assign xpb_primes[61] = 1026'h30fb3a3e01d46807c3eb389d464bcdbc68eeb6cc7e91b308cc29f8474807235d3c8e12baddbb69b19b6ab4170e2432920fd8222f56b38bbf33fa11cc6f559a72461e86fbab80176b2c1bff224c561bb7ef5cd14d67b2a940be325edc83bf3a5255d8a71a65e9b8562626acdbd0bab538037660cebd455eef553d4637e330d04;
assign xpb_primes[62] = 1026'h162dac772cdab73c61918bef68d8e1a050f3419c8628957fb5f8c9c1dfaead7ca246492e21b98035916f8be986db4e8d003df848a132170b6d8668fee255168d063b1bc88bb69dc37ba6e920bde58fa6e2077cafbade508bc1d8913e67121bebe0b9ace5f035d546753a661ef72477fc4d599e025f4e3b66d1d2af2bc99d70cb;
assign xpb_primes[63] = 1026'h68e5391c9c125643016fc0a3c9170c956d9dfac9b9a34c4578b05e836ffea09190743f5ae4675e96939a46c3d08ce0e86b8af8b01fd1ca7e673a218fb5343b8e110c3873aa216f094e161fc0fb05a5dbf5a20c7d35a930cd0f1ac70561b5644ac8370efcc63e8a9f80ccf63c1b53fdda83931789fb317406838a48c962f5a529;

    




    // xpb Outputs
    logic [NUM_XPB-1:0][BIT_LEN_XPB-1:0] xpb0[NUM_FLAG];
    logic [NUM_XPB-1:0][BIT_LEN_XPB-1:0] xpb1[NUM_FLAG];

    genvar i;
    generate;
        for (i=0; i<NUM_FLAG; i++) begin
            xpb #(
                .BIT_LEN_FLAG ( BIT_LEN_FLAG ),
                .BIT_LEN_XPB  ( BIT_LEN_XPB ),
                .NUM_XPB      ( NUM_XPB ))
                u_xpb (
                    .flag(xpb_flag[i]),
                    .xpb_prime(xpb_primes[i]),
                    .xpb0(xpb0[i]),
                    .xpb1(xpb1[i])
                    );
        end
    endgenerate




    // row_to_col parameter
    localparam INIT_NUMS_COLS = BIT_LEN_XPB*NUM_XPB;

    // row_to_col Intputs
    logic [INIT_NUMS_COLS-1:0] u_rtc0_in[NUM_FLAG+2];
    logic [INIT_NUMS_COLS-1:0] u_rtc1_in[NUM_FLAG];

    genvar i_0;
    generate;
        for (i_0=0; i_0<NUM_FLAG+2; i_0++)begin
            if (i_0 < NUM_FLAG)begin
                assign u_rtc0_in[i_0] = xpb0[i_0];
                assign u_rtc1_in[i_0] = xpb1[i_0];
            end else if(i_0 == NUM_FLAG)begin
                assign u_rtc0_in[i_0] = rest0;
            end else begin
                assign u_rtc0_in[i_0] = rest1;
            end
        end
    endgenerate

    // row_to_col Outputs
    logic [INIT_NUMS_COLS-1:0][NUM_FLAG+1:0] u_rtc0_out;
    logic [INIT_NUMS_COLS-1:0][NUM_FLAG-1:0] u_rtc1_out;


    genvar m,n;
    generate
        for ( m = 0; m < INIT_NUMS_COLS; m = m + 1)begin
            for ( n = 0; n < NUM_FLAG+2; n = n + 1)begin
                assign u_rtc0_out[m][n] = u_rtc0_in[n][m];
                if (n < NUM_FLAG) begin
                    assign u_rtc1_out[m][n] = u_rtc1_in[n][m];
                end
            end
        end
    endgenerate

    
    
    // compressor_array_reduction Parameter
    localparam NUM_ROWS = 66;

    // compressor_array_reduction Inputs
    logic [INIT_NUMS_COLS-1:0][NUM_ROWS-1:0] cols0;
    logic [INIT_NUMS_COLS-1:0][NUM_ROWS-1:0] cols1;

    genvar j;
    generate;
        for (j=0; j<INIT_NUMS_COLS; j++) begin
            assign cols0[j] = u_rtc0_out[j];
            assign cols1[j] = {u_rtc1_out[j], 2'b0};
        end
    endgenerate

    // compressor_array_reduction Outputs

    compressor_array_reduction #(
        .BIT_LEN_FLAG     ( BIT_LEN_FLAG   ),
        .BIT_LEN_XPB      ( BIT_LEN_XPB   ),
        .NUM_XPB          ( NUM_XPB   ),
        .NUM_ROWS         ( NUM_ROWS   ),
        .INIT_NUMS_COLS   ( INIT_NUMS_COLS ),
        .NUM_ELEMENTS_OUT ( NUM_ELEMENTS_OUT ))
        u_compressor_array_reduction (
            .cols0(cols0),
            .cols1(cols1),

            .C(C),
            .S(S)
        );

    
endmodule
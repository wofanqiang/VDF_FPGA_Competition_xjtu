module xpb_5_80
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'he844837d0ffafce16d93f03b5a9a26fc4ceb5ec239a14ec47558763a8bd6737ccc2c7b389b83028d3c3071e03ce6ddee17dbe9e90cceb9461d49d254bf539fcaa42bb265cc4626f90bd323c71ead7f73831ba23df8a9167e1d70274e1c1d952be0df405f42e30520b2784eea17482f1ade9739180b702cc87219ae0a954f3b4;
    5'b00010 : xpb = 1024'h1d08906fa1ff5f9c2db27e076b5344df899d6bd8473429d88eab0ec7517ace6f99858f6713706051a7860e3c079cdbbdc2fb7d3d2199d728c3a93a4a97ea73f95485764cb988c4df217a6478e3d5afee70637447bf1522cfc3ae04e9c383b2a57c1be80be85c60a4164f09dd42e905e35bd2e723016e05990e4335c152a9e768;
    5'b00011 : xpb = 1024'h2b8cd8a772ff0f6a448bbd0b20fce74f4e6c21c46ace3ec4d600962afa3835a76648571a9d28907a7b49155a0b6b499ca4793bdbb266c2bd257dd76fe3dfadf5fec83173164d274eb23796b555c087e5a8952e6b9e9fb437a585075ea5458bf83a29dc11dc8a90f621768ecbe45d88d509bc5ab4822508659564d0a1fbfedb1c;
    5'b00100 : xpb = 1024'h3a1120df43febf385b64fc0ed6a689bf133ad7b08e6853b11d561d8ea2f59cdf330b1ece26e0c0a34f0c1c780f39b77b85f6fa7a4333ae51875274952fd4e7f2a90aec99731189be42f4c8f1c7ab5fdce0c6e88f7e2a459f875c09d38707654af837d017d0b8c1482c9e13ba85d20bc6b7a5ce4602dc0b321c866b82a553ced0;
    5'b00101 : xpb = 1024'h4895691714fe6f06723e3b128c502c2ed8098d9cb202689d64aba4f24bb30416ffcde681b098f0cc22cf23961308255a6774b918d40099e5e92711ba7bca21ef534da7bfcfd5ec2dd3b1fb2e399637d418f8a2b35db4d70769330c4868c93e9db645c41dc4e6f19a37c598a927468eb8658f41d783930dfea3a806634ea8c284;
    5'b00110 : xpb = 1024'h5719b14ee5fe1ed489177a1641f9ce9e9cd84388d59c7d89ac012c55f4706b4ecc90ae353a5120f4f6922ab416d6933948f277b764cd857a4afbaedfc7bf5bebfd9062e62c9a4e9d646f2d6aab810fcb512a5cd73d3f686f4b0a0ebd4a8b17f07453b823b91521ec42ed1d97c8bb11aa1378b569044a10cb2ac9a143f7fdb638;
    5'b00111 : xpb = 1024'h659df986b6fdcea29ff0b919f7a3710e61a6f974f9369275f356b3b99d2dd286995375e8c409511dca5531d21aa501182a703655f59a710eacd04c0513b495e8a7d31e0c895eb10cf52c5fa71d6be7c2895c16fb1cc9f9d72ce111322c4cf1433261ac29ad43523e4e14a2866a2f949bc16228fa85011397b1eb3c24a152a9ec;
    5'b01000 : xpb = 1024'h742241be87fd7e70b6c9f81dad4d137e2675af611cd0a7623aac3b1d45eb39be66163d9c4dc181469e1838f01e736ef70bedf4f486675ca30ea4e92a5fa9cfe55215d932e623137c85e991e38f56bfb9c18dd11efc548b3f0eb813a70e0eca95f06fa02fa1718290593c27750ba4178d6f4b9c8c05b81664390cd7054aa79da0;
    5'b01001 : xpb = 1024'h82a689f658fd2e3ecda3372162f6b5edeb44654d406abc4e8201c280eea8a0f632d9054fd779b16f71db400e2241dcd5ed6bb393173448377079864fab9f09e1fc58945942e775ec16a6c420014197b0f9bf8b42dbdf1ca6f08f161befd0a3e8ae7d9435959fb2e26463ac63ad189a7f1d35101d866f1930c02e71e5f3fc9154;
    5'b01010 : xpb = 1024'h912ad22e29fcde0ce47c762518a0585db0131b396404d13ac95749e49766082dff9bcd036131e198459e472c26104ab4cee97231a80133cbd24e2374f79443dea69b4f7f9fabd85ba763f65c732c6fa831f14566bb69ae0ed2661890d1927d3b6c8b883b89cde3346f8b31524e8d1d70cb1e83af07261bfd47500cc69d518508;
    5'b01011 : xpb = 1024'h9faf1a65fafc8ddafb55b528ce49facd74e1d125879ee62710acd14840236f65cc5e94b6eaea11c119614e4a29deb893b06730d038ce1f603422c09a43897ddb50de0aa5fc703acb38212898e517479f6a22ff8a9af43f76b43d1b05b354568e2a997c417dfc13867ab2b640f001a0627907f74087dd1ec9ce71a7a746a678bc;
    5'b01100 : xpb = 1024'hae33629dcbfc3da9122ef42c83f39d3d39b08711ab38fb13580258abe8e0d69d99215c6a74a241e9ed2455682dad267291e4ef6ec99b0af495f75dbf8f7eb7d7fb20c5cc59349d3ac8de5ad557021f96a254b9ae7a7ed0de96141d7a95162fe0e8a77047722a43d885da3b2f9176235426f16ad20894219655934287effb6c70;
    5'b01101 : xpb = 1024'hc0a657fdb0db8ae5e02bb592942f85b8d0939ccf95b6f88217b26b9de9b90cd629ba6a53433f38421891d3f4e1d83870f48862737b5263d472cbb86a0a17d2331144c440668026547018a6f3011335ce6817a39cd833535c25e8df4bcad66a177add223b58f7b9d0a41d93f3b1a801c8600ff8138ffc73296456264106df9b9;
    5'b01110 : xpb = 1024'h1a8eadb7ac0d687c74dbfa5cdeec9acb51d7efb91cf5847468d0ae1d8758f8052f5e6e58bdec23acf54c245d51ebf165f0c644c5c88211d1a90158abec96b71fdb57076a632c64d4d7bebcaba1fc0b541eb3345dad0dc69da43590699e6f3ff435bbc629a9bdabef15695e2ddc8f030e33ea7312b9b6c9ff1d66fd44b9c2ed6d;
    5'b01111 : xpb = 1024'h2912f5ef7d0d184a8bb5396094963d3b16a6a5a5408f9960b026358130165f3cfc21360c47a453d5c90f2b7b55ba5f44d2440364594efd660ad5f5d1388bf11c8599c290bff0c744687beee813e6e34b56e4ee818c985805860c92de80311946f3c9ba2f9debdc412090e31c7e0385ffe1d3e6a43a6dcccba48898256317e121;
    5'b10000 : xpb = 1024'h37973e274e0cc818a28e78644a3fdfaadb755b916429ae4cf77bbce4d8d3c674c8e3fdbfd15c83fe9cd232995988cd23b3c1c202ea1be8fa6caa92f684812b192fdc7db71cb529b3f939212485d1bb428f16a8a56c22e96d67e3955361f2f299b1d7ae35921a0c932bb8680b1f7808f18fbd5a35bb24cf982baa33060c6cd4d5;
    5'b10001 : xpb = 1024'h461b865f1f0c77e6b967b767ffe9821aa044117d87c3c3393ed1444881912dac95a6c5735b14b427709539b75d573b02953f80a17ae8d48ece7f301bd0766515da1f38dd79798c2389f65360f7bc9339c74862c94bad7ad549ba97c843b4cbec6fe5a23b86483ce536dfecf9c0ec8be33da6cdc73bdbd264b2cbcde6b5c1c889;
    5'b10010 : xpb = 1024'h549fce96f00c27b4d040f66bb593248a6512c769ab5dd8258626cbac2a4e94e462698d26e4cce450445840d56125a8e176bd3f400bb5c0233053cd411c6b9f128461f403d63dee931ab3859d69a76b30ff7a1ced2b380c3d2b919a3d2576a53f2df396417a766d37420771e862610ed4eb904158bc92d53139ed68c75f16bc3d;
    5'b10011 : xpb = 1024'h632416cec10bd782e71a356f6b3cc6fa29e17d55cef7ed11cd7c530fd30bfc1c2f2c54da6e851479181b47f364f416c0583afdde9c82abb792286a666860d90f2ea4af2a33025102ab70b7d9db92432837abd7110ac29da50d689cb207387e91ec018a476ea49d894d2ef6d703d591c69979b4ea3d49d7fdc10f03a8086baff1;
    5'b10100 : xpb = 1024'h71a85f06920b8750fdf3747320e66969eeb03341f29201fe14d1da737bc96353fbef1c8df83d44a1ebde4f1168c2849f39b8bc7d2d4f974bf3fd078bb456130bd8e76a508fc6b3723c2dea164d7d1b1f6fdd9134ea4d2f0cef3f9f26e8fa57e4aa0f7e4d62d2cddb58567bc5a54a14b84763287bbe00daca48309e88b1c0a3a5;
    5'b10101 : xpb = 1024'h802ca73e630b371f14ccb376d6900bd9b37ee92e162c16ea5c2761d72486ca8bc8b1e44181f574cabfa1562f6c90f27e1b367b1bbe1c82e055d1a4b1004b4d08832a2576ec8b15e1cceb1c52bf67f316a80f4b58c9d7c074d116a19bcabc3137681d72535700fe2d637e00b446be97a9f54c9c0d3eb7dd96cf5239695b159759;
    5'b10110 : xpb = 1024'h8eb0ef76340ae6ed2ba5f27a8c39ae49784d9f1a39c62bd6a37ce93acd4431c39574abf50bada4f393645d4d705f605cfcb439ba4ee96e74b7a641d64c4087052d6ce09d494f78515da84e8f3152cb0de041057ca96251dcb2eda410ac7e0a8a262b66594b2f2e7f6ea585a2e8331a9ba3360f9ebf6ee0635673d44a046a8b0d;
    5'b10111 : xpb = 1024'h9d3537ae050a96bb427f317e41e350b93d1c55065d6040c2ead2709e760198fb623773a89565d51c6727646b742dce3bde31f858dfb65a09197adefb9835c101d7af9bc3a613dac0ee6580cba33da3051872bfa088ece34494c4a6858e3fe3dce4395a5f3f5d5ed179cd0a9189a79d8d511f83304025e32fdd956f2aadbf7ec1;
    5'b11000 : xpb = 1024'habb97fe5d60a468959587081f78cf32901eb0af280fa55af3227f8021ebf00332efa3b5c1f1e05453aea6b8977fc3c1abfafb6f77083459d7b4f7c20e42afafe81f256ea02d83d307f22b30815287afc50a479c4687774ac769ba8fa7001bd2fa2474e65338b8f2384f48f802b1c207eff08f6c1c0dce5fc64b70a0b57147275;
    5'b11001 : xpb = 1024'h99082c7e51bc18ea52c37ae9cdc4e475543bdadcf1cca23fba0c6101479ba62f8748596deafb6df6f4f3360986c992f3d134dafde9d60e62c84d9e7f54dc049b7e5dd61b00ba25afd45e2a1ee378ec294d13a4fbb7bd903a2e619749798f3f0314db04176f0c6e8095c2d8fd4c07d475e188b70f1488b98a56929e77786ffbe;
    5'b11010 : xpb = 1024'h1814caffb61b715cbc0576b25285f0b71a127399f2b6df1042f64d73bd37219ac5374d4a6867e70843123a7e9c3b070e1e910c4e6f6a4c7a8e59770d4142fa46622898880cd004ca8e0314de602266b9cd02f4739b066a6b84bd1be9795acd42ef5ba4476b1ef73a1483b27e763500390c01ff0271ff8e652c8ac4c820dbf372;
    5'b11011 : xpb = 1024'h26991337871b212ad2deb5b6082f9326dee129861650f3fc8a4bd4d765f488d291fa14fdf220173116d5419ca00974ed000ecaed0037380ef02e14328d3834430c6b53ae6994673a1ec0471ad20d3eb10534ae977a90fbd366941e5e5b1ca695ad69984d5f4d278c1fab376d17a9832ab9eb7293f2b69131b3ac5fa8ca30e726;
    5'b11100 : xpb = 1024'h351d5b6f581ad0f8e9b7f4b9bdd93596a3afdf7239eb08e8d1a15c3b0eb1f00a5ebcdcb17bd84759ea9848baa3d7e2cbe18c898b910423a35202b157d92d6e3fb6ae0ed4c658c9a9af7d795743f816a83d6668bb5a1b8d3b486b20d33cde7fe86b778c53537b57de2ad2bc5bb91e061c67d4e625736d93fe3acdfa897385dada;
    5'b11101 : xpb = 1024'h43a1a3a7291a80c7009133bd7382d806687e955e5d851dd518f6e39eb76f57422b7fa46505907782be5b4fd8a7a650aac30a482a21d10f37b3d74e7d2522a83c60f0c9fb231d2c19403aab93b5e2ee9f759822df39a61ea32a4223481ea0593b2985805947a9883035fa414a5a92890e15be59b6f42496cac1ef956a1cdace8e;
    5'b11110 : xpb = 1024'h5225ebdefa1a3095176a72c1292c7a762d4d4b4a811f32c1604c6b02602cbe79f8426c188f48a7ab921e56f6ab74be89a48806c8b29dfacc15abeba27117e2390b3385217fe18e88d0f7ddd027cdc696adc9dd031930b00b0c1925bd0062328de793745f3bd7b8824121c638fc070bffc3a7cd4874db99974911304ac62fc242;
    5'b11111 : xpb = 1024'h60aa3416cb19e0632e43b1c4ded61ce5f21c0136a4b947ada7a1f26608ea25b1c50533cc1900d7d465e15e14af432c688605c567436ae660778088c7bd0d1c35b5764047dca5f0f861b5100c99b89e8de5fb9726f8bb4172edf02831e2240be0a5a168653005e8d44c494b279d7b8ef1719140d9f5929c63d032cb2b6f84b5f6;
    endcase
end

endmodule
